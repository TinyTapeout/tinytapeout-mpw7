magic
tech sky130B
magscale 1 2
timestamp 1659434107
<< obsli1 >>
rect 17104 18159 547860 681425
<< obsm1 >>
rect 2774 3408 580506 700732
<< metal2 >>
rect 8546 703520 8658 704960
rect 24738 703520 24850 704960
rect 40930 703520 41042 704960
rect 57122 703520 57234 704960
rect 73314 703520 73426 704960
rect 89506 703520 89618 704960
rect 105698 703520 105810 704960
rect 121890 703520 122002 704960
rect 138082 703520 138194 704960
rect 154274 703520 154386 704960
rect 170466 703520 170578 704960
rect 186658 703520 186770 704960
rect 202850 703520 202962 704960
rect 219042 703520 219154 704960
rect 235234 703520 235346 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300002 703520 300114 704960
rect 316194 703520 316306 704960
rect 332386 703520 332498 704960
rect 348578 703520 348690 704960
rect 364770 703520 364882 704960
rect 380962 703520 381074 704960
rect 397154 703520 397266 704960
rect 413346 703520 413458 704960
rect 429538 703520 429650 704960
rect 445730 703520 445842 704960
rect 461922 703520 462034 704960
rect 478114 703520 478226 704960
rect 494306 703520 494418 704960
rect 510498 703520 510610 704960
rect 526690 703520 526802 704960
rect 542882 703520 542994 704960
rect 559074 703520 559186 704960
rect 575266 703520 575378 704960
rect 19770 -960 19882 480
rect 20874 -960 20986 480
rect 21978 -960 22090 480
rect 23082 -960 23194 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26394 -960 26506 480
rect 27498 -960 27610 480
rect 28602 -960 28714 480
rect 29706 -960 29818 480
rect 30810 -960 30922 480
rect 31914 -960 32026 480
rect 33018 -960 33130 480
rect 34122 -960 34234 480
rect 35226 -960 35338 480
rect 36330 -960 36442 480
rect 37434 -960 37546 480
rect 38538 -960 38650 480
rect 39642 -960 39754 480
rect 40746 -960 40858 480
rect 41850 -960 41962 480
rect 42954 -960 43066 480
rect 44058 -960 44170 480
rect 45162 -960 45274 480
rect 46266 -960 46378 480
rect 47370 -960 47482 480
rect 48474 -960 48586 480
rect 49578 -960 49690 480
rect 50682 -960 50794 480
rect 51786 -960 51898 480
rect 52890 -960 53002 480
rect 53994 -960 54106 480
rect 55098 -960 55210 480
rect 56202 -960 56314 480
rect 57306 -960 57418 480
rect 58410 -960 58522 480
rect 59514 -960 59626 480
rect 60618 -960 60730 480
rect 61722 -960 61834 480
rect 62826 -960 62938 480
rect 63930 -960 64042 480
rect 65034 -960 65146 480
rect 66138 -960 66250 480
rect 67242 -960 67354 480
rect 68346 -960 68458 480
rect 69450 -960 69562 480
rect 70554 -960 70666 480
rect 71658 -960 71770 480
rect 72762 -960 72874 480
rect 73866 -960 73978 480
rect 74970 -960 75082 480
rect 76074 -960 76186 480
rect 77178 -960 77290 480
rect 78282 -960 78394 480
rect 79386 -960 79498 480
rect 80490 -960 80602 480
rect 81594 -960 81706 480
rect 82698 -960 82810 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86010 -960 86122 480
rect 87114 -960 87226 480
rect 88218 -960 88330 480
rect 89322 -960 89434 480
rect 90426 -960 90538 480
rect 91530 -960 91642 480
rect 92634 -960 92746 480
rect 93738 -960 93850 480
rect 94842 -960 94954 480
rect 95946 -960 96058 480
rect 97050 -960 97162 480
rect 98154 -960 98266 480
rect 99258 -960 99370 480
rect 100362 -960 100474 480
rect 101466 -960 101578 480
rect 102570 -960 102682 480
rect 103674 -960 103786 480
rect 104778 -960 104890 480
rect 105882 -960 105994 480
rect 106986 -960 107098 480
rect 108090 -960 108202 480
rect 109194 -960 109306 480
rect 110298 -960 110410 480
rect 111402 -960 111514 480
rect 112506 -960 112618 480
rect 113610 -960 113722 480
rect 114714 -960 114826 480
rect 115818 -960 115930 480
rect 116922 -960 117034 480
rect 118026 -960 118138 480
rect 119130 -960 119242 480
rect 120234 -960 120346 480
rect 121338 -960 121450 480
rect 122442 -960 122554 480
rect 123546 -960 123658 480
rect 124650 -960 124762 480
rect 125754 -960 125866 480
rect 126858 -960 126970 480
rect 127962 -960 128074 480
rect 129066 -960 129178 480
rect 130170 -960 130282 480
rect 131274 -960 131386 480
rect 132378 -960 132490 480
rect 133482 -960 133594 480
rect 134586 -960 134698 480
rect 135690 -960 135802 480
rect 136794 -960 136906 480
rect 137898 -960 138010 480
rect 139002 -960 139114 480
rect 140106 -960 140218 480
rect 141210 -960 141322 480
rect 142314 -960 142426 480
rect 143418 -960 143530 480
rect 144522 -960 144634 480
rect 145626 -960 145738 480
rect 146730 -960 146842 480
rect 147834 -960 147946 480
rect 148938 -960 149050 480
rect 150042 -960 150154 480
rect 151146 -960 151258 480
rect 152250 -960 152362 480
rect 153354 -960 153466 480
rect 154458 -960 154570 480
rect 155562 -960 155674 480
rect 156666 -960 156778 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 159978 -960 160090 480
rect 161082 -960 161194 480
rect 162186 -960 162298 480
rect 163290 -960 163402 480
rect 164394 -960 164506 480
rect 165498 -960 165610 480
rect 166602 -960 166714 480
rect 167706 -960 167818 480
rect 168810 -960 168922 480
rect 169914 -960 170026 480
rect 171018 -960 171130 480
rect 172122 -960 172234 480
rect 173226 -960 173338 480
rect 174330 -960 174442 480
rect 175434 -960 175546 480
rect 176538 -960 176650 480
rect 177642 -960 177754 480
rect 178746 -960 178858 480
rect 179850 -960 179962 480
rect 180954 -960 181066 480
rect 182058 -960 182170 480
rect 183162 -960 183274 480
rect 184266 -960 184378 480
rect 185370 -960 185482 480
rect 186474 -960 186586 480
rect 187578 -960 187690 480
rect 188682 -960 188794 480
rect 189786 -960 189898 480
rect 190890 -960 191002 480
rect 191994 -960 192106 480
rect 193098 -960 193210 480
rect 194202 -960 194314 480
rect 195306 -960 195418 480
rect 196410 -960 196522 480
rect 197514 -960 197626 480
rect 198618 -960 198730 480
rect 199722 -960 199834 480
rect 200826 -960 200938 480
rect 201930 -960 202042 480
rect 203034 -960 203146 480
rect 204138 -960 204250 480
rect 205242 -960 205354 480
rect 206346 -960 206458 480
rect 207450 -960 207562 480
rect 208554 -960 208666 480
rect 209658 -960 209770 480
rect 210762 -960 210874 480
rect 211866 -960 211978 480
rect 212970 -960 213082 480
rect 214074 -960 214186 480
rect 215178 -960 215290 480
rect 216282 -960 216394 480
rect 217386 -960 217498 480
rect 218490 -960 218602 480
rect 219594 -960 219706 480
rect 220698 -960 220810 480
rect 221802 -960 221914 480
rect 222906 -960 223018 480
rect 224010 -960 224122 480
rect 225114 -960 225226 480
rect 226218 -960 226330 480
rect 227322 -960 227434 480
rect 228426 -960 228538 480
rect 229530 -960 229642 480
rect 230634 -960 230746 480
rect 231738 -960 231850 480
rect 232842 -960 232954 480
rect 233946 -960 234058 480
rect 235050 -960 235162 480
rect 236154 -960 236266 480
rect 237258 -960 237370 480
rect 238362 -960 238474 480
rect 239466 -960 239578 480
rect 240570 -960 240682 480
rect 241674 -960 241786 480
rect 242778 -960 242890 480
rect 243882 -960 243994 480
rect 244986 -960 245098 480
rect 246090 -960 246202 480
rect 247194 -960 247306 480
rect 248298 -960 248410 480
rect 249402 -960 249514 480
rect 250506 -960 250618 480
rect 251610 -960 251722 480
rect 252714 -960 252826 480
rect 253818 -960 253930 480
rect 254922 -960 255034 480
rect 256026 -960 256138 480
rect 257130 -960 257242 480
rect 258234 -960 258346 480
rect 259338 -960 259450 480
rect 260442 -960 260554 480
rect 261546 -960 261658 480
rect 262650 -960 262762 480
rect 263754 -960 263866 480
rect 264858 -960 264970 480
rect 265962 -960 266074 480
rect 267066 -960 267178 480
rect 268170 -960 268282 480
rect 269274 -960 269386 480
rect 270378 -960 270490 480
rect 271482 -960 271594 480
rect 272586 -960 272698 480
rect 273690 -960 273802 480
rect 274794 -960 274906 480
rect 275898 -960 276010 480
rect 277002 -960 277114 480
rect 278106 -960 278218 480
rect 279210 -960 279322 480
rect 280314 -960 280426 480
rect 281418 -960 281530 480
rect 282522 -960 282634 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285834 -960 285946 480
rect 286938 -960 287050 480
rect 288042 -960 288154 480
rect 289146 -960 289258 480
rect 290250 -960 290362 480
rect 291354 -960 291466 480
rect 292458 -960 292570 480
rect 293562 -960 293674 480
rect 294666 -960 294778 480
rect 295770 -960 295882 480
rect 296874 -960 296986 480
rect 297978 -960 298090 480
rect 299082 -960 299194 480
rect 300186 -960 300298 480
rect 301290 -960 301402 480
rect 302394 -960 302506 480
rect 303498 -960 303610 480
rect 304602 -960 304714 480
rect 305706 -960 305818 480
rect 306810 -960 306922 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310122 -960 310234 480
rect 311226 -960 311338 480
rect 312330 -960 312442 480
rect 313434 -960 313546 480
rect 314538 -960 314650 480
rect 315642 -960 315754 480
rect 316746 -960 316858 480
rect 317850 -960 317962 480
rect 318954 -960 319066 480
rect 320058 -960 320170 480
rect 321162 -960 321274 480
rect 322266 -960 322378 480
rect 323370 -960 323482 480
rect 324474 -960 324586 480
rect 325578 -960 325690 480
rect 326682 -960 326794 480
rect 327786 -960 327898 480
rect 328890 -960 329002 480
rect 329994 -960 330106 480
rect 331098 -960 331210 480
rect 332202 -960 332314 480
rect 333306 -960 333418 480
rect 334410 -960 334522 480
rect 335514 -960 335626 480
rect 336618 -960 336730 480
rect 337722 -960 337834 480
rect 338826 -960 338938 480
rect 339930 -960 340042 480
rect 341034 -960 341146 480
rect 342138 -960 342250 480
rect 343242 -960 343354 480
rect 344346 -960 344458 480
rect 345450 -960 345562 480
rect 346554 -960 346666 480
rect 347658 -960 347770 480
rect 348762 -960 348874 480
rect 349866 -960 349978 480
rect 350970 -960 351082 480
rect 352074 -960 352186 480
rect 353178 -960 353290 480
rect 354282 -960 354394 480
rect 355386 -960 355498 480
rect 356490 -960 356602 480
rect 357594 -960 357706 480
rect 358698 -960 358810 480
rect 359802 -960 359914 480
rect 360906 -960 361018 480
rect 362010 -960 362122 480
rect 363114 -960 363226 480
rect 364218 -960 364330 480
rect 365322 -960 365434 480
rect 366426 -960 366538 480
rect 367530 -960 367642 480
rect 368634 -960 368746 480
rect 369738 -960 369850 480
rect 370842 -960 370954 480
rect 371946 -960 372058 480
rect 373050 -960 373162 480
rect 374154 -960 374266 480
rect 375258 -960 375370 480
rect 376362 -960 376474 480
rect 377466 -960 377578 480
rect 378570 -960 378682 480
rect 379674 -960 379786 480
rect 380778 -960 380890 480
rect 381882 -960 381994 480
rect 382986 -960 383098 480
rect 384090 -960 384202 480
rect 385194 -960 385306 480
rect 386298 -960 386410 480
rect 387402 -960 387514 480
rect 388506 -960 388618 480
rect 389610 -960 389722 480
rect 390714 -960 390826 480
rect 391818 -960 391930 480
rect 392922 -960 393034 480
rect 394026 -960 394138 480
rect 395130 -960 395242 480
rect 396234 -960 396346 480
rect 397338 -960 397450 480
rect 398442 -960 398554 480
rect 399546 -960 399658 480
rect 400650 -960 400762 480
rect 401754 -960 401866 480
rect 402858 -960 402970 480
rect 403962 -960 404074 480
rect 405066 -960 405178 480
rect 406170 -960 406282 480
rect 407274 -960 407386 480
rect 408378 -960 408490 480
rect 409482 -960 409594 480
rect 410586 -960 410698 480
rect 411690 -960 411802 480
rect 412794 -960 412906 480
rect 413898 -960 414010 480
rect 415002 -960 415114 480
rect 416106 -960 416218 480
rect 417210 -960 417322 480
rect 418314 -960 418426 480
rect 419418 -960 419530 480
rect 420522 -960 420634 480
rect 421626 -960 421738 480
rect 422730 -960 422842 480
rect 423834 -960 423946 480
rect 424938 -960 425050 480
rect 426042 -960 426154 480
rect 427146 -960 427258 480
rect 428250 -960 428362 480
rect 429354 -960 429466 480
rect 430458 -960 430570 480
rect 431562 -960 431674 480
rect 432666 -960 432778 480
rect 433770 -960 433882 480
rect 434874 -960 434986 480
rect 435978 -960 436090 480
rect 437082 -960 437194 480
rect 438186 -960 438298 480
rect 439290 -960 439402 480
rect 440394 -960 440506 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443706 -960 443818 480
rect 444810 -960 444922 480
rect 445914 -960 446026 480
rect 447018 -960 447130 480
rect 448122 -960 448234 480
rect 449226 -960 449338 480
rect 450330 -960 450442 480
rect 451434 -960 451546 480
rect 452538 -960 452650 480
rect 453642 -960 453754 480
rect 454746 -960 454858 480
rect 455850 -960 455962 480
rect 456954 -960 457066 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460266 -960 460378 480
rect 461370 -960 461482 480
rect 462474 -960 462586 480
rect 463578 -960 463690 480
rect 464682 -960 464794 480
rect 465786 -960 465898 480
rect 466890 -960 467002 480
rect 467994 -960 468106 480
rect 469098 -960 469210 480
rect 470202 -960 470314 480
rect 471306 -960 471418 480
rect 472410 -960 472522 480
rect 473514 -960 473626 480
rect 474618 -960 474730 480
rect 475722 -960 475834 480
rect 476826 -960 476938 480
rect 477930 -960 478042 480
rect 479034 -960 479146 480
rect 480138 -960 480250 480
rect 481242 -960 481354 480
rect 482346 -960 482458 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485658 -960 485770 480
rect 486762 -960 486874 480
rect 487866 -960 487978 480
rect 488970 -960 489082 480
rect 490074 -960 490186 480
rect 491178 -960 491290 480
rect 492282 -960 492394 480
rect 493386 -960 493498 480
rect 494490 -960 494602 480
rect 495594 -960 495706 480
rect 496698 -960 496810 480
rect 497802 -960 497914 480
rect 498906 -960 499018 480
rect 500010 -960 500122 480
rect 501114 -960 501226 480
rect 502218 -960 502330 480
rect 503322 -960 503434 480
rect 504426 -960 504538 480
rect 505530 -960 505642 480
rect 506634 -960 506746 480
rect 507738 -960 507850 480
rect 508842 -960 508954 480
rect 509946 -960 510058 480
rect 511050 -960 511162 480
rect 512154 -960 512266 480
rect 513258 -960 513370 480
rect 514362 -960 514474 480
rect 515466 -960 515578 480
rect 516570 -960 516682 480
rect 517674 -960 517786 480
rect 518778 -960 518890 480
rect 519882 -960 519994 480
rect 520986 -960 521098 480
rect 522090 -960 522202 480
rect 523194 -960 523306 480
rect 524298 -960 524410 480
rect 525402 -960 525514 480
rect 526506 -960 526618 480
rect 527610 -960 527722 480
rect 528714 -960 528826 480
rect 529818 -960 529930 480
rect 530922 -960 531034 480
rect 532026 -960 532138 480
rect 533130 -960 533242 480
rect 534234 -960 534346 480
rect 535338 -960 535450 480
rect 536442 -960 536554 480
rect 537546 -960 537658 480
rect 538650 -960 538762 480
rect 539754 -960 539866 480
rect 540858 -960 540970 480
rect 541962 -960 542074 480
rect 543066 -960 543178 480
rect 544170 -960 544282 480
rect 545274 -960 545386 480
rect 546378 -960 546490 480
rect 547482 -960 547594 480
rect 548586 -960 548698 480
rect 549690 -960 549802 480
rect 550794 -960 550906 480
rect 551898 -960 552010 480
rect 553002 -960 553114 480
rect 554106 -960 554218 480
rect 555210 -960 555322 480
rect 556314 -960 556426 480
rect 557418 -960 557530 480
rect 558522 -960 558634 480
rect 559626 -960 559738 480
rect 560730 -960 560842 480
rect 561834 -960 561946 480
rect 562938 -960 563050 480
rect 564042 -960 564154 480
<< obsm2 >>
rect 2778 703464 8490 703520
rect 8714 703464 24682 703520
rect 24906 703464 40874 703520
rect 41098 703464 57066 703520
rect 57290 703464 73258 703520
rect 73482 703464 89450 703520
rect 89674 703464 105642 703520
rect 105866 703464 121834 703520
rect 122058 703464 138026 703520
rect 138250 703464 154218 703520
rect 154442 703464 170410 703520
rect 170634 703464 186602 703520
rect 186826 703464 202794 703520
rect 203018 703464 218986 703520
rect 219210 703464 235178 703520
rect 235402 703464 251370 703520
rect 251594 703464 267562 703520
rect 267786 703464 283754 703520
rect 283978 703464 299946 703520
rect 300170 703464 316138 703520
rect 316362 703464 332330 703520
rect 332554 703464 348522 703520
rect 348746 703464 364714 703520
rect 364938 703464 380906 703520
rect 381130 703464 397098 703520
rect 397322 703464 413290 703520
rect 413514 703464 429482 703520
rect 429706 703464 445674 703520
rect 445898 703464 461866 703520
rect 462090 703464 478058 703520
rect 478282 703464 494250 703520
rect 494474 703464 510442 703520
rect 510666 703464 526634 703520
rect 526858 703464 542826 703520
rect 543050 703464 559018 703520
rect 559242 703464 575210 703520
rect 575434 703464 580502 703520
rect 2778 536 580502 703464
rect 2778 480 19714 536
rect 19938 480 20818 536
rect 21042 480 21922 536
rect 22146 480 23026 536
rect 23250 480 24130 536
rect 24354 480 25234 536
rect 25458 480 26338 536
rect 26562 480 27442 536
rect 27666 480 28546 536
rect 28770 480 29650 536
rect 29874 480 30754 536
rect 30978 480 31858 536
rect 32082 480 32962 536
rect 33186 480 34066 536
rect 34290 480 35170 536
rect 35394 480 36274 536
rect 36498 480 37378 536
rect 37602 480 38482 536
rect 38706 480 39586 536
rect 39810 480 40690 536
rect 40914 480 41794 536
rect 42018 480 42898 536
rect 43122 480 44002 536
rect 44226 480 45106 536
rect 45330 480 46210 536
rect 46434 480 47314 536
rect 47538 480 48418 536
rect 48642 480 49522 536
rect 49746 480 50626 536
rect 50850 480 51730 536
rect 51954 480 52834 536
rect 53058 480 53938 536
rect 54162 480 55042 536
rect 55266 480 56146 536
rect 56370 480 57250 536
rect 57474 480 58354 536
rect 58578 480 59458 536
rect 59682 480 60562 536
rect 60786 480 61666 536
rect 61890 480 62770 536
rect 62994 480 63874 536
rect 64098 480 64978 536
rect 65202 480 66082 536
rect 66306 480 67186 536
rect 67410 480 68290 536
rect 68514 480 69394 536
rect 69618 480 70498 536
rect 70722 480 71602 536
rect 71826 480 72706 536
rect 72930 480 73810 536
rect 74034 480 74914 536
rect 75138 480 76018 536
rect 76242 480 77122 536
rect 77346 480 78226 536
rect 78450 480 79330 536
rect 79554 480 80434 536
rect 80658 480 81538 536
rect 81762 480 82642 536
rect 82866 480 83746 536
rect 83970 480 84850 536
rect 85074 480 85954 536
rect 86178 480 87058 536
rect 87282 480 88162 536
rect 88386 480 89266 536
rect 89490 480 90370 536
rect 90594 480 91474 536
rect 91698 480 92578 536
rect 92802 480 93682 536
rect 93906 480 94786 536
rect 95010 480 95890 536
rect 96114 480 96994 536
rect 97218 480 98098 536
rect 98322 480 99202 536
rect 99426 480 100306 536
rect 100530 480 101410 536
rect 101634 480 102514 536
rect 102738 480 103618 536
rect 103842 480 104722 536
rect 104946 480 105826 536
rect 106050 480 106930 536
rect 107154 480 108034 536
rect 108258 480 109138 536
rect 109362 480 110242 536
rect 110466 480 111346 536
rect 111570 480 112450 536
rect 112674 480 113554 536
rect 113778 480 114658 536
rect 114882 480 115762 536
rect 115986 480 116866 536
rect 117090 480 117970 536
rect 118194 480 119074 536
rect 119298 480 120178 536
rect 120402 480 121282 536
rect 121506 480 122386 536
rect 122610 480 123490 536
rect 123714 480 124594 536
rect 124818 480 125698 536
rect 125922 480 126802 536
rect 127026 480 127906 536
rect 128130 480 129010 536
rect 129234 480 130114 536
rect 130338 480 131218 536
rect 131442 480 132322 536
rect 132546 480 133426 536
rect 133650 480 134530 536
rect 134754 480 135634 536
rect 135858 480 136738 536
rect 136962 480 137842 536
rect 138066 480 138946 536
rect 139170 480 140050 536
rect 140274 480 141154 536
rect 141378 480 142258 536
rect 142482 480 143362 536
rect 143586 480 144466 536
rect 144690 480 145570 536
rect 145794 480 146674 536
rect 146898 480 147778 536
rect 148002 480 148882 536
rect 149106 480 149986 536
rect 150210 480 151090 536
rect 151314 480 152194 536
rect 152418 480 153298 536
rect 153522 480 154402 536
rect 154626 480 155506 536
rect 155730 480 156610 536
rect 156834 480 157714 536
rect 157938 480 158818 536
rect 159042 480 159922 536
rect 160146 480 161026 536
rect 161250 480 162130 536
rect 162354 480 163234 536
rect 163458 480 164338 536
rect 164562 480 165442 536
rect 165666 480 166546 536
rect 166770 480 167650 536
rect 167874 480 168754 536
rect 168978 480 169858 536
rect 170082 480 170962 536
rect 171186 480 172066 536
rect 172290 480 173170 536
rect 173394 480 174274 536
rect 174498 480 175378 536
rect 175602 480 176482 536
rect 176706 480 177586 536
rect 177810 480 178690 536
rect 178914 480 179794 536
rect 180018 480 180898 536
rect 181122 480 182002 536
rect 182226 480 183106 536
rect 183330 480 184210 536
rect 184434 480 185314 536
rect 185538 480 186418 536
rect 186642 480 187522 536
rect 187746 480 188626 536
rect 188850 480 189730 536
rect 189954 480 190834 536
rect 191058 480 191938 536
rect 192162 480 193042 536
rect 193266 480 194146 536
rect 194370 480 195250 536
rect 195474 480 196354 536
rect 196578 480 197458 536
rect 197682 480 198562 536
rect 198786 480 199666 536
rect 199890 480 200770 536
rect 200994 480 201874 536
rect 202098 480 202978 536
rect 203202 480 204082 536
rect 204306 480 205186 536
rect 205410 480 206290 536
rect 206514 480 207394 536
rect 207618 480 208498 536
rect 208722 480 209602 536
rect 209826 480 210706 536
rect 210930 480 211810 536
rect 212034 480 212914 536
rect 213138 480 214018 536
rect 214242 480 215122 536
rect 215346 480 216226 536
rect 216450 480 217330 536
rect 217554 480 218434 536
rect 218658 480 219538 536
rect 219762 480 220642 536
rect 220866 480 221746 536
rect 221970 480 222850 536
rect 223074 480 223954 536
rect 224178 480 225058 536
rect 225282 480 226162 536
rect 226386 480 227266 536
rect 227490 480 228370 536
rect 228594 480 229474 536
rect 229698 480 230578 536
rect 230802 480 231682 536
rect 231906 480 232786 536
rect 233010 480 233890 536
rect 234114 480 234994 536
rect 235218 480 236098 536
rect 236322 480 237202 536
rect 237426 480 238306 536
rect 238530 480 239410 536
rect 239634 480 240514 536
rect 240738 480 241618 536
rect 241842 480 242722 536
rect 242946 480 243826 536
rect 244050 480 244930 536
rect 245154 480 246034 536
rect 246258 480 247138 536
rect 247362 480 248242 536
rect 248466 480 249346 536
rect 249570 480 250450 536
rect 250674 480 251554 536
rect 251778 480 252658 536
rect 252882 480 253762 536
rect 253986 480 254866 536
rect 255090 480 255970 536
rect 256194 480 257074 536
rect 257298 480 258178 536
rect 258402 480 259282 536
rect 259506 480 260386 536
rect 260610 480 261490 536
rect 261714 480 262594 536
rect 262818 480 263698 536
rect 263922 480 264802 536
rect 265026 480 265906 536
rect 266130 480 267010 536
rect 267234 480 268114 536
rect 268338 480 269218 536
rect 269442 480 270322 536
rect 270546 480 271426 536
rect 271650 480 272530 536
rect 272754 480 273634 536
rect 273858 480 274738 536
rect 274962 480 275842 536
rect 276066 480 276946 536
rect 277170 480 278050 536
rect 278274 480 279154 536
rect 279378 480 280258 536
rect 280482 480 281362 536
rect 281586 480 282466 536
rect 282690 480 283570 536
rect 283794 480 284674 536
rect 284898 480 285778 536
rect 286002 480 286882 536
rect 287106 480 287986 536
rect 288210 480 289090 536
rect 289314 480 290194 536
rect 290418 480 291298 536
rect 291522 480 292402 536
rect 292626 480 293506 536
rect 293730 480 294610 536
rect 294834 480 295714 536
rect 295938 480 296818 536
rect 297042 480 297922 536
rect 298146 480 299026 536
rect 299250 480 300130 536
rect 300354 480 301234 536
rect 301458 480 302338 536
rect 302562 480 303442 536
rect 303666 480 304546 536
rect 304770 480 305650 536
rect 305874 480 306754 536
rect 306978 480 307858 536
rect 308082 480 308962 536
rect 309186 480 310066 536
rect 310290 480 311170 536
rect 311394 480 312274 536
rect 312498 480 313378 536
rect 313602 480 314482 536
rect 314706 480 315586 536
rect 315810 480 316690 536
rect 316914 480 317794 536
rect 318018 480 318898 536
rect 319122 480 320002 536
rect 320226 480 321106 536
rect 321330 480 322210 536
rect 322434 480 323314 536
rect 323538 480 324418 536
rect 324642 480 325522 536
rect 325746 480 326626 536
rect 326850 480 327730 536
rect 327954 480 328834 536
rect 329058 480 329938 536
rect 330162 480 331042 536
rect 331266 480 332146 536
rect 332370 480 333250 536
rect 333474 480 334354 536
rect 334578 480 335458 536
rect 335682 480 336562 536
rect 336786 480 337666 536
rect 337890 480 338770 536
rect 338994 480 339874 536
rect 340098 480 340978 536
rect 341202 480 342082 536
rect 342306 480 343186 536
rect 343410 480 344290 536
rect 344514 480 345394 536
rect 345618 480 346498 536
rect 346722 480 347602 536
rect 347826 480 348706 536
rect 348930 480 349810 536
rect 350034 480 350914 536
rect 351138 480 352018 536
rect 352242 480 353122 536
rect 353346 480 354226 536
rect 354450 480 355330 536
rect 355554 480 356434 536
rect 356658 480 357538 536
rect 357762 480 358642 536
rect 358866 480 359746 536
rect 359970 480 360850 536
rect 361074 480 361954 536
rect 362178 480 363058 536
rect 363282 480 364162 536
rect 364386 480 365266 536
rect 365490 480 366370 536
rect 366594 480 367474 536
rect 367698 480 368578 536
rect 368802 480 369682 536
rect 369906 480 370786 536
rect 371010 480 371890 536
rect 372114 480 372994 536
rect 373218 480 374098 536
rect 374322 480 375202 536
rect 375426 480 376306 536
rect 376530 480 377410 536
rect 377634 480 378514 536
rect 378738 480 379618 536
rect 379842 480 380722 536
rect 380946 480 381826 536
rect 382050 480 382930 536
rect 383154 480 384034 536
rect 384258 480 385138 536
rect 385362 480 386242 536
rect 386466 480 387346 536
rect 387570 480 388450 536
rect 388674 480 389554 536
rect 389778 480 390658 536
rect 390882 480 391762 536
rect 391986 480 392866 536
rect 393090 480 393970 536
rect 394194 480 395074 536
rect 395298 480 396178 536
rect 396402 480 397282 536
rect 397506 480 398386 536
rect 398610 480 399490 536
rect 399714 480 400594 536
rect 400818 480 401698 536
rect 401922 480 402802 536
rect 403026 480 403906 536
rect 404130 480 405010 536
rect 405234 480 406114 536
rect 406338 480 407218 536
rect 407442 480 408322 536
rect 408546 480 409426 536
rect 409650 480 410530 536
rect 410754 480 411634 536
rect 411858 480 412738 536
rect 412962 480 413842 536
rect 414066 480 414946 536
rect 415170 480 416050 536
rect 416274 480 417154 536
rect 417378 480 418258 536
rect 418482 480 419362 536
rect 419586 480 420466 536
rect 420690 480 421570 536
rect 421794 480 422674 536
rect 422898 480 423778 536
rect 424002 480 424882 536
rect 425106 480 425986 536
rect 426210 480 427090 536
rect 427314 480 428194 536
rect 428418 480 429298 536
rect 429522 480 430402 536
rect 430626 480 431506 536
rect 431730 480 432610 536
rect 432834 480 433714 536
rect 433938 480 434818 536
rect 435042 480 435922 536
rect 436146 480 437026 536
rect 437250 480 438130 536
rect 438354 480 439234 536
rect 439458 480 440338 536
rect 440562 480 441442 536
rect 441666 480 442546 536
rect 442770 480 443650 536
rect 443874 480 444754 536
rect 444978 480 445858 536
rect 446082 480 446962 536
rect 447186 480 448066 536
rect 448290 480 449170 536
rect 449394 480 450274 536
rect 450498 480 451378 536
rect 451602 480 452482 536
rect 452706 480 453586 536
rect 453810 480 454690 536
rect 454914 480 455794 536
rect 456018 480 456898 536
rect 457122 480 458002 536
rect 458226 480 459106 536
rect 459330 480 460210 536
rect 460434 480 461314 536
rect 461538 480 462418 536
rect 462642 480 463522 536
rect 463746 480 464626 536
rect 464850 480 465730 536
rect 465954 480 466834 536
rect 467058 480 467938 536
rect 468162 480 469042 536
rect 469266 480 470146 536
rect 470370 480 471250 536
rect 471474 480 472354 536
rect 472578 480 473458 536
rect 473682 480 474562 536
rect 474786 480 475666 536
rect 475890 480 476770 536
rect 476994 480 477874 536
rect 478098 480 478978 536
rect 479202 480 480082 536
rect 480306 480 481186 536
rect 481410 480 482290 536
rect 482514 480 483394 536
rect 483618 480 484498 536
rect 484722 480 485602 536
rect 485826 480 486706 536
rect 486930 480 487810 536
rect 488034 480 488914 536
rect 489138 480 490018 536
rect 490242 480 491122 536
rect 491346 480 492226 536
rect 492450 480 493330 536
rect 493554 480 494434 536
rect 494658 480 495538 536
rect 495762 480 496642 536
rect 496866 480 497746 536
rect 497970 480 498850 536
rect 499074 480 499954 536
rect 500178 480 501058 536
rect 501282 480 502162 536
rect 502386 480 503266 536
rect 503490 480 504370 536
rect 504594 480 505474 536
rect 505698 480 506578 536
rect 506802 480 507682 536
rect 507906 480 508786 536
rect 509010 480 509890 536
rect 510114 480 510994 536
rect 511218 480 512098 536
rect 512322 480 513202 536
rect 513426 480 514306 536
rect 514530 480 515410 536
rect 515634 480 516514 536
rect 516738 480 517618 536
rect 517842 480 518722 536
rect 518946 480 519826 536
rect 520050 480 520930 536
rect 521154 480 522034 536
rect 522258 480 523138 536
rect 523362 480 524242 536
rect 524466 480 525346 536
rect 525570 480 526450 536
rect 526674 480 527554 536
rect 527778 480 528658 536
rect 528882 480 529762 536
rect 529986 480 530866 536
rect 531090 480 531970 536
rect 532194 480 533074 536
rect 533298 480 534178 536
rect 534402 480 535282 536
rect 535506 480 536386 536
rect 536610 480 537490 536
rect 537714 480 538594 536
rect 538818 480 539698 536
rect 539922 480 540802 536
rect 541026 480 541906 536
rect 542130 480 543010 536
rect 543234 480 544114 536
rect 544338 480 545218 536
rect 545442 480 546322 536
rect 546546 480 547426 536
rect 547650 480 548530 536
rect 548754 480 549634 536
rect 549858 480 550738 536
rect 550962 480 551842 536
rect 552066 480 552946 536
rect 553170 480 554050 536
rect 554274 480 555154 536
rect 555378 480 556258 536
rect 556482 480 557362 536
rect 557586 480 558466 536
rect 558690 480 559570 536
rect 559794 480 560674 536
rect 560898 480 561778 536
rect 562002 480 562882 536
rect 563106 480 563986 536
rect 564210 480 580502 536
<< metal3 >>
rect 583520 694772 584960 695012
rect -960 694228 480 694468
rect 583520 681580 584960 681820
rect -960 681308 480 681548
rect -960 668388 480 668628
rect 583520 668388 584960 668628
rect -960 655468 480 655708
rect 583520 655196 584960 655436
rect -960 642548 480 642788
rect 583520 642004 584960 642244
rect -960 629628 480 629868
rect 583520 628812 584960 629052
rect -960 616708 480 616948
rect 583520 615620 584960 615860
rect -960 603788 480 604028
rect 583520 602428 584960 602668
rect -960 590868 480 591108
rect 583520 589236 584960 589476
rect -960 577948 480 578188
rect 583520 576044 584960 576284
rect -960 565028 480 565268
rect 583520 562852 584960 563092
rect -960 552108 480 552348
rect 583520 549660 584960 549900
rect -960 539188 480 539428
rect 583520 536468 584960 536708
rect -960 526268 480 526508
rect 583520 523276 584960 523516
rect -960 513348 480 513588
rect 583520 510084 584960 510324
rect -960 500428 480 500668
rect 583520 496892 584960 497132
rect -960 487508 480 487748
rect 583520 483700 584960 483940
rect -960 474588 480 474828
rect 583520 470508 584960 470748
rect -960 461668 480 461908
rect 583520 457316 584960 457556
rect -960 448748 480 448988
rect 583520 444124 584960 444364
rect -960 435828 480 436068
rect 583520 430932 584960 431172
rect -960 422908 480 423148
rect 583520 417740 584960 417980
rect -960 409988 480 410228
rect 583520 404548 584960 404788
rect -960 397068 480 397308
rect 583520 391356 584960 391596
rect -960 384148 480 384388
rect 583520 378164 584960 378404
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345388 480 345628
rect 583520 338588 584960 338828
rect -960 332468 480 332708
rect 583520 325396 584960 325636
rect -960 319548 480 319788
rect 583520 312204 584960 312444
rect -960 306628 480 306868
rect 583520 299012 584960 299252
rect -960 293708 480 293948
rect 583520 285820 584960 286060
rect -960 280788 480 281028
rect 583520 272628 584960 272868
rect -960 267868 480 268108
rect 583520 259436 584960 259676
rect -960 254948 480 255188
rect 583520 246244 584960 246484
rect -960 242028 480 242268
rect 583520 233052 584960 233292
rect -960 229108 480 229348
rect 583520 219860 584960 220100
rect -960 216188 480 216428
rect 583520 206668 584960 206908
rect -960 203268 480 203508
rect 583520 193476 584960 193716
rect -960 190348 480 190588
rect 583520 180284 584960 180524
rect -960 177428 480 177668
rect 583520 167092 584960 167332
rect -960 164508 480 164748
rect 583520 153900 584960 154140
rect -960 151588 480 151828
rect 583520 140708 584960 140948
rect -960 138668 480 138908
rect 583520 127516 584960 127756
rect -960 125748 480 125988
rect 583520 114324 584960 114564
rect -960 112828 480 113068
rect 583520 101132 584960 101372
rect -960 99908 480 100148
rect 583520 87940 584960 88180
rect -960 86988 480 87228
rect 583520 74748 584960 74988
rect -960 74068 480 74308
rect 583520 61556 584960 61796
rect -960 61148 480 61388
rect -960 48228 480 48468
rect 583520 48364 584960 48604
rect -960 35308 480 35548
rect 583520 35172 584960 35412
rect -960 22388 480 22628
rect 583520 21980 584960 22220
rect -960 9468 480 9708
rect 583520 8788 584960 9028
<< obsm3 >>
rect 560 681228 583520 681461
rect 480 668708 583520 681228
rect 560 668308 583440 668708
rect 480 655788 583520 668308
rect 560 655516 583520 655788
rect 560 655388 583440 655516
rect 480 655116 583440 655388
rect 480 642868 583520 655116
rect 560 642468 583520 642868
rect 480 642324 583520 642468
rect 480 641924 583440 642324
rect 480 629948 583520 641924
rect 560 629548 583520 629948
rect 480 629132 583520 629548
rect 480 628732 583440 629132
rect 480 617028 583520 628732
rect 560 616628 583520 617028
rect 480 615940 583520 616628
rect 480 615540 583440 615940
rect 480 604108 583520 615540
rect 560 603708 583520 604108
rect 480 602748 583520 603708
rect 480 602348 583440 602748
rect 480 591188 583520 602348
rect 560 590788 583520 591188
rect 480 589556 583520 590788
rect 480 589156 583440 589556
rect 480 578268 583520 589156
rect 560 577868 583520 578268
rect 480 576364 583520 577868
rect 480 575964 583440 576364
rect 480 565348 583520 575964
rect 560 564948 583520 565348
rect 480 563172 583520 564948
rect 480 562772 583440 563172
rect 480 552428 583520 562772
rect 560 552028 583520 552428
rect 480 549980 583520 552028
rect 480 549580 583440 549980
rect 480 539508 583520 549580
rect 560 539108 583520 539508
rect 480 536788 583520 539108
rect 480 536388 583440 536788
rect 480 526588 583520 536388
rect 560 526188 583520 526588
rect 480 523596 583520 526188
rect 480 523196 583440 523596
rect 480 513668 583520 523196
rect 560 513268 583520 513668
rect 480 510404 583520 513268
rect 480 510004 583440 510404
rect 480 500748 583520 510004
rect 560 500348 583520 500748
rect 480 497212 583520 500348
rect 480 496812 583440 497212
rect 480 487828 583520 496812
rect 560 487428 583520 487828
rect 480 484020 583520 487428
rect 480 483620 583440 484020
rect 480 474908 583520 483620
rect 560 474508 583520 474908
rect 480 470828 583520 474508
rect 480 470428 583440 470828
rect 480 461988 583520 470428
rect 560 461588 583520 461988
rect 480 457636 583520 461588
rect 480 457236 583440 457636
rect 480 449068 583520 457236
rect 560 448668 583520 449068
rect 480 444444 583520 448668
rect 480 444044 583440 444444
rect 480 436148 583520 444044
rect 560 435748 583520 436148
rect 480 431252 583520 435748
rect 480 430852 583440 431252
rect 480 423228 583520 430852
rect 560 422828 583520 423228
rect 480 418060 583520 422828
rect 480 417660 583440 418060
rect 480 410308 583520 417660
rect 560 409908 583520 410308
rect 480 404868 583520 409908
rect 480 404468 583440 404868
rect 480 397388 583520 404468
rect 560 396988 583520 397388
rect 480 391676 583520 396988
rect 480 391276 583440 391676
rect 480 384468 583520 391276
rect 560 384068 583520 384468
rect 480 378484 583520 384068
rect 480 378084 583440 378484
rect 480 371548 583520 378084
rect 560 371148 583520 371548
rect 480 365292 583520 371148
rect 480 364892 583440 365292
rect 480 358628 583520 364892
rect 560 358228 583520 358628
rect 480 352100 583520 358228
rect 480 351700 583440 352100
rect 480 345708 583520 351700
rect 560 345308 583520 345708
rect 480 338908 583520 345308
rect 480 338508 583440 338908
rect 480 332788 583520 338508
rect 560 332388 583520 332788
rect 480 325716 583520 332388
rect 480 325316 583440 325716
rect 480 319868 583520 325316
rect 560 319468 583520 319868
rect 480 312524 583520 319468
rect 480 312124 583440 312524
rect 480 306948 583520 312124
rect 560 306548 583520 306948
rect 480 299332 583520 306548
rect 480 298932 583440 299332
rect 480 294028 583520 298932
rect 560 293628 583520 294028
rect 480 286140 583520 293628
rect 480 285740 583440 286140
rect 480 281108 583520 285740
rect 560 280708 583520 281108
rect 480 272948 583520 280708
rect 480 272548 583440 272948
rect 480 268188 583520 272548
rect 560 267788 583520 268188
rect 480 259756 583520 267788
rect 480 259356 583440 259756
rect 480 255268 583520 259356
rect 560 254868 583520 255268
rect 480 246564 583520 254868
rect 480 246164 583440 246564
rect 480 242348 583520 246164
rect 560 241948 583520 242348
rect 480 233372 583520 241948
rect 480 232972 583440 233372
rect 480 229428 583520 232972
rect 560 229028 583520 229428
rect 480 220180 583520 229028
rect 480 219780 583440 220180
rect 480 216508 583520 219780
rect 560 216108 583520 216508
rect 480 206988 583520 216108
rect 480 206588 583440 206988
rect 480 203588 583520 206588
rect 560 203188 583520 203588
rect 480 193796 583520 203188
rect 480 193396 583440 193796
rect 480 190668 583520 193396
rect 560 190268 583520 190668
rect 480 180604 583520 190268
rect 480 180204 583440 180604
rect 480 177748 583520 180204
rect 560 177348 583520 177748
rect 480 167412 583520 177348
rect 480 167012 583440 167412
rect 480 164828 583520 167012
rect 560 164428 583520 164828
rect 480 154220 583520 164428
rect 480 153820 583440 154220
rect 480 151908 583520 153820
rect 560 151508 583520 151908
rect 480 141028 583520 151508
rect 480 140628 583440 141028
rect 480 138988 583520 140628
rect 560 138588 583520 138988
rect 480 127836 583520 138588
rect 480 127436 583440 127836
rect 480 126068 583520 127436
rect 560 125668 583520 126068
rect 480 114644 583520 125668
rect 480 114244 583440 114644
rect 480 113148 583520 114244
rect 560 112748 583520 113148
rect 480 101452 583520 112748
rect 480 101052 583440 101452
rect 480 100228 583520 101052
rect 560 99828 583520 100228
rect 480 88260 583520 99828
rect 480 87860 583440 88260
rect 480 87308 583520 87860
rect 560 86908 583520 87308
rect 480 75068 583520 86908
rect 480 74668 583440 75068
rect 480 74388 583520 74668
rect 560 73988 583520 74388
rect 480 61876 583520 73988
rect 480 61476 583440 61876
rect 480 61468 583520 61476
rect 560 61068 583520 61468
rect 480 48684 583520 61068
rect 480 48548 583440 48684
rect 560 48284 583440 48548
rect 560 48148 583520 48284
rect 480 35628 583520 48148
rect 560 35492 583520 35628
rect 560 35228 583440 35492
rect 480 35092 583440 35228
rect 480 22708 583520 35092
rect 560 22308 583520 22708
rect 480 22300 583520 22308
rect 480 21900 583440 22300
rect 480 9788 583520 21900
rect 560 9555 583520 9788
<< metal4 >>
rect -9036 -7964 -8416 711900
rect -8076 -7004 -7456 710940
rect -7116 -6044 -6496 709980
rect -6156 -5084 -5536 709020
rect -5196 -4124 -4576 708060
rect -4236 -3164 -3616 707100
rect -3276 -2204 -2656 706140
rect -2316 -1244 -1696 705180
rect 1794 -7964 2414 711900
rect 4044 -7964 4664 711900
rect 6294 -7964 6914 711900
rect 8544 -7964 9164 711900
rect 10794 -7964 11414 711900
rect 13044 -7964 13664 711900
rect 15294 686000 15914 711900
rect 19794 686000 20414 711900
rect 22044 686000 22664 711900
rect 24294 686000 24914 711900
rect 26544 686000 27164 711900
rect 28794 686000 29414 711900
rect 31044 686000 31664 711900
rect 33294 686000 33914 711900
rect 37794 686000 38414 711900
rect 40044 38000 40664 711900
rect 42294 686000 42914 711900
rect 44544 686000 45164 711900
rect 46794 686000 47414 711900
rect 49044 686000 49664 711900
rect 51294 686000 51914 711900
rect 55794 686000 56414 711900
rect 58044 686000 58664 711900
rect 60294 686000 60914 711900
rect 62544 686000 63164 711900
rect 64794 686000 65414 711900
rect 19794 -7964 20414 14000
rect 22044 -7964 22664 14000
rect 24294 -7964 24914 14000
rect 26544 -7964 27164 14000
rect 28794 -7964 29414 14000
rect 37794 -7964 38414 14000
rect 40044 -7964 40664 14000
rect 42294 -7964 42914 14000
rect 44544 -7964 45164 14000
rect 46794 -7964 47414 14000
rect 55794 -7964 56414 14000
rect 58044 -7964 58664 14000
rect 60294 -7964 60914 14000
rect 62544 -7964 63164 14000
rect 64794 -7964 65414 41000
rect 67044 -7964 67664 711900
rect 69294 686000 69914 711900
rect 73794 686000 74414 711900
rect 76044 686000 76664 711900
rect 78294 686000 78914 711900
rect 80544 686000 81164 711900
rect 82794 686000 83414 711900
rect 85044 686000 85664 711900
rect 87294 686000 87914 711900
rect 91794 686000 92414 711900
rect 73794 -7964 74414 14000
rect 76044 -7964 76664 14000
rect 78294 -7964 78914 14000
rect 80544 -7964 81164 14000
rect 82794 -7964 83414 14000
rect 91794 -7964 92414 14000
rect 94044 -7964 94664 711900
rect 96294 686000 96914 711900
rect 98544 686000 99164 711900
rect 100794 686000 101414 711900
rect 103044 686000 103664 711900
rect 105294 686000 105914 711900
rect 109794 686000 110414 711900
rect 112044 686000 112664 711900
rect 114294 686000 114914 711900
rect 116544 686000 117164 711900
rect 118794 686000 119414 711900
rect 96294 -7964 96914 14000
rect 98544 -7964 99164 14000
rect 100794 -7964 101414 14000
rect 109794 -7964 110414 14000
rect 112044 -7964 112664 14000
rect 114294 -7964 114914 14000
rect 116544 -7964 117164 14000
rect 118794 -7964 119414 14000
rect 121044 -7964 121664 711900
rect 123294 686000 123914 711900
rect 127794 686000 128414 711900
rect 130044 686000 130664 711900
rect 132294 686000 132914 711900
rect 134544 686000 135164 711900
rect 136794 686000 137414 711900
rect 139044 686000 139664 711900
rect 141294 686000 141914 711900
rect 145794 686000 146414 711900
rect 127794 -7964 128414 14000
rect 130044 -7964 130664 14000
rect 132294 -7964 132914 14000
rect 134544 -7964 135164 14000
rect 136794 -7964 137414 14000
rect 145794 -7964 146414 14000
rect 148044 -7964 148664 711900
rect 150294 686000 150914 711900
rect 152544 686000 153164 711900
rect 154794 686000 155414 711900
rect 157044 686000 157664 711900
rect 159294 686000 159914 711900
rect 163794 686000 164414 711900
rect 166044 686000 166664 711900
rect 168294 686000 168914 711900
rect 170544 686000 171164 711900
rect 172794 686000 173414 711900
rect 150294 -7964 150914 14000
rect 152544 -7964 153164 14000
rect 154794 -7964 155414 14000
rect 163794 -7964 164414 14000
rect 166044 -7964 166664 14000
rect 168294 -7964 168914 14000
rect 170544 -7964 171164 14000
rect 172794 -7964 173414 14000
rect 175044 -7964 175664 711900
rect 177294 686000 177914 711900
rect 181794 686000 182414 711900
rect 184044 686000 184664 711900
rect 186294 686000 186914 711900
rect 188544 686000 189164 711900
rect 190794 686000 191414 711900
rect 193044 686000 193664 711900
rect 195294 686000 195914 711900
rect 199794 686000 200414 711900
rect 181794 -7964 182414 14000
rect 184044 -7964 184664 14000
rect 186294 -7964 186914 14000
rect 188544 -7964 189164 14000
rect 190794 -7964 191414 14000
rect 199794 -7964 200414 14000
rect 202044 -7964 202664 711900
rect 204294 686000 204914 711900
rect 206544 686000 207164 711900
rect 208794 686000 209414 711900
rect 211044 686000 211664 711900
rect 213294 686000 213914 711900
rect 217794 686000 218414 711900
rect 220044 686000 220664 711900
rect 222294 686000 222914 711900
rect 224544 686000 225164 711900
rect 226794 686000 227414 711900
rect 204294 -7964 204914 14000
rect 206544 -7964 207164 14000
rect 208794 -7964 209414 14000
rect 217794 -7964 218414 14000
rect 220044 -7964 220664 14000
rect 222294 -7964 222914 14000
rect 224544 -7964 225164 14000
rect 226794 -7964 227414 14000
rect 229044 -7964 229664 711900
rect 231294 686000 231914 711900
rect 235794 686000 236414 711900
rect 238044 686000 238664 711900
rect 240294 686000 240914 711900
rect 242544 686000 243164 711900
rect 244794 686000 245414 711900
rect 247044 686000 247664 711900
rect 249294 686000 249914 711900
rect 253794 686000 254414 711900
rect 235794 -7964 236414 14000
rect 238044 -7964 238664 14000
rect 240294 -7964 240914 14000
rect 242544 -7964 243164 14000
rect 244794 -7964 245414 14000
rect 253794 -7964 254414 14000
rect 256044 -7964 256664 711900
rect 258294 686000 258914 711900
rect 260544 686000 261164 711900
rect 262794 686000 263414 711900
rect 265044 686000 265664 711900
rect 267294 686000 267914 711900
rect 271794 686000 272414 711900
rect 274044 686000 274664 711900
rect 276294 686000 276914 711900
rect 278544 686000 279164 711900
rect 280794 686000 281414 711900
rect 258294 -7964 258914 14000
rect 260544 -7964 261164 14000
rect 262794 -7964 263414 14000
rect 271794 -7964 272414 14000
rect 274044 -7964 274664 14000
rect 276294 -7964 276914 14000
rect 278544 -7964 279164 14000
rect 280794 -7964 281414 14000
rect 283044 -7964 283664 711900
rect 285294 686000 285914 711900
rect 289794 686000 290414 711900
rect 292044 686000 292664 711900
rect 294294 686000 294914 711900
rect 296544 686000 297164 711900
rect 298794 686000 299414 711900
rect 301044 686000 301664 711900
rect 303294 686000 303914 711900
rect 307794 686000 308414 711900
rect 289794 -7964 290414 14000
rect 292044 -7964 292664 14000
rect 294294 -7964 294914 14000
rect 296544 -7964 297164 14000
rect 298794 -7964 299414 14000
rect 307794 -7964 308414 14000
rect 310044 -7964 310664 711900
rect 312294 686000 312914 711900
rect 314544 686000 315164 711900
rect 316794 686000 317414 711900
rect 319044 686000 319664 711900
rect 321294 686000 321914 711900
rect 325794 686000 326414 711900
rect 328044 686000 328664 711900
rect 330294 686000 330914 711900
rect 332544 686000 333164 711900
rect 334794 686000 335414 711900
rect 312294 -7964 312914 14000
rect 314544 -7964 315164 14000
rect 316794 -7964 317414 14000
rect 325794 -7964 326414 14000
rect 328044 -7964 328664 14000
rect 330294 -7964 330914 14000
rect 332544 -7964 333164 14000
rect 334794 -7964 335414 14000
rect 337044 -7964 337664 711900
rect 339294 686000 339914 711900
rect 343794 686000 344414 711900
rect 346044 686000 346664 711900
rect 348294 686000 348914 711900
rect 350544 686000 351164 711900
rect 352794 686000 353414 711900
rect 355044 686000 355664 711900
rect 357294 686000 357914 711900
rect 361794 686000 362414 711900
rect 343794 -7964 344414 14000
rect 346044 -7964 346664 14000
rect 348294 -7964 348914 14000
rect 350544 -7964 351164 14000
rect 352794 -7964 353414 14000
rect 361794 -7964 362414 14000
rect 364044 -7964 364664 711900
rect 366294 686000 366914 711900
rect 368544 686000 369164 711900
rect 370794 686000 371414 711900
rect 373044 686000 373664 711900
rect 375294 686000 375914 711900
rect 379794 686000 380414 711900
rect 382044 686000 382664 711900
rect 384294 686000 384914 711900
rect 386544 686000 387164 711900
rect 388794 686000 389414 711900
rect 366294 -7964 366914 14000
rect 368544 -7964 369164 14000
rect 370794 -7964 371414 14000
rect 379794 -7964 380414 14000
rect 382044 -7964 382664 14000
rect 384294 -7964 384914 14000
rect 386544 -7964 387164 14000
rect 388794 -7964 389414 14000
rect 391044 -7964 391664 711900
rect 393294 686000 393914 711900
rect 397794 686000 398414 711900
rect 400044 686000 400664 711900
rect 402294 686000 402914 711900
rect 404544 686000 405164 711900
rect 406794 686000 407414 711900
rect 409044 686000 409664 711900
rect 411294 686000 411914 711900
rect 415794 686000 416414 711900
rect 397794 -7964 398414 14000
rect 400044 -7964 400664 14000
rect 402294 -7964 402914 14000
rect 404544 -7964 405164 14000
rect 406794 -7964 407414 14000
rect 415794 -7964 416414 14000
rect 418044 -7964 418664 711900
rect 420294 686000 420914 711900
rect 422544 686000 423164 711900
rect 424794 686000 425414 711900
rect 427044 686000 427664 711900
rect 429294 686000 429914 711900
rect 433794 686000 434414 711900
rect 436044 686000 436664 711900
rect 438294 686000 438914 711900
rect 440544 686000 441164 711900
rect 442794 686000 443414 711900
rect 420294 -7964 420914 14000
rect 422544 -7964 423164 14000
rect 424794 -7964 425414 14000
rect 433794 -7964 434414 14000
rect 436044 -7964 436664 14000
rect 438294 -7964 438914 14000
rect 440544 -7964 441164 14000
rect 442794 -7964 443414 14000
rect 445044 -7964 445664 711900
rect 447294 686000 447914 711900
rect 451794 686000 452414 711900
rect 454044 686000 454664 711900
rect 456294 686000 456914 711900
rect 458544 686000 459164 711900
rect 460794 686000 461414 711900
rect 463044 686000 463664 711900
rect 465294 686000 465914 711900
rect 469794 686000 470414 711900
rect 451794 -7964 452414 14000
rect 454044 -7964 454664 14000
rect 456294 -7964 456914 14000
rect 458544 -7964 459164 14000
rect 460794 -7964 461414 14000
rect 469794 -7964 470414 14000
rect 472044 -7964 472664 711900
rect 474294 686000 474914 711900
rect 476544 686000 477164 711900
rect 478794 686000 479414 711900
rect 481044 686000 481664 711900
rect 483294 686000 483914 711900
rect 487794 686000 488414 711900
rect 490044 686000 490664 711900
rect 492294 686000 492914 711900
rect 494544 686000 495164 711900
rect 496794 686000 497414 711900
rect 474294 -7964 474914 14000
rect 476544 -7964 477164 14000
rect 478794 -7964 479414 14000
rect 487794 -7964 488414 14000
rect 490044 -7964 490664 14000
rect 492294 -7964 492914 14000
rect 494544 -7964 495164 14000
rect 496794 -7964 497414 14000
rect 499044 -7964 499664 711900
rect 501294 686000 501914 711900
rect 505794 686000 506414 711900
rect 508044 686000 508664 711900
rect 510294 686000 510914 711900
rect 512544 686000 513164 711900
rect 514794 686000 515414 711900
rect 517044 686000 517664 711900
rect 519294 686000 519914 711900
rect 523794 686000 524414 711900
rect 505794 -7964 506414 14000
rect 508044 -7964 508664 14000
rect 510294 -7964 510914 14000
rect 512544 -7964 513164 14000
rect 514794 -7964 515414 14000
rect 523794 -7964 524414 14000
rect 526044 -7964 526664 711900
rect 528294 686000 528914 711900
rect 530544 686000 531164 711900
rect 532794 686000 533414 711900
rect 535044 686000 535664 711900
rect 537294 686000 537914 711900
rect 541794 686000 542414 711900
rect 544044 686000 544664 711900
rect 546294 686000 546914 711900
rect 548544 686000 549164 711900
rect 550794 686000 551414 711900
rect 528294 -7964 528914 14000
rect 530544 -7964 531164 14000
rect 532794 -7964 533414 14000
rect 541794 -7964 542414 14000
rect 544044 -7964 544664 14000
rect 546294 -7964 546914 14000
rect 548544 -7964 549164 14000
rect 550794 -7964 551414 14000
rect 553044 -7964 553664 711900
rect 555294 -7964 555914 711900
rect 557544 -7964 558164 711900
rect 559794 -7964 560414 711900
rect 562044 -7964 562664 711900
rect 564294 -7964 564914 711900
rect 566544 -7964 567164 711900
rect 568794 -7964 569414 711900
rect 571044 -7964 571664 711900
rect 573294 -7964 573914 711900
rect 575544 -7964 576164 711900
rect 577794 -7964 578414 711900
rect 580044 -7964 580664 711900
rect 582294 -7964 582914 711900
rect 585620 -1244 586240 705180
rect 586580 -2204 587200 706140
rect 587540 -3164 588160 707100
rect 588500 -4124 589120 708060
rect 589460 -5084 590080 709020
rect 590420 -6044 591040 709980
rect 591380 -7004 592000 710940
rect 592340 -7964 592960 711900
<< obsm4 >>
rect 19910 37920 39964 681456
rect 40744 41080 66964 681456
rect 40744 37920 64714 41080
rect 19910 18128 64714 37920
rect 65494 18128 66964 41080
rect 67744 18128 93964 681456
rect 94744 18128 120964 681456
rect 121744 18128 147964 681456
rect 148744 18128 174964 681456
rect 175744 18128 201964 681456
rect 202744 18128 228964 681456
rect 229744 18128 255964 681456
rect 256744 18128 282964 681456
rect 283744 18128 309964 681456
rect 310744 18128 336964 681456
rect 337744 18128 363964 681456
rect 364744 18128 390964 681456
rect 391744 18128 417964 681456
rect 418744 18128 444964 681456
rect 445744 18128 471964 681456
rect 472744 18128 498964 681456
rect 499744 18128 525964 681456
rect 526744 18128 545091 681456
<< metal5 >>
rect -9036 711280 592960 711900
rect -8076 710320 592000 710940
rect -7116 709360 591040 709980
rect -6156 708400 590080 709020
rect -5196 707440 589120 708060
rect -4236 706480 588160 707100
rect -3276 705520 587200 706140
rect -2316 704560 586240 705180
rect -9036 700366 592960 700986
rect -9036 698116 592960 698736
rect -9036 695866 592960 696486
rect -9036 693616 592960 694236
rect -9036 691366 592960 691986
rect -9036 689116 592960 689736
rect -9036 686866 592960 687486
rect -9036 684616 592960 685236
rect -9036 682366 592960 682986
rect -9036 680116 592960 680736
rect -9036 677866 592960 678486
rect -9036 675616 592960 676236
rect -9036 673366 592960 673986
rect -9036 671116 592960 671736
rect -9036 668866 592960 669486
rect -9036 666616 592960 667236
rect -9036 664366 592960 664986
rect -9036 662116 592960 662736
rect -9036 659866 592960 660486
rect -9036 657616 592960 658236
rect -9036 655366 592960 655986
rect -9036 653116 592960 653736
rect -9036 650866 592960 651486
rect -9036 648616 592960 649236
rect -9036 646366 592960 646986
rect -9036 644116 592960 644736
rect -9036 641866 592960 642486
rect -9036 639616 592960 640236
rect -9036 637366 592960 637986
rect -9036 635116 592960 635736
rect -9036 632866 592960 633486
rect -9036 630616 592960 631236
rect -9036 628366 592960 628986
rect -9036 626116 592960 626736
rect -9036 623866 592960 624486
rect -9036 621616 592960 622236
rect -9036 619366 592960 619986
rect -9036 617116 592960 617736
rect -9036 614866 592960 615486
rect -9036 612616 592960 613236
rect -9036 610366 592960 610986
rect -9036 608116 592960 608736
rect -9036 605866 592960 606486
rect -9036 603616 592960 604236
rect -9036 601366 592960 601986
rect -9036 599116 592960 599736
rect -9036 596866 592960 597486
rect -9036 594616 592960 595236
rect -9036 592366 592960 592986
rect -9036 590116 592960 590736
rect -9036 587866 592960 588486
rect -9036 585616 592960 586236
rect -9036 583366 592960 583986
rect -9036 581116 592960 581736
rect -9036 578866 592960 579486
rect -9036 576616 592960 577236
rect -9036 574366 592960 574986
rect -9036 572116 592960 572736
rect -9036 569866 592960 570486
rect -9036 567616 592960 568236
rect -9036 565366 592960 565986
rect -9036 563116 592960 563736
rect -9036 560866 592960 561486
rect -9036 558616 592960 559236
rect -9036 556366 592960 556986
rect -9036 554116 592960 554736
rect -9036 551866 592960 552486
rect -9036 549616 592960 550236
rect -9036 547366 592960 547986
rect -9036 545116 592960 545736
rect -9036 542866 592960 543486
rect -9036 540616 592960 541236
rect -9036 538366 592960 538986
rect -9036 536116 592960 536736
rect -9036 533866 592960 534486
rect -9036 531616 592960 532236
rect -9036 529366 592960 529986
rect -9036 527116 592960 527736
rect -9036 524866 592960 525486
rect -9036 522616 592960 523236
rect -9036 520366 592960 520986
rect -9036 518116 592960 518736
rect -9036 515866 592960 516486
rect -9036 513616 592960 514236
rect -9036 511366 592960 511986
rect -9036 509116 592960 509736
rect -9036 506866 592960 507486
rect -9036 504616 592960 505236
rect -9036 502366 592960 502986
rect -9036 500116 592960 500736
rect -9036 497866 592960 498486
rect -9036 495616 592960 496236
rect -9036 493366 592960 493986
rect -9036 491116 592960 491736
rect -9036 488866 592960 489486
rect -9036 486616 592960 487236
rect -9036 484366 592960 484986
rect -9036 482116 592960 482736
rect -9036 479866 592960 480486
rect -9036 477616 592960 478236
rect -9036 475366 592960 475986
rect -9036 473116 592960 473736
rect -9036 470866 592960 471486
rect -9036 468616 592960 469236
rect -9036 466366 592960 466986
rect -9036 464116 592960 464736
rect -9036 461866 592960 462486
rect -9036 459616 592960 460236
rect -9036 457366 592960 457986
rect -9036 455116 592960 455736
rect -9036 452866 592960 453486
rect -9036 450616 592960 451236
rect -9036 448366 592960 448986
rect -9036 446116 592960 446736
rect -9036 443866 592960 444486
rect -9036 441616 592960 442236
rect -9036 439366 592960 439986
rect -9036 437116 592960 437736
rect -9036 434866 592960 435486
rect -9036 432616 592960 433236
rect -9036 430366 592960 430986
rect -9036 428116 592960 428736
rect -9036 425866 592960 426486
rect -9036 423616 592960 424236
rect -9036 421366 592960 421986
rect -9036 419116 592960 419736
rect -9036 416866 592960 417486
rect -9036 414616 592960 415236
rect -9036 412366 592960 412986
rect -9036 410116 592960 410736
rect -9036 407866 592960 408486
rect -9036 405616 592960 406236
rect -9036 403366 592960 403986
rect -9036 401116 592960 401736
rect -9036 398866 592960 399486
rect -9036 396616 592960 397236
rect -9036 394366 592960 394986
rect -9036 392116 592960 392736
rect -9036 389866 592960 390486
rect -9036 387616 592960 388236
rect -9036 385366 592960 385986
rect -9036 383116 592960 383736
rect -9036 380866 592960 381486
rect -9036 378616 592960 379236
rect -9036 376366 592960 376986
rect -9036 374116 592960 374736
rect -9036 371866 592960 372486
rect -9036 369616 592960 370236
rect -9036 367366 592960 367986
rect -9036 365116 592960 365736
rect -9036 362866 592960 363486
rect -9036 360616 592960 361236
rect -9036 358366 592960 358986
rect -9036 356116 592960 356736
rect -9036 353866 592960 354486
rect -9036 351616 592960 352236
rect -9036 349366 592960 349986
rect -9036 347116 592960 347736
rect -9036 344866 592960 345486
rect -9036 342616 592960 343236
rect -9036 340366 592960 340986
rect -9036 338116 592960 338736
rect -9036 335866 592960 336486
rect -9036 333616 592960 334236
rect -9036 331366 592960 331986
rect -9036 329116 592960 329736
rect -9036 326866 592960 327486
rect -9036 324616 592960 325236
rect -9036 322366 592960 322986
rect -9036 320116 592960 320736
rect -9036 317866 592960 318486
rect -9036 315616 592960 316236
rect -9036 313366 592960 313986
rect -9036 311116 592960 311736
rect -9036 308866 592960 309486
rect -9036 306616 592960 307236
rect -9036 304366 592960 304986
rect -9036 302116 592960 302736
rect -9036 299866 592960 300486
rect -9036 297616 592960 298236
rect -9036 295366 592960 295986
rect -9036 293116 592960 293736
rect -9036 290866 592960 291486
rect -9036 288616 592960 289236
rect -9036 286366 592960 286986
rect -9036 284116 592960 284736
rect -9036 281866 592960 282486
rect -9036 279616 592960 280236
rect -9036 277366 592960 277986
rect -9036 275116 592960 275736
rect -9036 272866 592960 273486
rect -9036 270616 592960 271236
rect -9036 268366 592960 268986
rect -9036 266116 592960 266736
rect -9036 263866 592960 264486
rect -9036 261616 592960 262236
rect -9036 259366 592960 259986
rect -9036 257116 592960 257736
rect -9036 254866 592960 255486
rect -9036 252616 592960 253236
rect -9036 250366 592960 250986
rect -9036 248116 592960 248736
rect -9036 245866 592960 246486
rect -9036 243616 592960 244236
rect -9036 241366 592960 241986
rect -9036 239116 592960 239736
rect -9036 236866 592960 237486
rect -9036 234616 592960 235236
rect -9036 232366 592960 232986
rect -9036 230116 592960 230736
rect -9036 227866 592960 228486
rect -9036 225616 592960 226236
rect -9036 223366 592960 223986
rect -9036 221116 592960 221736
rect -9036 218866 592960 219486
rect -9036 216616 592960 217236
rect -9036 214366 592960 214986
rect -9036 212116 592960 212736
rect -9036 209866 592960 210486
rect -9036 207616 592960 208236
rect -9036 205366 592960 205986
rect -9036 203116 592960 203736
rect -9036 200866 592960 201486
rect -9036 198616 592960 199236
rect -9036 196366 592960 196986
rect -9036 194116 592960 194736
rect -9036 191866 592960 192486
rect -9036 189616 592960 190236
rect -9036 187366 592960 187986
rect -9036 185116 592960 185736
rect -9036 182866 592960 183486
rect -9036 180616 592960 181236
rect -9036 178366 592960 178986
rect -9036 176116 592960 176736
rect -9036 173866 592960 174486
rect -9036 171616 592960 172236
rect -9036 169366 592960 169986
rect -9036 167116 592960 167736
rect -9036 164866 592960 165486
rect -9036 162616 592960 163236
rect -9036 160366 592960 160986
rect -9036 158116 592960 158736
rect -9036 155866 592960 156486
rect -9036 153616 592960 154236
rect -9036 151366 592960 151986
rect -9036 149116 592960 149736
rect -9036 146866 592960 147486
rect -9036 144616 592960 145236
rect -9036 142366 592960 142986
rect -9036 140116 592960 140736
rect -9036 137866 592960 138486
rect -9036 135616 592960 136236
rect -9036 133366 592960 133986
rect -9036 131116 592960 131736
rect -9036 128866 592960 129486
rect -9036 126616 592960 127236
rect -9036 124366 592960 124986
rect -9036 122116 592960 122736
rect -9036 119866 592960 120486
rect -9036 117616 592960 118236
rect -9036 115366 592960 115986
rect -9036 113116 592960 113736
rect -9036 110866 592960 111486
rect -9036 108616 592960 109236
rect -9036 106366 592960 106986
rect -9036 104116 592960 104736
rect -9036 101866 592960 102486
rect -9036 99616 592960 100236
rect -9036 97366 592960 97986
rect -9036 95116 592960 95736
rect -9036 92866 592960 93486
rect -9036 90616 592960 91236
rect -9036 88366 592960 88986
rect -9036 86116 592960 86736
rect -9036 83866 592960 84486
rect -9036 81616 592960 82236
rect -9036 79366 592960 79986
rect -9036 77116 592960 77736
rect -9036 74866 592960 75486
rect -9036 72616 592960 73236
rect -9036 70366 592960 70986
rect -9036 68116 592960 68736
rect -9036 65866 592960 66486
rect -9036 63616 592960 64236
rect -9036 61366 592960 61986
rect -9036 59116 592960 59736
rect -9036 56866 592960 57486
rect -9036 54616 592960 55236
rect -9036 52366 592960 52986
rect -9036 50116 592960 50736
rect -9036 47866 592960 48486
rect -9036 45616 592960 46236
rect -9036 43366 592960 43986
rect -9036 41116 592960 41736
rect -9036 38866 592960 39486
rect -9036 36616 592960 37236
rect -9036 34366 592960 34986
rect -9036 32116 592960 32736
rect -9036 29866 592960 30486
rect -9036 27616 592960 28236
rect -9036 25366 592960 25986
rect -9036 23116 592960 23736
rect -9036 20866 592960 21486
rect -9036 18616 592960 19236
rect -9036 16366 592960 16986
rect -9036 14116 592960 14736
rect -9036 11866 592960 12486
rect -9036 9616 592960 10236
rect -9036 7366 592960 7986
rect -9036 5116 592960 5736
rect -9036 2866 592960 3486
rect -2316 -1244 586240 -624
rect -3276 -2204 587200 -1584
rect -4236 -3164 588160 -2544
rect -5196 -4124 589120 -3504
rect -6156 -5084 590080 -4464
rect -7116 -6044 591040 -5424
rect -8076 -7004 592000 -6384
rect -9036 -7964 592960 -7344
<< labels >>
rlabel metal3 s 583520 285820 584960 286060 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 445730 703520 445842 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 380962 703520 381074 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316194 703520 316306 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186658 703520 186770 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121890 703520 122002 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 57122 703520 57234 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 694228 480 694468 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 642548 480 642788 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 590868 480 591108 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338588 584960 338828 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 539188 480 539428 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 487508 480 487748 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 435828 480 436068 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384148 480 384388 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332468 480 332708 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 280788 480 281028 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 229108 480 229348 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 177428 480 177668 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 125748 480 125988 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391356 584960 391596 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444124 584960 444364 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 496892 584960 497132 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 549660 584960 549900 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 602428 584960 602668 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 655196 584960 655436 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575266 703520 575378 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510498 703520 510610 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 8788 584960 9028 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457316 584960 457556 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 510084 584960 510324 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 562852 584960 563092 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 615620 584960 615860 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 668388 584960 668628 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559074 703520 559186 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494306 703520 494418 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429538 703520 429650 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364770 703520 364882 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300002 703520 300114 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 48364 584960 48604 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235234 703520 235346 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170466 703520 170578 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105698 703520 105810 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40930 703520 41042 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 681308 480 681548 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 629628 480 629868 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 577948 480 578188 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 526268 480 526508 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 474588 480 474828 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 422908 480 423148 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 87940 584960 88180 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319548 480 319788 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267868 480 268108 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 216188 480 216428 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 164508 480 164748 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 112828 480 113068 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 74068 480 74308 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 35308 480 35548 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 127516 584960 127756 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 167092 584960 167332 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 206668 584960 206908 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 246244 584960 246484 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404548 584960 404788 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 35172 584960 35412 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 483700 584960 483940 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 536468 584960 536708 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 589236 584960 589476 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 642004 584960 642244 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 694772 584960 695012 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 526690 703520 526802 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 461922 703520 462034 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397154 703520 397266 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332386 703520 332498 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 74748 584960 74988 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202850 703520 202962 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 138082 703520 138194 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 73314 703520 73426 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8546 703520 8658 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 655468 480 655708 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 603788 480 604028 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 552108 480 552348 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 500428 480 500668 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 448748 480 448988 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397068 480 397308 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 114324 584960 114564 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345388 480 345628 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293708 480 293948 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 242028 480 242268 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 190348 480 190588 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 138668 480 138908 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 86988 480 87228 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 48228 480 48468 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 9468 480 9708 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 153900 584960 154140 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 193476 584960 193716 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 233052 584960 233292 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272628 584960 272868 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325396 584960 325636 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378164 584960 378404 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 430932 584960 431172 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 21980 584960 22220 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 470508 584960 470748 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 523276 584960 523516 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 576044 584960 576284 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 628812 584960 629052 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 681580 584960 681820 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 542882 703520 542994 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478114 703520 478226 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413346 703520 413458 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348578 703520 348690 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 61556 584960 61796 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 219042 703520 219154 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154274 703520 154386 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89506 703520 89618 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24738 703520 24850 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 668388 480 668628 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 616708 480 616948 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 565028 480 565268 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 513348 480 513588 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 461668 480 461908 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 409988 480 410228 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 101132 584960 101372 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306628 480 306868 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 254948 480 255188 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 203268 480 203508 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 151588 480 151828 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 99908 480 100148 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 61148 480 61388 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 22388 480 22628 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 140708 584960 140948 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 180284 584960 180524 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 219860 584960 220100 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 259436 584960 259676 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 312204 584960 312444 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 417740 584960 417980 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 136794 -960 136906 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 467994 -960 468106 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 471306 -960 471418 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 474618 -960 474730 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 477930 -960 478042 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 481242 -960 481354 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 484554 -960 484666 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 487866 -960 487978 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 491178 -960 491290 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 494490 -960 494602 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 497802 -960 497914 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 169914 -960 170026 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 501114 -960 501226 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 504426 -960 504538 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 507738 -960 507850 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 511050 -960 511162 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 514362 -960 514474 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 517674 -960 517786 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 520986 -960 521098 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 524298 -960 524410 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 527610 -960 527722 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 530922 -960 531034 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 173226 -960 173338 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 534234 -960 534346 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 537546 -960 537658 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 540858 -960 540970 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 544170 -960 544282 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 547482 -960 547594 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 550794 -960 550906 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 554106 -960 554218 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 557418 -960 557530 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 179850 -960 179962 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 183162 -960 183274 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 186474 -960 186586 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 189786 -960 189898 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 193098 -960 193210 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 196410 -960 196522 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 199722 -960 199834 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 140106 -960 140218 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 203034 -960 203146 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 206346 -960 206458 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 209658 -960 209770 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 212970 -960 213082 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 216282 -960 216394 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 219594 -960 219706 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 226218 -960 226330 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 229530 -960 229642 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 232842 -960 232954 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 143418 -960 143530 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 236154 -960 236266 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 239466 -960 239578 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 242778 -960 242890 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 246090 -960 246202 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 249402 -960 249514 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 252714 -960 252826 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 256026 -960 256138 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 259338 -960 259450 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 262650 -960 262762 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 265962 -960 266074 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 146730 -960 146842 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 272586 -960 272698 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 275898 -960 276010 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 279210 -960 279322 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 282522 -960 282634 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285834 -960 285946 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 289146 -960 289258 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292458 -960 292570 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 295770 -960 295882 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299082 -960 299194 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 150042 -960 150154 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 302394 -960 302506 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 305706 -960 305818 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 312330 -960 312442 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 315642 -960 315754 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 318954 -960 319066 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 322266 -960 322378 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 325578 -960 325690 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 328890 -960 329002 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 332202 -960 332314 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 153354 -960 153466 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 335514 -960 335626 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 338826 -960 338938 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 345450 -960 345562 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 348762 -960 348874 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 352074 -960 352186 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 355386 -960 355498 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 362010 -960 362122 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 365322 -960 365434 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 156666 -960 156778 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 368634 -960 368746 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 371946 -960 372058 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 375258 -960 375370 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 378570 -960 378682 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 381882 -960 381994 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 385194 -960 385306 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 388506 -960 388618 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 395130 -960 395242 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 398442 -960 398554 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 159978 -960 160090 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 401754 -960 401866 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 405066 -960 405178 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 411690 -960 411802 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 415002 -960 415114 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 418314 -960 418426 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 421626 -960 421738 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 424938 -960 425050 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 428250 -960 428362 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 431562 -960 431674 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 163290 -960 163402 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 434874 -960 434986 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 438186 -960 438298 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 444810 -960 444922 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 448122 -960 448234 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 451434 -960 451546 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 454746 -960 454858 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 461370 -960 461482 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 464682 -960 464794 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 166602 -960 166714 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 137898 -960 138010 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 469098 -960 469210 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 472410 -960 472522 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 475722 -960 475834 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 479034 -960 479146 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 482346 -960 482458 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 485658 -960 485770 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 488970 -960 489082 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 495594 -960 495706 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 171018 -960 171130 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 502218 -960 502330 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 505530 -960 505642 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 508842 -960 508954 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 512154 -960 512266 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 515466 -960 515578 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 518778 -960 518890 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 522090 -960 522202 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 525402 -960 525514 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 528714 -960 528826 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 532026 -960 532138 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 174330 -960 174442 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 535338 -960 535450 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 538650 -960 538762 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 548586 -960 548698 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 551898 -960 552010 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 555210 -960 555322 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 558522 -960 558634 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 177642 -960 177754 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 180954 -960 181066 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 184266 -960 184378 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 187578 -960 187690 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 190890 -960 191002 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 194202 -960 194314 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 197514 -960 197626 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 200826 -960 200938 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 204138 -960 204250 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 207450 -960 207562 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 210762 -960 210874 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 214074 -960 214186 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 217386 -960 217498 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 220698 -960 220810 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 224010 -960 224122 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 227322 -960 227434 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 230634 -960 230746 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 233946 -960 234058 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 144522 -960 144634 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 237258 -960 237370 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 240570 -960 240682 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 243882 -960 243994 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 247194 -960 247306 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 250506 -960 250618 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 253818 -960 253930 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 257130 -960 257242 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 260442 -960 260554 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 263754 -960 263866 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 267066 -960 267178 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 147834 -960 147946 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 270378 -960 270490 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 273690 -960 273802 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 277002 -960 277114 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 280314 -960 280426 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283626 -960 283738 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286938 -960 287050 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290250 -960 290362 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293562 -960 293674 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 296874 -960 296986 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300186 -960 300298 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 151146 -960 151258 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 303498 -960 303610 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 306810 -960 306922 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 310122 -960 310234 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 313434 -960 313546 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 316746 -960 316858 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 320058 -960 320170 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 323370 -960 323482 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 326682 -960 326794 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 329994 -960 330106 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 333306 -960 333418 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 154458 -960 154570 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 336618 -960 336730 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 339930 -960 340042 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 343242 -960 343354 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 346554 -960 346666 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 349866 -960 349978 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 353178 -960 353290 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 356490 -960 356602 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 359802 -960 359914 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 363114 -960 363226 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 366426 -960 366538 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 157770 -960 157882 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 369738 -960 369850 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 373050 -960 373162 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 376362 -960 376474 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 379674 -960 379786 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 382986 -960 383098 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 386298 -960 386410 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 389610 -960 389722 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 392922 -960 393034 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 396234 -960 396346 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 399546 -960 399658 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 161082 -960 161194 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 402858 -960 402970 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 406170 -960 406282 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 409482 -960 409594 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 412794 -960 412906 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 416106 -960 416218 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 419418 -960 419530 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 422730 -960 422842 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 426042 -960 426154 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 429354 -960 429466 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 432666 -960 432778 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 164394 -960 164506 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 435978 -960 436090 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 439290 -960 439402 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 445914 -960 446026 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 449226 -960 449338 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 452538 -960 452650 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 455850 -960 455962 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 459162 -960 459274 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 462474 -960 462586 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 465786 -960 465898 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 167706 -960 167818 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 139002 -960 139114 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 470202 -960 470314 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 473514 -960 473626 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 476826 -960 476938 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 480138 -960 480250 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 483450 -960 483562 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 486762 -960 486874 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 490074 -960 490186 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 493386 -960 493498 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 496698 -960 496810 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 500010 -960 500122 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 172122 -960 172234 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 503322 -960 503434 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 506634 -960 506746 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 509946 -960 510058 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 513258 -960 513370 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 516570 -960 516682 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 519882 -960 519994 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 523194 -960 523306 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 526506 -960 526618 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 529818 -960 529930 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 533130 -960 533242 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 536442 -960 536554 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 539754 -960 539866 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 543066 -960 543178 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 546378 -960 546490 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 549690 -960 549802 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 553002 -960 553114 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 556314 -960 556426 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 559626 -960 559738 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 178746 -960 178858 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 182058 -960 182170 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 185370 -960 185482 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 188682 -960 188794 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 195306 -960 195418 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 198618 -960 198730 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 201930 -960 202042 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 142314 -960 142426 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 205242 -960 205354 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 208554 -960 208666 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 211866 -960 211978 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 215178 -960 215290 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 218490 -960 218602 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 221802 -960 221914 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 228426 -960 228538 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 231738 -960 231850 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 235050 -960 235162 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 145626 -960 145738 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 238362 -960 238474 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 244986 -960 245098 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 248298 -960 248410 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 251610 -960 251722 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 254922 -960 255034 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 258234 -960 258346 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 261546 -960 261658 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 264858 -960 264970 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 268170 -960 268282 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 148938 -960 149050 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 271482 -960 271594 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 278106 -960 278218 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 281418 -960 281530 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284730 -960 284842 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 288042 -960 288154 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294666 -960 294778 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 297978 -960 298090 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301290 -960 301402 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 152250 -960 152362 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 304602 -960 304714 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 307914 -960 308026 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 311226 -960 311338 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 314538 -960 314650 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 317850 -960 317962 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 321162 -960 321274 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 324474 -960 324586 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 327786 -960 327898 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 331098 -960 331210 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 334410 -960 334522 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 155562 -960 155674 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 337722 -960 337834 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 341034 -960 341146 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 344346 -960 344458 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 347658 -960 347770 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 350970 -960 351082 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 354282 -960 354394 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 357594 -960 357706 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 360906 -960 361018 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 364218 -960 364330 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 367530 -960 367642 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 158874 -960 158986 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 370842 -960 370954 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 374154 -960 374266 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 377466 -960 377578 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 380778 -960 380890 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 384090 -960 384202 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 387402 -960 387514 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 390714 -960 390826 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 394026 -960 394138 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 397338 -960 397450 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 400650 -960 400762 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 162186 -960 162298 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 403962 -960 404074 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 407274 -960 407386 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 410586 -960 410698 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 413898 -960 414010 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 417210 -960 417322 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 420522 -960 420634 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 423834 -960 423946 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 427146 -960 427258 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 430458 -960 430570 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 433770 -960 433882 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 165498 -960 165610 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 437082 -960 437194 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 440394 -960 440506 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 443706 -960 443818 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 447018 -960 447130 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 450330 -960 450442 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 453642 -960 453754 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 456954 -960 457066 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 460266 -960 460378 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 463578 -960 463690 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 466890 -960 467002 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 168810 -960 168922 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 560730 -960 560842 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 561834 -960 561946 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 562938 -960 563050 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 564042 -960 564154 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal4 s -2316 -1244 -1696 705180 4 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2316 -1244 586240 -624 8 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2316 704560 586240 705180 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 585620 -1244 586240 705180 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 1794 -7964 2414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 19794 -7964 20414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 19794 686000 20414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 37794 -7964 38414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 37794 686000 38414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 55794 -7964 56414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 55794 686000 56414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 -7964 74414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 686000 74414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 91794 -7964 92414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 91794 686000 92414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 -7964 110414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 686000 110414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127794 -7964 128414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127794 686000 128414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 -7964 146414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 686000 146414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 163794 -7964 164414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 163794 686000 164414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 -7964 182414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 686000 182414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 199794 -7964 200414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 199794 686000 200414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 217794 -7964 218414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 217794 686000 218414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 235794 -7964 236414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 235794 686000 236414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253794 -7964 254414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253794 686000 254414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 271794 -7964 272414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 271794 686000 272414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 289794 -7964 290414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 289794 686000 290414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 307794 -7964 308414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 307794 686000 308414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 325794 -7964 326414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 325794 686000 326414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 343794 -7964 344414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 343794 686000 344414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 361794 -7964 362414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 361794 686000 362414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 379794 -7964 380414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 379794 686000 380414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 -7964 398414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 686000 398414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 415794 -7964 416414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 415794 686000 416414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 -7964 434414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 686000 434414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 451794 -7964 452414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 451794 686000 452414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 -7964 470414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 686000 470414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 487794 -7964 488414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 487794 686000 488414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 -7964 506414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 686000 506414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 523794 -7964 524414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 523794 686000 524414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 541794 -7964 542414 14000 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 541794 686000 542414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 559794 -7964 560414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 577794 -7964 578414 711900 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 2866 592960 3486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 20866 592960 21486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 38866 592960 39486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 56866 592960 57486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 74866 592960 75486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 92866 592960 93486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 110866 592960 111486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 128866 592960 129486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 146866 592960 147486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 164866 592960 165486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 182866 592960 183486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 200866 592960 201486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 218866 592960 219486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 236866 592960 237486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 254866 592960 255486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 272866 592960 273486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 290866 592960 291486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 308866 592960 309486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 326866 592960 327486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 344866 592960 345486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 362866 592960 363486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 380866 592960 381486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 398866 592960 399486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 416866 592960 417486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 434866 592960 435486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 452866 592960 453486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 470866 592960 471486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 488866 592960 489486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 506866 592960 507486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 524866 592960 525486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 542866 592960 543486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 560866 592960 561486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 578866 592960 579486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 596866 592960 597486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 614866 592960 615486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 632866 592960 633486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 650866 592960 651486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 668866 592960 669486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -9036 686866 592960 687486 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s -4236 -3164 -3616 707100 4 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4236 -3164 588160 -2544 8 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -4236 706480 588160 707100 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 587540 -3164 588160 707100 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 6294 -7964 6914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 24294 -7964 24914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 24294 686000 24914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 42294 -7964 42914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 42294 686000 42914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 60294 -7964 60914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 60294 686000 60914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 78294 -7964 78914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 78294 686000 78914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 96294 -7964 96914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 96294 686000 96914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 114294 -7964 114914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 114294 686000 114914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 132294 -7964 132914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 132294 686000 132914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 150294 -7964 150914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 150294 686000 150914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 168294 -7964 168914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 168294 686000 168914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 186294 -7964 186914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 186294 686000 186914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 204294 -7964 204914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 204294 686000 204914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 222294 -7964 222914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 222294 686000 222914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 240294 -7964 240914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 240294 686000 240914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 258294 -7964 258914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 258294 686000 258914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 276294 -7964 276914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 276294 686000 276914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 294294 -7964 294914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 294294 686000 294914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 312294 -7964 312914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 312294 686000 312914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 330294 -7964 330914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 330294 686000 330914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 348294 -7964 348914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 348294 686000 348914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 366294 -7964 366914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 366294 686000 366914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 384294 -7964 384914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 384294 686000 384914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 402294 -7964 402914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 402294 686000 402914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 420294 -7964 420914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 420294 686000 420914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 438294 -7964 438914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 438294 686000 438914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 456294 -7964 456914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 456294 686000 456914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 474294 -7964 474914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 474294 686000 474914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 492294 -7964 492914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 492294 686000 492914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 510294 -7964 510914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 510294 686000 510914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 528294 -7964 528914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 528294 686000 528914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 546294 -7964 546914 14000 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 546294 686000 546914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 564294 -7964 564914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 582294 -7964 582914 711900 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 7366 592960 7986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 25366 592960 25986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 43366 592960 43986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 61366 592960 61986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 79366 592960 79986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 97366 592960 97986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 115366 592960 115986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 133366 592960 133986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 151366 592960 151986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 169366 592960 169986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 187366 592960 187986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 205366 592960 205986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 223366 592960 223986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 241366 592960 241986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 259366 592960 259986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 277366 592960 277986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 295366 592960 295986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 313366 592960 313986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 331366 592960 331986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 349366 592960 349986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 367366 592960 367986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 385366 592960 385986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 403366 592960 403986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 421366 592960 421986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 439366 592960 439986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 457366 592960 457986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 475366 592960 475986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 493366 592960 493986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 511366 592960 511986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 529366 592960 529986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 547366 592960 547986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 565366 592960 565986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 583366 592960 583986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 601366 592960 601986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 619366 592960 619986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 637366 592960 637986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 655366 592960 655986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 673366 592960 673986 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -9036 691366 592960 691986 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s -6156 -5084 -5536 709020 4 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -6156 -5084 590080 -4464 8 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -6156 708400 590080 709020 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 589460 -5084 590080 709020 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 10794 -7964 11414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 28794 -7964 29414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 28794 686000 29414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 46794 -7964 47414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 46794 686000 47414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 64794 -7964 65414 41000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 64794 686000 65414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 82794 -7964 83414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 82794 686000 83414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 100794 -7964 101414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 100794 686000 101414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 118794 -7964 119414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 118794 686000 119414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 136794 -7964 137414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 136794 686000 137414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 154794 -7964 155414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 154794 686000 155414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 172794 -7964 173414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 172794 686000 173414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 190794 -7964 191414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 190794 686000 191414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 208794 -7964 209414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 208794 686000 209414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 226794 -7964 227414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 226794 686000 227414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 244794 -7964 245414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 244794 686000 245414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 262794 -7964 263414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 262794 686000 263414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 280794 -7964 281414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 280794 686000 281414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 298794 -7964 299414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 298794 686000 299414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 316794 -7964 317414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 316794 686000 317414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 334794 -7964 335414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 334794 686000 335414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 352794 -7964 353414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 352794 686000 353414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 370794 -7964 371414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 370794 686000 371414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 388794 -7964 389414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 388794 686000 389414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 406794 -7964 407414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 406794 686000 407414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 424794 -7964 425414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 424794 686000 425414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 442794 -7964 443414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 442794 686000 443414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 460794 -7964 461414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 460794 686000 461414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 478794 -7964 479414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 478794 686000 479414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 496794 -7964 497414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 496794 686000 497414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 514794 -7964 515414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 514794 686000 515414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 532794 -7964 533414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 532794 686000 533414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 550794 -7964 551414 14000 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 550794 686000 551414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 568794 -7964 569414 711900 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 11866 592960 12486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 29866 592960 30486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 47866 592960 48486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 65866 592960 66486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 83866 592960 84486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 101866 592960 102486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 119866 592960 120486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 137866 592960 138486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 155866 592960 156486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 173866 592960 174486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 191866 592960 192486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 209866 592960 210486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 227866 592960 228486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 245866 592960 246486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 263866 592960 264486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 281866 592960 282486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 299866 592960 300486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 317866 592960 318486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 335866 592960 336486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 353866 592960 354486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 371866 592960 372486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 389866 592960 390486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 407866 592960 408486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 425866 592960 426486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 443866 592960 444486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 461866 592960 462486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 479866 592960 480486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 497866 592960 498486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 515866 592960 516486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 533866 592960 534486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 551866 592960 552486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 569866 592960 570486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 587866 592960 588486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 605866 592960 606486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 623866 592960 624486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 641866 592960 642486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 659866 592960 660486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 677866 592960 678486 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -9036 695866 592960 696486 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s -8076 -7004 -7456 710940 4 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8076 -7004 592000 -6384 8 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8076 710320 592000 710940 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 591380 -7004 592000 710940 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 15294 686000 15914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 33294 686000 33914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 51294 686000 51914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 69294 686000 69914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 87294 686000 87914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 105294 686000 105914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 123294 686000 123914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 141294 686000 141914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 159294 686000 159914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 177294 686000 177914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 195294 686000 195914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 213294 686000 213914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 231294 686000 231914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 249294 686000 249914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 267294 686000 267914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 285294 686000 285914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 303294 686000 303914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 321294 686000 321914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 339294 686000 339914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 357294 686000 357914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 375294 686000 375914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 393294 686000 393914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 411294 686000 411914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 429294 686000 429914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 447294 686000 447914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 465294 686000 465914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 483294 686000 483914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 501294 686000 501914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 519294 686000 519914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 537294 686000 537914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 555294 -7964 555914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 573294 -7964 573914 711900 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 16366 592960 16986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 34366 592960 34986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 52366 592960 52986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 70366 592960 70986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 88366 592960 88986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 106366 592960 106986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 124366 592960 124986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 142366 592960 142986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 160366 592960 160986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 178366 592960 178986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 196366 592960 196986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 214366 592960 214986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 232366 592960 232986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 250366 592960 250986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 268366 592960 268986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 286366 592960 286986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 304366 592960 304986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 322366 592960 322986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 340366 592960 340986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 358366 592960 358986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 376366 592960 376986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 394366 592960 394986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 412366 592960 412986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 430366 592960 430986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 448366 592960 448986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 466366 592960 466986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 484366 592960 484986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 502366 592960 502986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 520366 592960 520986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 538366 592960 538986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 556366 592960 556986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 574366 592960 574986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 592366 592960 592986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 610366 592960 610986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 628366 592960 628986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 646366 592960 646986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 664366 592960 664986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 682366 592960 682986 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -9036 700366 592960 700986 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s -7116 -6044 -6496 709980 4 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -7116 -6044 591040 -5424 8 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -7116 709360 591040 709980 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 590420 -6044 591040 709980 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 13044 -7964 13664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 31044 686000 31664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 49044 686000 49664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 67044 -7964 67664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 85044 686000 85664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 103044 686000 103664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 121044 -7964 121664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 139044 686000 139664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 157044 686000 157664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 175044 -7964 175664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 193044 686000 193664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 211044 686000 211664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 229044 -7964 229664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 247044 686000 247664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 265044 686000 265664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 283044 -7964 283664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 301044 686000 301664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 319044 686000 319664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 337044 -7964 337664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 355044 686000 355664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 373044 686000 373664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 391044 -7964 391664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 409044 686000 409664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 427044 686000 427664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 445044 -7964 445664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 463044 686000 463664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 481044 686000 481664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 499044 -7964 499664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 517044 686000 517664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 535044 686000 535664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 553044 -7964 553664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 571044 -7964 571664 711900 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 14116 592960 14736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 32116 592960 32736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 50116 592960 50736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 68116 592960 68736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 86116 592960 86736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 104116 592960 104736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 122116 592960 122736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 140116 592960 140736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 158116 592960 158736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 176116 592960 176736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 194116 592960 194736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 212116 592960 212736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 230116 592960 230736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 248116 592960 248736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 266116 592960 266736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 284116 592960 284736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 302116 592960 302736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 320116 592960 320736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 338116 592960 338736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 356116 592960 356736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 374116 592960 374736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 392116 592960 392736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 410116 592960 410736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 428116 592960 428736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 446116 592960 446736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 464116 592960 464736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 482116 592960 482736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 500116 592960 500736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 518116 592960 518736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 536116 592960 536736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 554116 592960 554736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 572116 592960 572736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 590116 592960 590736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 608116 592960 608736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 626116 592960 626736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 644116 592960 644736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 662116 592960 662736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 680116 592960 680736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -9036 698116 592960 698736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s -9036 -7964 -8416 711900 4 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 -7964 592960 -7344 8 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 711280 592960 711900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 592340 -7964 592960 711900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 557544 -7964 558164 711900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 575544 -7964 576164 711900 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 18616 592960 19236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 36616 592960 37236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 54616 592960 55236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 72616 592960 73236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 90616 592960 91236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 108616 592960 109236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 126616 592960 127236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 144616 592960 145236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 162616 592960 163236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 180616 592960 181236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 198616 592960 199236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 216616 592960 217236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 234616 592960 235236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 252616 592960 253236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 270616 592960 271236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 288616 592960 289236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 306616 592960 307236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 324616 592960 325236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 342616 592960 343236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 360616 592960 361236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 378616 592960 379236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 396616 592960 397236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 414616 592960 415236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 432616 592960 433236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 450616 592960 451236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 468616 592960 469236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 486616 592960 487236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 504616 592960 505236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 522616 592960 523236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 540616 592960 541236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 558616 592960 559236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 576616 592960 577236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 594616 592960 595236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 612616 592960 613236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 630616 592960 631236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 648616 592960 649236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 666616 592960 667236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -9036 684616 592960 685236 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s -3276 -2204 -2656 706140 4 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -3276 -2204 587200 -1584 8 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -3276 705520 587200 706140 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 586580 -2204 587200 706140 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 4044 -7964 4664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 22044 -7964 22664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 22044 686000 22664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 40044 -7964 40664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 40044 38000 40664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 58044 -7964 58664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 58044 686000 58664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 76044 -7964 76664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 76044 686000 76664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 94044 -7964 94664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 112044 -7964 112664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 112044 686000 112664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 130044 -7964 130664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 130044 686000 130664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 148044 -7964 148664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 166044 -7964 166664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 166044 686000 166664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 184044 -7964 184664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 184044 686000 184664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 202044 -7964 202664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 220044 -7964 220664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 220044 686000 220664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 238044 -7964 238664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 238044 686000 238664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 256044 -7964 256664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 274044 -7964 274664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 274044 686000 274664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 292044 -7964 292664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 292044 686000 292664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 310044 -7964 310664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 328044 -7964 328664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 328044 686000 328664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 346044 -7964 346664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 346044 686000 346664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 364044 -7964 364664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382044 -7964 382664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 382044 686000 382664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 400044 -7964 400664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 400044 686000 400664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 418044 -7964 418664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 436044 -7964 436664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 436044 686000 436664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 454044 -7964 454664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 454044 686000 454664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 472044 -7964 472664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 490044 -7964 490664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 490044 686000 490664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 508044 -7964 508664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 508044 686000 508664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 526044 -7964 526664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 544044 -7964 544664 14000 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 544044 686000 544664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 562044 -7964 562664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 580044 -7964 580664 711900 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 5116 592960 5736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 23116 592960 23736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 41116 592960 41736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 59116 592960 59736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 77116 592960 77736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 95116 592960 95736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 113116 592960 113736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 131116 592960 131736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 149116 592960 149736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 167116 592960 167736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 185116 592960 185736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 203116 592960 203736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 221116 592960 221736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 239116 592960 239736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 257116 592960 257736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 275116 592960 275736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 293116 592960 293736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 311116 592960 311736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 329116 592960 329736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 347116 592960 347736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 365116 592960 365736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 383116 592960 383736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 401116 592960 401736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 419116 592960 419736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 437116 592960 437736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 455116 592960 455736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 473116 592960 473736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 491116 592960 491736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 509116 592960 509736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 527116 592960 527736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 545116 592960 545736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 563116 592960 563736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 581116 592960 581736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 599116 592960 599736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 617116 592960 617736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 635116 592960 635736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 653116 592960 653736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 671116 592960 671736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -9036 689116 592960 689736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s -5196 -4124 -4576 708060 4 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5196 -4124 589120 -3504 8 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5196 707440 589120 708060 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 588500 -4124 589120 708060 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 8544 -7964 9164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 26544 -7964 27164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 26544 686000 27164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 44544 -7964 45164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 44544 686000 45164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 62544 -7964 63164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 62544 686000 63164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 80544 -7964 81164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 80544 686000 81164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 98544 -7964 99164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 98544 686000 99164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 116544 -7964 117164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 116544 686000 117164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 134544 -7964 135164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 134544 686000 135164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 152544 -7964 153164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 152544 686000 153164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 170544 -7964 171164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 170544 686000 171164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 188544 -7964 189164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 188544 686000 189164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 206544 -7964 207164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 206544 686000 207164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 224544 -7964 225164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 224544 686000 225164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 242544 -7964 243164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 242544 686000 243164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 260544 -7964 261164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 260544 686000 261164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 278544 -7964 279164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 278544 686000 279164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 296544 -7964 297164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 296544 686000 297164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 314544 -7964 315164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 314544 686000 315164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 332544 -7964 333164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 332544 686000 333164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 350544 -7964 351164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 350544 686000 351164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 368544 -7964 369164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 368544 686000 369164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 386544 -7964 387164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 386544 686000 387164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 404544 -7964 405164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 404544 686000 405164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 422544 -7964 423164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 422544 686000 423164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 440544 -7964 441164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 440544 686000 441164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 458544 -7964 459164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 458544 686000 459164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 476544 -7964 477164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 476544 686000 477164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 494544 -7964 495164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 494544 686000 495164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 512544 -7964 513164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 512544 686000 513164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 530544 -7964 531164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 530544 686000 531164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 548544 -7964 549164 14000 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 548544 686000 549164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 566544 -7964 567164 711900 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 9616 592960 10236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 27616 592960 28236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 45616 592960 46236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 63616 592960 64236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 81616 592960 82236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 99616 592960 100236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 117616 592960 118236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 135616 592960 136236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 153616 592960 154236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 171616 592960 172236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 189616 592960 190236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 207616 592960 208236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 225616 592960 226236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 243616 592960 244236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 261616 592960 262236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 279616 592960 280236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 297616 592960 298236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 315616 592960 316236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 333616 592960 334236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 351616 592960 352236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 369616 592960 370236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 387616 592960 388236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 405616 592960 406236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 423616 592960 424236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 441616 592960 442236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 459616 592960 460236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 477616 592960 478236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 495616 592960 496236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 513616 592960 514236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 531616 592960 532236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 549616 592960 550236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 567616 592960 568236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 585616 592960 586236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 603616 592960 604236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 621616 592960 622236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 639616 592960 640236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 657616 592960 658236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 675616 592960 676236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -9036 693616 592960 694236 6 vssd2
port 539 nsew ground bidirectional
rlabel metal2 s 19770 -960 19882 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 20874 -960 20986 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 21978 -960 22090 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 26394 -960 26506 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 63930 -960 64042 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 67242 -960 67354 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 70554 -960 70666 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 73866 -960 73978 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 77178 -960 77290 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 80490 -960 80602 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 87114 -960 87226 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 90426 -960 90538 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 93738 -960 93850 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 30810 -960 30922 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 97050 -960 97162 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 100362 -960 100474 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 103674 -960 103786 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 106986 -960 107098 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 110298 -960 110410 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 113610 -960 113722 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 116922 -960 117034 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 120234 -960 120346 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 123546 -960 123658 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 126858 -960 126970 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 35226 -960 35338 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 130170 -960 130282 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 133482 -960 133594 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 39642 -960 39754 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 44058 -960 44170 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 47370 -960 47482 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 50682 -960 50794 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 53994 -960 54106 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 57306 -960 57418 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 60618 -960 60730 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 23082 -960 23194 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 27498 -960 27610 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 65034 -960 65146 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 68346 -960 68458 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 71658 -960 71770 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 78282 -960 78394 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 81594 -960 81706 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 88218 -960 88330 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 94842 -960 94954 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 31914 -960 32026 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 98154 -960 98266 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 101466 -960 101578 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 104778 -960 104890 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 111402 -960 111514 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 118026 -960 118138 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 121338 -960 121450 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 127962 -960 128074 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 36330 -960 36442 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 131274 -960 131386 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 134586 -960 134698 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 40746 -960 40858 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 45162 -960 45274 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 48474 -960 48586 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 51786 -960 51898 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 55098 -960 55210 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 61722 -960 61834 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 28602 -960 28714 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 66138 -960 66250 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 69450 -960 69562 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 72762 -960 72874 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 76074 -960 76186 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 79386 -960 79498 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 82698 -960 82810 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 86010 -960 86122 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 89322 -960 89434 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 92634 -960 92746 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 95946 -960 96058 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 33018 -960 33130 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 102570 -960 102682 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 105882 -960 105994 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 109194 -960 109306 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 112506 -960 112618 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 115818 -960 115930 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 119130 -960 119242 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 122442 -960 122554 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 125754 -960 125866 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 129066 -960 129178 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 37434 -960 37546 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 132378 -960 132490 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 135690 -960 135802 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 46266 -960 46378 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 49578 -960 49690 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 52890 -960 53002 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 56202 -960 56314 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 59514 -960 59626 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 62826 -960 62938 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 29706 -960 29818 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 34122 -960 34234 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 38538 -960 38650 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 42954 -960 43066 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 24186 -960 24298 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5368500
string GDS_FILE /home/matt/work/asic-workshop/shuttle7/tiny-tapeout/openlane/user_project_wrapper/runs/22_08_02_11_52/results/signoff/user_project_wrapper.magic.gds
string GDS_START 1457838
<< end >>

