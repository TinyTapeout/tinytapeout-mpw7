* NGSPICE file created from user_project_wrapper.ext - technology: sky130B

* Black-box entry subcircuit for scan_wrapper_334445762078310996 abstract view
.subckt scan_wrapper_334445762078310996 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_335404063203000914 abstract view
.subckt scan_wrapper_335404063203000914 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_controller abstract view
.subckt scan_controller active_select[0] active_select[1] active_select[2] active_select[3]
+ active_select[4] active_select[5] active_select[6] active_select[7] active_select[8]
+ clk inputs[0] inputs[1] inputs[2] inputs[3] inputs[4] inputs[5] inputs[6] inputs[7]
+ oeb[0] oeb[1] oeb[2] oeb[3] oeb[4] oeb[5] oeb[6] oeb[7] oeb[8] outputs[0] outputs[1]
+ outputs[2] outputs[3] outputs[4] outputs[5] outputs[6] outputs[7] ready reset scan_clk
+ scan_data_in scan_data_out scan_latch_enable scan_select vccd1 vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xscan_wrapper_334445762078310996_397 scan_wrapper_334445762078310996_397/clk_in scan_wrapper_334445762078310996_398/clk_in
+ scan_wrapper_334445762078310996_397/data_in scan_wrapper_334445762078310996_398/data_in
+ scan_wrapper_334445762078310996_397/latch_enable_in scan_wrapper_334445762078310996_398/latch_enable_in
+ scan_wrapper_334445762078310996_397/scan_select_in scan_wrapper_334445762078310996_398/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_386 scan_wrapper_334445762078310996_386/clk_in scan_wrapper_334445762078310996_387/clk_in
+ scan_wrapper_334445762078310996_386/data_in scan_wrapper_334445762078310996_387/data_in
+ scan_wrapper_334445762078310996_386/latch_enable_in scan_wrapper_334445762078310996_387/latch_enable_in
+ scan_wrapper_334445762078310996_386/scan_select_in scan_wrapper_334445762078310996_387/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_320 scan_wrapper_334445762078310996_320/clk_in scan_wrapper_334445762078310996_321/clk_in
+ scan_wrapper_334445762078310996_320/data_in scan_wrapper_334445762078310996_321/data_in
+ scan_wrapper_334445762078310996_320/latch_enable_in scan_wrapper_334445762078310996_321/latch_enable_in
+ scan_wrapper_334445762078310996_320/scan_select_in scan_wrapper_334445762078310996_321/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_331 scan_wrapper_334445762078310996_331/clk_in scan_wrapper_334445762078310996_332/clk_in
+ scan_wrapper_334445762078310996_331/data_in scan_wrapper_334445762078310996_332/data_in
+ scan_wrapper_334445762078310996_331/latch_enable_in scan_wrapper_334445762078310996_332/latch_enable_in
+ scan_wrapper_334445762078310996_331/scan_select_in scan_wrapper_334445762078310996_332/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_342 scan_wrapper_334445762078310996_342/clk_in scan_wrapper_334445762078310996_343/clk_in
+ scan_wrapper_334445762078310996_342/data_in scan_wrapper_334445762078310996_343/data_in
+ scan_wrapper_334445762078310996_342/latch_enable_in scan_wrapper_334445762078310996_343/latch_enable_in
+ scan_wrapper_334445762078310996_342/scan_select_in scan_wrapper_334445762078310996_343/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_353 scan_wrapper_334445762078310996_353/clk_in scan_wrapper_334445762078310996_354/clk_in
+ scan_wrapper_334445762078310996_353/data_in scan_wrapper_334445762078310996_354/data_in
+ scan_wrapper_334445762078310996_353/latch_enable_in scan_wrapper_334445762078310996_354/latch_enable_in
+ scan_wrapper_334445762078310996_353/scan_select_in scan_wrapper_334445762078310996_354/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_364 scan_wrapper_334445762078310996_364/clk_in scan_wrapper_334445762078310996_365/clk_in
+ scan_wrapper_334445762078310996_364/data_in scan_wrapper_334445762078310996_365/data_in
+ scan_wrapper_334445762078310996_364/latch_enable_in scan_wrapper_334445762078310996_365/latch_enable_in
+ scan_wrapper_334445762078310996_364/scan_select_in scan_wrapper_334445762078310996_365/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_375 scan_wrapper_334445762078310996_375/clk_in scan_wrapper_334445762078310996_376/clk_in
+ scan_wrapper_334445762078310996_375/data_in scan_wrapper_334445762078310996_376/data_in
+ scan_wrapper_334445762078310996_375/latch_enable_in scan_wrapper_334445762078310996_376/latch_enable_in
+ scan_wrapper_334445762078310996_375/scan_select_in scan_wrapper_334445762078310996_376/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_150 scan_wrapper_334445762078310996_150/clk_in scan_wrapper_334445762078310996_151/clk_in
+ scan_wrapper_334445762078310996_150/data_in scan_wrapper_334445762078310996_151/data_in
+ scan_wrapper_334445762078310996_150/latch_enable_in scan_wrapper_334445762078310996_151/latch_enable_in
+ scan_wrapper_334445762078310996_150/scan_select_in scan_wrapper_334445762078310996_151/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_161 scan_wrapper_334445762078310996_161/clk_in scan_wrapper_334445762078310996_162/clk_in
+ scan_wrapper_334445762078310996_161/data_in scan_wrapper_334445762078310996_162/data_in
+ scan_wrapper_334445762078310996_161/latch_enable_in scan_wrapper_334445762078310996_162/latch_enable_in
+ scan_wrapper_334445762078310996_161/scan_select_in scan_wrapper_334445762078310996_162/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_172 scan_wrapper_334445762078310996_172/clk_in scan_wrapper_334445762078310996_173/clk_in
+ scan_wrapper_334445762078310996_172/data_in scan_wrapper_334445762078310996_173/data_in
+ scan_wrapper_334445762078310996_172/latch_enable_in scan_wrapper_334445762078310996_173/latch_enable_in
+ scan_wrapper_334445762078310996_172/scan_select_in scan_wrapper_334445762078310996_173/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_183 scan_wrapper_334445762078310996_183/clk_in scan_wrapper_334445762078310996_184/clk_in
+ scan_wrapper_334445762078310996_183/data_in scan_wrapper_334445762078310996_184/data_in
+ scan_wrapper_334445762078310996_183/latch_enable_in scan_wrapper_334445762078310996_184/latch_enable_in
+ scan_wrapper_334445762078310996_183/scan_select_in scan_wrapper_334445762078310996_184/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_194 scan_wrapper_334445762078310996_194/clk_in scan_wrapper_334445762078310996_195/clk_in
+ scan_wrapper_334445762078310996_194/data_in scan_wrapper_334445762078310996_195/data_in
+ scan_wrapper_334445762078310996_194/latch_enable_in scan_wrapper_334445762078310996_195/latch_enable_in
+ scan_wrapper_334445762078310996_194/scan_select_in scan_wrapper_334445762078310996_195/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_398 scan_wrapper_334445762078310996_398/clk_in scan_wrapper_334445762078310996_399/clk_in
+ scan_wrapper_334445762078310996_398/data_in scan_wrapper_334445762078310996_399/data_in
+ scan_wrapper_334445762078310996_398/latch_enable_in scan_wrapper_334445762078310996_399/latch_enable_in
+ scan_wrapper_334445762078310996_398/scan_select_in scan_wrapper_334445762078310996_399/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_387 scan_wrapper_334445762078310996_387/clk_in scan_wrapper_334445762078310996_388/clk_in
+ scan_wrapper_334445762078310996_387/data_in scan_wrapper_334445762078310996_388/data_in
+ scan_wrapper_334445762078310996_387/latch_enable_in scan_wrapper_334445762078310996_388/latch_enable_in
+ scan_wrapper_334445762078310996_387/scan_select_in scan_wrapper_334445762078310996_388/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_90 scan_wrapper_334445762078310996_90/clk_in scan_wrapper_334445762078310996_91/clk_in
+ scan_wrapper_334445762078310996_90/data_in scan_wrapper_334445762078310996_91/data_in
+ scan_wrapper_334445762078310996_90/latch_enable_in scan_wrapper_334445762078310996_91/latch_enable_in
+ scan_wrapper_334445762078310996_90/scan_select_in scan_wrapper_334445762078310996_91/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_310 scan_wrapper_334445762078310996_310/clk_in scan_wrapper_334445762078310996_311/clk_in
+ scan_wrapper_334445762078310996_310/data_in scan_wrapper_334445762078310996_311/data_in
+ scan_wrapper_334445762078310996_310/latch_enable_in scan_wrapper_334445762078310996_311/latch_enable_in
+ scan_wrapper_334445762078310996_310/scan_select_in scan_wrapper_334445762078310996_311/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_321 scan_wrapper_334445762078310996_321/clk_in scan_wrapper_334445762078310996_322/clk_in
+ scan_wrapper_334445762078310996_321/data_in scan_wrapper_334445762078310996_322/data_in
+ scan_wrapper_334445762078310996_321/latch_enable_in scan_wrapper_334445762078310996_322/latch_enable_in
+ scan_wrapper_334445762078310996_321/scan_select_in scan_wrapper_334445762078310996_322/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_332 scan_wrapper_334445762078310996_332/clk_in scan_wrapper_334445762078310996_333/clk_in
+ scan_wrapper_334445762078310996_332/data_in scan_wrapper_334445762078310996_333/data_in
+ scan_wrapper_334445762078310996_332/latch_enable_in scan_wrapper_334445762078310996_333/latch_enable_in
+ scan_wrapper_334445762078310996_332/scan_select_in scan_wrapper_334445762078310996_333/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_343 scan_wrapper_334445762078310996_343/clk_in scan_wrapper_334445762078310996_344/clk_in
+ scan_wrapper_334445762078310996_343/data_in scan_wrapper_334445762078310996_344/data_in
+ scan_wrapper_334445762078310996_343/latch_enable_in scan_wrapper_334445762078310996_344/latch_enable_in
+ scan_wrapper_334445762078310996_343/scan_select_in scan_wrapper_334445762078310996_344/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_354 scan_wrapper_334445762078310996_354/clk_in scan_wrapper_334445762078310996_355/clk_in
+ scan_wrapper_334445762078310996_354/data_in scan_wrapper_334445762078310996_355/data_in
+ scan_wrapper_334445762078310996_354/latch_enable_in scan_wrapper_334445762078310996_355/latch_enable_in
+ scan_wrapper_334445762078310996_354/scan_select_in scan_wrapper_334445762078310996_355/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_365 scan_wrapper_334445762078310996_365/clk_in scan_wrapper_334445762078310996_366/clk_in
+ scan_wrapper_334445762078310996_365/data_in scan_wrapper_334445762078310996_366/data_in
+ scan_wrapper_334445762078310996_365/latch_enable_in scan_wrapper_334445762078310996_366/latch_enable_in
+ scan_wrapper_334445762078310996_365/scan_select_in scan_wrapper_334445762078310996_366/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_376 scan_wrapper_334445762078310996_376/clk_in scan_wrapper_334445762078310996_377/clk_in
+ scan_wrapper_334445762078310996_376/data_in scan_wrapper_334445762078310996_377/data_in
+ scan_wrapper_334445762078310996_376/latch_enable_in scan_wrapper_334445762078310996_377/latch_enable_in
+ scan_wrapper_334445762078310996_376/scan_select_in scan_wrapper_334445762078310996_377/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_140 scan_wrapper_334445762078310996_140/clk_in scan_wrapper_334445762078310996_141/clk_in
+ scan_wrapper_334445762078310996_140/data_in scan_wrapper_334445762078310996_141/data_in
+ scan_wrapper_334445762078310996_140/latch_enable_in scan_wrapper_334445762078310996_141/latch_enable_in
+ scan_wrapper_334445762078310996_140/scan_select_in scan_wrapper_334445762078310996_141/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_151 scan_wrapper_334445762078310996_151/clk_in scan_wrapper_334445762078310996_152/clk_in
+ scan_wrapper_334445762078310996_151/data_in scan_wrapper_334445762078310996_152/data_in
+ scan_wrapper_334445762078310996_151/latch_enable_in scan_wrapper_334445762078310996_152/latch_enable_in
+ scan_wrapper_334445762078310996_151/scan_select_in scan_wrapper_334445762078310996_152/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_162 scan_wrapper_334445762078310996_162/clk_in scan_wrapper_334445762078310996_163/clk_in
+ scan_wrapper_334445762078310996_162/data_in scan_wrapper_334445762078310996_163/data_in
+ scan_wrapper_334445762078310996_162/latch_enable_in scan_wrapper_334445762078310996_163/latch_enable_in
+ scan_wrapper_334445762078310996_162/scan_select_in scan_wrapper_334445762078310996_163/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_173 scan_wrapper_334445762078310996_173/clk_in scan_wrapper_334445762078310996_174/clk_in
+ scan_wrapper_334445762078310996_173/data_in scan_wrapper_334445762078310996_174/data_in
+ scan_wrapper_334445762078310996_173/latch_enable_in scan_wrapper_334445762078310996_174/latch_enable_in
+ scan_wrapper_334445762078310996_173/scan_select_in scan_wrapper_334445762078310996_174/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_184 scan_wrapper_334445762078310996_184/clk_in scan_wrapper_334445762078310996_185/clk_in
+ scan_wrapper_334445762078310996_184/data_in scan_wrapper_334445762078310996_185/data_in
+ scan_wrapper_334445762078310996_184/latch_enable_in scan_wrapper_334445762078310996_185/latch_enable_in
+ scan_wrapper_334445762078310996_184/scan_select_in scan_wrapper_334445762078310996_185/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_195 scan_wrapper_334445762078310996_195/clk_in scan_wrapper_334445762078310996_196/clk_in
+ scan_wrapper_334445762078310996_195/data_in scan_wrapper_334445762078310996_196/data_in
+ scan_wrapper_334445762078310996_195/latch_enable_in scan_wrapper_334445762078310996_196/latch_enable_in
+ scan_wrapper_334445762078310996_195/scan_select_in scan_wrapper_334445762078310996_196/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_399 scan_wrapper_334445762078310996_399/clk_in scan_wrapper_334445762078310996_400/clk_in
+ scan_wrapper_334445762078310996_399/data_in scan_wrapper_334445762078310996_400/data_in
+ scan_wrapper_334445762078310996_399/latch_enable_in scan_wrapper_334445762078310996_400/latch_enable_in
+ scan_wrapper_334445762078310996_399/scan_select_in scan_wrapper_334445762078310996_400/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_388 scan_wrapper_334445762078310996_388/clk_in scan_wrapper_334445762078310996_389/clk_in
+ scan_wrapper_334445762078310996_388/data_in scan_wrapper_334445762078310996_389/data_in
+ scan_wrapper_334445762078310996_388/latch_enable_in scan_wrapper_334445762078310996_389/latch_enable_in
+ scan_wrapper_334445762078310996_388/scan_select_in scan_wrapper_334445762078310996_389/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_91 scan_wrapper_334445762078310996_91/clk_in scan_wrapper_334445762078310996_92/clk_in
+ scan_wrapper_334445762078310996_91/data_in scan_wrapper_334445762078310996_92/data_in
+ scan_wrapper_334445762078310996_91/latch_enable_in scan_wrapper_334445762078310996_92/latch_enable_in
+ scan_wrapper_334445762078310996_91/scan_select_in scan_wrapper_334445762078310996_92/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_80 scan_wrapper_334445762078310996_80/clk_in scan_wrapper_334445762078310996_81/clk_in
+ scan_wrapper_334445762078310996_80/data_in scan_wrapper_334445762078310996_81/data_in
+ scan_wrapper_334445762078310996_80/latch_enable_in scan_wrapper_334445762078310996_81/latch_enable_in
+ scan_wrapper_334445762078310996_80/scan_select_in scan_wrapper_334445762078310996_81/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_300 scan_wrapper_334445762078310996_300/clk_in scan_wrapper_334445762078310996_301/clk_in
+ scan_wrapper_334445762078310996_300/data_in scan_wrapper_334445762078310996_301/data_in
+ scan_wrapper_334445762078310996_300/latch_enable_in scan_wrapper_334445762078310996_301/latch_enable_in
+ scan_wrapper_334445762078310996_300/scan_select_in scan_wrapper_334445762078310996_301/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_311 scan_wrapper_334445762078310996_311/clk_in scan_wrapper_334445762078310996_312/clk_in
+ scan_wrapper_334445762078310996_311/data_in scan_wrapper_334445762078310996_312/data_in
+ scan_wrapper_334445762078310996_311/latch_enable_in scan_wrapper_334445762078310996_312/latch_enable_in
+ scan_wrapper_334445762078310996_311/scan_select_in scan_wrapper_334445762078310996_312/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_322 scan_wrapper_334445762078310996_322/clk_in scan_wrapper_334445762078310996_323/clk_in
+ scan_wrapper_334445762078310996_322/data_in scan_wrapper_334445762078310996_323/data_in
+ scan_wrapper_334445762078310996_322/latch_enable_in scan_wrapper_334445762078310996_323/latch_enable_in
+ scan_wrapper_334445762078310996_322/scan_select_in scan_wrapper_334445762078310996_323/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_333 scan_wrapper_334445762078310996_333/clk_in scan_wrapper_334445762078310996_334/clk_in
+ scan_wrapper_334445762078310996_333/data_in scan_wrapper_334445762078310996_334/data_in
+ scan_wrapper_334445762078310996_333/latch_enable_in scan_wrapper_334445762078310996_334/latch_enable_in
+ scan_wrapper_334445762078310996_333/scan_select_in scan_wrapper_334445762078310996_334/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_344 scan_wrapper_334445762078310996_344/clk_in scan_wrapper_334445762078310996_345/clk_in
+ scan_wrapper_334445762078310996_344/data_in scan_wrapper_334445762078310996_345/data_in
+ scan_wrapper_334445762078310996_344/latch_enable_in scan_wrapper_334445762078310996_345/latch_enable_in
+ scan_wrapper_334445762078310996_344/scan_select_in scan_wrapper_334445762078310996_345/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_355 scan_wrapper_334445762078310996_355/clk_in scan_wrapper_334445762078310996_356/clk_in
+ scan_wrapper_334445762078310996_355/data_in scan_wrapper_334445762078310996_356/data_in
+ scan_wrapper_334445762078310996_355/latch_enable_in scan_wrapper_334445762078310996_356/latch_enable_in
+ scan_wrapper_334445762078310996_355/scan_select_in scan_wrapper_334445762078310996_356/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_366 scan_wrapper_334445762078310996_366/clk_in scan_wrapper_334445762078310996_367/clk_in
+ scan_wrapper_334445762078310996_366/data_in scan_wrapper_334445762078310996_367/data_in
+ scan_wrapper_334445762078310996_366/latch_enable_in scan_wrapper_334445762078310996_367/latch_enable_in
+ scan_wrapper_334445762078310996_366/scan_select_in scan_wrapper_334445762078310996_367/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_377 scan_wrapper_334445762078310996_377/clk_in scan_wrapper_334445762078310996_378/clk_in
+ scan_wrapper_334445762078310996_377/data_in scan_wrapper_334445762078310996_378/data_in
+ scan_wrapper_334445762078310996_377/latch_enable_in scan_wrapper_334445762078310996_378/latch_enable_in
+ scan_wrapper_334445762078310996_377/scan_select_in scan_wrapper_334445762078310996_378/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_130 scan_wrapper_334445762078310996_130/clk_in scan_wrapper_334445762078310996_131/clk_in
+ scan_wrapper_334445762078310996_130/data_in scan_wrapper_334445762078310996_131/data_in
+ scan_wrapper_334445762078310996_130/latch_enable_in scan_wrapper_334445762078310996_131/latch_enable_in
+ scan_wrapper_334445762078310996_130/scan_select_in scan_wrapper_334445762078310996_131/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_141 scan_wrapper_334445762078310996_141/clk_in scan_wrapper_334445762078310996_142/clk_in
+ scan_wrapper_334445762078310996_141/data_in scan_wrapper_334445762078310996_142/data_in
+ scan_wrapper_334445762078310996_141/latch_enable_in scan_wrapper_334445762078310996_142/latch_enable_in
+ scan_wrapper_334445762078310996_141/scan_select_in scan_wrapper_334445762078310996_142/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_152 scan_wrapper_334445762078310996_152/clk_in scan_wrapper_334445762078310996_153/clk_in
+ scan_wrapper_334445762078310996_152/data_in scan_wrapper_334445762078310996_153/data_in
+ scan_wrapper_334445762078310996_152/latch_enable_in scan_wrapper_334445762078310996_153/latch_enable_in
+ scan_wrapper_334445762078310996_152/scan_select_in scan_wrapper_334445762078310996_153/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_163 scan_wrapper_334445762078310996_163/clk_in scan_wrapper_334445762078310996_164/clk_in
+ scan_wrapper_334445762078310996_163/data_in scan_wrapper_334445762078310996_164/data_in
+ scan_wrapper_334445762078310996_163/latch_enable_in scan_wrapper_334445762078310996_164/latch_enable_in
+ scan_wrapper_334445762078310996_163/scan_select_in scan_wrapper_334445762078310996_164/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_174 scan_wrapper_334445762078310996_174/clk_in scan_wrapper_334445762078310996_175/clk_in
+ scan_wrapper_334445762078310996_174/data_in scan_wrapper_334445762078310996_175/data_in
+ scan_wrapper_334445762078310996_174/latch_enable_in scan_wrapper_334445762078310996_175/latch_enable_in
+ scan_wrapper_334445762078310996_174/scan_select_in scan_wrapper_334445762078310996_175/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_185 scan_wrapper_334445762078310996_185/clk_in scan_wrapper_334445762078310996_186/clk_in
+ scan_wrapper_334445762078310996_185/data_in scan_wrapper_334445762078310996_186/data_in
+ scan_wrapper_334445762078310996_185/latch_enable_in scan_wrapper_334445762078310996_186/latch_enable_in
+ scan_wrapper_334445762078310996_185/scan_select_in scan_wrapper_334445762078310996_186/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_196 scan_wrapper_334445762078310996_196/clk_in scan_wrapper_334445762078310996_197/clk_in
+ scan_wrapper_334445762078310996_196/data_in scan_wrapper_334445762078310996_197/data_in
+ scan_wrapper_334445762078310996_196/latch_enable_in scan_wrapper_334445762078310996_197/latch_enable_in
+ scan_wrapper_334445762078310996_196/scan_select_in scan_wrapper_334445762078310996_197/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_92 scan_wrapper_334445762078310996_92/clk_in scan_wrapper_334445762078310996_93/clk_in
+ scan_wrapper_334445762078310996_92/data_in scan_wrapper_334445762078310996_93/data_in
+ scan_wrapper_334445762078310996_92/latch_enable_in scan_wrapper_334445762078310996_93/latch_enable_in
+ scan_wrapper_334445762078310996_92/scan_select_in scan_wrapper_334445762078310996_93/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_81 scan_wrapper_334445762078310996_81/clk_in scan_wrapper_334445762078310996_82/clk_in
+ scan_wrapper_334445762078310996_81/data_in scan_wrapper_334445762078310996_82/data_in
+ scan_wrapper_334445762078310996_81/latch_enable_in scan_wrapper_334445762078310996_82/latch_enable_in
+ scan_wrapper_334445762078310996_81/scan_select_in scan_wrapper_334445762078310996_82/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_70 scan_wrapper_334445762078310996_70/clk_in scan_wrapper_334445762078310996_71/clk_in
+ scan_wrapper_334445762078310996_70/data_in scan_wrapper_334445762078310996_71/data_in
+ scan_wrapper_334445762078310996_70/latch_enable_in scan_wrapper_334445762078310996_71/latch_enable_in
+ scan_wrapper_334445762078310996_70/scan_select_in scan_wrapper_334445762078310996_71/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_301 scan_wrapper_334445762078310996_301/clk_in scan_wrapper_334445762078310996_302/clk_in
+ scan_wrapper_334445762078310996_301/data_in scan_wrapper_334445762078310996_302/data_in
+ scan_wrapper_334445762078310996_301/latch_enable_in scan_wrapper_334445762078310996_302/latch_enable_in
+ scan_wrapper_334445762078310996_301/scan_select_in scan_wrapper_334445762078310996_302/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_312 scan_wrapper_334445762078310996_312/clk_in scan_wrapper_334445762078310996_313/clk_in
+ scan_wrapper_334445762078310996_312/data_in scan_wrapper_334445762078310996_313/data_in
+ scan_wrapper_334445762078310996_312/latch_enable_in scan_wrapper_334445762078310996_313/latch_enable_in
+ scan_wrapper_334445762078310996_312/scan_select_in scan_wrapper_334445762078310996_313/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_323 scan_wrapper_334445762078310996_323/clk_in scan_wrapper_334445762078310996_324/clk_in
+ scan_wrapper_334445762078310996_323/data_in scan_wrapper_334445762078310996_324/data_in
+ scan_wrapper_334445762078310996_323/latch_enable_in scan_wrapper_334445762078310996_324/latch_enable_in
+ scan_wrapper_334445762078310996_323/scan_select_in scan_wrapper_334445762078310996_324/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_389 scan_wrapper_334445762078310996_389/clk_in scan_wrapper_334445762078310996_390/clk_in
+ scan_wrapper_334445762078310996_389/data_in scan_wrapper_334445762078310996_390/data_in
+ scan_wrapper_334445762078310996_389/latch_enable_in scan_wrapper_334445762078310996_390/latch_enable_in
+ scan_wrapper_334445762078310996_389/scan_select_in scan_wrapper_334445762078310996_390/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_334 scan_wrapper_334445762078310996_334/clk_in scan_wrapper_334445762078310996_335/clk_in
+ scan_wrapper_334445762078310996_334/data_in scan_wrapper_334445762078310996_335/data_in
+ scan_wrapper_334445762078310996_334/latch_enable_in scan_wrapper_334445762078310996_335/latch_enable_in
+ scan_wrapper_334445762078310996_334/scan_select_in scan_wrapper_334445762078310996_335/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_345 scan_wrapper_334445762078310996_345/clk_in scan_wrapper_334445762078310996_346/clk_in
+ scan_wrapper_334445762078310996_345/data_in scan_wrapper_334445762078310996_346/data_in
+ scan_wrapper_334445762078310996_345/latch_enable_in scan_wrapper_334445762078310996_346/latch_enable_in
+ scan_wrapper_334445762078310996_345/scan_select_in scan_wrapper_334445762078310996_346/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_356 scan_wrapper_334445762078310996_356/clk_in scan_wrapper_334445762078310996_357/clk_in
+ scan_wrapper_334445762078310996_356/data_in scan_wrapper_334445762078310996_357/data_in
+ scan_wrapper_334445762078310996_356/latch_enable_in scan_wrapper_334445762078310996_357/latch_enable_in
+ scan_wrapper_334445762078310996_356/scan_select_in scan_wrapper_334445762078310996_357/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_367 scan_wrapper_334445762078310996_367/clk_in scan_wrapper_334445762078310996_368/clk_in
+ scan_wrapper_334445762078310996_367/data_in scan_wrapper_334445762078310996_368/data_in
+ scan_wrapper_334445762078310996_367/latch_enable_in scan_wrapper_334445762078310996_368/latch_enable_in
+ scan_wrapper_334445762078310996_367/scan_select_in scan_wrapper_334445762078310996_368/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_378 scan_wrapper_334445762078310996_378/clk_in scan_wrapper_334445762078310996_379/clk_in
+ scan_wrapper_334445762078310996_378/data_in scan_wrapper_334445762078310996_379/data_in
+ scan_wrapper_334445762078310996_378/latch_enable_in scan_wrapper_334445762078310996_379/latch_enable_in
+ scan_wrapper_334445762078310996_378/scan_select_in scan_wrapper_334445762078310996_379/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_120 scan_wrapper_334445762078310996_120/clk_in scan_wrapper_334445762078310996_121/clk_in
+ scan_wrapper_334445762078310996_120/data_in scan_wrapper_334445762078310996_121/data_in
+ scan_wrapper_334445762078310996_120/latch_enable_in scan_wrapper_334445762078310996_121/latch_enable_in
+ scan_wrapper_334445762078310996_120/scan_select_in scan_wrapper_334445762078310996_121/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_131 scan_wrapper_334445762078310996_131/clk_in scan_wrapper_334445762078310996_132/clk_in
+ scan_wrapper_334445762078310996_131/data_in scan_wrapper_334445762078310996_132/data_in
+ scan_wrapper_334445762078310996_131/latch_enable_in scan_wrapper_334445762078310996_132/latch_enable_in
+ scan_wrapper_334445762078310996_131/scan_select_in scan_wrapper_334445762078310996_132/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_142 scan_wrapper_334445762078310996_142/clk_in scan_wrapper_334445762078310996_143/clk_in
+ scan_wrapper_334445762078310996_142/data_in scan_wrapper_334445762078310996_143/data_in
+ scan_wrapper_334445762078310996_142/latch_enable_in scan_wrapper_334445762078310996_143/latch_enable_in
+ scan_wrapper_334445762078310996_142/scan_select_in scan_wrapper_334445762078310996_143/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_153 scan_wrapper_334445762078310996_153/clk_in scan_wrapper_334445762078310996_154/clk_in
+ scan_wrapper_334445762078310996_153/data_in scan_wrapper_334445762078310996_154/data_in
+ scan_wrapper_334445762078310996_153/latch_enable_in scan_wrapper_334445762078310996_154/latch_enable_in
+ scan_wrapper_334445762078310996_153/scan_select_in scan_wrapper_334445762078310996_154/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_164 scan_wrapper_334445762078310996_164/clk_in scan_wrapper_334445762078310996_165/clk_in
+ scan_wrapper_334445762078310996_164/data_in scan_wrapper_334445762078310996_165/data_in
+ scan_wrapper_334445762078310996_164/latch_enable_in scan_wrapper_334445762078310996_165/latch_enable_in
+ scan_wrapper_334445762078310996_164/scan_select_in scan_wrapper_334445762078310996_165/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_175 scan_wrapper_334445762078310996_175/clk_in scan_wrapper_334445762078310996_176/clk_in
+ scan_wrapper_334445762078310996_175/data_in scan_wrapper_334445762078310996_176/data_in
+ scan_wrapper_334445762078310996_175/latch_enable_in scan_wrapper_334445762078310996_176/latch_enable_in
+ scan_wrapper_334445762078310996_175/scan_select_in scan_wrapper_334445762078310996_176/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_186 scan_wrapper_334445762078310996_186/clk_in scan_wrapper_334445762078310996_187/clk_in
+ scan_wrapper_334445762078310996_186/data_in scan_wrapper_334445762078310996_187/data_in
+ scan_wrapper_334445762078310996_186/latch_enable_in scan_wrapper_334445762078310996_187/latch_enable_in
+ scan_wrapper_334445762078310996_186/scan_select_in scan_wrapper_334445762078310996_187/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_197 scan_wrapper_334445762078310996_197/clk_in scan_wrapper_334445762078310996_198/clk_in
+ scan_wrapper_334445762078310996_197/data_in scan_wrapper_334445762078310996_198/data_in
+ scan_wrapper_334445762078310996_197/latch_enable_in scan_wrapper_334445762078310996_198/latch_enable_in
+ scan_wrapper_334445762078310996_197/scan_select_in scan_wrapper_334445762078310996_198/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_93 scan_wrapper_334445762078310996_93/clk_in scan_wrapper_334445762078310996_94/clk_in
+ scan_wrapper_334445762078310996_93/data_in scan_wrapper_334445762078310996_94/data_in
+ scan_wrapper_334445762078310996_93/latch_enable_in scan_wrapper_334445762078310996_94/latch_enable_in
+ scan_wrapper_334445762078310996_93/scan_select_in scan_wrapper_334445762078310996_94/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_82 scan_wrapper_334445762078310996_82/clk_in scan_wrapper_334445762078310996_83/clk_in
+ scan_wrapper_334445762078310996_82/data_in scan_wrapper_334445762078310996_83/data_in
+ scan_wrapper_334445762078310996_82/latch_enable_in scan_wrapper_334445762078310996_83/latch_enable_in
+ scan_wrapper_334445762078310996_82/scan_select_in scan_wrapper_334445762078310996_83/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_71 scan_wrapper_334445762078310996_71/clk_in scan_wrapper_334445762078310996_72/clk_in
+ scan_wrapper_334445762078310996_71/data_in scan_wrapper_334445762078310996_72/data_in
+ scan_wrapper_334445762078310996_71/latch_enable_in scan_wrapper_334445762078310996_72/latch_enable_in
+ scan_wrapper_334445762078310996_71/scan_select_in scan_wrapper_334445762078310996_72/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_60 scan_wrapper_334445762078310996_60/clk_in scan_wrapper_334445762078310996_61/clk_in
+ scan_wrapper_334445762078310996_60/data_in scan_wrapper_334445762078310996_61/data_in
+ scan_wrapper_334445762078310996_60/latch_enable_in scan_wrapper_334445762078310996_61/latch_enable_in
+ scan_wrapper_334445762078310996_60/scan_select_in scan_wrapper_334445762078310996_61/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_302 scan_wrapper_334445762078310996_302/clk_in scan_wrapper_334445762078310996_303/clk_in
+ scan_wrapper_334445762078310996_302/data_in scan_wrapper_334445762078310996_303/data_in
+ scan_wrapper_334445762078310996_302/latch_enable_in scan_wrapper_334445762078310996_303/latch_enable_in
+ scan_wrapper_334445762078310996_302/scan_select_in scan_wrapper_334445762078310996_303/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_313 scan_wrapper_334445762078310996_313/clk_in scan_wrapper_334445762078310996_314/clk_in
+ scan_wrapper_334445762078310996_313/data_in scan_wrapper_334445762078310996_314/data_in
+ scan_wrapper_334445762078310996_313/latch_enable_in scan_wrapper_334445762078310996_314/latch_enable_in
+ scan_wrapper_334445762078310996_313/scan_select_in scan_wrapper_334445762078310996_314/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_324 scan_wrapper_334445762078310996_324/clk_in scan_wrapper_334445762078310996_325/clk_in
+ scan_wrapper_334445762078310996_324/data_in scan_wrapper_334445762078310996_325/data_in
+ scan_wrapper_334445762078310996_324/latch_enable_in scan_wrapper_334445762078310996_325/latch_enable_in
+ scan_wrapper_334445762078310996_324/scan_select_in scan_wrapper_334445762078310996_325/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_335 scan_wrapper_334445762078310996_335/clk_in scan_wrapper_334445762078310996_336/clk_in
+ scan_wrapper_334445762078310996_335/data_in scan_wrapper_334445762078310996_336/data_in
+ scan_wrapper_334445762078310996_335/latch_enable_in scan_wrapper_334445762078310996_336/latch_enable_in
+ scan_wrapper_334445762078310996_335/scan_select_in scan_wrapper_334445762078310996_336/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_346 scan_wrapper_334445762078310996_346/clk_in scan_wrapper_334445762078310996_347/clk_in
+ scan_wrapper_334445762078310996_346/data_in scan_wrapper_334445762078310996_347/data_in
+ scan_wrapper_334445762078310996_346/latch_enable_in scan_wrapper_334445762078310996_347/latch_enable_in
+ scan_wrapper_334445762078310996_346/scan_select_in scan_wrapper_334445762078310996_347/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_357 scan_wrapper_334445762078310996_357/clk_in scan_wrapper_334445762078310996_358/clk_in
+ scan_wrapper_334445762078310996_357/data_in scan_wrapper_334445762078310996_358/data_in
+ scan_wrapper_334445762078310996_357/latch_enable_in scan_wrapper_334445762078310996_358/latch_enable_in
+ scan_wrapper_334445762078310996_357/scan_select_in scan_wrapper_334445762078310996_358/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_368 scan_wrapper_334445762078310996_368/clk_in scan_wrapper_334445762078310996_369/clk_in
+ scan_wrapper_334445762078310996_368/data_in scan_wrapper_334445762078310996_369/data_in
+ scan_wrapper_334445762078310996_368/latch_enable_in scan_wrapper_334445762078310996_369/latch_enable_in
+ scan_wrapper_334445762078310996_368/scan_select_in scan_wrapper_334445762078310996_369/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_379 scan_wrapper_334445762078310996_379/clk_in scan_wrapper_334445762078310996_380/clk_in
+ scan_wrapper_334445762078310996_379/data_in scan_wrapper_334445762078310996_380/data_in
+ scan_wrapper_334445762078310996_379/latch_enable_in scan_wrapper_334445762078310996_380/latch_enable_in
+ scan_wrapper_334445762078310996_379/scan_select_in scan_wrapper_334445762078310996_380/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_110 scan_wrapper_334445762078310996_110/clk_in scan_wrapper_334445762078310996_111/clk_in
+ scan_wrapper_334445762078310996_110/data_in scan_wrapper_334445762078310996_111/data_in
+ scan_wrapper_334445762078310996_110/latch_enable_in scan_wrapper_334445762078310996_111/latch_enable_in
+ scan_wrapper_334445762078310996_110/scan_select_in scan_wrapper_334445762078310996_111/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_121 scan_wrapper_334445762078310996_121/clk_in scan_wrapper_334445762078310996_122/clk_in
+ scan_wrapper_334445762078310996_121/data_in scan_wrapper_334445762078310996_122/data_in
+ scan_wrapper_334445762078310996_121/latch_enable_in scan_wrapper_334445762078310996_122/latch_enable_in
+ scan_wrapper_334445762078310996_121/scan_select_in scan_wrapper_334445762078310996_122/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_132 scan_wrapper_334445762078310996_132/clk_in scan_wrapper_334445762078310996_133/clk_in
+ scan_wrapper_334445762078310996_132/data_in scan_wrapper_334445762078310996_133/data_in
+ scan_wrapper_334445762078310996_132/latch_enable_in scan_wrapper_334445762078310996_133/latch_enable_in
+ scan_wrapper_334445762078310996_132/scan_select_in scan_wrapper_334445762078310996_133/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_143 scan_wrapper_334445762078310996_143/clk_in scan_wrapper_334445762078310996_144/clk_in
+ scan_wrapper_334445762078310996_143/data_in scan_wrapper_334445762078310996_144/data_in
+ scan_wrapper_334445762078310996_143/latch_enable_in scan_wrapper_334445762078310996_144/latch_enable_in
+ scan_wrapper_334445762078310996_143/scan_select_in scan_wrapper_334445762078310996_144/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_154 scan_wrapper_334445762078310996_154/clk_in scan_wrapper_334445762078310996_155/clk_in
+ scan_wrapper_334445762078310996_154/data_in scan_wrapper_334445762078310996_155/data_in
+ scan_wrapper_334445762078310996_154/latch_enable_in scan_wrapper_334445762078310996_155/latch_enable_in
+ scan_wrapper_334445762078310996_154/scan_select_in scan_wrapper_334445762078310996_155/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_165 scan_wrapper_334445762078310996_165/clk_in scan_wrapper_334445762078310996_166/clk_in
+ scan_wrapper_334445762078310996_165/data_in scan_wrapper_334445762078310996_166/data_in
+ scan_wrapper_334445762078310996_165/latch_enable_in scan_wrapper_334445762078310996_166/latch_enable_in
+ scan_wrapper_334445762078310996_165/scan_select_in scan_wrapper_334445762078310996_166/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_176 scan_wrapper_334445762078310996_176/clk_in scan_wrapper_334445762078310996_177/clk_in
+ scan_wrapper_334445762078310996_176/data_in scan_wrapper_334445762078310996_177/data_in
+ scan_wrapper_334445762078310996_176/latch_enable_in scan_wrapper_334445762078310996_177/latch_enable_in
+ scan_wrapper_334445762078310996_176/scan_select_in scan_wrapper_334445762078310996_177/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_187 scan_wrapper_334445762078310996_187/clk_in scan_wrapper_334445762078310996_188/clk_in
+ scan_wrapper_334445762078310996_187/data_in scan_wrapper_334445762078310996_188/data_in
+ scan_wrapper_334445762078310996_187/latch_enable_in scan_wrapper_334445762078310996_188/latch_enable_in
+ scan_wrapper_334445762078310996_187/scan_select_in scan_wrapper_334445762078310996_188/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_198 scan_wrapper_334445762078310996_198/clk_in scan_wrapper_334445762078310996_199/clk_in
+ scan_wrapper_334445762078310996_198/data_in scan_wrapper_334445762078310996_199/data_in
+ scan_wrapper_334445762078310996_198/latch_enable_in scan_wrapper_334445762078310996_199/latch_enable_in
+ scan_wrapper_334445762078310996_198/scan_select_in scan_wrapper_334445762078310996_199/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_94 scan_wrapper_334445762078310996_94/clk_in scan_wrapper_334445762078310996_95/clk_in
+ scan_wrapper_334445762078310996_94/data_in scan_wrapper_334445762078310996_95/data_in
+ scan_wrapper_334445762078310996_94/latch_enable_in scan_wrapper_334445762078310996_95/latch_enable_in
+ scan_wrapper_334445762078310996_94/scan_select_in scan_wrapper_334445762078310996_95/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_83 scan_wrapper_334445762078310996_83/clk_in scan_wrapper_334445762078310996_84/clk_in
+ scan_wrapper_334445762078310996_83/data_in scan_wrapper_334445762078310996_84/data_in
+ scan_wrapper_334445762078310996_83/latch_enable_in scan_wrapper_334445762078310996_84/latch_enable_in
+ scan_wrapper_334445762078310996_83/scan_select_in scan_wrapper_334445762078310996_84/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_72 scan_wrapper_334445762078310996_72/clk_in scan_wrapper_334445762078310996_73/clk_in
+ scan_wrapper_334445762078310996_72/data_in scan_wrapper_334445762078310996_73/data_in
+ scan_wrapper_334445762078310996_72/latch_enable_in scan_wrapper_334445762078310996_73/latch_enable_in
+ scan_wrapper_334445762078310996_72/scan_select_in scan_wrapper_334445762078310996_73/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_61 scan_wrapper_334445762078310996_61/clk_in scan_wrapper_334445762078310996_62/clk_in
+ scan_wrapper_334445762078310996_61/data_in scan_wrapper_334445762078310996_62/data_in
+ scan_wrapper_334445762078310996_61/latch_enable_in scan_wrapper_334445762078310996_62/latch_enable_in
+ scan_wrapper_334445762078310996_61/scan_select_in scan_wrapper_334445762078310996_62/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_50 scan_wrapper_334445762078310996_50/clk_in scan_wrapper_334445762078310996_51/clk_in
+ scan_wrapper_334445762078310996_50/data_in scan_wrapper_334445762078310996_51/data_in
+ scan_wrapper_334445762078310996_50/latch_enable_in scan_wrapper_334445762078310996_51/latch_enable_in
+ scan_wrapper_334445762078310996_50/scan_select_in scan_wrapper_334445762078310996_51/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_303 scan_wrapper_334445762078310996_303/clk_in scan_wrapper_334445762078310996_304/clk_in
+ scan_wrapper_334445762078310996_303/data_in scan_wrapper_334445762078310996_304/data_in
+ scan_wrapper_334445762078310996_303/latch_enable_in scan_wrapper_334445762078310996_304/latch_enable_in
+ scan_wrapper_334445762078310996_303/scan_select_in scan_wrapper_334445762078310996_304/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_314 scan_wrapper_334445762078310996_314/clk_in scan_wrapper_334445762078310996_315/clk_in
+ scan_wrapper_334445762078310996_314/data_in scan_wrapper_334445762078310996_315/data_in
+ scan_wrapper_334445762078310996_314/latch_enable_in scan_wrapper_334445762078310996_315/latch_enable_in
+ scan_wrapper_334445762078310996_314/scan_select_in scan_wrapper_334445762078310996_315/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_325 scan_wrapper_334445762078310996_325/clk_in scan_wrapper_334445762078310996_326/clk_in
+ scan_wrapper_334445762078310996_325/data_in scan_wrapper_334445762078310996_326/data_in
+ scan_wrapper_334445762078310996_325/latch_enable_in scan_wrapper_334445762078310996_326/latch_enable_in
+ scan_wrapper_334445762078310996_325/scan_select_in scan_wrapper_334445762078310996_326/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_336 scan_wrapper_334445762078310996_336/clk_in scan_wrapper_334445762078310996_337/clk_in
+ scan_wrapper_334445762078310996_336/data_in scan_wrapper_334445762078310996_337/data_in
+ scan_wrapper_334445762078310996_336/latch_enable_in scan_wrapper_334445762078310996_337/latch_enable_in
+ scan_wrapper_334445762078310996_336/scan_select_in scan_wrapper_334445762078310996_337/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_347 scan_wrapper_334445762078310996_347/clk_in scan_wrapper_334445762078310996_348/clk_in
+ scan_wrapper_334445762078310996_347/data_in scan_wrapper_334445762078310996_348/data_in
+ scan_wrapper_334445762078310996_347/latch_enable_in scan_wrapper_334445762078310996_348/latch_enable_in
+ scan_wrapper_334445762078310996_347/scan_select_in scan_wrapper_334445762078310996_348/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_358 scan_wrapper_334445762078310996_358/clk_in scan_wrapper_334445762078310996_359/clk_in
+ scan_wrapper_334445762078310996_358/data_in scan_wrapper_334445762078310996_359/data_in
+ scan_wrapper_334445762078310996_358/latch_enable_in scan_wrapper_334445762078310996_359/latch_enable_in
+ scan_wrapper_334445762078310996_358/scan_select_in scan_wrapper_334445762078310996_359/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_369 scan_wrapper_334445762078310996_369/clk_in scan_wrapper_334445762078310996_370/clk_in
+ scan_wrapper_334445762078310996_369/data_in scan_wrapper_334445762078310996_370/data_in
+ scan_wrapper_334445762078310996_369/latch_enable_in scan_wrapper_334445762078310996_370/latch_enable_in
+ scan_wrapper_334445762078310996_369/scan_select_in scan_wrapper_334445762078310996_370/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_100 scan_wrapper_334445762078310996_99/clk_out scan_wrapper_334445762078310996_101/clk_in
+ scan_wrapper_334445762078310996_99/data_out scan_wrapper_334445762078310996_101/data_in
+ scan_wrapper_334445762078310996_99/latch_enable_out scan_wrapper_334445762078310996_101/latch_enable_in
+ scan_wrapper_334445762078310996_99/scan_select_out scan_wrapper_334445762078310996_101/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_111 scan_wrapper_334445762078310996_111/clk_in scan_wrapper_334445762078310996_112/clk_in
+ scan_wrapper_334445762078310996_111/data_in scan_wrapper_334445762078310996_112/data_in
+ scan_wrapper_334445762078310996_111/latch_enable_in scan_wrapper_334445762078310996_112/latch_enable_in
+ scan_wrapper_334445762078310996_111/scan_select_in scan_wrapper_334445762078310996_112/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_122 scan_wrapper_334445762078310996_122/clk_in scan_wrapper_334445762078310996_123/clk_in
+ scan_wrapper_334445762078310996_122/data_in scan_wrapper_334445762078310996_123/data_in
+ scan_wrapper_334445762078310996_122/latch_enable_in scan_wrapper_334445762078310996_123/latch_enable_in
+ scan_wrapper_334445762078310996_122/scan_select_in scan_wrapper_334445762078310996_123/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_133 scan_wrapper_334445762078310996_133/clk_in scan_wrapper_334445762078310996_134/clk_in
+ scan_wrapper_334445762078310996_133/data_in scan_wrapper_334445762078310996_134/data_in
+ scan_wrapper_334445762078310996_133/latch_enable_in scan_wrapper_334445762078310996_134/latch_enable_in
+ scan_wrapper_334445762078310996_133/scan_select_in scan_wrapper_334445762078310996_134/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_144 scan_wrapper_334445762078310996_144/clk_in scan_wrapper_334445762078310996_145/clk_in
+ scan_wrapper_334445762078310996_144/data_in scan_wrapper_334445762078310996_145/data_in
+ scan_wrapper_334445762078310996_144/latch_enable_in scan_wrapper_334445762078310996_145/latch_enable_in
+ scan_wrapper_334445762078310996_144/scan_select_in scan_wrapper_334445762078310996_145/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_155 scan_wrapper_334445762078310996_155/clk_in scan_wrapper_334445762078310996_156/clk_in
+ scan_wrapper_334445762078310996_155/data_in scan_wrapper_334445762078310996_156/data_in
+ scan_wrapper_334445762078310996_155/latch_enable_in scan_wrapper_334445762078310996_156/latch_enable_in
+ scan_wrapper_334445762078310996_155/scan_select_in scan_wrapper_334445762078310996_156/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_166 scan_wrapper_334445762078310996_166/clk_in scan_wrapper_334445762078310996_167/clk_in
+ scan_wrapper_334445762078310996_166/data_in scan_wrapper_334445762078310996_167/data_in
+ scan_wrapper_334445762078310996_166/latch_enable_in scan_wrapper_334445762078310996_167/latch_enable_in
+ scan_wrapper_334445762078310996_166/scan_select_in scan_wrapper_334445762078310996_167/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_177 scan_wrapper_334445762078310996_177/clk_in scan_wrapper_334445762078310996_178/clk_in
+ scan_wrapper_334445762078310996_177/data_in scan_wrapper_334445762078310996_178/data_in
+ scan_wrapper_334445762078310996_177/latch_enable_in scan_wrapper_334445762078310996_178/latch_enable_in
+ scan_wrapper_334445762078310996_177/scan_select_in scan_wrapper_334445762078310996_178/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_188 scan_wrapper_334445762078310996_188/clk_in scan_wrapper_334445762078310996_189/clk_in
+ scan_wrapper_334445762078310996_188/data_in scan_wrapper_334445762078310996_189/data_in
+ scan_wrapper_334445762078310996_188/latch_enable_in scan_wrapper_334445762078310996_189/latch_enable_in
+ scan_wrapper_334445762078310996_188/scan_select_in scan_wrapper_334445762078310996_189/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_199 scan_wrapper_334445762078310996_199/clk_in scan_wrapper_334445762078310996_200/clk_in
+ scan_wrapper_334445762078310996_199/data_in scan_wrapper_334445762078310996_200/data_in
+ scan_wrapper_334445762078310996_199/latch_enable_in scan_wrapper_334445762078310996_200/latch_enable_in
+ scan_wrapper_334445762078310996_199/scan_select_in scan_wrapper_334445762078310996_200/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_84 scan_wrapper_334445762078310996_84/clk_in scan_wrapper_334445762078310996_85/clk_in
+ scan_wrapper_334445762078310996_84/data_in scan_wrapper_334445762078310996_85/data_in
+ scan_wrapper_334445762078310996_84/latch_enable_in scan_wrapper_334445762078310996_85/latch_enable_in
+ scan_wrapper_334445762078310996_84/scan_select_in scan_wrapper_334445762078310996_85/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_73 scan_wrapper_334445762078310996_73/clk_in scan_wrapper_334445762078310996_74/clk_in
+ scan_wrapper_334445762078310996_73/data_in scan_wrapper_334445762078310996_74/data_in
+ scan_wrapper_334445762078310996_73/latch_enable_in scan_wrapper_334445762078310996_74/latch_enable_in
+ scan_wrapper_334445762078310996_73/scan_select_in scan_wrapper_334445762078310996_74/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_62 scan_wrapper_334445762078310996_62/clk_in scan_wrapper_334445762078310996_63/clk_in
+ scan_wrapper_334445762078310996_62/data_in scan_wrapper_334445762078310996_63/data_in
+ scan_wrapper_334445762078310996_62/latch_enable_in scan_wrapper_334445762078310996_63/latch_enable_in
+ scan_wrapper_334445762078310996_62/scan_select_in scan_wrapper_334445762078310996_63/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_51 scan_wrapper_334445762078310996_51/clk_in scan_wrapper_334445762078310996_52/clk_in
+ scan_wrapper_334445762078310996_51/data_in scan_wrapper_334445762078310996_52/data_in
+ scan_wrapper_334445762078310996_51/latch_enable_in scan_wrapper_334445762078310996_52/latch_enable_in
+ scan_wrapper_334445762078310996_51/scan_select_in scan_wrapper_334445762078310996_52/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_40 scan_wrapper_334445762078310996_40/clk_in scan_wrapper_334445762078310996_41/clk_in
+ scan_wrapper_334445762078310996_40/data_in scan_wrapper_334445762078310996_41/data_in
+ scan_wrapper_334445762078310996_40/latch_enable_in scan_wrapper_334445762078310996_41/latch_enable_in
+ scan_wrapper_334445762078310996_40/scan_select_in scan_wrapper_334445762078310996_41/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_95 scan_wrapper_334445762078310996_95/clk_in scan_wrapper_334445762078310996_96/clk_in
+ scan_wrapper_334445762078310996_95/data_in scan_wrapper_334445762078310996_96/data_in
+ scan_wrapper_334445762078310996_95/latch_enable_in scan_wrapper_334445762078310996_96/latch_enable_in
+ scan_wrapper_334445762078310996_95/scan_select_in scan_wrapper_334445762078310996_96/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_304 scan_wrapper_334445762078310996_304/clk_in scan_wrapper_334445762078310996_305/clk_in
+ scan_wrapper_334445762078310996_304/data_in scan_wrapper_334445762078310996_305/data_in
+ scan_wrapper_334445762078310996_304/latch_enable_in scan_wrapper_334445762078310996_305/latch_enable_in
+ scan_wrapper_334445762078310996_304/scan_select_in scan_wrapper_334445762078310996_305/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_315 scan_wrapper_334445762078310996_315/clk_in scan_wrapper_334445762078310996_316/clk_in
+ scan_wrapper_334445762078310996_315/data_in scan_wrapper_334445762078310996_316/data_in
+ scan_wrapper_334445762078310996_315/latch_enable_in scan_wrapper_334445762078310996_316/latch_enable_in
+ scan_wrapper_334445762078310996_315/scan_select_in scan_wrapper_334445762078310996_316/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_326 scan_wrapper_334445762078310996_326/clk_in scan_wrapper_334445762078310996_327/clk_in
+ scan_wrapper_334445762078310996_326/data_in scan_wrapper_334445762078310996_327/data_in
+ scan_wrapper_334445762078310996_326/latch_enable_in scan_wrapper_334445762078310996_327/latch_enable_in
+ scan_wrapper_334445762078310996_326/scan_select_in scan_wrapper_334445762078310996_327/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_337 scan_wrapper_334445762078310996_337/clk_in scan_wrapper_334445762078310996_338/clk_in
+ scan_wrapper_334445762078310996_337/data_in scan_wrapper_334445762078310996_338/data_in
+ scan_wrapper_334445762078310996_337/latch_enable_in scan_wrapper_334445762078310996_338/latch_enable_in
+ scan_wrapper_334445762078310996_337/scan_select_in scan_wrapper_334445762078310996_338/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_348 scan_wrapper_334445762078310996_348/clk_in scan_wrapper_334445762078310996_349/clk_in
+ scan_wrapper_334445762078310996_348/data_in scan_wrapper_334445762078310996_349/data_in
+ scan_wrapper_334445762078310996_348/latch_enable_in scan_wrapper_334445762078310996_349/latch_enable_in
+ scan_wrapper_334445762078310996_348/scan_select_in scan_wrapper_334445762078310996_349/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_359 scan_wrapper_334445762078310996_359/clk_in scan_wrapper_334445762078310996_360/clk_in
+ scan_wrapper_334445762078310996_359/data_in scan_wrapper_334445762078310996_360/data_in
+ scan_wrapper_334445762078310996_359/latch_enable_in scan_wrapper_334445762078310996_360/latch_enable_in
+ scan_wrapper_334445762078310996_359/scan_select_in scan_wrapper_334445762078310996_360/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_101 scan_wrapper_334445762078310996_101/clk_in scan_wrapper_334445762078310996_102/clk_in
+ scan_wrapper_334445762078310996_101/data_in scan_wrapper_334445762078310996_102/data_in
+ scan_wrapper_334445762078310996_101/latch_enable_in scan_wrapper_334445762078310996_102/latch_enable_in
+ scan_wrapper_334445762078310996_101/scan_select_in scan_wrapper_334445762078310996_102/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_112 scan_wrapper_334445762078310996_112/clk_in scan_wrapper_334445762078310996_113/clk_in
+ scan_wrapper_334445762078310996_112/data_in scan_wrapper_334445762078310996_113/data_in
+ scan_wrapper_334445762078310996_112/latch_enable_in scan_wrapper_334445762078310996_113/latch_enable_in
+ scan_wrapper_334445762078310996_112/scan_select_in scan_wrapper_334445762078310996_113/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_123 scan_wrapper_334445762078310996_123/clk_in scan_wrapper_334445762078310996_124/clk_in
+ scan_wrapper_334445762078310996_123/data_in scan_wrapper_334445762078310996_124/data_in
+ scan_wrapper_334445762078310996_123/latch_enable_in scan_wrapper_334445762078310996_124/latch_enable_in
+ scan_wrapper_334445762078310996_123/scan_select_in scan_wrapper_334445762078310996_124/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_134 scan_wrapper_334445762078310996_134/clk_in scan_wrapper_334445762078310996_135/clk_in
+ scan_wrapper_334445762078310996_134/data_in scan_wrapper_334445762078310996_135/data_in
+ scan_wrapper_334445762078310996_134/latch_enable_in scan_wrapper_334445762078310996_135/latch_enable_in
+ scan_wrapper_334445762078310996_134/scan_select_in scan_wrapper_334445762078310996_135/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_145 scan_wrapper_334445762078310996_145/clk_in scan_wrapper_334445762078310996_146/clk_in
+ scan_wrapper_334445762078310996_145/data_in scan_wrapper_334445762078310996_146/data_in
+ scan_wrapper_334445762078310996_145/latch_enable_in scan_wrapper_334445762078310996_146/latch_enable_in
+ scan_wrapper_334445762078310996_145/scan_select_in scan_wrapper_334445762078310996_146/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_156 scan_wrapper_334445762078310996_156/clk_in scan_wrapper_334445762078310996_157/clk_in
+ scan_wrapper_334445762078310996_156/data_in scan_wrapper_334445762078310996_157/data_in
+ scan_wrapper_334445762078310996_156/latch_enable_in scan_wrapper_334445762078310996_157/latch_enable_in
+ scan_wrapper_334445762078310996_156/scan_select_in scan_wrapper_334445762078310996_157/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_167 scan_wrapper_334445762078310996_167/clk_in scan_wrapper_334445762078310996_168/clk_in
+ scan_wrapper_334445762078310996_167/data_in scan_wrapper_334445762078310996_168/data_in
+ scan_wrapper_334445762078310996_167/latch_enable_in scan_wrapper_334445762078310996_168/latch_enable_in
+ scan_wrapper_334445762078310996_167/scan_select_in scan_wrapper_334445762078310996_168/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_178 scan_wrapper_334445762078310996_178/clk_in scan_wrapper_334445762078310996_179/clk_in
+ scan_wrapper_334445762078310996_178/data_in scan_wrapper_334445762078310996_179/data_in
+ scan_wrapper_334445762078310996_178/latch_enable_in scan_wrapper_334445762078310996_179/latch_enable_in
+ scan_wrapper_334445762078310996_178/scan_select_in scan_wrapper_334445762078310996_179/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_189 scan_wrapper_334445762078310996_189/clk_in scan_wrapper_334445762078310996_190/clk_in
+ scan_wrapper_334445762078310996_189/data_in scan_wrapper_334445762078310996_190/data_in
+ scan_wrapper_334445762078310996_189/latch_enable_in scan_wrapper_334445762078310996_190/latch_enable_in
+ scan_wrapper_334445762078310996_189/scan_select_in scan_wrapper_334445762078310996_190/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_85 scan_wrapper_334445762078310996_85/clk_in scan_wrapper_334445762078310996_86/clk_in
+ scan_wrapper_334445762078310996_85/data_in scan_wrapper_334445762078310996_86/data_in
+ scan_wrapper_334445762078310996_85/latch_enable_in scan_wrapper_334445762078310996_86/latch_enable_in
+ scan_wrapper_334445762078310996_85/scan_select_in scan_wrapper_334445762078310996_86/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_74 scan_wrapper_334445762078310996_74/clk_in scan_wrapper_334445762078310996_75/clk_in
+ scan_wrapper_334445762078310996_74/data_in scan_wrapper_334445762078310996_75/data_in
+ scan_wrapper_334445762078310996_74/latch_enable_in scan_wrapper_334445762078310996_75/latch_enable_in
+ scan_wrapper_334445762078310996_74/scan_select_in scan_wrapper_334445762078310996_75/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_63 scan_wrapper_334445762078310996_63/clk_in scan_wrapper_334445762078310996_64/clk_in
+ scan_wrapper_334445762078310996_63/data_in scan_wrapper_334445762078310996_64/data_in
+ scan_wrapper_334445762078310996_63/latch_enable_in scan_wrapper_334445762078310996_64/latch_enable_in
+ scan_wrapper_334445762078310996_63/scan_select_in scan_wrapper_334445762078310996_64/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_52 scan_wrapper_334445762078310996_52/clk_in scan_wrapper_334445762078310996_53/clk_in
+ scan_wrapper_334445762078310996_52/data_in scan_wrapper_334445762078310996_53/data_in
+ scan_wrapper_334445762078310996_52/latch_enable_in scan_wrapper_334445762078310996_53/latch_enable_in
+ scan_wrapper_334445762078310996_52/scan_select_in scan_wrapper_334445762078310996_53/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_41 scan_wrapper_334445762078310996_41/clk_in scan_wrapper_334445762078310996_42/clk_in
+ scan_wrapper_334445762078310996_41/data_in scan_wrapper_334445762078310996_42/data_in
+ scan_wrapper_334445762078310996_41/latch_enable_in scan_wrapper_334445762078310996_42/latch_enable_in
+ scan_wrapper_334445762078310996_41/scan_select_in scan_wrapper_334445762078310996_42/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_30 scan_wrapper_334445762078310996_30/clk_in scan_wrapper_334445762078310996_31/clk_in
+ scan_wrapper_334445762078310996_30/data_in scan_wrapper_334445762078310996_31/data_in
+ scan_wrapper_334445762078310996_30/latch_enable_in scan_wrapper_334445762078310996_31/latch_enable_in
+ scan_wrapper_334445762078310996_30/scan_select_in scan_wrapper_334445762078310996_31/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_96 scan_wrapper_334445762078310996_96/clk_in scan_wrapper_334445762078310996_97/clk_in
+ scan_wrapper_334445762078310996_96/data_in scan_wrapper_334445762078310996_97/data_in
+ scan_wrapper_334445762078310996_96/latch_enable_in scan_wrapper_334445762078310996_97/latch_enable_in
+ scan_wrapper_334445762078310996_96/scan_select_in scan_wrapper_334445762078310996_97/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_305 scan_wrapper_334445762078310996_305/clk_in scan_wrapper_334445762078310996_306/clk_in
+ scan_wrapper_334445762078310996_305/data_in scan_wrapper_334445762078310996_306/data_in
+ scan_wrapper_334445762078310996_305/latch_enable_in scan_wrapper_334445762078310996_306/latch_enable_in
+ scan_wrapper_334445762078310996_305/scan_select_in scan_wrapper_334445762078310996_306/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_316 scan_wrapper_334445762078310996_316/clk_in scan_wrapper_334445762078310996_317/clk_in
+ scan_wrapper_334445762078310996_316/data_in scan_wrapper_334445762078310996_317/data_in
+ scan_wrapper_334445762078310996_316/latch_enable_in scan_wrapper_334445762078310996_317/latch_enable_in
+ scan_wrapper_334445762078310996_316/scan_select_in scan_wrapper_334445762078310996_317/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_327 scan_wrapper_334445762078310996_327/clk_in scan_wrapper_334445762078310996_328/clk_in
+ scan_wrapper_334445762078310996_327/data_in scan_wrapper_334445762078310996_328/data_in
+ scan_wrapper_334445762078310996_327/latch_enable_in scan_wrapper_334445762078310996_328/latch_enable_in
+ scan_wrapper_334445762078310996_327/scan_select_in scan_wrapper_334445762078310996_328/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_338 scan_wrapper_334445762078310996_338/clk_in scan_wrapper_334445762078310996_339/clk_in
+ scan_wrapper_334445762078310996_338/data_in scan_wrapper_334445762078310996_339/data_in
+ scan_wrapper_334445762078310996_338/latch_enable_in scan_wrapper_334445762078310996_339/latch_enable_in
+ scan_wrapper_334445762078310996_338/scan_select_in scan_wrapper_334445762078310996_339/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_349 scan_wrapper_334445762078310996_349/clk_in scan_wrapper_334445762078310996_350/clk_in
+ scan_wrapper_334445762078310996_349/data_in scan_wrapper_334445762078310996_350/data_in
+ scan_wrapper_334445762078310996_349/latch_enable_in scan_wrapper_334445762078310996_350/latch_enable_in
+ scan_wrapper_334445762078310996_349/scan_select_in scan_wrapper_334445762078310996_350/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_102 scan_wrapper_334445762078310996_102/clk_in scan_wrapper_334445762078310996_103/clk_in
+ scan_wrapper_334445762078310996_102/data_in scan_wrapper_334445762078310996_103/data_in
+ scan_wrapper_334445762078310996_102/latch_enable_in scan_wrapper_334445762078310996_103/latch_enable_in
+ scan_wrapper_334445762078310996_102/scan_select_in scan_wrapper_334445762078310996_103/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_113 scan_wrapper_334445762078310996_113/clk_in scan_wrapper_334445762078310996_114/clk_in
+ scan_wrapper_334445762078310996_113/data_in scan_wrapper_334445762078310996_114/data_in
+ scan_wrapper_334445762078310996_113/latch_enable_in scan_wrapper_334445762078310996_114/latch_enable_in
+ scan_wrapper_334445762078310996_113/scan_select_in scan_wrapper_334445762078310996_114/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_124 scan_wrapper_334445762078310996_124/clk_in scan_wrapper_334445762078310996_125/clk_in
+ scan_wrapper_334445762078310996_124/data_in scan_wrapper_334445762078310996_125/data_in
+ scan_wrapper_334445762078310996_124/latch_enable_in scan_wrapper_334445762078310996_125/latch_enable_in
+ scan_wrapper_334445762078310996_124/scan_select_in scan_wrapper_334445762078310996_125/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_135 scan_wrapper_334445762078310996_135/clk_in scan_wrapper_334445762078310996_136/clk_in
+ scan_wrapper_334445762078310996_135/data_in scan_wrapper_334445762078310996_136/data_in
+ scan_wrapper_334445762078310996_135/latch_enable_in scan_wrapper_334445762078310996_136/latch_enable_in
+ scan_wrapper_334445762078310996_135/scan_select_in scan_wrapper_334445762078310996_136/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_146 scan_wrapper_334445762078310996_146/clk_in scan_wrapper_334445762078310996_147/clk_in
+ scan_wrapper_334445762078310996_146/data_in scan_wrapper_334445762078310996_147/data_in
+ scan_wrapper_334445762078310996_146/latch_enable_in scan_wrapper_334445762078310996_147/latch_enable_in
+ scan_wrapper_334445762078310996_146/scan_select_in scan_wrapper_334445762078310996_147/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_157 scan_wrapper_334445762078310996_157/clk_in scan_wrapper_334445762078310996_158/clk_in
+ scan_wrapper_334445762078310996_157/data_in scan_wrapper_334445762078310996_158/data_in
+ scan_wrapper_334445762078310996_157/latch_enable_in scan_wrapper_334445762078310996_158/latch_enable_in
+ scan_wrapper_334445762078310996_157/scan_select_in scan_wrapper_334445762078310996_158/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_168 scan_wrapper_334445762078310996_168/clk_in scan_wrapper_334445762078310996_169/clk_in
+ scan_wrapper_334445762078310996_168/data_in scan_wrapper_334445762078310996_169/data_in
+ scan_wrapper_334445762078310996_168/latch_enable_in scan_wrapper_334445762078310996_169/latch_enable_in
+ scan_wrapper_334445762078310996_168/scan_select_in scan_wrapper_334445762078310996_169/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_179 scan_wrapper_334445762078310996_179/clk_in scan_wrapper_334445762078310996_180/clk_in
+ scan_wrapper_334445762078310996_179/data_in scan_wrapper_334445762078310996_180/data_in
+ scan_wrapper_334445762078310996_179/latch_enable_in scan_wrapper_334445762078310996_180/latch_enable_in
+ scan_wrapper_334445762078310996_179/scan_select_in scan_wrapper_334445762078310996_180/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_86 scan_wrapper_334445762078310996_86/clk_in scan_wrapper_334445762078310996_87/clk_in
+ scan_wrapper_334445762078310996_86/data_in scan_wrapper_334445762078310996_87/data_in
+ scan_wrapper_334445762078310996_86/latch_enable_in scan_wrapper_334445762078310996_87/latch_enable_in
+ scan_wrapper_334445762078310996_86/scan_select_in scan_wrapper_334445762078310996_87/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_75 scan_wrapper_334445762078310996_75/clk_in scan_wrapper_334445762078310996_76/clk_in
+ scan_wrapper_334445762078310996_75/data_in scan_wrapper_334445762078310996_76/data_in
+ scan_wrapper_334445762078310996_75/latch_enable_in scan_wrapper_334445762078310996_76/latch_enable_in
+ scan_wrapper_334445762078310996_75/scan_select_in scan_wrapper_334445762078310996_76/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_64 scan_wrapper_334445762078310996_64/clk_in scan_wrapper_334445762078310996_65/clk_in
+ scan_wrapper_334445762078310996_64/data_in scan_wrapper_334445762078310996_65/data_in
+ scan_wrapper_334445762078310996_64/latch_enable_in scan_wrapper_334445762078310996_65/latch_enable_in
+ scan_wrapper_334445762078310996_64/scan_select_in scan_wrapper_334445762078310996_65/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_53 scan_wrapper_334445762078310996_53/clk_in scan_wrapper_334445762078310996_54/clk_in
+ scan_wrapper_334445762078310996_53/data_in scan_wrapper_334445762078310996_54/data_in
+ scan_wrapper_334445762078310996_53/latch_enable_in scan_wrapper_334445762078310996_54/latch_enable_in
+ scan_wrapper_334445762078310996_53/scan_select_in scan_wrapper_334445762078310996_54/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_42 scan_wrapper_334445762078310996_42/clk_in scan_wrapper_334445762078310996_43/clk_in
+ scan_wrapper_334445762078310996_42/data_in scan_wrapper_334445762078310996_43/data_in
+ scan_wrapper_334445762078310996_42/latch_enable_in scan_wrapper_334445762078310996_43/latch_enable_in
+ scan_wrapper_334445762078310996_42/scan_select_in scan_wrapper_334445762078310996_43/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_31 scan_wrapper_334445762078310996_31/clk_in scan_wrapper_334445762078310996_32/clk_in
+ scan_wrapper_334445762078310996_31/data_in scan_wrapper_334445762078310996_32/data_in
+ scan_wrapper_334445762078310996_31/latch_enable_in scan_wrapper_334445762078310996_32/latch_enable_in
+ scan_wrapper_334445762078310996_31/scan_select_in scan_wrapper_334445762078310996_32/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_20 scan_wrapper_334445762078310996_20/clk_in scan_wrapper_334445762078310996_21/clk_in
+ scan_wrapper_334445762078310996_20/data_in scan_wrapper_334445762078310996_21/data_in
+ scan_wrapper_334445762078310996_20/latch_enable_in scan_wrapper_334445762078310996_21/latch_enable_in
+ scan_wrapper_334445762078310996_20/scan_select_in scan_wrapper_334445762078310996_21/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_97 scan_wrapper_334445762078310996_97/clk_in scan_wrapper_334445762078310996_98/clk_in
+ scan_wrapper_334445762078310996_97/data_in scan_wrapper_334445762078310996_98/data_in
+ scan_wrapper_334445762078310996_97/latch_enable_in scan_wrapper_334445762078310996_98/latch_enable_in
+ scan_wrapper_334445762078310996_97/scan_select_in scan_wrapper_334445762078310996_98/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_306 scan_wrapper_334445762078310996_306/clk_in scan_wrapper_334445762078310996_307/clk_in
+ scan_wrapper_334445762078310996_306/data_in scan_wrapper_334445762078310996_307/data_in
+ scan_wrapper_334445762078310996_306/latch_enable_in scan_wrapper_334445762078310996_307/latch_enable_in
+ scan_wrapper_334445762078310996_306/scan_select_in scan_wrapper_334445762078310996_307/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_317 scan_wrapper_334445762078310996_317/clk_in scan_wrapper_334445762078310996_318/clk_in
+ scan_wrapper_334445762078310996_317/data_in scan_wrapper_334445762078310996_318/data_in
+ scan_wrapper_334445762078310996_317/latch_enable_in scan_wrapper_334445762078310996_318/latch_enable_in
+ scan_wrapper_334445762078310996_317/scan_select_in scan_wrapper_334445762078310996_318/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_328 scan_wrapper_334445762078310996_328/clk_in scan_wrapper_334445762078310996_329/clk_in
+ scan_wrapper_334445762078310996_328/data_in scan_wrapper_334445762078310996_329/data_in
+ scan_wrapper_334445762078310996_328/latch_enable_in scan_wrapper_334445762078310996_329/latch_enable_in
+ scan_wrapper_334445762078310996_328/scan_select_in scan_wrapper_334445762078310996_329/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_339 scan_wrapper_334445762078310996_339/clk_in scan_wrapper_334445762078310996_340/clk_in
+ scan_wrapper_334445762078310996_339/data_in scan_wrapper_334445762078310996_340/data_in
+ scan_wrapper_334445762078310996_339/latch_enable_in scan_wrapper_334445762078310996_340/latch_enable_in
+ scan_wrapper_334445762078310996_339/scan_select_in scan_wrapper_334445762078310996_340/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_103 scan_wrapper_334445762078310996_103/clk_in scan_wrapper_334445762078310996_104/clk_in
+ scan_wrapper_334445762078310996_103/data_in scan_wrapper_334445762078310996_104/data_in
+ scan_wrapper_334445762078310996_103/latch_enable_in scan_wrapper_334445762078310996_104/latch_enable_in
+ scan_wrapper_334445762078310996_103/scan_select_in scan_wrapper_334445762078310996_104/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_114 scan_wrapper_334445762078310996_114/clk_in scan_wrapper_334445762078310996_115/clk_in
+ scan_wrapper_334445762078310996_114/data_in scan_wrapper_334445762078310996_115/data_in
+ scan_wrapper_334445762078310996_114/latch_enable_in scan_wrapper_334445762078310996_115/latch_enable_in
+ scan_wrapper_334445762078310996_114/scan_select_in scan_wrapper_334445762078310996_115/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_125 scan_wrapper_334445762078310996_125/clk_in scan_wrapper_334445762078310996_126/clk_in
+ scan_wrapper_334445762078310996_125/data_in scan_wrapper_334445762078310996_126/data_in
+ scan_wrapper_334445762078310996_125/latch_enable_in scan_wrapper_334445762078310996_126/latch_enable_in
+ scan_wrapper_334445762078310996_125/scan_select_in scan_wrapper_334445762078310996_126/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_136 scan_wrapper_334445762078310996_136/clk_in scan_wrapper_334445762078310996_137/clk_in
+ scan_wrapper_334445762078310996_136/data_in scan_wrapper_334445762078310996_137/data_in
+ scan_wrapper_334445762078310996_136/latch_enable_in scan_wrapper_334445762078310996_137/latch_enable_in
+ scan_wrapper_334445762078310996_136/scan_select_in scan_wrapper_334445762078310996_137/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_147 scan_wrapper_334445762078310996_147/clk_in scan_wrapper_334445762078310996_148/clk_in
+ scan_wrapper_334445762078310996_147/data_in scan_wrapper_334445762078310996_148/data_in
+ scan_wrapper_334445762078310996_147/latch_enable_in scan_wrapper_334445762078310996_148/latch_enable_in
+ scan_wrapper_334445762078310996_147/scan_select_in scan_wrapper_334445762078310996_148/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_158 scan_wrapper_334445762078310996_158/clk_in scan_wrapper_334445762078310996_159/clk_in
+ scan_wrapper_334445762078310996_158/data_in scan_wrapper_334445762078310996_159/data_in
+ scan_wrapper_334445762078310996_158/latch_enable_in scan_wrapper_334445762078310996_159/latch_enable_in
+ scan_wrapper_334445762078310996_158/scan_select_in scan_wrapper_334445762078310996_159/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_169 scan_wrapper_334445762078310996_169/clk_in scan_wrapper_334445762078310996_170/clk_in
+ scan_wrapper_334445762078310996_169/data_in scan_wrapper_334445762078310996_170/data_in
+ scan_wrapper_334445762078310996_169/latch_enable_in scan_wrapper_334445762078310996_170/latch_enable_in
+ scan_wrapper_334445762078310996_169/scan_select_in scan_wrapper_334445762078310996_170/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_87 scan_wrapper_334445762078310996_87/clk_in scan_wrapper_334445762078310996_88/clk_in
+ scan_wrapper_334445762078310996_87/data_in scan_wrapper_334445762078310996_88/data_in
+ scan_wrapper_334445762078310996_87/latch_enable_in scan_wrapper_334445762078310996_88/latch_enable_in
+ scan_wrapper_334445762078310996_87/scan_select_in scan_wrapper_334445762078310996_88/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_76 scan_wrapper_334445762078310996_76/clk_in scan_wrapper_334445762078310996_77/clk_in
+ scan_wrapper_334445762078310996_76/data_in scan_wrapper_334445762078310996_77/data_in
+ scan_wrapper_334445762078310996_76/latch_enable_in scan_wrapper_334445762078310996_77/latch_enable_in
+ scan_wrapper_334445762078310996_76/scan_select_in scan_wrapper_334445762078310996_77/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_65 scan_wrapper_334445762078310996_65/clk_in scan_wrapper_334445762078310996_66/clk_in
+ scan_wrapper_334445762078310996_65/data_in scan_wrapper_334445762078310996_66/data_in
+ scan_wrapper_334445762078310996_65/latch_enable_in scan_wrapper_334445762078310996_66/latch_enable_in
+ scan_wrapper_334445762078310996_65/scan_select_in scan_wrapper_334445762078310996_66/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_54 scan_wrapper_334445762078310996_54/clk_in scan_wrapper_334445762078310996_55/clk_in
+ scan_wrapper_334445762078310996_54/data_in scan_wrapper_334445762078310996_55/data_in
+ scan_wrapper_334445762078310996_54/latch_enable_in scan_wrapper_334445762078310996_55/latch_enable_in
+ scan_wrapper_334445762078310996_54/scan_select_in scan_wrapper_334445762078310996_55/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_43 scan_wrapper_334445762078310996_43/clk_in scan_wrapper_334445762078310996_44/clk_in
+ scan_wrapper_334445762078310996_43/data_in scan_wrapper_334445762078310996_44/data_in
+ scan_wrapper_334445762078310996_43/latch_enable_in scan_wrapper_334445762078310996_44/latch_enable_in
+ scan_wrapper_334445762078310996_43/scan_select_in scan_wrapper_334445762078310996_44/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_32 scan_wrapper_334445762078310996_32/clk_in scan_wrapper_334445762078310996_33/clk_in
+ scan_wrapper_334445762078310996_32/data_in scan_wrapper_334445762078310996_33/data_in
+ scan_wrapper_334445762078310996_32/latch_enable_in scan_wrapper_334445762078310996_33/latch_enable_in
+ scan_wrapper_334445762078310996_32/scan_select_in scan_wrapper_334445762078310996_33/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_21 scan_wrapper_334445762078310996_21/clk_in scan_wrapper_334445762078310996_22/clk_in
+ scan_wrapper_334445762078310996_21/data_in scan_wrapper_334445762078310996_22/data_in
+ scan_wrapper_334445762078310996_21/latch_enable_in scan_wrapper_334445762078310996_22/latch_enable_in
+ scan_wrapper_334445762078310996_21/scan_select_in scan_wrapper_334445762078310996_22/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_10 scan_wrapper_334445762078310996_9/clk_out scan_wrapper_334445762078310996_11/clk_in
+ scan_wrapper_334445762078310996_9/data_out scan_wrapper_334445762078310996_11/data_in
+ scan_wrapper_334445762078310996_9/latch_enable_out scan_wrapper_334445762078310996_11/latch_enable_in
+ scan_wrapper_334445762078310996_9/scan_select_out scan_wrapper_334445762078310996_11/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_98 scan_wrapper_334445762078310996_98/clk_in scan_wrapper_334445762078310996_99/clk_in
+ scan_wrapper_334445762078310996_98/data_in scan_wrapper_334445762078310996_99/data_in
+ scan_wrapper_334445762078310996_98/latch_enable_in scan_wrapper_334445762078310996_99/latch_enable_in
+ scan_wrapper_334445762078310996_98/scan_select_in scan_wrapper_334445762078310996_99/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_307 scan_wrapper_334445762078310996_307/clk_in scan_wrapper_334445762078310996_308/clk_in
+ scan_wrapper_334445762078310996_307/data_in scan_wrapper_334445762078310996_308/data_in
+ scan_wrapper_334445762078310996_307/latch_enable_in scan_wrapper_334445762078310996_308/latch_enable_in
+ scan_wrapper_334445762078310996_307/scan_select_in scan_wrapper_334445762078310996_308/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_318 scan_wrapper_334445762078310996_318/clk_in scan_wrapper_334445762078310996_319/clk_in
+ scan_wrapper_334445762078310996_318/data_in scan_wrapper_334445762078310996_319/data_in
+ scan_wrapper_334445762078310996_318/latch_enable_in scan_wrapper_334445762078310996_319/latch_enable_in
+ scan_wrapper_334445762078310996_318/scan_select_in scan_wrapper_334445762078310996_319/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_329 scan_wrapper_334445762078310996_329/clk_in scan_wrapper_334445762078310996_330/clk_in
+ scan_wrapper_334445762078310996_329/data_in scan_wrapper_334445762078310996_330/data_in
+ scan_wrapper_334445762078310996_329/latch_enable_in scan_wrapper_334445762078310996_330/latch_enable_in
+ scan_wrapper_334445762078310996_329/scan_select_in scan_wrapper_334445762078310996_330/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_104 scan_wrapper_334445762078310996_104/clk_in scan_wrapper_334445762078310996_105/clk_in
+ scan_wrapper_334445762078310996_104/data_in scan_wrapper_334445762078310996_105/data_in
+ scan_wrapper_334445762078310996_104/latch_enable_in scan_wrapper_334445762078310996_105/latch_enable_in
+ scan_wrapper_334445762078310996_104/scan_select_in scan_wrapper_334445762078310996_105/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_115 scan_wrapper_334445762078310996_115/clk_in scan_wrapper_334445762078310996_116/clk_in
+ scan_wrapper_334445762078310996_115/data_in scan_wrapper_334445762078310996_116/data_in
+ scan_wrapper_334445762078310996_115/latch_enable_in scan_wrapper_334445762078310996_116/latch_enable_in
+ scan_wrapper_334445762078310996_115/scan_select_in scan_wrapper_334445762078310996_116/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_126 scan_wrapper_334445762078310996_126/clk_in scan_wrapper_334445762078310996_127/clk_in
+ scan_wrapper_334445762078310996_126/data_in scan_wrapper_334445762078310996_127/data_in
+ scan_wrapper_334445762078310996_126/latch_enable_in scan_wrapper_334445762078310996_127/latch_enable_in
+ scan_wrapper_334445762078310996_126/scan_select_in scan_wrapper_334445762078310996_127/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_137 scan_wrapper_334445762078310996_137/clk_in scan_wrapper_334445762078310996_138/clk_in
+ scan_wrapper_334445762078310996_137/data_in scan_wrapper_334445762078310996_138/data_in
+ scan_wrapper_334445762078310996_137/latch_enable_in scan_wrapper_334445762078310996_138/latch_enable_in
+ scan_wrapper_334445762078310996_137/scan_select_in scan_wrapper_334445762078310996_138/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_148 scan_wrapper_334445762078310996_148/clk_in scan_wrapper_334445762078310996_149/clk_in
+ scan_wrapper_334445762078310996_148/data_in scan_wrapper_334445762078310996_149/data_in
+ scan_wrapper_334445762078310996_148/latch_enable_in scan_wrapper_334445762078310996_149/latch_enable_in
+ scan_wrapper_334445762078310996_148/scan_select_in scan_wrapper_334445762078310996_149/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_159 scan_wrapper_334445762078310996_159/clk_in scan_wrapper_334445762078310996_160/clk_in
+ scan_wrapper_334445762078310996_159/data_in scan_wrapper_334445762078310996_160/data_in
+ scan_wrapper_334445762078310996_159/latch_enable_in scan_wrapper_334445762078310996_160/latch_enable_in
+ scan_wrapper_334445762078310996_159/scan_select_in scan_wrapper_334445762078310996_160/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_490 scan_wrapper_334445762078310996_490/clk_in scan_wrapper_334445762078310996_491/clk_in
+ scan_wrapper_334445762078310996_490/data_in scan_wrapper_334445762078310996_491/data_in
+ scan_wrapper_334445762078310996_490/latch_enable_in scan_wrapper_334445762078310996_491/latch_enable_in
+ scan_wrapper_334445762078310996_490/scan_select_in scan_wrapper_334445762078310996_491/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_88 scan_wrapper_334445762078310996_88/clk_in scan_wrapper_334445762078310996_89/clk_in
+ scan_wrapper_334445762078310996_88/data_in scan_wrapper_334445762078310996_89/data_in
+ scan_wrapper_334445762078310996_88/latch_enable_in scan_wrapper_334445762078310996_89/latch_enable_in
+ scan_wrapper_334445762078310996_88/scan_select_in scan_wrapper_334445762078310996_89/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_77 scan_wrapper_334445762078310996_77/clk_in scan_wrapper_334445762078310996_78/clk_in
+ scan_wrapper_334445762078310996_77/data_in scan_wrapper_334445762078310996_78/data_in
+ scan_wrapper_334445762078310996_77/latch_enable_in scan_wrapper_334445762078310996_78/latch_enable_in
+ scan_wrapper_334445762078310996_77/scan_select_in scan_wrapper_334445762078310996_78/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_66 scan_wrapper_334445762078310996_66/clk_in scan_wrapper_334445762078310996_67/clk_in
+ scan_wrapper_334445762078310996_66/data_in scan_wrapper_334445762078310996_67/data_in
+ scan_wrapper_334445762078310996_66/latch_enable_in scan_wrapper_334445762078310996_67/latch_enable_in
+ scan_wrapper_334445762078310996_66/scan_select_in scan_wrapper_334445762078310996_67/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_55 scan_wrapper_334445762078310996_55/clk_in scan_wrapper_334445762078310996_56/clk_in
+ scan_wrapper_334445762078310996_55/data_in scan_wrapper_334445762078310996_56/data_in
+ scan_wrapper_334445762078310996_55/latch_enable_in scan_wrapper_334445762078310996_56/latch_enable_in
+ scan_wrapper_334445762078310996_55/scan_select_in scan_wrapper_334445762078310996_56/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_44 scan_wrapper_334445762078310996_44/clk_in scan_wrapper_334445762078310996_45/clk_in
+ scan_wrapper_334445762078310996_44/data_in scan_wrapper_334445762078310996_45/data_in
+ scan_wrapper_334445762078310996_44/latch_enable_in scan_wrapper_334445762078310996_45/latch_enable_in
+ scan_wrapper_334445762078310996_44/scan_select_in scan_wrapper_334445762078310996_45/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_33 scan_wrapper_334445762078310996_33/clk_in scan_wrapper_334445762078310996_34/clk_in
+ scan_wrapper_334445762078310996_33/data_in scan_wrapper_334445762078310996_34/data_in
+ scan_wrapper_334445762078310996_33/latch_enable_in scan_wrapper_334445762078310996_34/latch_enable_in
+ scan_wrapper_334445762078310996_33/scan_select_in scan_wrapper_334445762078310996_34/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_22 scan_wrapper_334445762078310996_22/clk_in scan_wrapper_334445762078310996_23/clk_in
+ scan_wrapper_334445762078310996_22/data_in scan_wrapper_334445762078310996_23/data_in
+ scan_wrapper_334445762078310996_22/latch_enable_in scan_wrapper_334445762078310996_23/latch_enable_in
+ scan_wrapper_334445762078310996_22/scan_select_in scan_wrapper_334445762078310996_23/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_11 scan_wrapper_334445762078310996_11/clk_in scan_wrapper_334445762078310996_12/clk_in
+ scan_wrapper_334445762078310996_11/data_in scan_wrapper_334445762078310996_12/data_in
+ scan_wrapper_334445762078310996_11/latch_enable_in scan_wrapper_334445762078310996_12/latch_enable_in
+ scan_wrapper_334445762078310996_11/scan_select_in scan_wrapper_334445762078310996_12/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_99 scan_wrapper_334445762078310996_99/clk_in scan_wrapper_334445762078310996_99/clk_out
+ scan_wrapper_334445762078310996_99/data_in scan_wrapper_334445762078310996_99/data_out
+ scan_wrapper_334445762078310996_99/latch_enable_in scan_wrapper_334445762078310996_99/latch_enable_out
+ scan_wrapper_334445762078310996_99/scan_select_in scan_wrapper_334445762078310996_99/scan_select_out
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_308 scan_wrapper_334445762078310996_308/clk_in scan_wrapper_334445762078310996_309/clk_in
+ scan_wrapper_334445762078310996_308/data_in scan_wrapper_334445762078310996_309/data_in
+ scan_wrapper_334445762078310996_308/latch_enable_in scan_wrapper_334445762078310996_309/latch_enable_in
+ scan_wrapper_334445762078310996_308/scan_select_in scan_wrapper_334445762078310996_309/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_319 scan_wrapper_334445762078310996_319/clk_in scan_wrapper_334445762078310996_320/clk_in
+ scan_wrapper_334445762078310996_319/data_in scan_wrapper_334445762078310996_320/data_in
+ scan_wrapper_334445762078310996_319/latch_enable_in scan_wrapper_334445762078310996_320/latch_enable_in
+ scan_wrapper_334445762078310996_319/scan_select_in scan_wrapper_334445762078310996_320/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_105 scan_wrapper_334445762078310996_105/clk_in scan_wrapper_334445762078310996_106/clk_in
+ scan_wrapper_334445762078310996_105/data_in scan_wrapper_334445762078310996_106/data_in
+ scan_wrapper_334445762078310996_105/latch_enable_in scan_wrapper_334445762078310996_106/latch_enable_in
+ scan_wrapper_334445762078310996_105/scan_select_in scan_wrapper_334445762078310996_106/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_116 scan_wrapper_334445762078310996_116/clk_in scan_wrapper_334445762078310996_117/clk_in
+ scan_wrapper_334445762078310996_116/data_in scan_wrapper_334445762078310996_117/data_in
+ scan_wrapper_334445762078310996_116/latch_enable_in scan_wrapper_334445762078310996_117/latch_enable_in
+ scan_wrapper_334445762078310996_116/scan_select_in scan_wrapper_334445762078310996_117/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_127 scan_wrapper_334445762078310996_127/clk_in scan_wrapper_334445762078310996_128/clk_in
+ scan_wrapper_334445762078310996_127/data_in scan_wrapper_334445762078310996_128/data_in
+ scan_wrapper_334445762078310996_127/latch_enable_in scan_wrapper_334445762078310996_128/latch_enable_in
+ scan_wrapper_334445762078310996_127/scan_select_in scan_wrapper_334445762078310996_128/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_138 scan_wrapper_334445762078310996_138/clk_in scan_wrapper_334445762078310996_139/clk_in
+ scan_wrapper_334445762078310996_138/data_in scan_wrapper_334445762078310996_139/data_in
+ scan_wrapper_334445762078310996_138/latch_enable_in scan_wrapper_334445762078310996_139/latch_enable_in
+ scan_wrapper_334445762078310996_138/scan_select_in scan_wrapper_334445762078310996_139/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_149 scan_wrapper_334445762078310996_149/clk_in scan_wrapper_334445762078310996_150/clk_in
+ scan_wrapper_334445762078310996_149/data_in scan_wrapper_334445762078310996_150/data_in
+ scan_wrapper_334445762078310996_149/latch_enable_in scan_wrapper_334445762078310996_150/latch_enable_in
+ scan_wrapper_334445762078310996_149/scan_select_in scan_wrapper_334445762078310996_150/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_491 scan_wrapper_334445762078310996_491/clk_in scan_wrapper_334445762078310996_492/clk_in
+ scan_wrapper_334445762078310996_491/data_in scan_wrapper_334445762078310996_492/data_in
+ scan_wrapper_334445762078310996_491/latch_enable_in scan_wrapper_334445762078310996_492/latch_enable_in
+ scan_wrapper_334445762078310996_491/scan_select_in scan_wrapper_334445762078310996_492/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_480 scan_wrapper_334445762078310996_480/clk_in scan_wrapper_334445762078310996_481/clk_in
+ scan_wrapper_334445762078310996_480/data_in scan_wrapper_334445762078310996_481/data_in
+ scan_wrapper_334445762078310996_480/latch_enable_in scan_wrapper_334445762078310996_481/latch_enable_in
+ scan_wrapper_334445762078310996_480/scan_select_in scan_wrapper_334445762078310996_481/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_89 scan_wrapper_334445762078310996_89/clk_in scan_wrapper_334445762078310996_90/clk_in
+ scan_wrapper_334445762078310996_89/data_in scan_wrapper_334445762078310996_90/data_in
+ scan_wrapper_334445762078310996_89/latch_enable_in scan_wrapper_334445762078310996_90/latch_enable_in
+ scan_wrapper_334445762078310996_89/scan_select_in scan_wrapper_334445762078310996_90/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_78 scan_wrapper_334445762078310996_78/clk_in scan_wrapper_334445762078310996_79/clk_in
+ scan_wrapper_334445762078310996_78/data_in scan_wrapper_334445762078310996_79/data_in
+ scan_wrapper_334445762078310996_78/latch_enable_in scan_wrapper_334445762078310996_79/latch_enable_in
+ scan_wrapper_334445762078310996_78/scan_select_in scan_wrapper_334445762078310996_79/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_67 scan_wrapper_334445762078310996_67/clk_in scan_wrapper_334445762078310996_68/clk_in
+ scan_wrapper_334445762078310996_67/data_in scan_wrapper_334445762078310996_68/data_in
+ scan_wrapper_334445762078310996_67/latch_enable_in scan_wrapper_334445762078310996_68/latch_enable_in
+ scan_wrapper_334445762078310996_67/scan_select_in scan_wrapper_334445762078310996_68/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_56 scan_wrapper_334445762078310996_56/clk_in scan_wrapper_334445762078310996_57/clk_in
+ scan_wrapper_334445762078310996_56/data_in scan_wrapper_334445762078310996_57/data_in
+ scan_wrapper_334445762078310996_56/latch_enable_in scan_wrapper_334445762078310996_57/latch_enable_in
+ scan_wrapper_334445762078310996_56/scan_select_in scan_wrapper_334445762078310996_57/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_45 scan_wrapper_334445762078310996_45/clk_in scan_wrapper_334445762078310996_46/clk_in
+ scan_wrapper_334445762078310996_45/data_in scan_wrapper_334445762078310996_46/data_in
+ scan_wrapper_334445762078310996_45/latch_enable_in scan_wrapper_334445762078310996_46/latch_enable_in
+ scan_wrapper_334445762078310996_45/scan_select_in scan_wrapper_334445762078310996_46/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_34 scan_wrapper_334445762078310996_34/clk_in scan_wrapper_334445762078310996_35/clk_in
+ scan_wrapper_334445762078310996_34/data_in scan_wrapper_334445762078310996_35/data_in
+ scan_wrapper_334445762078310996_34/latch_enable_in scan_wrapper_334445762078310996_35/latch_enable_in
+ scan_wrapper_334445762078310996_34/scan_select_in scan_wrapper_334445762078310996_35/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_23 scan_wrapper_334445762078310996_23/clk_in scan_wrapper_334445762078310996_24/clk_in
+ scan_wrapper_334445762078310996_23/data_in scan_wrapper_334445762078310996_24/data_in
+ scan_wrapper_334445762078310996_23/latch_enable_in scan_wrapper_334445762078310996_24/latch_enable_in
+ scan_wrapper_334445762078310996_23/scan_select_in scan_wrapper_334445762078310996_24/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_12 scan_wrapper_334445762078310996_12/clk_in scan_wrapper_334445762078310996_13/clk_in
+ scan_wrapper_334445762078310996_12/data_in scan_wrapper_334445762078310996_13/data_in
+ scan_wrapper_334445762078310996_12/latch_enable_in scan_wrapper_334445762078310996_13/latch_enable_in
+ scan_wrapper_334445762078310996_12/scan_select_in scan_wrapper_334445762078310996_13/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_309 scan_wrapper_334445762078310996_309/clk_in scan_wrapper_334445762078310996_310/clk_in
+ scan_wrapper_334445762078310996_309/data_in scan_wrapper_334445762078310996_310/data_in
+ scan_wrapper_334445762078310996_309/latch_enable_in scan_wrapper_334445762078310996_310/latch_enable_in
+ scan_wrapper_334445762078310996_309/scan_select_in scan_wrapper_334445762078310996_310/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_106 scan_wrapper_334445762078310996_106/clk_in scan_wrapper_334445762078310996_107/clk_in
+ scan_wrapper_334445762078310996_106/data_in scan_wrapper_334445762078310996_107/data_in
+ scan_wrapper_334445762078310996_106/latch_enable_in scan_wrapper_334445762078310996_107/latch_enable_in
+ scan_wrapper_334445762078310996_106/scan_select_in scan_wrapper_334445762078310996_107/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_117 scan_wrapper_334445762078310996_117/clk_in scan_wrapper_334445762078310996_118/clk_in
+ scan_wrapper_334445762078310996_117/data_in scan_wrapper_334445762078310996_118/data_in
+ scan_wrapper_334445762078310996_117/latch_enable_in scan_wrapper_334445762078310996_118/latch_enable_in
+ scan_wrapper_334445762078310996_117/scan_select_in scan_wrapper_334445762078310996_118/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_128 scan_wrapper_334445762078310996_128/clk_in scan_wrapper_334445762078310996_129/clk_in
+ scan_wrapper_334445762078310996_128/data_in scan_wrapper_334445762078310996_129/data_in
+ scan_wrapper_334445762078310996_128/latch_enable_in scan_wrapper_334445762078310996_129/latch_enable_in
+ scan_wrapper_334445762078310996_128/scan_select_in scan_wrapper_334445762078310996_129/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_139 scan_wrapper_334445762078310996_139/clk_in scan_wrapper_334445762078310996_140/clk_in
+ scan_wrapper_334445762078310996_139/data_in scan_wrapper_334445762078310996_140/data_in
+ scan_wrapper_334445762078310996_139/latch_enable_in scan_wrapper_334445762078310996_140/latch_enable_in
+ scan_wrapper_334445762078310996_139/scan_select_in scan_wrapper_334445762078310996_140/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_492 scan_wrapper_334445762078310996_492/clk_in scan_wrapper_334445762078310996_493/clk_in
+ scan_wrapper_334445762078310996_492/data_in scan_wrapper_334445762078310996_493/data_in
+ scan_wrapper_334445762078310996_492/latch_enable_in scan_wrapper_334445762078310996_493/latch_enable_in
+ scan_wrapper_334445762078310996_492/scan_select_in scan_wrapper_334445762078310996_493/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_481 scan_wrapper_334445762078310996_481/clk_in scan_wrapper_334445762078310996_482/clk_in
+ scan_wrapper_334445762078310996_481/data_in scan_wrapper_334445762078310996_482/data_in
+ scan_wrapper_334445762078310996_481/latch_enable_in scan_wrapper_334445762078310996_482/latch_enable_in
+ scan_wrapper_334445762078310996_481/scan_select_in scan_wrapper_334445762078310996_482/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_470 scan_wrapper_334445762078310996_470/clk_in scan_wrapper_334445762078310996_471/clk_in
+ scan_wrapper_334445762078310996_470/data_in scan_wrapper_334445762078310996_471/data_in
+ scan_wrapper_334445762078310996_470/latch_enable_in scan_wrapper_334445762078310996_471/latch_enable_in
+ scan_wrapper_334445762078310996_470/scan_select_in scan_wrapper_334445762078310996_471/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_79 scan_wrapper_334445762078310996_79/clk_in scan_wrapper_334445762078310996_80/clk_in
+ scan_wrapper_334445762078310996_79/data_in scan_wrapper_334445762078310996_80/data_in
+ scan_wrapper_334445762078310996_79/latch_enable_in scan_wrapper_334445762078310996_80/latch_enable_in
+ scan_wrapper_334445762078310996_79/scan_select_in scan_wrapper_334445762078310996_80/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_68 scan_wrapper_334445762078310996_68/clk_in scan_wrapper_334445762078310996_69/clk_in
+ scan_wrapper_334445762078310996_68/data_in scan_wrapper_334445762078310996_69/data_in
+ scan_wrapper_334445762078310996_68/latch_enable_in scan_wrapper_334445762078310996_69/latch_enable_in
+ scan_wrapper_334445762078310996_68/scan_select_in scan_wrapper_334445762078310996_69/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_57 scan_wrapper_334445762078310996_57/clk_in scan_wrapper_334445762078310996_58/clk_in
+ scan_wrapper_334445762078310996_57/data_in scan_wrapper_334445762078310996_58/data_in
+ scan_wrapper_334445762078310996_57/latch_enable_in scan_wrapper_334445762078310996_58/latch_enable_in
+ scan_wrapper_334445762078310996_57/scan_select_in scan_wrapper_334445762078310996_58/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_46 scan_wrapper_334445762078310996_46/clk_in scan_wrapper_334445762078310996_47/clk_in
+ scan_wrapper_334445762078310996_46/data_in scan_wrapper_334445762078310996_47/data_in
+ scan_wrapper_334445762078310996_46/latch_enable_in scan_wrapper_334445762078310996_47/latch_enable_in
+ scan_wrapper_334445762078310996_46/scan_select_in scan_wrapper_334445762078310996_47/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_35 scan_wrapper_334445762078310996_35/clk_in scan_wrapper_334445762078310996_36/clk_in
+ scan_wrapper_334445762078310996_35/data_in scan_wrapper_334445762078310996_36/data_in
+ scan_wrapper_334445762078310996_35/latch_enable_in scan_wrapper_334445762078310996_36/latch_enable_in
+ scan_wrapper_334445762078310996_35/scan_select_in scan_wrapper_334445762078310996_36/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_24 scan_wrapper_334445762078310996_24/clk_in scan_wrapper_334445762078310996_25/clk_in
+ scan_wrapper_334445762078310996_24/data_in scan_wrapper_334445762078310996_25/data_in
+ scan_wrapper_334445762078310996_24/latch_enable_in scan_wrapper_334445762078310996_25/latch_enable_in
+ scan_wrapper_334445762078310996_24/scan_select_in scan_wrapper_334445762078310996_25/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_13 scan_wrapper_334445762078310996_13/clk_in scan_wrapper_334445762078310996_14/clk_in
+ scan_wrapper_334445762078310996_13/data_in scan_wrapper_334445762078310996_14/data_in
+ scan_wrapper_334445762078310996_13/latch_enable_in scan_wrapper_334445762078310996_14/latch_enable_in
+ scan_wrapper_334445762078310996_13/scan_select_in scan_wrapper_334445762078310996_14/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_107 scan_wrapper_334445762078310996_107/clk_in scan_wrapper_334445762078310996_108/clk_in
+ scan_wrapper_334445762078310996_107/data_in scan_wrapper_334445762078310996_108/data_in
+ scan_wrapper_334445762078310996_107/latch_enable_in scan_wrapper_334445762078310996_108/latch_enable_in
+ scan_wrapper_334445762078310996_107/scan_select_in scan_wrapper_334445762078310996_108/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_118 scan_wrapper_334445762078310996_118/clk_in scan_wrapper_334445762078310996_119/clk_in
+ scan_wrapper_334445762078310996_118/data_in scan_wrapper_334445762078310996_119/data_in
+ scan_wrapper_334445762078310996_118/latch_enable_in scan_wrapper_334445762078310996_119/latch_enable_in
+ scan_wrapper_334445762078310996_118/scan_select_in scan_wrapper_334445762078310996_119/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_129 scan_wrapper_334445762078310996_129/clk_in scan_wrapper_334445762078310996_130/clk_in
+ scan_wrapper_334445762078310996_129/data_in scan_wrapper_334445762078310996_130/data_in
+ scan_wrapper_334445762078310996_129/latch_enable_in scan_wrapper_334445762078310996_130/latch_enable_in
+ scan_wrapper_334445762078310996_129/scan_select_in scan_wrapper_334445762078310996_130/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_493 scan_wrapper_334445762078310996_493/clk_in scan_wrapper_334445762078310996_494/clk_in
+ scan_wrapper_334445762078310996_493/data_in scan_wrapper_334445762078310996_494/data_in
+ scan_wrapper_334445762078310996_493/latch_enable_in scan_wrapper_334445762078310996_494/latch_enable_in
+ scan_wrapper_334445762078310996_493/scan_select_in scan_wrapper_334445762078310996_494/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_482 scan_wrapper_334445762078310996_482/clk_in scan_wrapper_334445762078310996_483/clk_in
+ scan_wrapper_334445762078310996_482/data_in scan_wrapper_334445762078310996_483/data_in
+ scan_wrapper_334445762078310996_482/latch_enable_in scan_wrapper_334445762078310996_483/latch_enable_in
+ scan_wrapper_334445762078310996_482/scan_select_in scan_wrapper_334445762078310996_483/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_471 scan_wrapper_334445762078310996_471/clk_in scan_wrapper_334445762078310996_472/clk_in
+ scan_wrapper_334445762078310996_471/data_in scan_wrapper_334445762078310996_472/data_in
+ scan_wrapper_334445762078310996_471/latch_enable_in scan_wrapper_334445762078310996_472/latch_enable_in
+ scan_wrapper_334445762078310996_471/scan_select_in scan_wrapper_334445762078310996_472/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_460 scan_wrapper_334445762078310996_460/clk_in scan_wrapper_334445762078310996_461/clk_in
+ scan_wrapper_334445762078310996_460/data_in scan_wrapper_334445762078310996_461/data_in
+ scan_wrapper_334445762078310996_460/latch_enable_in scan_wrapper_334445762078310996_461/latch_enable_in
+ scan_wrapper_334445762078310996_460/scan_select_in scan_wrapper_334445762078310996_461/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_290 scan_wrapper_334445762078310996_290/clk_in scan_wrapper_334445762078310996_291/clk_in
+ scan_wrapper_334445762078310996_290/data_in scan_wrapper_334445762078310996_291/data_in
+ scan_wrapper_334445762078310996_290/latch_enable_in scan_wrapper_334445762078310996_291/latch_enable_in
+ scan_wrapper_334445762078310996_290/scan_select_in scan_wrapper_334445762078310996_291/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_69 scan_wrapper_334445762078310996_69/clk_in scan_wrapper_334445762078310996_70/clk_in
+ scan_wrapper_334445762078310996_69/data_in scan_wrapper_334445762078310996_70/data_in
+ scan_wrapper_334445762078310996_69/latch_enable_in scan_wrapper_334445762078310996_70/latch_enable_in
+ scan_wrapper_334445762078310996_69/scan_select_in scan_wrapper_334445762078310996_70/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_58 scan_wrapper_334445762078310996_58/clk_in scan_wrapper_334445762078310996_59/clk_in
+ scan_wrapper_334445762078310996_58/data_in scan_wrapper_334445762078310996_59/data_in
+ scan_wrapper_334445762078310996_58/latch_enable_in scan_wrapper_334445762078310996_59/latch_enable_in
+ scan_wrapper_334445762078310996_58/scan_select_in scan_wrapper_334445762078310996_59/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_47 scan_wrapper_334445762078310996_47/clk_in scan_wrapper_334445762078310996_48/clk_in
+ scan_wrapper_334445762078310996_47/data_in scan_wrapper_334445762078310996_48/data_in
+ scan_wrapper_334445762078310996_47/latch_enable_in scan_wrapper_334445762078310996_48/latch_enable_in
+ scan_wrapper_334445762078310996_47/scan_select_in scan_wrapper_334445762078310996_48/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_36 scan_wrapper_334445762078310996_36/clk_in scan_wrapper_334445762078310996_37/clk_in
+ scan_wrapper_334445762078310996_36/data_in scan_wrapper_334445762078310996_37/data_in
+ scan_wrapper_334445762078310996_36/latch_enable_in scan_wrapper_334445762078310996_37/latch_enable_in
+ scan_wrapper_334445762078310996_36/scan_select_in scan_wrapper_334445762078310996_37/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_25 scan_wrapper_334445762078310996_25/clk_in scan_wrapper_334445762078310996_26/clk_in
+ scan_wrapper_334445762078310996_25/data_in scan_wrapper_334445762078310996_26/data_in
+ scan_wrapper_334445762078310996_25/latch_enable_in scan_wrapper_334445762078310996_26/latch_enable_in
+ scan_wrapper_334445762078310996_25/scan_select_in scan_wrapper_334445762078310996_26/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_14 scan_wrapper_334445762078310996_14/clk_in scan_wrapper_334445762078310996_15/clk_in
+ scan_wrapper_334445762078310996_14/data_in scan_wrapper_334445762078310996_15/data_in
+ scan_wrapper_334445762078310996_14/latch_enable_in scan_wrapper_334445762078310996_15/latch_enable_in
+ scan_wrapper_334445762078310996_14/scan_select_in scan_wrapper_334445762078310996_15/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_108 scan_wrapper_334445762078310996_108/clk_in scan_wrapper_334445762078310996_109/clk_in
+ scan_wrapper_334445762078310996_108/data_in scan_wrapper_334445762078310996_109/data_in
+ scan_wrapper_334445762078310996_108/latch_enable_in scan_wrapper_334445762078310996_109/latch_enable_in
+ scan_wrapper_334445762078310996_108/scan_select_in scan_wrapper_334445762078310996_109/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_119 scan_wrapper_334445762078310996_119/clk_in scan_wrapper_334445762078310996_120/clk_in
+ scan_wrapper_334445762078310996_119/data_in scan_wrapper_334445762078310996_120/data_in
+ scan_wrapper_334445762078310996_119/latch_enable_in scan_wrapper_334445762078310996_120/latch_enable_in
+ scan_wrapper_334445762078310996_119/scan_select_in scan_wrapper_334445762078310996_120/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_494 scan_wrapper_334445762078310996_494/clk_in scan_wrapper_334445762078310996_495/clk_in
+ scan_wrapper_334445762078310996_494/data_in scan_wrapper_334445762078310996_495/data_in
+ scan_wrapper_334445762078310996_494/latch_enable_in scan_wrapper_334445762078310996_495/latch_enable_in
+ scan_wrapper_334445762078310996_494/scan_select_in scan_wrapper_334445762078310996_495/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_483 scan_wrapper_334445762078310996_483/clk_in scan_wrapper_334445762078310996_484/clk_in
+ scan_wrapper_334445762078310996_483/data_in scan_wrapper_334445762078310996_484/data_in
+ scan_wrapper_334445762078310996_483/latch_enable_in scan_wrapper_334445762078310996_484/latch_enable_in
+ scan_wrapper_334445762078310996_483/scan_select_in scan_wrapper_334445762078310996_484/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_472 scan_wrapper_334445762078310996_472/clk_in scan_wrapper_334445762078310996_473/clk_in
+ scan_wrapper_334445762078310996_472/data_in scan_wrapper_334445762078310996_473/data_in
+ scan_wrapper_334445762078310996_472/latch_enable_in scan_wrapper_334445762078310996_473/latch_enable_in
+ scan_wrapper_334445762078310996_472/scan_select_in scan_wrapper_334445762078310996_473/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_461 scan_wrapper_334445762078310996_461/clk_in scan_wrapper_334445762078310996_462/clk_in
+ scan_wrapper_334445762078310996_461/data_in scan_wrapper_334445762078310996_462/data_in
+ scan_wrapper_334445762078310996_461/latch_enable_in scan_wrapper_334445762078310996_462/latch_enable_in
+ scan_wrapper_334445762078310996_461/scan_select_in scan_wrapper_334445762078310996_462/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_450 scan_wrapper_334445762078310996_450/clk_in scan_wrapper_334445762078310996_451/clk_in
+ scan_wrapper_334445762078310996_450/data_in scan_wrapper_334445762078310996_451/data_in
+ scan_wrapper_334445762078310996_450/latch_enable_in scan_wrapper_334445762078310996_451/latch_enable_in
+ scan_wrapper_334445762078310996_450/scan_select_in scan_wrapper_334445762078310996_451/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_280 scan_wrapper_334445762078310996_280/clk_in scan_wrapper_334445762078310996_281/clk_in
+ scan_wrapper_334445762078310996_280/data_in scan_wrapper_334445762078310996_281/data_in
+ scan_wrapper_334445762078310996_280/latch_enable_in scan_wrapper_334445762078310996_281/latch_enable_in
+ scan_wrapper_334445762078310996_280/scan_select_in scan_wrapper_334445762078310996_281/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_291 scan_wrapper_334445762078310996_291/clk_in scan_wrapper_334445762078310996_292/clk_in
+ scan_wrapper_334445762078310996_291/data_in scan_wrapper_334445762078310996_292/data_in
+ scan_wrapper_334445762078310996_291/latch_enable_in scan_wrapper_334445762078310996_292/latch_enable_in
+ scan_wrapper_334445762078310996_291/scan_select_in scan_wrapper_334445762078310996_292/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_59 scan_wrapper_334445762078310996_59/clk_in scan_wrapper_334445762078310996_60/clk_in
+ scan_wrapper_334445762078310996_59/data_in scan_wrapper_334445762078310996_60/data_in
+ scan_wrapper_334445762078310996_59/latch_enable_in scan_wrapper_334445762078310996_60/latch_enable_in
+ scan_wrapper_334445762078310996_59/scan_select_in scan_wrapper_334445762078310996_60/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_48 scan_wrapper_334445762078310996_48/clk_in scan_wrapper_334445762078310996_49/clk_in
+ scan_wrapper_334445762078310996_48/data_in scan_wrapper_334445762078310996_49/data_in
+ scan_wrapper_334445762078310996_48/latch_enable_in scan_wrapper_334445762078310996_49/latch_enable_in
+ scan_wrapper_334445762078310996_48/scan_select_in scan_wrapper_334445762078310996_49/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_37 scan_wrapper_334445762078310996_37/clk_in scan_wrapper_334445762078310996_38/clk_in
+ scan_wrapper_334445762078310996_37/data_in scan_wrapper_334445762078310996_38/data_in
+ scan_wrapper_334445762078310996_37/latch_enable_in scan_wrapper_334445762078310996_38/latch_enable_in
+ scan_wrapper_334445762078310996_37/scan_select_in scan_wrapper_334445762078310996_38/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_26 scan_wrapper_334445762078310996_26/clk_in scan_wrapper_334445762078310996_27/clk_in
+ scan_wrapper_334445762078310996_26/data_in scan_wrapper_334445762078310996_27/data_in
+ scan_wrapper_334445762078310996_26/latch_enable_in scan_wrapper_334445762078310996_27/latch_enable_in
+ scan_wrapper_334445762078310996_26/scan_select_in scan_wrapper_334445762078310996_27/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_15 scan_wrapper_334445762078310996_15/clk_in scan_wrapper_334445762078310996_16/clk_in
+ scan_wrapper_334445762078310996_15/data_in scan_wrapper_334445762078310996_16/data_in
+ scan_wrapper_334445762078310996_15/latch_enable_in scan_wrapper_334445762078310996_16/latch_enable_in
+ scan_wrapper_334445762078310996_15/scan_select_in scan_wrapper_334445762078310996_16/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_109 scan_wrapper_334445762078310996_109/clk_in scan_wrapper_334445762078310996_110/clk_in
+ scan_wrapper_334445762078310996_109/data_in scan_wrapper_334445762078310996_110/data_in
+ scan_wrapper_334445762078310996_109/latch_enable_in scan_wrapper_334445762078310996_110/latch_enable_in
+ scan_wrapper_334445762078310996_109/scan_select_in scan_wrapper_334445762078310996_110/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_495 scan_wrapper_334445762078310996_495/clk_in scan_wrapper_334445762078310996_496/clk_in
+ scan_wrapper_334445762078310996_495/data_in scan_wrapper_334445762078310996_496/data_in
+ scan_wrapper_334445762078310996_495/latch_enable_in scan_wrapper_334445762078310996_496/latch_enable_in
+ scan_wrapper_334445762078310996_495/scan_select_in scan_wrapper_334445762078310996_496/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_484 scan_wrapper_334445762078310996_484/clk_in scan_wrapper_334445762078310996_485/clk_in
+ scan_wrapper_334445762078310996_484/data_in scan_wrapper_334445762078310996_485/data_in
+ scan_wrapper_334445762078310996_484/latch_enable_in scan_wrapper_334445762078310996_485/latch_enable_in
+ scan_wrapper_334445762078310996_484/scan_select_in scan_wrapper_334445762078310996_485/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_473 scan_wrapper_334445762078310996_473/clk_in scan_wrapper_334445762078310996_474/clk_in
+ scan_wrapper_334445762078310996_473/data_in scan_wrapper_334445762078310996_474/data_in
+ scan_wrapper_334445762078310996_473/latch_enable_in scan_wrapper_334445762078310996_474/latch_enable_in
+ scan_wrapper_334445762078310996_473/scan_select_in scan_wrapper_334445762078310996_474/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_462 scan_wrapper_334445762078310996_462/clk_in scan_wrapper_334445762078310996_463/clk_in
+ scan_wrapper_334445762078310996_462/data_in scan_wrapper_334445762078310996_463/data_in
+ scan_wrapper_334445762078310996_462/latch_enable_in scan_wrapper_334445762078310996_463/latch_enable_in
+ scan_wrapper_334445762078310996_462/scan_select_in scan_wrapper_334445762078310996_463/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_451 scan_wrapper_334445762078310996_451/clk_in scan_wrapper_334445762078310996_452/clk_in
+ scan_wrapper_334445762078310996_451/data_in scan_wrapper_334445762078310996_452/data_in
+ scan_wrapper_334445762078310996_451/latch_enable_in scan_wrapper_334445762078310996_452/latch_enable_in
+ scan_wrapper_334445762078310996_451/scan_select_in scan_wrapper_334445762078310996_452/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_440 scan_wrapper_334445762078310996_440/clk_in scan_wrapper_334445762078310996_441/clk_in
+ scan_wrapper_334445762078310996_440/data_in scan_wrapper_334445762078310996_441/data_in
+ scan_wrapper_334445762078310996_440/latch_enable_in scan_wrapper_334445762078310996_441/latch_enable_in
+ scan_wrapper_334445762078310996_440/scan_select_in scan_wrapper_334445762078310996_441/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_270 scan_wrapper_334445762078310996_270/clk_in scan_wrapper_334445762078310996_271/clk_in
+ scan_wrapper_334445762078310996_270/data_in scan_wrapper_334445762078310996_271/data_in
+ scan_wrapper_334445762078310996_270/latch_enable_in scan_wrapper_334445762078310996_271/latch_enable_in
+ scan_wrapper_334445762078310996_270/scan_select_in scan_wrapper_334445762078310996_271/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_281 scan_wrapper_334445762078310996_281/clk_in scan_wrapper_334445762078310996_282/clk_in
+ scan_wrapper_334445762078310996_281/data_in scan_wrapper_334445762078310996_282/data_in
+ scan_wrapper_334445762078310996_281/latch_enable_in scan_wrapper_334445762078310996_282/latch_enable_in
+ scan_wrapper_334445762078310996_281/scan_select_in scan_wrapper_334445762078310996_282/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_292 scan_wrapper_334445762078310996_292/clk_in scan_wrapper_334445762078310996_293/clk_in
+ scan_wrapper_334445762078310996_292/data_in scan_wrapper_334445762078310996_293/data_in
+ scan_wrapper_334445762078310996_292/latch_enable_in scan_wrapper_334445762078310996_293/latch_enable_in
+ scan_wrapper_334445762078310996_292/scan_select_in scan_wrapper_334445762078310996_293/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_49 scan_wrapper_334445762078310996_49/clk_in scan_wrapper_334445762078310996_50/clk_in
+ scan_wrapper_334445762078310996_49/data_in scan_wrapper_334445762078310996_50/data_in
+ scan_wrapper_334445762078310996_49/latch_enable_in scan_wrapper_334445762078310996_50/latch_enable_in
+ scan_wrapper_334445762078310996_49/scan_select_in scan_wrapper_334445762078310996_50/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_38 scan_wrapper_334445762078310996_38/clk_in scan_wrapper_334445762078310996_39/clk_in
+ scan_wrapper_334445762078310996_38/data_in scan_wrapper_334445762078310996_39/data_in
+ scan_wrapper_334445762078310996_38/latch_enable_in scan_wrapper_334445762078310996_39/latch_enable_in
+ scan_wrapper_334445762078310996_38/scan_select_in scan_wrapper_334445762078310996_39/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_27 scan_wrapper_334445762078310996_27/clk_in scan_wrapper_334445762078310996_28/clk_in
+ scan_wrapper_334445762078310996_27/data_in scan_wrapper_334445762078310996_28/data_in
+ scan_wrapper_334445762078310996_27/latch_enable_in scan_wrapper_334445762078310996_28/latch_enable_in
+ scan_wrapper_334445762078310996_27/scan_select_in scan_wrapper_334445762078310996_28/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_16 scan_wrapper_334445762078310996_16/clk_in scan_wrapper_334445762078310996_17/clk_in
+ scan_wrapper_334445762078310996_16/data_in scan_wrapper_334445762078310996_17/data_in
+ scan_wrapper_334445762078310996_16/latch_enable_in scan_wrapper_334445762078310996_17/latch_enable_in
+ scan_wrapper_334445762078310996_16/scan_select_in scan_wrapper_334445762078310996_17/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_496 scan_wrapper_334445762078310996_496/clk_in scan_wrapper_334445762078310996_497/clk_in
+ scan_wrapper_334445762078310996_496/data_in scan_wrapper_334445762078310996_497/data_in
+ scan_wrapper_334445762078310996_496/latch_enable_in scan_wrapper_334445762078310996_497/latch_enable_in
+ scan_wrapper_334445762078310996_496/scan_select_in scan_wrapper_334445762078310996_497/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_485 scan_wrapper_334445762078310996_485/clk_in scan_wrapper_334445762078310996_486/clk_in
+ scan_wrapper_334445762078310996_485/data_in scan_wrapper_334445762078310996_486/data_in
+ scan_wrapper_334445762078310996_485/latch_enable_in scan_wrapper_334445762078310996_486/latch_enable_in
+ scan_wrapper_334445762078310996_485/scan_select_in scan_wrapper_334445762078310996_486/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_474 scan_wrapper_334445762078310996_474/clk_in scan_wrapper_334445762078310996_475/clk_in
+ scan_wrapper_334445762078310996_474/data_in scan_wrapper_334445762078310996_475/data_in
+ scan_wrapper_334445762078310996_474/latch_enable_in scan_wrapper_334445762078310996_475/latch_enable_in
+ scan_wrapper_334445762078310996_474/scan_select_in scan_wrapper_334445762078310996_475/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_463 scan_wrapper_334445762078310996_463/clk_in scan_wrapper_334445762078310996_464/clk_in
+ scan_wrapper_334445762078310996_463/data_in scan_wrapper_334445762078310996_464/data_in
+ scan_wrapper_334445762078310996_463/latch_enable_in scan_wrapper_334445762078310996_464/latch_enable_in
+ scan_wrapper_334445762078310996_463/scan_select_in scan_wrapper_334445762078310996_464/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_452 scan_wrapper_334445762078310996_452/clk_in scan_wrapper_334445762078310996_453/clk_in
+ scan_wrapper_334445762078310996_452/data_in scan_wrapper_334445762078310996_453/data_in
+ scan_wrapper_334445762078310996_452/latch_enable_in scan_wrapper_334445762078310996_453/latch_enable_in
+ scan_wrapper_334445762078310996_452/scan_select_in scan_wrapper_334445762078310996_453/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_441 scan_wrapper_334445762078310996_441/clk_in scan_wrapper_334445762078310996_442/clk_in
+ scan_wrapper_334445762078310996_441/data_in scan_wrapper_334445762078310996_442/data_in
+ scan_wrapper_334445762078310996_441/latch_enable_in scan_wrapper_334445762078310996_442/latch_enable_in
+ scan_wrapper_334445762078310996_441/scan_select_in scan_wrapper_334445762078310996_442/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_430 scan_wrapper_334445762078310996_430/clk_in scan_wrapper_334445762078310996_431/clk_in
+ scan_wrapper_334445762078310996_430/data_in scan_wrapper_334445762078310996_431/data_in
+ scan_wrapper_334445762078310996_430/latch_enable_in scan_wrapper_334445762078310996_431/latch_enable_in
+ scan_wrapper_334445762078310996_430/scan_select_in scan_wrapper_334445762078310996_431/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_260 scan_wrapper_334445762078310996_260/clk_in scan_wrapper_334445762078310996_261/clk_in
+ scan_wrapper_334445762078310996_260/data_in scan_wrapper_334445762078310996_261/data_in
+ scan_wrapper_334445762078310996_260/latch_enable_in scan_wrapper_334445762078310996_261/latch_enable_in
+ scan_wrapper_334445762078310996_260/scan_select_in scan_wrapper_334445762078310996_261/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_271 scan_wrapper_334445762078310996_271/clk_in scan_wrapper_334445762078310996_272/clk_in
+ scan_wrapper_334445762078310996_271/data_in scan_wrapper_334445762078310996_272/data_in
+ scan_wrapper_334445762078310996_271/latch_enable_in scan_wrapper_334445762078310996_272/latch_enable_in
+ scan_wrapper_334445762078310996_271/scan_select_in scan_wrapper_334445762078310996_272/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_282 scan_wrapper_334445762078310996_282/clk_in scan_wrapper_334445762078310996_283/clk_in
+ scan_wrapper_334445762078310996_282/data_in scan_wrapper_334445762078310996_283/data_in
+ scan_wrapper_334445762078310996_282/latch_enable_in scan_wrapper_334445762078310996_283/latch_enable_in
+ scan_wrapper_334445762078310996_282/scan_select_in scan_wrapper_334445762078310996_283/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_293 scan_wrapper_334445762078310996_293/clk_in scan_wrapper_334445762078310996_294/clk_in
+ scan_wrapper_334445762078310996_293/data_in scan_wrapper_334445762078310996_294/data_in
+ scan_wrapper_334445762078310996_293/latch_enable_in scan_wrapper_334445762078310996_294/latch_enable_in
+ scan_wrapper_334445762078310996_293/scan_select_in scan_wrapper_334445762078310996_294/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_39 scan_wrapper_334445762078310996_39/clk_in scan_wrapper_334445762078310996_40/clk_in
+ scan_wrapper_334445762078310996_39/data_in scan_wrapper_334445762078310996_40/data_in
+ scan_wrapper_334445762078310996_39/latch_enable_in scan_wrapper_334445762078310996_40/latch_enable_in
+ scan_wrapper_334445762078310996_39/scan_select_in scan_wrapper_334445762078310996_40/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_28 scan_wrapper_334445762078310996_28/clk_in scan_wrapper_334445762078310996_29/clk_in
+ scan_wrapper_334445762078310996_28/data_in scan_wrapper_334445762078310996_29/data_in
+ scan_wrapper_334445762078310996_28/latch_enable_in scan_wrapper_334445762078310996_29/latch_enable_in
+ scan_wrapper_334445762078310996_28/scan_select_in scan_wrapper_334445762078310996_29/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_17 scan_wrapper_334445762078310996_17/clk_in scan_wrapper_334445762078310996_18/clk_in
+ scan_wrapper_334445762078310996_17/data_in scan_wrapper_334445762078310996_18/data_in
+ scan_wrapper_334445762078310996_17/latch_enable_in scan_wrapper_334445762078310996_18/latch_enable_in
+ scan_wrapper_334445762078310996_17/scan_select_in scan_wrapper_334445762078310996_18/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_497 scan_wrapper_334445762078310996_497/clk_in scan_wrapper_334445762078310996_497/clk_out
+ scan_wrapper_334445762078310996_497/data_in scan_controller/scan_data_in scan_wrapper_334445762078310996_497/latch_enable_in
+ scan_wrapper_334445762078310996_497/latch_enable_out scan_wrapper_334445762078310996_497/scan_select_in
+ scan_wrapper_334445762078310996_497/scan_select_out vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_486 scan_wrapper_334445762078310996_486/clk_in scan_wrapper_334445762078310996_487/clk_in
+ scan_wrapper_334445762078310996_486/data_in scan_wrapper_334445762078310996_487/data_in
+ scan_wrapper_334445762078310996_486/latch_enable_in scan_wrapper_334445762078310996_487/latch_enable_in
+ scan_wrapper_334445762078310996_486/scan_select_in scan_wrapper_334445762078310996_487/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_475 scan_wrapper_334445762078310996_475/clk_in scan_wrapper_334445762078310996_476/clk_in
+ scan_wrapper_334445762078310996_475/data_in scan_wrapper_334445762078310996_476/data_in
+ scan_wrapper_334445762078310996_475/latch_enable_in scan_wrapper_334445762078310996_476/latch_enable_in
+ scan_wrapper_334445762078310996_475/scan_select_in scan_wrapper_334445762078310996_476/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_464 scan_wrapper_334445762078310996_464/clk_in scan_wrapper_334445762078310996_465/clk_in
+ scan_wrapper_334445762078310996_464/data_in scan_wrapper_334445762078310996_465/data_in
+ scan_wrapper_334445762078310996_464/latch_enable_in scan_wrapper_334445762078310996_465/latch_enable_in
+ scan_wrapper_334445762078310996_464/scan_select_in scan_wrapper_334445762078310996_465/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_453 scan_wrapper_334445762078310996_453/clk_in scan_wrapper_334445762078310996_454/clk_in
+ scan_wrapper_334445762078310996_453/data_in scan_wrapper_334445762078310996_454/data_in
+ scan_wrapper_334445762078310996_453/latch_enable_in scan_wrapper_334445762078310996_454/latch_enable_in
+ scan_wrapper_334445762078310996_453/scan_select_in scan_wrapper_334445762078310996_454/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_442 scan_wrapper_334445762078310996_442/clk_in scan_wrapper_334445762078310996_443/clk_in
+ scan_wrapper_334445762078310996_442/data_in scan_wrapper_334445762078310996_443/data_in
+ scan_wrapper_334445762078310996_442/latch_enable_in scan_wrapper_334445762078310996_443/latch_enable_in
+ scan_wrapper_334445762078310996_442/scan_select_in scan_wrapper_334445762078310996_443/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_431 scan_wrapper_334445762078310996_431/clk_in scan_wrapper_334445762078310996_432/clk_in
+ scan_wrapper_334445762078310996_431/data_in scan_wrapper_334445762078310996_432/data_in
+ scan_wrapper_334445762078310996_431/latch_enable_in scan_wrapper_334445762078310996_432/latch_enable_in
+ scan_wrapper_334445762078310996_431/scan_select_in scan_wrapper_334445762078310996_432/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_420 scan_wrapper_334445762078310996_420/clk_in scan_wrapper_334445762078310996_421/clk_in
+ scan_wrapper_334445762078310996_420/data_in scan_wrapper_334445762078310996_421/data_in
+ scan_wrapper_334445762078310996_420/latch_enable_in scan_wrapper_334445762078310996_421/latch_enable_in
+ scan_wrapper_334445762078310996_420/scan_select_in scan_wrapper_334445762078310996_421/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_250 scan_wrapper_334445762078310996_250/clk_in scan_wrapper_334445762078310996_251/clk_in
+ scan_wrapper_334445762078310996_250/data_in scan_wrapper_334445762078310996_251/data_in
+ scan_wrapper_334445762078310996_250/latch_enable_in scan_wrapper_334445762078310996_251/latch_enable_in
+ scan_wrapper_334445762078310996_250/scan_select_in scan_wrapper_334445762078310996_251/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_261 scan_wrapper_334445762078310996_261/clk_in scan_wrapper_334445762078310996_262/clk_in
+ scan_wrapper_334445762078310996_261/data_in scan_wrapper_334445762078310996_262/data_in
+ scan_wrapper_334445762078310996_261/latch_enable_in scan_wrapper_334445762078310996_262/latch_enable_in
+ scan_wrapper_334445762078310996_261/scan_select_in scan_wrapper_334445762078310996_262/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_272 scan_wrapper_334445762078310996_272/clk_in scan_wrapper_334445762078310996_273/clk_in
+ scan_wrapper_334445762078310996_272/data_in scan_wrapper_334445762078310996_273/data_in
+ scan_wrapper_334445762078310996_272/latch_enable_in scan_wrapper_334445762078310996_273/latch_enable_in
+ scan_wrapper_334445762078310996_272/scan_select_in scan_wrapper_334445762078310996_273/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_283 scan_wrapper_334445762078310996_283/clk_in scan_wrapper_334445762078310996_284/clk_in
+ scan_wrapper_334445762078310996_283/data_in scan_wrapper_334445762078310996_284/data_in
+ scan_wrapper_334445762078310996_283/latch_enable_in scan_wrapper_334445762078310996_284/latch_enable_in
+ scan_wrapper_334445762078310996_283/scan_select_in scan_wrapper_334445762078310996_284/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_294 scan_wrapper_334445762078310996_294/clk_in scan_wrapper_334445762078310996_295/clk_in
+ scan_wrapper_334445762078310996_294/data_in scan_wrapper_334445762078310996_295/data_in
+ scan_wrapper_334445762078310996_294/latch_enable_in scan_wrapper_334445762078310996_295/latch_enable_in
+ scan_wrapper_334445762078310996_294/scan_select_in scan_wrapper_334445762078310996_295/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_29 scan_wrapper_334445762078310996_29/clk_in scan_wrapper_334445762078310996_30/clk_in
+ scan_wrapper_334445762078310996_29/data_in scan_wrapper_334445762078310996_30/data_in
+ scan_wrapper_334445762078310996_29/latch_enable_in scan_wrapper_334445762078310996_30/latch_enable_in
+ scan_wrapper_334445762078310996_29/scan_select_in scan_wrapper_334445762078310996_30/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_18 scan_wrapper_334445762078310996_18/clk_in scan_wrapper_334445762078310996_19/clk_in
+ scan_wrapper_334445762078310996_18/data_in scan_wrapper_334445762078310996_19/data_in
+ scan_wrapper_334445762078310996_18/latch_enable_in scan_wrapper_334445762078310996_19/latch_enable_in
+ scan_wrapper_334445762078310996_18/scan_select_in scan_wrapper_334445762078310996_19/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_0 scan_controller/scan_clk scan_wrapper_335404063203000914_1/clk_in
+ scan_controller/scan_data_out scan_wrapper_335404063203000914_1/data_in scan_controller/scan_latch_enable
+ scan_wrapper_335404063203000914_1/latch_enable_in scan_controller/scan_select scan_wrapper_335404063203000914_1/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_432 scan_wrapper_334445762078310996_432/clk_in scan_wrapper_334445762078310996_433/clk_in
+ scan_wrapper_334445762078310996_432/data_in scan_wrapper_334445762078310996_433/data_in
+ scan_wrapper_334445762078310996_432/latch_enable_in scan_wrapper_334445762078310996_433/latch_enable_in
+ scan_wrapper_334445762078310996_432/scan_select_in scan_wrapper_334445762078310996_433/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_421 scan_wrapper_334445762078310996_421/clk_in scan_wrapper_334445762078310996_422/clk_in
+ scan_wrapper_334445762078310996_421/data_in scan_wrapper_334445762078310996_422/data_in
+ scan_wrapper_334445762078310996_421/latch_enable_in scan_wrapper_334445762078310996_422/latch_enable_in
+ scan_wrapper_334445762078310996_421/scan_select_in scan_wrapper_334445762078310996_422/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_410 scan_wrapper_334445762078310996_410/clk_in scan_wrapper_334445762078310996_411/clk_in
+ scan_wrapper_334445762078310996_410/data_in scan_wrapper_334445762078310996_411/data_in
+ scan_wrapper_334445762078310996_410/latch_enable_in scan_wrapper_334445762078310996_411/latch_enable_in
+ scan_wrapper_334445762078310996_410/scan_select_in scan_wrapper_334445762078310996_411/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_487 scan_wrapper_334445762078310996_487/clk_in scan_wrapper_334445762078310996_488/clk_in
+ scan_wrapper_334445762078310996_487/data_in scan_wrapper_334445762078310996_488/data_in
+ scan_wrapper_334445762078310996_487/latch_enable_in scan_wrapper_334445762078310996_488/latch_enable_in
+ scan_wrapper_334445762078310996_487/scan_select_in scan_wrapper_334445762078310996_488/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_476 scan_wrapper_334445762078310996_476/clk_in scan_wrapper_334445762078310996_477/clk_in
+ scan_wrapper_334445762078310996_476/data_in scan_wrapper_334445762078310996_477/data_in
+ scan_wrapper_334445762078310996_476/latch_enable_in scan_wrapper_334445762078310996_477/latch_enable_in
+ scan_wrapper_334445762078310996_476/scan_select_in scan_wrapper_334445762078310996_477/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_465 scan_wrapper_334445762078310996_465/clk_in scan_wrapper_334445762078310996_466/clk_in
+ scan_wrapper_334445762078310996_465/data_in scan_wrapper_334445762078310996_466/data_in
+ scan_wrapper_334445762078310996_465/latch_enable_in scan_wrapper_334445762078310996_466/latch_enable_in
+ scan_wrapper_334445762078310996_465/scan_select_in scan_wrapper_334445762078310996_466/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_454 scan_wrapper_334445762078310996_454/clk_in scan_wrapper_334445762078310996_455/clk_in
+ scan_wrapper_334445762078310996_454/data_in scan_wrapper_334445762078310996_455/data_in
+ scan_wrapper_334445762078310996_454/latch_enable_in scan_wrapper_334445762078310996_455/latch_enable_in
+ scan_wrapper_334445762078310996_454/scan_select_in scan_wrapper_334445762078310996_455/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_443 scan_wrapper_334445762078310996_443/clk_in scan_wrapper_334445762078310996_444/clk_in
+ scan_wrapper_334445762078310996_443/data_in scan_wrapper_334445762078310996_444/data_in
+ scan_wrapper_334445762078310996_443/latch_enable_in scan_wrapper_334445762078310996_444/latch_enable_in
+ scan_wrapper_334445762078310996_443/scan_select_in scan_wrapper_334445762078310996_444/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_240 scan_wrapper_334445762078310996_240/clk_in scan_wrapper_334445762078310996_241/clk_in
+ scan_wrapper_334445762078310996_240/data_in scan_wrapper_334445762078310996_241/data_in
+ scan_wrapper_334445762078310996_240/latch_enable_in scan_wrapper_334445762078310996_241/latch_enable_in
+ scan_wrapper_334445762078310996_240/scan_select_in scan_wrapper_334445762078310996_241/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_251 scan_wrapper_334445762078310996_251/clk_in scan_wrapper_334445762078310996_252/clk_in
+ scan_wrapper_334445762078310996_251/data_in scan_wrapper_334445762078310996_252/data_in
+ scan_wrapper_334445762078310996_251/latch_enable_in scan_wrapper_334445762078310996_252/latch_enable_in
+ scan_wrapper_334445762078310996_251/scan_select_in scan_wrapper_334445762078310996_252/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_262 scan_wrapper_334445762078310996_262/clk_in scan_wrapper_334445762078310996_263/clk_in
+ scan_wrapper_334445762078310996_262/data_in scan_wrapper_334445762078310996_263/data_in
+ scan_wrapper_334445762078310996_262/latch_enable_in scan_wrapper_334445762078310996_263/latch_enable_in
+ scan_wrapper_334445762078310996_262/scan_select_in scan_wrapper_334445762078310996_263/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_273 scan_wrapper_334445762078310996_273/clk_in scan_wrapper_334445762078310996_274/clk_in
+ scan_wrapper_334445762078310996_273/data_in scan_wrapper_334445762078310996_274/data_in
+ scan_wrapper_334445762078310996_273/latch_enable_in scan_wrapper_334445762078310996_274/latch_enable_in
+ scan_wrapper_334445762078310996_273/scan_select_in scan_wrapper_334445762078310996_274/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_284 scan_wrapper_334445762078310996_284/clk_in scan_wrapper_334445762078310996_285/clk_in
+ scan_wrapper_334445762078310996_284/data_in scan_wrapper_334445762078310996_285/data_in
+ scan_wrapper_334445762078310996_284/latch_enable_in scan_wrapper_334445762078310996_285/latch_enable_in
+ scan_wrapper_334445762078310996_284/scan_select_in scan_wrapper_334445762078310996_285/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_295 scan_wrapper_334445762078310996_295/clk_in scan_wrapper_334445762078310996_296/clk_in
+ scan_wrapper_334445762078310996_295/data_in scan_wrapper_334445762078310996_296/data_in
+ scan_wrapper_334445762078310996_295/latch_enable_in scan_wrapper_334445762078310996_296/latch_enable_in
+ scan_wrapper_334445762078310996_295/scan_select_in scan_wrapper_334445762078310996_296/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_19 scan_wrapper_334445762078310996_19/clk_in scan_wrapper_334445762078310996_20/clk_in
+ scan_wrapper_334445762078310996_19/data_in scan_wrapper_334445762078310996_20/data_in
+ scan_wrapper_334445762078310996_19/latch_enable_in scan_wrapper_334445762078310996_20/latch_enable_in
+ scan_wrapper_334445762078310996_19/scan_select_in scan_wrapper_334445762078310996_20/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_488 scan_wrapper_334445762078310996_488/clk_in scan_wrapper_334445762078310996_489/clk_in
+ scan_wrapper_334445762078310996_488/data_in scan_wrapper_334445762078310996_489/data_in
+ scan_wrapper_334445762078310996_488/latch_enable_in scan_wrapper_334445762078310996_489/latch_enable_in
+ scan_wrapper_334445762078310996_488/scan_select_in scan_wrapper_334445762078310996_489/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_477 scan_wrapper_334445762078310996_477/clk_in scan_wrapper_334445762078310996_478/clk_in
+ scan_wrapper_334445762078310996_477/data_in scan_wrapper_334445762078310996_478/data_in
+ scan_wrapper_334445762078310996_477/latch_enable_in scan_wrapper_334445762078310996_478/latch_enable_in
+ scan_wrapper_334445762078310996_477/scan_select_in scan_wrapper_334445762078310996_478/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_466 scan_wrapper_334445762078310996_466/clk_in scan_wrapper_334445762078310996_467/clk_in
+ scan_wrapper_334445762078310996_466/data_in scan_wrapper_334445762078310996_467/data_in
+ scan_wrapper_334445762078310996_466/latch_enable_in scan_wrapper_334445762078310996_467/latch_enable_in
+ scan_wrapper_334445762078310996_466/scan_select_in scan_wrapper_334445762078310996_467/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_455 scan_wrapper_334445762078310996_455/clk_in scan_wrapper_334445762078310996_456/clk_in
+ scan_wrapper_334445762078310996_455/data_in scan_wrapper_334445762078310996_456/data_in
+ scan_wrapper_334445762078310996_455/latch_enable_in scan_wrapper_334445762078310996_456/latch_enable_in
+ scan_wrapper_334445762078310996_455/scan_select_in scan_wrapper_334445762078310996_456/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_444 scan_wrapper_334445762078310996_444/clk_in scan_wrapper_334445762078310996_445/clk_in
+ scan_wrapper_334445762078310996_444/data_in scan_wrapper_334445762078310996_445/data_in
+ scan_wrapper_334445762078310996_444/latch_enable_in scan_wrapper_334445762078310996_445/latch_enable_in
+ scan_wrapper_334445762078310996_444/scan_select_in scan_wrapper_334445762078310996_445/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_433 scan_wrapper_334445762078310996_433/clk_in scan_wrapper_334445762078310996_434/clk_in
+ scan_wrapper_334445762078310996_433/data_in scan_wrapper_334445762078310996_434/data_in
+ scan_wrapper_334445762078310996_433/latch_enable_in scan_wrapper_334445762078310996_434/latch_enable_in
+ scan_wrapper_334445762078310996_433/scan_select_in scan_wrapper_334445762078310996_434/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_422 scan_wrapper_334445762078310996_422/clk_in scan_wrapper_334445762078310996_423/clk_in
+ scan_wrapper_334445762078310996_422/data_in scan_wrapper_334445762078310996_423/data_in
+ scan_wrapper_334445762078310996_422/latch_enable_in scan_wrapper_334445762078310996_423/latch_enable_in
+ scan_wrapper_334445762078310996_422/scan_select_in scan_wrapper_334445762078310996_423/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_411 scan_wrapper_334445762078310996_411/clk_in scan_wrapper_334445762078310996_412/clk_in
+ scan_wrapper_334445762078310996_411/data_in scan_wrapper_334445762078310996_412/data_in
+ scan_wrapper_334445762078310996_411/latch_enable_in scan_wrapper_334445762078310996_412/latch_enable_in
+ scan_wrapper_334445762078310996_411/scan_select_in scan_wrapper_334445762078310996_412/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_400 scan_wrapper_334445762078310996_400/clk_in scan_wrapper_334445762078310996_401/clk_in
+ scan_wrapper_334445762078310996_400/data_in scan_wrapper_334445762078310996_401/data_in
+ scan_wrapper_334445762078310996_400/latch_enable_in scan_wrapper_334445762078310996_401/latch_enable_in
+ scan_wrapper_334445762078310996_400/scan_select_in scan_wrapper_334445762078310996_401/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_230 scan_wrapper_334445762078310996_230/clk_in scan_wrapper_334445762078310996_231/clk_in
+ scan_wrapper_334445762078310996_230/data_in scan_wrapper_334445762078310996_231/data_in
+ scan_wrapper_334445762078310996_230/latch_enable_in scan_wrapper_334445762078310996_231/latch_enable_in
+ scan_wrapper_334445762078310996_230/scan_select_in scan_wrapper_334445762078310996_231/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_241 scan_wrapper_334445762078310996_241/clk_in scan_wrapper_334445762078310996_242/clk_in
+ scan_wrapper_334445762078310996_241/data_in scan_wrapper_334445762078310996_242/data_in
+ scan_wrapper_334445762078310996_241/latch_enable_in scan_wrapper_334445762078310996_242/latch_enable_in
+ scan_wrapper_334445762078310996_241/scan_select_in scan_wrapper_334445762078310996_242/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_252 scan_wrapper_334445762078310996_252/clk_in scan_wrapper_334445762078310996_253/clk_in
+ scan_wrapper_334445762078310996_252/data_in scan_wrapper_334445762078310996_253/data_in
+ scan_wrapper_334445762078310996_252/latch_enable_in scan_wrapper_334445762078310996_253/latch_enable_in
+ scan_wrapper_334445762078310996_252/scan_select_in scan_wrapper_334445762078310996_253/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_263 scan_wrapper_334445762078310996_263/clk_in scan_wrapper_334445762078310996_264/clk_in
+ scan_wrapper_334445762078310996_263/data_in scan_wrapper_334445762078310996_264/data_in
+ scan_wrapper_334445762078310996_263/latch_enable_in scan_wrapper_334445762078310996_264/latch_enable_in
+ scan_wrapper_334445762078310996_263/scan_select_in scan_wrapper_334445762078310996_264/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_274 scan_wrapper_334445762078310996_274/clk_in scan_wrapper_334445762078310996_275/clk_in
+ scan_wrapper_334445762078310996_274/data_in scan_wrapper_334445762078310996_275/data_in
+ scan_wrapper_334445762078310996_274/latch_enable_in scan_wrapper_334445762078310996_275/latch_enable_in
+ scan_wrapper_334445762078310996_274/scan_select_in scan_wrapper_334445762078310996_275/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_285 scan_wrapper_334445762078310996_285/clk_in scan_wrapper_334445762078310996_286/clk_in
+ scan_wrapper_334445762078310996_285/data_in scan_wrapper_334445762078310996_286/data_in
+ scan_wrapper_334445762078310996_285/latch_enable_in scan_wrapper_334445762078310996_286/latch_enable_in
+ scan_wrapper_334445762078310996_285/scan_select_in scan_wrapper_334445762078310996_286/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_296 scan_wrapper_334445762078310996_296/clk_in scan_wrapper_334445762078310996_297/clk_in
+ scan_wrapper_334445762078310996_296/data_in scan_wrapper_334445762078310996_297/data_in
+ scan_wrapper_334445762078310996_296/latch_enable_in scan_wrapper_334445762078310996_297/latch_enable_in
+ scan_wrapper_334445762078310996_296/scan_select_in scan_wrapper_334445762078310996_297/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_2 scan_wrapper_334445762078310996_2/clk_in scan_wrapper_334445762078310996_3/clk_in
+ scan_wrapper_334445762078310996_2/data_in scan_wrapper_334445762078310996_3/data_in
+ scan_wrapper_334445762078310996_2/latch_enable_in scan_wrapper_334445762078310996_3/latch_enable_in
+ scan_wrapper_334445762078310996_2/scan_select_in scan_wrapper_334445762078310996_3/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_489 scan_wrapper_334445762078310996_489/clk_in scan_wrapper_334445762078310996_490/clk_in
+ scan_wrapper_334445762078310996_489/data_in scan_wrapper_334445762078310996_490/data_in
+ scan_wrapper_334445762078310996_489/latch_enable_in scan_wrapper_334445762078310996_490/latch_enable_in
+ scan_wrapper_334445762078310996_489/scan_select_in scan_wrapper_334445762078310996_490/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_478 scan_wrapper_334445762078310996_478/clk_in scan_wrapper_334445762078310996_479/clk_in
+ scan_wrapper_334445762078310996_478/data_in scan_wrapper_334445762078310996_479/data_in
+ scan_wrapper_334445762078310996_478/latch_enable_in scan_wrapper_334445762078310996_479/latch_enable_in
+ scan_wrapper_334445762078310996_478/scan_select_in scan_wrapper_334445762078310996_479/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_467 scan_wrapper_334445762078310996_467/clk_in scan_wrapper_334445762078310996_468/clk_in
+ scan_wrapper_334445762078310996_467/data_in scan_wrapper_334445762078310996_468/data_in
+ scan_wrapper_334445762078310996_467/latch_enable_in scan_wrapper_334445762078310996_468/latch_enable_in
+ scan_wrapper_334445762078310996_467/scan_select_in scan_wrapper_334445762078310996_468/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_456 scan_wrapper_334445762078310996_456/clk_in scan_wrapper_334445762078310996_457/clk_in
+ scan_wrapper_334445762078310996_456/data_in scan_wrapper_334445762078310996_457/data_in
+ scan_wrapper_334445762078310996_456/latch_enable_in scan_wrapper_334445762078310996_457/latch_enable_in
+ scan_wrapper_334445762078310996_456/scan_select_in scan_wrapper_334445762078310996_457/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_445 scan_wrapper_334445762078310996_445/clk_in scan_wrapper_334445762078310996_446/clk_in
+ scan_wrapper_334445762078310996_445/data_in scan_wrapper_334445762078310996_446/data_in
+ scan_wrapper_334445762078310996_445/latch_enable_in scan_wrapper_334445762078310996_446/latch_enable_in
+ scan_wrapper_334445762078310996_445/scan_select_in scan_wrapper_334445762078310996_446/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_434 scan_wrapper_334445762078310996_434/clk_in scan_wrapper_334445762078310996_435/clk_in
+ scan_wrapper_334445762078310996_434/data_in scan_wrapper_334445762078310996_435/data_in
+ scan_wrapper_334445762078310996_434/latch_enable_in scan_wrapper_334445762078310996_435/latch_enable_in
+ scan_wrapper_334445762078310996_434/scan_select_in scan_wrapper_334445762078310996_435/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_423 scan_wrapper_334445762078310996_423/clk_in scan_wrapper_334445762078310996_424/clk_in
+ scan_wrapper_334445762078310996_423/data_in scan_wrapper_334445762078310996_424/data_in
+ scan_wrapper_334445762078310996_423/latch_enable_in scan_wrapper_334445762078310996_424/latch_enable_in
+ scan_wrapper_334445762078310996_423/scan_select_in scan_wrapper_334445762078310996_424/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_412 scan_wrapper_334445762078310996_412/clk_in scan_wrapper_334445762078310996_413/clk_in
+ scan_wrapper_334445762078310996_412/data_in scan_wrapper_334445762078310996_413/data_in
+ scan_wrapper_334445762078310996_412/latch_enable_in scan_wrapper_334445762078310996_413/latch_enable_in
+ scan_wrapper_334445762078310996_412/scan_select_in scan_wrapper_334445762078310996_413/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_401 scan_wrapper_334445762078310996_401/clk_in scan_wrapper_334445762078310996_402/clk_in
+ scan_wrapper_334445762078310996_401/data_in scan_wrapper_334445762078310996_402/data_in
+ scan_wrapper_334445762078310996_401/latch_enable_in scan_wrapper_334445762078310996_402/latch_enable_in
+ scan_wrapper_334445762078310996_401/scan_select_in scan_wrapper_334445762078310996_402/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_220 scan_wrapper_334445762078310996_220/clk_in scan_wrapper_334445762078310996_221/clk_in
+ scan_wrapper_334445762078310996_220/data_in scan_wrapper_334445762078310996_221/data_in
+ scan_wrapper_334445762078310996_220/latch_enable_in scan_wrapper_334445762078310996_221/latch_enable_in
+ scan_wrapper_334445762078310996_220/scan_select_in scan_wrapper_334445762078310996_221/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_231 scan_wrapper_334445762078310996_231/clk_in scan_wrapper_334445762078310996_232/clk_in
+ scan_wrapper_334445762078310996_231/data_in scan_wrapper_334445762078310996_232/data_in
+ scan_wrapper_334445762078310996_231/latch_enable_in scan_wrapper_334445762078310996_232/latch_enable_in
+ scan_wrapper_334445762078310996_231/scan_select_in scan_wrapper_334445762078310996_232/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_242 scan_wrapper_334445762078310996_242/clk_in scan_wrapper_334445762078310996_243/clk_in
+ scan_wrapper_334445762078310996_242/data_in scan_wrapper_334445762078310996_243/data_in
+ scan_wrapper_334445762078310996_242/latch_enable_in scan_wrapper_334445762078310996_243/latch_enable_in
+ scan_wrapper_334445762078310996_242/scan_select_in scan_wrapper_334445762078310996_243/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_253 scan_wrapper_334445762078310996_253/clk_in scan_wrapper_334445762078310996_254/clk_in
+ scan_wrapper_334445762078310996_253/data_in scan_wrapper_334445762078310996_254/data_in
+ scan_wrapper_334445762078310996_253/latch_enable_in scan_wrapper_334445762078310996_254/latch_enable_in
+ scan_wrapper_334445762078310996_253/scan_select_in scan_wrapper_334445762078310996_254/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_264 scan_wrapper_334445762078310996_264/clk_in scan_wrapper_334445762078310996_265/clk_in
+ scan_wrapper_334445762078310996_264/data_in scan_wrapper_334445762078310996_265/data_in
+ scan_wrapper_334445762078310996_264/latch_enable_in scan_wrapper_334445762078310996_265/latch_enable_in
+ scan_wrapper_334445762078310996_264/scan_select_in scan_wrapper_334445762078310996_265/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_275 scan_wrapper_334445762078310996_275/clk_in scan_wrapper_334445762078310996_276/clk_in
+ scan_wrapper_334445762078310996_275/data_in scan_wrapper_334445762078310996_276/data_in
+ scan_wrapper_334445762078310996_275/latch_enable_in scan_wrapper_334445762078310996_276/latch_enable_in
+ scan_wrapper_334445762078310996_275/scan_select_in scan_wrapper_334445762078310996_276/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_286 scan_wrapper_334445762078310996_286/clk_in scan_wrapper_334445762078310996_287/clk_in
+ scan_wrapper_334445762078310996_286/data_in scan_wrapper_334445762078310996_287/data_in
+ scan_wrapper_334445762078310996_286/latch_enable_in scan_wrapper_334445762078310996_287/latch_enable_in
+ scan_wrapper_334445762078310996_286/scan_select_in scan_wrapper_334445762078310996_287/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_297 scan_wrapper_334445762078310996_297/clk_in scan_wrapper_334445762078310996_298/clk_in
+ scan_wrapper_334445762078310996_297/data_in scan_wrapper_334445762078310996_298/data_in
+ scan_wrapper_334445762078310996_297/latch_enable_in scan_wrapper_334445762078310996_298/latch_enable_in
+ scan_wrapper_334445762078310996_297/scan_select_in scan_wrapper_334445762078310996_298/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_3 scan_wrapper_334445762078310996_3/clk_in scan_wrapper_334445762078310996_4/clk_in
+ scan_wrapper_334445762078310996_3/data_in scan_wrapper_334445762078310996_4/data_in
+ scan_wrapper_334445762078310996_3/latch_enable_in scan_wrapper_334445762078310996_4/latch_enable_in
+ scan_wrapper_334445762078310996_3/scan_select_in scan_wrapper_334445762078310996_4/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_479 scan_wrapper_334445762078310996_479/clk_in scan_wrapper_334445762078310996_480/clk_in
+ scan_wrapper_334445762078310996_479/data_in scan_wrapper_334445762078310996_480/data_in
+ scan_wrapper_334445762078310996_479/latch_enable_in scan_wrapper_334445762078310996_480/latch_enable_in
+ scan_wrapper_334445762078310996_479/scan_select_in scan_wrapper_334445762078310996_480/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_468 scan_wrapper_334445762078310996_468/clk_in scan_wrapper_334445762078310996_469/clk_in
+ scan_wrapper_334445762078310996_468/data_in scan_wrapper_334445762078310996_469/data_in
+ scan_wrapper_334445762078310996_468/latch_enable_in scan_wrapper_334445762078310996_469/latch_enable_in
+ scan_wrapper_334445762078310996_468/scan_select_in scan_wrapper_334445762078310996_469/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_457 scan_wrapper_334445762078310996_457/clk_in scan_wrapper_334445762078310996_458/clk_in
+ scan_wrapper_334445762078310996_457/data_in scan_wrapper_334445762078310996_458/data_in
+ scan_wrapper_334445762078310996_457/latch_enable_in scan_wrapper_334445762078310996_458/latch_enable_in
+ scan_wrapper_334445762078310996_457/scan_select_in scan_wrapper_334445762078310996_458/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_446 scan_wrapper_334445762078310996_446/clk_in scan_wrapper_334445762078310996_447/clk_in
+ scan_wrapper_334445762078310996_446/data_in scan_wrapper_334445762078310996_447/data_in
+ scan_wrapper_334445762078310996_446/latch_enable_in scan_wrapper_334445762078310996_447/latch_enable_in
+ scan_wrapper_334445762078310996_446/scan_select_in scan_wrapper_334445762078310996_447/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_435 scan_wrapper_334445762078310996_435/clk_in scan_wrapper_334445762078310996_436/clk_in
+ scan_wrapper_334445762078310996_435/data_in scan_wrapper_334445762078310996_436/data_in
+ scan_wrapper_334445762078310996_435/latch_enable_in scan_wrapper_334445762078310996_436/latch_enable_in
+ scan_wrapper_334445762078310996_435/scan_select_in scan_wrapper_334445762078310996_436/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_424 scan_wrapper_334445762078310996_424/clk_in scan_wrapper_334445762078310996_425/clk_in
+ scan_wrapper_334445762078310996_424/data_in scan_wrapper_334445762078310996_425/data_in
+ scan_wrapper_334445762078310996_424/latch_enable_in scan_wrapper_334445762078310996_425/latch_enable_in
+ scan_wrapper_334445762078310996_424/scan_select_in scan_wrapper_334445762078310996_425/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_413 scan_wrapper_334445762078310996_413/clk_in scan_wrapper_334445762078310996_414/clk_in
+ scan_wrapper_334445762078310996_413/data_in scan_wrapper_334445762078310996_414/data_in
+ scan_wrapper_334445762078310996_413/latch_enable_in scan_wrapper_334445762078310996_414/latch_enable_in
+ scan_wrapper_334445762078310996_413/scan_select_in scan_wrapper_334445762078310996_414/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_402 scan_wrapper_334445762078310996_402/clk_in scan_wrapper_334445762078310996_403/clk_in
+ scan_wrapper_334445762078310996_402/data_in scan_wrapper_334445762078310996_403/data_in
+ scan_wrapper_334445762078310996_402/latch_enable_in scan_wrapper_334445762078310996_403/latch_enable_in
+ scan_wrapper_334445762078310996_402/scan_select_in scan_wrapper_334445762078310996_403/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_210 scan_wrapper_334445762078310996_210/clk_in scan_wrapper_334445762078310996_211/clk_in
+ scan_wrapper_334445762078310996_210/data_in scan_wrapper_334445762078310996_211/data_in
+ scan_wrapper_334445762078310996_210/latch_enable_in scan_wrapper_334445762078310996_211/latch_enable_in
+ scan_wrapper_334445762078310996_210/scan_select_in scan_wrapper_334445762078310996_211/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_221 scan_wrapper_334445762078310996_221/clk_in scan_wrapper_334445762078310996_222/clk_in
+ scan_wrapper_334445762078310996_221/data_in scan_wrapper_334445762078310996_222/data_in
+ scan_wrapper_334445762078310996_221/latch_enable_in scan_wrapper_334445762078310996_222/latch_enable_in
+ scan_wrapper_334445762078310996_221/scan_select_in scan_wrapper_334445762078310996_222/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_232 scan_wrapper_334445762078310996_232/clk_in scan_wrapper_334445762078310996_233/clk_in
+ scan_wrapper_334445762078310996_232/data_in scan_wrapper_334445762078310996_233/data_in
+ scan_wrapper_334445762078310996_232/latch_enable_in scan_wrapper_334445762078310996_233/latch_enable_in
+ scan_wrapper_334445762078310996_232/scan_select_in scan_wrapper_334445762078310996_233/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_243 scan_wrapper_334445762078310996_243/clk_in scan_wrapper_334445762078310996_244/clk_in
+ scan_wrapper_334445762078310996_243/data_in scan_wrapper_334445762078310996_244/data_in
+ scan_wrapper_334445762078310996_243/latch_enable_in scan_wrapper_334445762078310996_244/latch_enable_in
+ scan_wrapper_334445762078310996_243/scan_select_in scan_wrapper_334445762078310996_244/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_254 scan_wrapper_334445762078310996_254/clk_in scan_wrapper_334445762078310996_255/clk_in
+ scan_wrapper_334445762078310996_254/data_in scan_wrapper_334445762078310996_255/data_in
+ scan_wrapper_334445762078310996_254/latch_enable_in scan_wrapper_334445762078310996_255/latch_enable_in
+ scan_wrapper_334445762078310996_254/scan_select_in scan_wrapper_334445762078310996_255/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_265 scan_wrapper_334445762078310996_265/clk_in scan_wrapper_334445762078310996_266/clk_in
+ scan_wrapper_334445762078310996_265/data_in scan_wrapper_334445762078310996_266/data_in
+ scan_wrapper_334445762078310996_265/latch_enable_in scan_wrapper_334445762078310996_266/latch_enable_in
+ scan_wrapper_334445762078310996_265/scan_select_in scan_wrapper_334445762078310996_266/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_276 scan_wrapper_334445762078310996_276/clk_in scan_wrapper_334445762078310996_277/clk_in
+ scan_wrapper_334445762078310996_276/data_in scan_wrapper_334445762078310996_277/data_in
+ scan_wrapper_334445762078310996_276/latch_enable_in scan_wrapper_334445762078310996_277/latch_enable_in
+ scan_wrapper_334445762078310996_276/scan_select_in scan_wrapper_334445762078310996_277/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_287 scan_wrapper_334445762078310996_287/clk_in scan_wrapper_334445762078310996_288/clk_in
+ scan_wrapper_334445762078310996_287/data_in scan_wrapper_334445762078310996_288/data_in
+ scan_wrapper_334445762078310996_287/latch_enable_in scan_wrapper_334445762078310996_288/latch_enable_in
+ scan_wrapper_334445762078310996_287/scan_select_in scan_wrapper_334445762078310996_288/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_298 scan_wrapper_334445762078310996_298/clk_in scan_wrapper_334445762078310996_299/clk_in
+ scan_wrapper_334445762078310996_298/data_in scan_wrapper_334445762078310996_299/data_in
+ scan_wrapper_334445762078310996_298/latch_enable_in scan_wrapper_334445762078310996_299/latch_enable_in
+ scan_wrapper_334445762078310996_298/scan_select_in scan_wrapper_334445762078310996_299/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_335404063203000914_1 scan_wrapper_335404063203000914_1/clk_in scan_wrapper_334445762078310996_2/clk_in
+ scan_wrapper_335404063203000914_1/data_in scan_wrapper_334445762078310996_2/data_in
+ scan_wrapper_335404063203000914_1/latch_enable_in scan_wrapper_334445762078310996_2/latch_enable_in
+ scan_wrapper_335404063203000914_1/scan_select_in scan_wrapper_334445762078310996_2/scan_select_in
+ vccd1 vssd1 scan_wrapper_335404063203000914
Xscan_wrapper_334445762078310996_4 scan_wrapper_334445762078310996_4/clk_in scan_wrapper_334445762078310996_5/clk_in
+ scan_wrapper_334445762078310996_4/data_in scan_wrapper_334445762078310996_5/data_in
+ scan_wrapper_334445762078310996_4/latch_enable_in scan_wrapper_334445762078310996_5/latch_enable_in
+ scan_wrapper_334445762078310996_4/scan_select_in scan_wrapper_334445762078310996_5/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_469 scan_wrapper_334445762078310996_469/clk_in scan_wrapper_334445762078310996_470/clk_in
+ scan_wrapper_334445762078310996_469/data_in scan_wrapper_334445762078310996_470/data_in
+ scan_wrapper_334445762078310996_469/latch_enable_in scan_wrapper_334445762078310996_470/latch_enable_in
+ scan_wrapper_334445762078310996_469/scan_select_in scan_wrapper_334445762078310996_470/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_458 scan_wrapper_334445762078310996_458/clk_in scan_wrapper_334445762078310996_459/clk_in
+ scan_wrapper_334445762078310996_458/data_in scan_wrapper_334445762078310996_459/data_in
+ scan_wrapper_334445762078310996_458/latch_enable_in scan_wrapper_334445762078310996_459/latch_enable_in
+ scan_wrapper_334445762078310996_458/scan_select_in scan_wrapper_334445762078310996_459/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_447 scan_wrapper_334445762078310996_447/clk_in scan_wrapper_334445762078310996_448/clk_in
+ scan_wrapper_334445762078310996_447/data_in scan_wrapper_334445762078310996_448/data_in
+ scan_wrapper_334445762078310996_447/latch_enable_in scan_wrapper_334445762078310996_448/latch_enable_in
+ scan_wrapper_334445762078310996_447/scan_select_in scan_wrapper_334445762078310996_448/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_436 scan_wrapper_334445762078310996_436/clk_in scan_wrapper_334445762078310996_437/clk_in
+ scan_wrapper_334445762078310996_436/data_in scan_wrapper_334445762078310996_437/data_in
+ scan_wrapper_334445762078310996_436/latch_enable_in scan_wrapper_334445762078310996_437/latch_enable_in
+ scan_wrapper_334445762078310996_436/scan_select_in scan_wrapper_334445762078310996_437/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_425 scan_wrapper_334445762078310996_425/clk_in scan_wrapper_334445762078310996_426/clk_in
+ scan_wrapper_334445762078310996_425/data_in scan_wrapper_334445762078310996_426/data_in
+ scan_wrapper_334445762078310996_425/latch_enable_in scan_wrapper_334445762078310996_426/latch_enable_in
+ scan_wrapper_334445762078310996_425/scan_select_in scan_wrapper_334445762078310996_426/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_414 scan_wrapper_334445762078310996_414/clk_in scan_wrapper_334445762078310996_415/clk_in
+ scan_wrapper_334445762078310996_414/data_in scan_wrapper_334445762078310996_415/data_in
+ scan_wrapper_334445762078310996_414/latch_enable_in scan_wrapper_334445762078310996_415/latch_enable_in
+ scan_wrapper_334445762078310996_414/scan_select_in scan_wrapper_334445762078310996_415/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_403 scan_wrapper_334445762078310996_403/clk_in scan_wrapper_334445762078310996_404/clk_in
+ scan_wrapper_334445762078310996_403/data_in scan_wrapper_334445762078310996_404/data_in
+ scan_wrapper_334445762078310996_403/latch_enable_in scan_wrapper_334445762078310996_404/latch_enable_in
+ scan_wrapper_334445762078310996_403/scan_select_in scan_wrapper_334445762078310996_404/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_200 scan_wrapper_334445762078310996_200/clk_in scan_wrapper_334445762078310996_201/clk_in
+ scan_wrapper_334445762078310996_200/data_in scan_wrapper_334445762078310996_201/data_in
+ scan_wrapper_334445762078310996_200/latch_enable_in scan_wrapper_334445762078310996_201/latch_enable_in
+ scan_wrapper_334445762078310996_200/scan_select_in scan_wrapper_334445762078310996_201/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_211 scan_wrapper_334445762078310996_211/clk_in scan_wrapper_334445762078310996_212/clk_in
+ scan_wrapper_334445762078310996_211/data_in scan_wrapper_334445762078310996_212/data_in
+ scan_wrapper_334445762078310996_211/latch_enable_in scan_wrapper_334445762078310996_212/latch_enable_in
+ scan_wrapper_334445762078310996_211/scan_select_in scan_wrapper_334445762078310996_212/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_222 scan_wrapper_334445762078310996_222/clk_in scan_wrapper_334445762078310996_223/clk_in
+ scan_wrapper_334445762078310996_222/data_in scan_wrapper_334445762078310996_223/data_in
+ scan_wrapper_334445762078310996_222/latch_enable_in scan_wrapper_334445762078310996_223/latch_enable_in
+ scan_wrapper_334445762078310996_222/scan_select_in scan_wrapper_334445762078310996_223/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_233 scan_wrapper_334445762078310996_233/clk_in scan_wrapper_334445762078310996_234/clk_in
+ scan_wrapper_334445762078310996_233/data_in scan_wrapper_334445762078310996_234/data_in
+ scan_wrapper_334445762078310996_233/latch_enable_in scan_wrapper_334445762078310996_234/latch_enable_in
+ scan_wrapper_334445762078310996_233/scan_select_in scan_wrapper_334445762078310996_234/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_244 scan_wrapper_334445762078310996_244/clk_in scan_wrapper_334445762078310996_245/clk_in
+ scan_wrapper_334445762078310996_244/data_in scan_wrapper_334445762078310996_245/data_in
+ scan_wrapper_334445762078310996_244/latch_enable_in scan_wrapper_334445762078310996_245/latch_enable_in
+ scan_wrapper_334445762078310996_244/scan_select_in scan_wrapper_334445762078310996_245/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_255 scan_wrapper_334445762078310996_255/clk_in scan_wrapper_334445762078310996_256/clk_in
+ scan_wrapper_334445762078310996_255/data_in scan_wrapper_334445762078310996_256/data_in
+ scan_wrapper_334445762078310996_255/latch_enable_in scan_wrapper_334445762078310996_256/latch_enable_in
+ scan_wrapper_334445762078310996_255/scan_select_in scan_wrapper_334445762078310996_256/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_266 scan_wrapper_334445762078310996_266/clk_in scan_wrapper_334445762078310996_267/clk_in
+ scan_wrapper_334445762078310996_266/data_in scan_wrapper_334445762078310996_267/data_in
+ scan_wrapper_334445762078310996_266/latch_enable_in scan_wrapper_334445762078310996_267/latch_enable_in
+ scan_wrapper_334445762078310996_266/scan_select_in scan_wrapper_334445762078310996_267/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_277 scan_wrapper_334445762078310996_277/clk_in scan_wrapper_334445762078310996_278/clk_in
+ scan_wrapper_334445762078310996_277/data_in scan_wrapper_334445762078310996_278/data_in
+ scan_wrapper_334445762078310996_277/latch_enable_in scan_wrapper_334445762078310996_278/latch_enable_in
+ scan_wrapper_334445762078310996_277/scan_select_in scan_wrapper_334445762078310996_278/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_288 scan_wrapper_334445762078310996_288/clk_in scan_wrapper_334445762078310996_289/clk_in
+ scan_wrapper_334445762078310996_288/data_in scan_wrapper_334445762078310996_289/data_in
+ scan_wrapper_334445762078310996_288/latch_enable_in scan_wrapper_334445762078310996_289/latch_enable_in
+ scan_wrapper_334445762078310996_288/scan_select_in scan_wrapper_334445762078310996_289/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_299 scan_wrapper_334445762078310996_299/clk_in scan_wrapper_334445762078310996_300/clk_in
+ scan_wrapper_334445762078310996_299/data_in scan_wrapper_334445762078310996_300/data_in
+ scan_wrapper_334445762078310996_299/latch_enable_in scan_wrapper_334445762078310996_300/latch_enable_in
+ scan_wrapper_334445762078310996_299/scan_select_in scan_wrapper_334445762078310996_300/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_5 scan_wrapper_334445762078310996_5/clk_in scan_wrapper_334445762078310996_6/clk_in
+ scan_wrapper_334445762078310996_5/data_in scan_wrapper_334445762078310996_6/data_in
+ scan_wrapper_334445762078310996_5/latch_enable_in scan_wrapper_334445762078310996_6/latch_enable_in
+ scan_wrapper_334445762078310996_5/scan_select_in scan_wrapper_334445762078310996_6/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_448 scan_wrapper_334445762078310996_448/clk_in scan_wrapper_334445762078310996_449/clk_in
+ scan_wrapper_334445762078310996_448/data_in scan_wrapper_334445762078310996_449/data_in
+ scan_wrapper_334445762078310996_448/latch_enable_in scan_wrapper_334445762078310996_449/latch_enable_in
+ scan_wrapper_334445762078310996_448/scan_select_in scan_wrapper_334445762078310996_449/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_437 scan_wrapper_334445762078310996_437/clk_in scan_wrapper_334445762078310996_438/clk_in
+ scan_wrapper_334445762078310996_437/data_in scan_wrapper_334445762078310996_438/data_in
+ scan_wrapper_334445762078310996_437/latch_enable_in scan_wrapper_334445762078310996_438/latch_enable_in
+ scan_wrapper_334445762078310996_437/scan_select_in scan_wrapper_334445762078310996_438/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_426 scan_wrapper_334445762078310996_426/clk_in scan_wrapper_334445762078310996_427/clk_in
+ scan_wrapper_334445762078310996_426/data_in scan_wrapper_334445762078310996_427/data_in
+ scan_wrapper_334445762078310996_426/latch_enable_in scan_wrapper_334445762078310996_427/latch_enable_in
+ scan_wrapper_334445762078310996_426/scan_select_in scan_wrapper_334445762078310996_427/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_415 scan_wrapper_334445762078310996_415/clk_in scan_wrapper_334445762078310996_416/clk_in
+ scan_wrapper_334445762078310996_415/data_in scan_wrapper_334445762078310996_416/data_in
+ scan_wrapper_334445762078310996_415/latch_enable_in scan_wrapper_334445762078310996_416/latch_enable_in
+ scan_wrapper_334445762078310996_415/scan_select_in scan_wrapper_334445762078310996_416/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_404 scan_wrapper_334445762078310996_404/clk_in scan_wrapper_334445762078310996_405/clk_in
+ scan_wrapper_334445762078310996_404/data_in scan_wrapper_334445762078310996_405/data_in
+ scan_wrapper_334445762078310996_404/latch_enable_in scan_wrapper_334445762078310996_405/latch_enable_in
+ scan_wrapper_334445762078310996_404/scan_select_in scan_wrapper_334445762078310996_405/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_459 scan_wrapper_334445762078310996_459/clk_in scan_wrapper_334445762078310996_460/clk_in
+ scan_wrapper_334445762078310996_459/data_in scan_wrapper_334445762078310996_460/data_in
+ scan_wrapper_334445762078310996_459/latch_enable_in scan_wrapper_334445762078310996_460/latch_enable_in
+ scan_wrapper_334445762078310996_459/scan_select_in scan_wrapper_334445762078310996_460/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_201 scan_wrapper_334445762078310996_201/clk_in scan_wrapper_334445762078310996_202/clk_in
+ scan_wrapper_334445762078310996_201/data_in scan_wrapper_334445762078310996_202/data_in
+ scan_wrapper_334445762078310996_201/latch_enable_in scan_wrapper_334445762078310996_202/latch_enable_in
+ scan_wrapper_334445762078310996_201/scan_select_in scan_wrapper_334445762078310996_202/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_212 scan_wrapper_334445762078310996_212/clk_in scan_wrapper_334445762078310996_213/clk_in
+ scan_wrapper_334445762078310996_212/data_in scan_wrapper_334445762078310996_213/data_in
+ scan_wrapper_334445762078310996_212/latch_enable_in scan_wrapper_334445762078310996_213/latch_enable_in
+ scan_wrapper_334445762078310996_212/scan_select_in scan_wrapper_334445762078310996_213/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_223 scan_wrapper_334445762078310996_223/clk_in scan_wrapper_334445762078310996_224/clk_in
+ scan_wrapper_334445762078310996_223/data_in scan_wrapper_334445762078310996_224/data_in
+ scan_wrapper_334445762078310996_223/latch_enable_in scan_wrapper_334445762078310996_224/latch_enable_in
+ scan_wrapper_334445762078310996_223/scan_select_in scan_wrapper_334445762078310996_224/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_234 scan_wrapper_334445762078310996_234/clk_in scan_wrapper_334445762078310996_235/clk_in
+ scan_wrapper_334445762078310996_234/data_in scan_wrapper_334445762078310996_235/data_in
+ scan_wrapper_334445762078310996_234/latch_enable_in scan_wrapper_334445762078310996_235/latch_enable_in
+ scan_wrapper_334445762078310996_234/scan_select_in scan_wrapper_334445762078310996_235/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_245 scan_wrapper_334445762078310996_245/clk_in scan_wrapper_334445762078310996_246/clk_in
+ scan_wrapper_334445762078310996_245/data_in scan_wrapper_334445762078310996_246/data_in
+ scan_wrapper_334445762078310996_245/latch_enable_in scan_wrapper_334445762078310996_246/latch_enable_in
+ scan_wrapper_334445762078310996_245/scan_select_in scan_wrapper_334445762078310996_246/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_256 scan_wrapper_334445762078310996_256/clk_in scan_wrapper_334445762078310996_257/clk_in
+ scan_wrapper_334445762078310996_256/data_in scan_wrapper_334445762078310996_257/data_in
+ scan_wrapper_334445762078310996_256/latch_enable_in scan_wrapper_334445762078310996_257/latch_enable_in
+ scan_wrapper_334445762078310996_256/scan_select_in scan_wrapper_334445762078310996_257/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_267 scan_wrapper_334445762078310996_267/clk_in scan_wrapper_334445762078310996_268/clk_in
+ scan_wrapper_334445762078310996_267/data_in scan_wrapper_334445762078310996_268/data_in
+ scan_wrapper_334445762078310996_267/latch_enable_in scan_wrapper_334445762078310996_268/latch_enable_in
+ scan_wrapper_334445762078310996_267/scan_select_in scan_wrapper_334445762078310996_268/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_278 scan_wrapper_334445762078310996_278/clk_in scan_wrapper_334445762078310996_279/clk_in
+ scan_wrapper_334445762078310996_278/data_in scan_wrapper_334445762078310996_279/data_in
+ scan_wrapper_334445762078310996_278/latch_enable_in scan_wrapper_334445762078310996_279/latch_enable_in
+ scan_wrapper_334445762078310996_278/scan_select_in scan_wrapper_334445762078310996_279/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_289 scan_wrapper_334445762078310996_289/clk_in scan_wrapper_334445762078310996_290/clk_in
+ scan_wrapper_334445762078310996_289/data_in scan_wrapper_334445762078310996_290/data_in
+ scan_wrapper_334445762078310996_289/latch_enable_in scan_wrapper_334445762078310996_290/latch_enable_in
+ scan_wrapper_334445762078310996_289/scan_select_in scan_wrapper_334445762078310996_290/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_6 scan_wrapper_334445762078310996_6/clk_in scan_wrapper_334445762078310996_7/clk_in
+ scan_wrapper_334445762078310996_6/data_in scan_wrapper_334445762078310996_7/data_in
+ scan_wrapper_334445762078310996_6/latch_enable_in scan_wrapper_334445762078310996_7/latch_enable_in
+ scan_wrapper_334445762078310996_6/scan_select_in scan_wrapper_334445762078310996_7/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_449 scan_wrapper_334445762078310996_449/clk_in scan_wrapper_334445762078310996_450/clk_in
+ scan_wrapper_334445762078310996_449/data_in scan_wrapper_334445762078310996_450/data_in
+ scan_wrapper_334445762078310996_449/latch_enable_in scan_wrapper_334445762078310996_450/latch_enable_in
+ scan_wrapper_334445762078310996_449/scan_select_in scan_wrapper_334445762078310996_450/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_438 scan_wrapper_334445762078310996_438/clk_in scan_wrapper_334445762078310996_439/clk_in
+ scan_wrapper_334445762078310996_438/data_in scan_wrapper_334445762078310996_439/data_in
+ scan_wrapper_334445762078310996_438/latch_enable_in scan_wrapper_334445762078310996_439/latch_enable_in
+ scan_wrapper_334445762078310996_438/scan_select_in scan_wrapper_334445762078310996_439/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_427 scan_wrapper_334445762078310996_427/clk_in scan_wrapper_334445762078310996_428/clk_in
+ scan_wrapper_334445762078310996_427/data_in scan_wrapper_334445762078310996_428/data_in
+ scan_wrapper_334445762078310996_427/latch_enable_in scan_wrapper_334445762078310996_428/latch_enable_in
+ scan_wrapper_334445762078310996_427/scan_select_in scan_wrapper_334445762078310996_428/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_416 scan_wrapper_334445762078310996_416/clk_in scan_wrapper_334445762078310996_417/clk_in
+ scan_wrapper_334445762078310996_416/data_in scan_wrapper_334445762078310996_417/data_in
+ scan_wrapper_334445762078310996_416/latch_enable_in scan_wrapper_334445762078310996_417/latch_enable_in
+ scan_wrapper_334445762078310996_416/scan_select_in scan_wrapper_334445762078310996_417/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_405 scan_wrapper_334445762078310996_405/clk_in scan_wrapper_334445762078310996_406/clk_in
+ scan_wrapper_334445762078310996_405/data_in scan_wrapper_334445762078310996_406/data_in
+ scan_wrapper_334445762078310996_405/latch_enable_in scan_wrapper_334445762078310996_406/latch_enable_in
+ scan_wrapper_334445762078310996_405/scan_select_in scan_wrapper_334445762078310996_406/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_202 scan_wrapper_334445762078310996_202/clk_in scan_wrapper_334445762078310996_203/clk_in
+ scan_wrapper_334445762078310996_202/data_in scan_wrapper_334445762078310996_203/data_in
+ scan_wrapper_334445762078310996_202/latch_enable_in scan_wrapper_334445762078310996_203/latch_enable_in
+ scan_wrapper_334445762078310996_202/scan_select_in scan_wrapper_334445762078310996_203/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_213 scan_wrapper_334445762078310996_213/clk_in scan_wrapper_334445762078310996_214/clk_in
+ scan_wrapper_334445762078310996_213/data_in scan_wrapper_334445762078310996_214/data_in
+ scan_wrapper_334445762078310996_213/latch_enable_in scan_wrapper_334445762078310996_214/latch_enable_in
+ scan_wrapper_334445762078310996_213/scan_select_in scan_wrapper_334445762078310996_214/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_224 scan_wrapper_334445762078310996_224/clk_in scan_wrapper_334445762078310996_225/clk_in
+ scan_wrapper_334445762078310996_224/data_in scan_wrapper_334445762078310996_225/data_in
+ scan_wrapper_334445762078310996_224/latch_enable_in scan_wrapper_334445762078310996_225/latch_enable_in
+ scan_wrapper_334445762078310996_224/scan_select_in scan_wrapper_334445762078310996_225/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_235 scan_wrapper_334445762078310996_235/clk_in scan_wrapper_334445762078310996_236/clk_in
+ scan_wrapper_334445762078310996_235/data_in scan_wrapper_334445762078310996_236/data_in
+ scan_wrapper_334445762078310996_235/latch_enable_in scan_wrapper_334445762078310996_236/latch_enable_in
+ scan_wrapper_334445762078310996_235/scan_select_in scan_wrapper_334445762078310996_236/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_246 scan_wrapper_334445762078310996_246/clk_in scan_wrapper_334445762078310996_247/clk_in
+ scan_wrapper_334445762078310996_246/data_in scan_wrapper_334445762078310996_247/data_in
+ scan_wrapper_334445762078310996_246/latch_enable_in scan_wrapper_334445762078310996_247/latch_enable_in
+ scan_wrapper_334445762078310996_246/scan_select_in scan_wrapper_334445762078310996_247/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_257 scan_wrapper_334445762078310996_257/clk_in scan_wrapper_334445762078310996_258/clk_in
+ scan_wrapper_334445762078310996_257/data_in scan_wrapper_334445762078310996_258/data_in
+ scan_wrapper_334445762078310996_257/latch_enable_in scan_wrapper_334445762078310996_258/latch_enable_in
+ scan_wrapper_334445762078310996_257/scan_select_in scan_wrapper_334445762078310996_258/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_268 scan_wrapper_334445762078310996_268/clk_in scan_wrapper_334445762078310996_269/clk_in
+ scan_wrapper_334445762078310996_268/data_in scan_wrapper_334445762078310996_269/data_in
+ scan_wrapper_334445762078310996_268/latch_enable_in scan_wrapper_334445762078310996_269/latch_enable_in
+ scan_wrapper_334445762078310996_268/scan_select_in scan_wrapper_334445762078310996_269/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_279 scan_wrapper_334445762078310996_279/clk_in scan_wrapper_334445762078310996_280/clk_in
+ scan_wrapper_334445762078310996_279/data_in scan_wrapper_334445762078310996_280/data_in
+ scan_wrapper_334445762078310996_279/latch_enable_in scan_wrapper_334445762078310996_280/latch_enable_in
+ scan_wrapper_334445762078310996_279/scan_select_in scan_wrapper_334445762078310996_280/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_7 scan_wrapper_334445762078310996_7/clk_in scan_wrapper_334445762078310996_8/clk_in
+ scan_wrapper_334445762078310996_7/data_in scan_wrapper_334445762078310996_8/data_in
+ scan_wrapper_334445762078310996_7/latch_enable_in scan_wrapper_334445762078310996_8/latch_enable_in
+ scan_wrapper_334445762078310996_7/scan_select_in scan_wrapper_334445762078310996_8/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_439 scan_wrapper_334445762078310996_439/clk_in scan_wrapper_334445762078310996_440/clk_in
+ scan_wrapper_334445762078310996_439/data_in scan_wrapper_334445762078310996_440/data_in
+ scan_wrapper_334445762078310996_439/latch_enable_in scan_wrapper_334445762078310996_440/latch_enable_in
+ scan_wrapper_334445762078310996_439/scan_select_in scan_wrapper_334445762078310996_440/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_428 scan_wrapper_334445762078310996_428/clk_in scan_wrapper_334445762078310996_429/clk_in
+ scan_wrapper_334445762078310996_428/data_in scan_wrapper_334445762078310996_429/data_in
+ scan_wrapper_334445762078310996_428/latch_enable_in scan_wrapper_334445762078310996_429/latch_enable_in
+ scan_wrapper_334445762078310996_428/scan_select_in scan_wrapper_334445762078310996_429/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_417 scan_wrapper_334445762078310996_417/clk_in scan_wrapper_334445762078310996_418/clk_in
+ scan_wrapper_334445762078310996_417/data_in scan_wrapper_334445762078310996_418/data_in
+ scan_wrapper_334445762078310996_417/latch_enable_in scan_wrapper_334445762078310996_418/latch_enable_in
+ scan_wrapper_334445762078310996_417/scan_select_in scan_wrapper_334445762078310996_418/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_406 scan_wrapper_334445762078310996_406/clk_in scan_wrapper_334445762078310996_407/clk_in
+ scan_wrapper_334445762078310996_406/data_in scan_wrapper_334445762078310996_407/data_in
+ scan_wrapper_334445762078310996_406/latch_enable_in scan_wrapper_334445762078310996_407/latch_enable_in
+ scan_wrapper_334445762078310996_406/scan_select_in scan_wrapper_334445762078310996_407/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_203 scan_wrapper_334445762078310996_203/clk_in scan_wrapper_334445762078310996_204/clk_in
+ scan_wrapper_334445762078310996_203/data_in scan_wrapper_334445762078310996_204/data_in
+ scan_wrapper_334445762078310996_203/latch_enable_in scan_wrapper_334445762078310996_204/latch_enable_in
+ scan_wrapper_334445762078310996_203/scan_select_in scan_wrapper_334445762078310996_204/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_214 scan_wrapper_334445762078310996_214/clk_in scan_wrapper_334445762078310996_215/clk_in
+ scan_wrapper_334445762078310996_214/data_in scan_wrapper_334445762078310996_215/data_in
+ scan_wrapper_334445762078310996_214/latch_enable_in scan_wrapper_334445762078310996_215/latch_enable_in
+ scan_wrapper_334445762078310996_214/scan_select_in scan_wrapper_334445762078310996_215/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_225 scan_wrapper_334445762078310996_225/clk_in scan_wrapper_334445762078310996_226/clk_in
+ scan_wrapper_334445762078310996_225/data_in scan_wrapper_334445762078310996_226/data_in
+ scan_wrapper_334445762078310996_225/latch_enable_in scan_wrapper_334445762078310996_226/latch_enable_in
+ scan_wrapper_334445762078310996_225/scan_select_in scan_wrapper_334445762078310996_226/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_236 scan_wrapper_334445762078310996_236/clk_in scan_wrapper_334445762078310996_237/clk_in
+ scan_wrapper_334445762078310996_236/data_in scan_wrapper_334445762078310996_237/data_in
+ scan_wrapper_334445762078310996_236/latch_enable_in scan_wrapper_334445762078310996_237/latch_enable_in
+ scan_wrapper_334445762078310996_236/scan_select_in scan_wrapper_334445762078310996_237/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_247 scan_wrapper_334445762078310996_247/clk_in scan_wrapper_334445762078310996_248/clk_in
+ scan_wrapper_334445762078310996_247/data_in scan_wrapper_334445762078310996_248/data_in
+ scan_wrapper_334445762078310996_247/latch_enable_in scan_wrapper_334445762078310996_248/latch_enable_in
+ scan_wrapper_334445762078310996_247/scan_select_in scan_wrapper_334445762078310996_248/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_258 scan_wrapper_334445762078310996_258/clk_in scan_wrapper_334445762078310996_259/clk_in
+ scan_wrapper_334445762078310996_258/data_in scan_wrapper_334445762078310996_259/data_in
+ scan_wrapper_334445762078310996_258/latch_enable_in scan_wrapper_334445762078310996_259/latch_enable_in
+ scan_wrapper_334445762078310996_258/scan_select_in scan_wrapper_334445762078310996_259/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_269 scan_wrapper_334445762078310996_269/clk_in scan_wrapper_334445762078310996_270/clk_in
+ scan_wrapper_334445762078310996_269/data_in scan_wrapper_334445762078310996_270/data_in
+ scan_wrapper_334445762078310996_269/latch_enable_in scan_wrapper_334445762078310996_270/latch_enable_in
+ scan_wrapper_334445762078310996_269/scan_select_in scan_wrapper_334445762078310996_270/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_8 scan_wrapper_334445762078310996_8/clk_in scan_wrapper_334445762078310996_9/clk_in
+ scan_wrapper_334445762078310996_8/data_in scan_wrapper_334445762078310996_9/data_in
+ scan_wrapper_334445762078310996_8/latch_enable_in scan_wrapper_334445762078310996_9/latch_enable_in
+ scan_wrapper_334445762078310996_8/scan_select_in scan_wrapper_334445762078310996_9/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_429 scan_wrapper_334445762078310996_429/clk_in scan_wrapper_334445762078310996_430/clk_in
+ scan_wrapper_334445762078310996_429/data_in scan_wrapper_334445762078310996_430/data_in
+ scan_wrapper_334445762078310996_429/latch_enable_in scan_wrapper_334445762078310996_430/latch_enable_in
+ scan_wrapper_334445762078310996_429/scan_select_in scan_wrapper_334445762078310996_430/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_418 scan_wrapper_334445762078310996_418/clk_in scan_wrapper_334445762078310996_419/clk_in
+ scan_wrapper_334445762078310996_418/data_in scan_wrapper_334445762078310996_419/data_in
+ scan_wrapper_334445762078310996_418/latch_enable_in scan_wrapper_334445762078310996_419/latch_enable_in
+ scan_wrapper_334445762078310996_418/scan_select_in scan_wrapper_334445762078310996_419/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_407 scan_wrapper_334445762078310996_407/clk_in scan_wrapper_334445762078310996_408/clk_in
+ scan_wrapper_334445762078310996_407/data_in scan_wrapper_334445762078310996_408/data_in
+ scan_wrapper_334445762078310996_407/latch_enable_in scan_wrapper_334445762078310996_408/latch_enable_in
+ scan_wrapper_334445762078310996_407/scan_select_in scan_wrapper_334445762078310996_408/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_204 scan_wrapper_334445762078310996_204/clk_in scan_wrapper_334445762078310996_205/clk_in
+ scan_wrapper_334445762078310996_204/data_in scan_wrapper_334445762078310996_205/data_in
+ scan_wrapper_334445762078310996_204/latch_enable_in scan_wrapper_334445762078310996_205/latch_enable_in
+ scan_wrapper_334445762078310996_204/scan_select_in scan_wrapper_334445762078310996_205/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_215 scan_wrapper_334445762078310996_215/clk_in scan_wrapper_334445762078310996_216/clk_in
+ scan_wrapper_334445762078310996_215/data_in scan_wrapper_334445762078310996_216/data_in
+ scan_wrapper_334445762078310996_215/latch_enable_in scan_wrapper_334445762078310996_216/latch_enable_in
+ scan_wrapper_334445762078310996_215/scan_select_in scan_wrapper_334445762078310996_216/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_226 scan_wrapper_334445762078310996_226/clk_in scan_wrapper_334445762078310996_227/clk_in
+ scan_wrapper_334445762078310996_226/data_in scan_wrapper_334445762078310996_227/data_in
+ scan_wrapper_334445762078310996_226/latch_enable_in scan_wrapper_334445762078310996_227/latch_enable_in
+ scan_wrapper_334445762078310996_226/scan_select_in scan_wrapper_334445762078310996_227/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_237 scan_wrapper_334445762078310996_237/clk_in scan_wrapper_334445762078310996_238/clk_in
+ scan_wrapper_334445762078310996_237/data_in scan_wrapper_334445762078310996_238/data_in
+ scan_wrapper_334445762078310996_237/latch_enable_in scan_wrapper_334445762078310996_238/latch_enable_in
+ scan_wrapper_334445762078310996_237/scan_select_in scan_wrapper_334445762078310996_238/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_248 scan_wrapper_334445762078310996_248/clk_in scan_wrapper_334445762078310996_249/clk_in
+ scan_wrapper_334445762078310996_248/data_in scan_wrapper_334445762078310996_249/data_in
+ scan_wrapper_334445762078310996_248/latch_enable_in scan_wrapper_334445762078310996_249/latch_enable_in
+ scan_wrapper_334445762078310996_248/scan_select_in scan_wrapper_334445762078310996_249/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_259 scan_wrapper_334445762078310996_259/clk_in scan_wrapper_334445762078310996_260/clk_in
+ scan_wrapper_334445762078310996_259/data_in scan_wrapper_334445762078310996_260/data_in
+ scan_wrapper_334445762078310996_259/latch_enable_in scan_wrapper_334445762078310996_260/latch_enable_in
+ scan_wrapper_334445762078310996_259/scan_select_in scan_wrapper_334445762078310996_260/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_9 scan_wrapper_334445762078310996_9/clk_in scan_wrapper_334445762078310996_9/clk_out
+ scan_wrapper_334445762078310996_9/data_in scan_wrapper_334445762078310996_9/data_out
+ scan_wrapper_334445762078310996_9/latch_enable_in scan_wrapper_334445762078310996_9/latch_enable_out
+ scan_wrapper_334445762078310996_9/scan_select_in scan_wrapper_334445762078310996_9/scan_select_out
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_419 scan_wrapper_334445762078310996_419/clk_in scan_wrapper_334445762078310996_420/clk_in
+ scan_wrapper_334445762078310996_419/data_in scan_wrapper_334445762078310996_420/data_in
+ scan_wrapper_334445762078310996_419/latch_enable_in scan_wrapper_334445762078310996_420/latch_enable_in
+ scan_wrapper_334445762078310996_419/scan_select_in scan_wrapper_334445762078310996_420/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_408 scan_wrapper_334445762078310996_408/clk_in scan_wrapper_334445762078310996_409/clk_in
+ scan_wrapper_334445762078310996_408/data_in scan_wrapper_334445762078310996_409/data_in
+ scan_wrapper_334445762078310996_408/latch_enable_in scan_wrapper_334445762078310996_409/latch_enable_in
+ scan_wrapper_334445762078310996_408/scan_select_in scan_wrapper_334445762078310996_409/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_205 scan_wrapper_334445762078310996_205/clk_in scan_wrapper_334445762078310996_206/clk_in
+ scan_wrapper_334445762078310996_205/data_in scan_wrapper_334445762078310996_206/data_in
+ scan_wrapper_334445762078310996_205/latch_enable_in scan_wrapper_334445762078310996_206/latch_enable_in
+ scan_wrapper_334445762078310996_205/scan_select_in scan_wrapper_334445762078310996_206/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_216 scan_wrapper_334445762078310996_216/clk_in scan_wrapper_334445762078310996_217/clk_in
+ scan_wrapper_334445762078310996_216/data_in scan_wrapper_334445762078310996_217/data_in
+ scan_wrapper_334445762078310996_216/latch_enable_in scan_wrapper_334445762078310996_217/latch_enable_in
+ scan_wrapper_334445762078310996_216/scan_select_in scan_wrapper_334445762078310996_217/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_227 scan_wrapper_334445762078310996_227/clk_in scan_wrapper_334445762078310996_228/clk_in
+ scan_wrapper_334445762078310996_227/data_in scan_wrapper_334445762078310996_228/data_in
+ scan_wrapper_334445762078310996_227/latch_enable_in scan_wrapper_334445762078310996_228/latch_enable_in
+ scan_wrapper_334445762078310996_227/scan_select_in scan_wrapper_334445762078310996_228/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_238 scan_wrapper_334445762078310996_238/clk_in scan_wrapper_334445762078310996_239/clk_in
+ scan_wrapper_334445762078310996_238/data_in scan_wrapper_334445762078310996_239/data_in
+ scan_wrapper_334445762078310996_238/latch_enable_in scan_wrapper_334445762078310996_239/latch_enable_in
+ scan_wrapper_334445762078310996_238/scan_select_in scan_wrapper_334445762078310996_239/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_249 scan_wrapper_334445762078310996_249/clk_in scan_wrapper_334445762078310996_250/clk_in
+ scan_wrapper_334445762078310996_249/data_in scan_wrapper_334445762078310996_250/data_in
+ scan_wrapper_334445762078310996_249/latch_enable_in scan_wrapper_334445762078310996_250/latch_enable_in
+ scan_wrapper_334445762078310996_249/scan_select_in scan_wrapper_334445762078310996_250/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_409 scan_wrapper_334445762078310996_409/clk_in scan_wrapper_334445762078310996_410/clk_in
+ scan_wrapper_334445762078310996_409/data_in scan_wrapper_334445762078310996_410/data_in
+ scan_wrapper_334445762078310996_409/latch_enable_in scan_wrapper_334445762078310996_410/latch_enable_in
+ scan_wrapper_334445762078310996_409/scan_select_in scan_wrapper_334445762078310996_410/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_206 scan_wrapper_334445762078310996_206/clk_in scan_wrapper_334445762078310996_207/clk_in
+ scan_wrapper_334445762078310996_206/data_in scan_wrapper_334445762078310996_207/data_in
+ scan_wrapper_334445762078310996_206/latch_enable_in scan_wrapper_334445762078310996_207/latch_enable_in
+ scan_wrapper_334445762078310996_206/scan_select_in scan_wrapper_334445762078310996_207/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_217 scan_wrapper_334445762078310996_217/clk_in scan_wrapper_334445762078310996_218/clk_in
+ scan_wrapper_334445762078310996_217/data_in scan_wrapper_334445762078310996_218/data_in
+ scan_wrapper_334445762078310996_217/latch_enable_in scan_wrapper_334445762078310996_218/latch_enable_in
+ scan_wrapper_334445762078310996_217/scan_select_in scan_wrapper_334445762078310996_218/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_228 scan_wrapper_334445762078310996_228/clk_in scan_wrapper_334445762078310996_229/clk_in
+ scan_wrapper_334445762078310996_228/data_in scan_wrapper_334445762078310996_229/data_in
+ scan_wrapper_334445762078310996_228/latch_enable_in scan_wrapper_334445762078310996_229/latch_enable_in
+ scan_wrapper_334445762078310996_228/scan_select_in scan_wrapper_334445762078310996_229/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_239 scan_wrapper_334445762078310996_239/clk_in scan_wrapper_334445762078310996_240/clk_in
+ scan_wrapper_334445762078310996_239/data_in scan_wrapper_334445762078310996_240/data_in
+ scan_wrapper_334445762078310996_239/latch_enable_in scan_wrapper_334445762078310996_240/latch_enable_in
+ scan_wrapper_334445762078310996_239/scan_select_in scan_wrapper_334445762078310996_240/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_207 scan_wrapper_334445762078310996_207/clk_in scan_wrapper_334445762078310996_208/clk_in
+ scan_wrapper_334445762078310996_207/data_in scan_wrapper_334445762078310996_208/data_in
+ scan_wrapper_334445762078310996_207/latch_enable_in scan_wrapper_334445762078310996_208/latch_enable_in
+ scan_wrapper_334445762078310996_207/scan_select_in scan_wrapper_334445762078310996_208/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_218 scan_wrapper_334445762078310996_218/clk_in scan_wrapper_334445762078310996_219/clk_in
+ scan_wrapper_334445762078310996_218/data_in scan_wrapper_334445762078310996_219/data_in
+ scan_wrapper_334445762078310996_218/latch_enable_in scan_wrapper_334445762078310996_219/latch_enable_in
+ scan_wrapper_334445762078310996_218/scan_select_in scan_wrapper_334445762078310996_219/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_229 scan_wrapper_334445762078310996_229/clk_in scan_wrapper_334445762078310996_230/clk_in
+ scan_wrapper_334445762078310996_229/data_in scan_wrapper_334445762078310996_230/data_in
+ scan_wrapper_334445762078310996_229/latch_enable_in scan_wrapper_334445762078310996_230/latch_enable_in
+ scan_wrapper_334445762078310996_229/scan_select_in scan_wrapper_334445762078310996_230/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_390 scan_wrapper_334445762078310996_390/clk_in scan_wrapper_334445762078310996_391/clk_in
+ scan_wrapper_334445762078310996_390/data_in scan_wrapper_334445762078310996_391/data_in
+ scan_wrapper_334445762078310996_390/latch_enable_in scan_wrapper_334445762078310996_391/latch_enable_in
+ scan_wrapper_334445762078310996_390/scan_select_in scan_wrapper_334445762078310996_391/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_208 scan_wrapper_334445762078310996_208/clk_in scan_wrapper_334445762078310996_209/clk_in
+ scan_wrapper_334445762078310996_208/data_in scan_wrapper_334445762078310996_209/data_in
+ scan_wrapper_334445762078310996_208/latch_enable_in scan_wrapper_334445762078310996_209/latch_enable_in
+ scan_wrapper_334445762078310996_208/scan_select_in scan_wrapper_334445762078310996_209/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_219 scan_wrapper_334445762078310996_219/clk_in scan_wrapper_334445762078310996_220/clk_in
+ scan_wrapper_334445762078310996_219/data_in scan_wrapper_334445762078310996_220/data_in
+ scan_wrapper_334445762078310996_219/latch_enable_in scan_wrapper_334445762078310996_220/latch_enable_in
+ scan_wrapper_334445762078310996_219/scan_select_in scan_wrapper_334445762078310996_220/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_391 scan_wrapper_334445762078310996_391/clk_in scan_wrapper_334445762078310996_392/clk_in
+ scan_wrapper_334445762078310996_391/data_in scan_wrapper_334445762078310996_392/data_in
+ scan_wrapper_334445762078310996_391/latch_enable_in scan_wrapper_334445762078310996_392/latch_enable_in
+ scan_wrapper_334445762078310996_391/scan_select_in scan_wrapper_334445762078310996_392/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_380 scan_wrapper_334445762078310996_380/clk_in scan_wrapper_334445762078310996_381/clk_in
+ scan_wrapper_334445762078310996_380/data_in scan_wrapper_334445762078310996_381/data_in
+ scan_wrapper_334445762078310996_380/latch_enable_in scan_wrapper_334445762078310996_381/latch_enable_in
+ scan_wrapper_334445762078310996_380/scan_select_in scan_wrapper_334445762078310996_381/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_209 scan_wrapper_334445762078310996_209/clk_in scan_wrapper_334445762078310996_210/clk_in
+ scan_wrapper_334445762078310996_209/data_in scan_wrapper_334445762078310996_210/data_in
+ scan_wrapper_334445762078310996_209/latch_enable_in scan_wrapper_334445762078310996_210/latch_enable_in
+ scan_wrapper_334445762078310996_209/scan_select_in scan_wrapper_334445762078310996_210/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_392 scan_wrapper_334445762078310996_392/clk_in scan_wrapper_334445762078310996_393/clk_in
+ scan_wrapper_334445762078310996_392/data_in scan_wrapper_334445762078310996_393/data_in
+ scan_wrapper_334445762078310996_392/latch_enable_in scan_wrapper_334445762078310996_393/latch_enable_in
+ scan_wrapper_334445762078310996_392/scan_select_in scan_wrapper_334445762078310996_393/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_370 scan_wrapper_334445762078310996_370/clk_in scan_wrapper_334445762078310996_371/clk_in
+ scan_wrapper_334445762078310996_370/data_in scan_wrapper_334445762078310996_371/data_in
+ scan_wrapper_334445762078310996_370/latch_enable_in scan_wrapper_334445762078310996_371/latch_enable_in
+ scan_wrapper_334445762078310996_370/scan_select_in scan_wrapper_334445762078310996_371/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_381 scan_wrapper_334445762078310996_381/clk_in scan_wrapper_334445762078310996_382/clk_in
+ scan_wrapper_334445762078310996_381/data_in scan_wrapper_334445762078310996_382/data_in
+ scan_wrapper_334445762078310996_381/latch_enable_in scan_wrapper_334445762078310996_382/latch_enable_in
+ scan_wrapper_334445762078310996_381/scan_select_in scan_wrapper_334445762078310996_382/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_controller io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18]
+ io_in[19] io_in[20] wb_clk_i io_in[21] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26]
+ io_in[27] io_in[28] io_oeb[29] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_out[29] io_out[30] io_out[31] io_out[32] io_out[33]
+ io_out[34] io_out[35] io_out[36] io_out[37] wb_rst_i scan_controller/scan_clk scan_controller/scan_data_in
+ scan_controller/scan_data_out scan_controller/scan_latch_enable scan_controller/scan_select
+ vccd1 vssd1 scan_controller
Xscan_wrapper_334445762078310996_393 scan_wrapper_334445762078310996_393/clk_in scan_wrapper_334445762078310996_394/clk_in
+ scan_wrapper_334445762078310996_393/data_in scan_wrapper_334445762078310996_394/data_in
+ scan_wrapper_334445762078310996_393/latch_enable_in scan_wrapper_334445762078310996_394/latch_enable_in
+ scan_wrapper_334445762078310996_393/scan_select_in scan_wrapper_334445762078310996_394/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_360 scan_wrapper_334445762078310996_360/clk_in scan_wrapper_334445762078310996_361/clk_in
+ scan_wrapper_334445762078310996_360/data_in scan_wrapper_334445762078310996_361/data_in
+ scan_wrapper_334445762078310996_360/latch_enable_in scan_wrapper_334445762078310996_361/latch_enable_in
+ scan_wrapper_334445762078310996_360/scan_select_in scan_wrapper_334445762078310996_361/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_371 scan_wrapper_334445762078310996_371/clk_in scan_wrapper_334445762078310996_372/clk_in
+ scan_wrapper_334445762078310996_371/data_in scan_wrapper_334445762078310996_372/data_in
+ scan_wrapper_334445762078310996_371/latch_enable_in scan_wrapper_334445762078310996_372/latch_enable_in
+ scan_wrapper_334445762078310996_371/scan_select_in scan_wrapper_334445762078310996_372/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_382 scan_wrapper_334445762078310996_382/clk_in scan_wrapper_334445762078310996_383/clk_in
+ scan_wrapper_334445762078310996_382/data_in scan_wrapper_334445762078310996_383/data_in
+ scan_wrapper_334445762078310996_382/latch_enable_in scan_wrapper_334445762078310996_383/latch_enable_in
+ scan_wrapper_334445762078310996_382/scan_select_in scan_wrapper_334445762078310996_383/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_190 scan_wrapper_334445762078310996_190/clk_in scan_wrapper_334445762078310996_191/clk_in
+ scan_wrapper_334445762078310996_190/data_in scan_wrapper_334445762078310996_191/data_in
+ scan_wrapper_334445762078310996_190/latch_enable_in scan_wrapper_334445762078310996_191/latch_enable_in
+ scan_wrapper_334445762078310996_190/scan_select_in scan_wrapper_334445762078310996_191/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_394 scan_wrapper_334445762078310996_394/clk_in scan_wrapper_334445762078310996_395/clk_in
+ scan_wrapper_334445762078310996_394/data_in scan_wrapper_334445762078310996_395/data_in
+ scan_wrapper_334445762078310996_394/latch_enable_in scan_wrapper_334445762078310996_395/latch_enable_in
+ scan_wrapper_334445762078310996_394/scan_select_in scan_wrapper_334445762078310996_395/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_383 scan_wrapper_334445762078310996_383/clk_in scan_wrapper_334445762078310996_384/clk_in
+ scan_wrapper_334445762078310996_383/data_in scan_wrapper_334445762078310996_384/data_in
+ scan_wrapper_334445762078310996_383/latch_enable_in scan_wrapper_334445762078310996_384/latch_enable_in
+ scan_wrapper_334445762078310996_383/scan_select_in scan_wrapper_334445762078310996_384/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_350 scan_wrapper_334445762078310996_350/clk_in scan_wrapper_334445762078310996_351/clk_in
+ scan_wrapper_334445762078310996_350/data_in scan_wrapper_334445762078310996_351/data_in
+ scan_wrapper_334445762078310996_350/latch_enable_in scan_wrapper_334445762078310996_351/latch_enable_in
+ scan_wrapper_334445762078310996_350/scan_select_in scan_wrapper_334445762078310996_351/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_361 scan_wrapper_334445762078310996_361/clk_in scan_wrapper_334445762078310996_362/clk_in
+ scan_wrapper_334445762078310996_361/data_in scan_wrapper_334445762078310996_362/data_in
+ scan_wrapper_334445762078310996_361/latch_enable_in scan_wrapper_334445762078310996_362/latch_enable_in
+ scan_wrapper_334445762078310996_361/scan_select_in scan_wrapper_334445762078310996_362/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_372 scan_wrapper_334445762078310996_372/clk_in scan_wrapper_334445762078310996_373/clk_in
+ scan_wrapper_334445762078310996_372/data_in scan_wrapper_334445762078310996_373/data_in
+ scan_wrapper_334445762078310996_372/latch_enable_in scan_wrapper_334445762078310996_373/latch_enable_in
+ scan_wrapper_334445762078310996_372/scan_select_in scan_wrapper_334445762078310996_373/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_180 scan_wrapper_334445762078310996_180/clk_in scan_wrapper_334445762078310996_181/clk_in
+ scan_wrapper_334445762078310996_180/data_in scan_wrapper_334445762078310996_181/data_in
+ scan_wrapper_334445762078310996_180/latch_enable_in scan_wrapper_334445762078310996_181/latch_enable_in
+ scan_wrapper_334445762078310996_180/scan_select_in scan_wrapper_334445762078310996_181/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_191 scan_wrapper_334445762078310996_191/clk_in scan_wrapper_334445762078310996_192/clk_in
+ scan_wrapper_334445762078310996_191/data_in scan_wrapper_334445762078310996_192/data_in
+ scan_wrapper_334445762078310996_191/latch_enable_in scan_wrapper_334445762078310996_192/latch_enable_in
+ scan_wrapper_334445762078310996_191/scan_select_in scan_wrapper_334445762078310996_192/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_395 scan_wrapper_334445762078310996_395/clk_in scan_wrapper_334445762078310996_396/clk_in
+ scan_wrapper_334445762078310996_395/data_in scan_wrapper_334445762078310996_396/data_in
+ scan_wrapper_334445762078310996_395/latch_enable_in scan_wrapper_334445762078310996_396/latch_enable_in
+ scan_wrapper_334445762078310996_395/scan_select_in scan_wrapper_334445762078310996_396/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_384 scan_wrapper_334445762078310996_384/clk_in scan_wrapper_334445762078310996_385/clk_in
+ scan_wrapper_334445762078310996_384/data_in scan_wrapper_334445762078310996_385/data_in
+ scan_wrapper_334445762078310996_384/latch_enable_in scan_wrapper_334445762078310996_385/latch_enable_in
+ scan_wrapper_334445762078310996_384/scan_select_in scan_wrapper_334445762078310996_385/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_340 scan_wrapper_334445762078310996_340/clk_in scan_wrapper_334445762078310996_341/clk_in
+ scan_wrapper_334445762078310996_340/data_in scan_wrapper_334445762078310996_341/data_in
+ scan_wrapper_334445762078310996_340/latch_enable_in scan_wrapper_334445762078310996_341/latch_enable_in
+ scan_wrapper_334445762078310996_340/scan_select_in scan_wrapper_334445762078310996_341/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_351 scan_wrapper_334445762078310996_351/clk_in scan_wrapper_334445762078310996_352/clk_in
+ scan_wrapper_334445762078310996_351/data_in scan_wrapper_334445762078310996_352/data_in
+ scan_wrapper_334445762078310996_351/latch_enable_in scan_wrapper_334445762078310996_352/latch_enable_in
+ scan_wrapper_334445762078310996_351/scan_select_in scan_wrapper_334445762078310996_352/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_362 scan_wrapper_334445762078310996_362/clk_in scan_wrapper_334445762078310996_363/clk_in
+ scan_wrapper_334445762078310996_362/data_in scan_wrapper_334445762078310996_363/data_in
+ scan_wrapper_334445762078310996_362/latch_enable_in scan_wrapper_334445762078310996_363/latch_enable_in
+ scan_wrapper_334445762078310996_362/scan_select_in scan_wrapper_334445762078310996_363/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_373 scan_wrapper_334445762078310996_373/clk_in scan_wrapper_334445762078310996_374/clk_in
+ scan_wrapper_334445762078310996_373/data_in scan_wrapper_334445762078310996_374/data_in
+ scan_wrapper_334445762078310996_373/latch_enable_in scan_wrapper_334445762078310996_374/latch_enable_in
+ scan_wrapper_334445762078310996_373/scan_select_in scan_wrapper_334445762078310996_374/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_170 scan_wrapper_334445762078310996_170/clk_in scan_wrapper_334445762078310996_171/clk_in
+ scan_wrapper_334445762078310996_170/data_in scan_wrapper_334445762078310996_171/data_in
+ scan_wrapper_334445762078310996_170/latch_enable_in scan_wrapper_334445762078310996_171/latch_enable_in
+ scan_wrapper_334445762078310996_170/scan_select_in scan_wrapper_334445762078310996_171/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_181 scan_wrapper_334445762078310996_181/clk_in scan_wrapper_334445762078310996_182/clk_in
+ scan_wrapper_334445762078310996_181/data_in scan_wrapper_334445762078310996_182/data_in
+ scan_wrapper_334445762078310996_181/latch_enable_in scan_wrapper_334445762078310996_182/latch_enable_in
+ scan_wrapper_334445762078310996_181/scan_select_in scan_wrapper_334445762078310996_182/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_192 scan_wrapper_334445762078310996_192/clk_in scan_wrapper_334445762078310996_193/clk_in
+ scan_wrapper_334445762078310996_192/data_in scan_wrapper_334445762078310996_193/data_in
+ scan_wrapper_334445762078310996_192/latch_enable_in scan_wrapper_334445762078310996_193/latch_enable_in
+ scan_wrapper_334445762078310996_192/scan_select_in scan_wrapper_334445762078310996_193/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_396 scan_wrapper_334445762078310996_396/clk_in scan_wrapper_334445762078310996_397/clk_in
+ scan_wrapper_334445762078310996_396/data_in scan_wrapper_334445762078310996_397/data_in
+ scan_wrapper_334445762078310996_396/latch_enable_in scan_wrapper_334445762078310996_397/latch_enable_in
+ scan_wrapper_334445762078310996_396/scan_select_in scan_wrapper_334445762078310996_397/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_385 scan_wrapper_334445762078310996_385/clk_in scan_wrapper_334445762078310996_386/clk_in
+ scan_wrapper_334445762078310996_385/data_in scan_wrapper_334445762078310996_386/data_in
+ scan_wrapper_334445762078310996_385/latch_enable_in scan_wrapper_334445762078310996_386/latch_enable_in
+ scan_wrapper_334445762078310996_385/scan_select_in scan_wrapper_334445762078310996_386/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_330 scan_wrapper_334445762078310996_330/clk_in scan_wrapper_334445762078310996_331/clk_in
+ scan_wrapper_334445762078310996_330/data_in scan_wrapper_334445762078310996_331/data_in
+ scan_wrapper_334445762078310996_330/latch_enable_in scan_wrapper_334445762078310996_331/latch_enable_in
+ scan_wrapper_334445762078310996_330/scan_select_in scan_wrapper_334445762078310996_331/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_341 scan_wrapper_334445762078310996_341/clk_in scan_wrapper_334445762078310996_342/clk_in
+ scan_wrapper_334445762078310996_341/data_in scan_wrapper_334445762078310996_342/data_in
+ scan_wrapper_334445762078310996_341/latch_enable_in scan_wrapper_334445762078310996_342/latch_enable_in
+ scan_wrapper_334445762078310996_341/scan_select_in scan_wrapper_334445762078310996_342/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_352 scan_wrapper_334445762078310996_352/clk_in scan_wrapper_334445762078310996_353/clk_in
+ scan_wrapper_334445762078310996_352/data_in scan_wrapper_334445762078310996_353/data_in
+ scan_wrapper_334445762078310996_352/latch_enable_in scan_wrapper_334445762078310996_353/latch_enable_in
+ scan_wrapper_334445762078310996_352/scan_select_in scan_wrapper_334445762078310996_353/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_363 scan_wrapper_334445762078310996_363/clk_in scan_wrapper_334445762078310996_364/clk_in
+ scan_wrapper_334445762078310996_363/data_in scan_wrapper_334445762078310996_364/data_in
+ scan_wrapper_334445762078310996_363/latch_enable_in scan_wrapper_334445762078310996_364/latch_enable_in
+ scan_wrapper_334445762078310996_363/scan_select_in scan_wrapper_334445762078310996_364/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_374 scan_wrapper_334445762078310996_374/clk_in scan_wrapper_334445762078310996_375/clk_in
+ scan_wrapper_334445762078310996_374/data_in scan_wrapper_334445762078310996_375/data_in
+ scan_wrapper_334445762078310996_374/latch_enable_in scan_wrapper_334445762078310996_375/latch_enable_in
+ scan_wrapper_334445762078310996_374/scan_select_in scan_wrapper_334445762078310996_375/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_160 scan_wrapper_334445762078310996_160/clk_in scan_wrapper_334445762078310996_161/clk_in
+ scan_wrapper_334445762078310996_160/data_in scan_wrapper_334445762078310996_161/data_in
+ scan_wrapper_334445762078310996_160/latch_enable_in scan_wrapper_334445762078310996_161/latch_enable_in
+ scan_wrapper_334445762078310996_160/scan_select_in scan_wrapper_334445762078310996_161/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_171 scan_wrapper_334445762078310996_171/clk_in scan_wrapper_334445762078310996_172/clk_in
+ scan_wrapper_334445762078310996_171/data_in scan_wrapper_334445762078310996_172/data_in
+ scan_wrapper_334445762078310996_171/latch_enable_in scan_wrapper_334445762078310996_172/latch_enable_in
+ scan_wrapper_334445762078310996_171/scan_select_in scan_wrapper_334445762078310996_172/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_182 scan_wrapper_334445762078310996_182/clk_in scan_wrapper_334445762078310996_183/clk_in
+ scan_wrapper_334445762078310996_182/data_in scan_wrapper_334445762078310996_183/data_in
+ scan_wrapper_334445762078310996_182/latch_enable_in scan_wrapper_334445762078310996_183/latch_enable_in
+ scan_wrapper_334445762078310996_182/scan_select_in scan_wrapper_334445762078310996_183/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
Xscan_wrapper_334445762078310996_193 scan_wrapper_334445762078310996_193/clk_in scan_wrapper_334445762078310996_194/clk_in
+ scan_wrapper_334445762078310996_193/data_in scan_wrapper_334445762078310996_194/data_in
+ scan_wrapper_334445762078310996_193/latch_enable_in scan_wrapper_334445762078310996_194/latch_enable_in
+ scan_wrapper_334445762078310996_193/scan_select_in scan_wrapper_334445762078310996_194/scan_select_in
+ vccd1 vssd1 scan_wrapper_334445762078310996
.ends

