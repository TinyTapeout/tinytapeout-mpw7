module scan_wrapper_341438392303616596 (clk_in,
    clk_out,
    data_in,
    data_out,
    latch_enable_in,
    latch_enable_out,
    scan_select_in,
    scan_select_out,
    vccd1,
    vssd1);
 input clk_in;
 output clk_out;
 input data_in;
 output data_out;
 input latch_enable_in;
 output latch_enable_out;
 input scan_select_in;
 output scan_select_out;
 input vccd1;
 input vssd1;

 wire clk;
 wire data_out_i;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire \scan_data_in[1] ;
 wire \scan_data_in[2] ;
 wire \scan_data_in[3] ;
 wire \scan_data_in[4] ;
 wire \scan_data_in[5] ;
 wire \scan_data_in[6] ;
 wire \scan_data_in[7] ;
 wire \scan_data_out[7] ;
 wire \user_module.net1 ;
 wire \user_module.net10 ;
 wire \user_module.net11 ;
 wire \user_module.net12 ;
 wire \user_module.net2 ;
 wire \user_module.net3 ;
 wire \user_module.net4 ;
 wire \user_module.net5 ;
 wire \user_module.net6 ;
 wire \user_module.net7 ;
 wire \user_module.net8 ;
 wire \user_module.net9 ;

 sky130_fd_sc_hd__decap_3 FILLER_0_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_13 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_111 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_123 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_11_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_11_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_119 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_12_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_12_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_12_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_133 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_145 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_13_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_13_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_13_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_14_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_49 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_14_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_14_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_15_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_146 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_15_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_127 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_16_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_17_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_119 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_18_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_18_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_18_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_19_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_1_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_21_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_23_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_24_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_24_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_24_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_25_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_26_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_174 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_26_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_18 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_27_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_27_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_30 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_42 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_27_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_28_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_28_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_28_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_29_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_29_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_29_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_29_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_29_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_2_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_2_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_2_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_2_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_3_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_3_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_3_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_5_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_7_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_9_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _45_ (.A(\user_module.net1 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.net9 ));
 sky130_fd_sc_hd__clkinv_2 _46_ (.A(\user_module.net4 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.net12 ));
 sky130_fd_sc_hd__clkinv_2 _47_ (.A(\user_module.net3 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.net11 ));
 sky130_fd_sc_hd__clkinv_2 _48_ (.A(\user_module.net2 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.net10 ));
 sky130_fd_sc_hd__conb_1 _58__4 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net4));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(data_in),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(latch_enable_in),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(scan_select_in),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input_buf_clk (.A(clk_in),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clk));
 sky130_fd_sc_hd__dlxtp_1 \latch[0]  (.D(\scan_data_in[1] ),
    .GATE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.net1 ));
 sky130_fd_sc_hd__dlxtp_1 \latch[1]  (.D(\scan_data_in[2] ),
    .GATE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.net2 ));
 sky130_fd_sc_hd__dlxtp_1 \latch[2]  (.D(\scan_data_in[3] ),
    .GATE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.net3 ));
 sky130_fd_sc_hd__dlxtp_1 \latch[3]  (.D(\scan_data_in[4] ),
    .GATE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.net4 ));
 sky130_fd_sc_hd__dlxtp_1 \latch[4]  (.D(\scan_data_in[5] ),
    .GATE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.net5 ));
 sky130_fd_sc_hd__dlxtp_1 \latch[5]  (.D(\scan_data_in[6] ),
    .GATE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.net6 ));
 sky130_fd_sc_hd__dlxtp_1 \latch[6]  (.D(\scan_data_in[7] ),
    .GATE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.net7 ));
 sky130_fd_sc_hd__dlxtp_1 \latch[7]  (.D(\scan_data_out[7] ),
    .GATE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.net8 ));
 sky130_fd_sc_hd__dfrtn_1 out_flop (.CLK_N(clk),
    .D(\scan_data_out[7] ),
    .RESET_B(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(data_out_i));
 sky130_fd_sc_hd__buf_4 \output_buffers[0]  (.A(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(latch_enable_out));
 sky130_fd_sc_hd__buf_4 \output_buffers[1]  (.A(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(scan_select_out));
 sky130_fd_sc_hd__buf_4 \output_buffers[2]  (.A(data_out_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(data_out));
 sky130_fd_sc_hd__buf_4 \output_buffers[3]  (.A(clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clk_out));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[0]  (.CLK(clk),
    .D(net1),
    .SCD(\user_module.net9 ),
    .SCE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\scan_data_in[1] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[1]  (.CLK(clk),
    .D(\scan_data_in[1] ),
    .SCD(\user_module.net10 ),
    .SCE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\scan_data_in[2] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[2]  (.CLK(clk),
    .D(\scan_data_in[2] ),
    .SCD(\user_module.net11 ),
    .SCE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\scan_data_in[3] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[3]  (.CLK(clk),
    .D(\scan_data_in[3] ),
    .SCD(\user_module.net12 ),
    .SCE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\scan_data_in[4] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[4]  (.CLK(clk),
    .D(\scan_data_in[4] ),
    .SCD(\user_module.net5 ),
    .SCE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\scan_data_in[5] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[5]  (.CLK(clk),
    .D(\scan_data_in[5] ),
    .SCD(\user_module.net6 ),
    .SCE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\scan_data_in[6] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[6]  (.CLK(clk),
    .D(\scan_data_in[6] ),
    .SCD(\user_module.net7 ),
    .SCE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\scan_data_in[7] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[7]  (.CLK(clk),
    .D(\scan_data_in[7] ),
    .SCD(\user_module.net8 ),
    .SCE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\scan_data_out[7] ));
endmodule
