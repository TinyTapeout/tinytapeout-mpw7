module scan_wrapper_341263346544149074 (clk_in,
    clk_out,
    data_in,
    data_out,
    latch_enable_in,
    latch_enable_out,
    scan_select_in,
    scan_select_out,
    vccd1,
    vssd1);
 input clk_in;
 output clk_out;
 input data_in;
 output data_out;
 input latch_enable_in;
 output latch_enable_out;
 input scan_select_in;
 output scan_select_out;
 input vccd1;
 input vssd1;

 wire clk;
 wire data_out_i;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire \scan_data_in[1] ;
 wire \scan_data_in[2] ;
 wire \scan_data_in[3] ;
 wire \scan_data_in[4] ;
 wire \scan_data_in[5] ;
 wire \scan_data_in[6] ;
 wire \scan_data_in[7] ;
 wire \scan_data_out[7] ;
 wire \user_module.clk ;
 wire \user_module.data[10][0] ;
 wire \user_module.data[10][1] ;
 wire \user_module.data[10][2] ;
 wire \user_module.data[10][3] ;
 wire \user_module.data[11][0] ;
 wire \user_module.data[11][1] ;
 wire \user_module.data[11][2] ;
 wire \user_module.data[11][3] ;
 wire \user_module.data[12][0] ;
 wire \user_module.data[12][1] ;
 wire \user_module.data[12][2] ;
 wire \user_module.data[12][3] ;
 wire \user_module.data[13][0] ;
 wire \user_module.data[13][1] ;
 wire \user_module.data[13][2] ;
 wire \user_module.data[13][3] ;
 wire \user_module.data[14][0] ;
 wire \user_module.data[14][1] ;
 wire \user_module.data[14][2] ;
 wire \user_module.data[14][3] ;
 wire \user_module.data[15][0] ;
 wire \user_module.data[15][1] ;
 wire \user_module.data[15][2] ;
 wire \user_module.data[15][3] ;
 wire \user_module.data[16][0] ;
 wire \user_module.data[16][1] ;
 wire \user_module.data[16][2] ;
 wire \user_module.data[16][3] ;
 wire \user_module.data[17][0] ;
 wire \user_module.data[17][1] ;
 wire \user_module.data[17][2] ;
 wire \user_module.data[17][3] ;
 wire \user_module.data[18][0] ;
 wire \user_module.data[18][1] ;
 wire \user_module.data[18][2] ;
 wire \user_module.data[18][3] ;
 wire \user_module.data[19][0] ;
 wire \user_module.data[19][1] ;
 wire \user_module.data[19][2] ;
 wire \user_module.data[19][3] ;
 wire \user_module.data[1][0] ;
 wire \user_module.data[1][1] ;
 wire \user_module.data[1][2] ;
 wire \user_module.data[1][3] ;
 wire \user_module.data[20][0] ;
 wire \user_module.data[20][1] ;
 wire \user_module.data[20][2] ;
 wire \user_module.data[20][3] ;
 wire \user_module.data[21][0] ;
 wire \user_module.data[21][1] ;
 wire \user_module.data[21][2] ;
 wire \user_module.data[21][3] ;
 wire \user_module.data[22][0] ;
 wire \user_module.data[22][1] ;
 wire \user_module.data[22][2] ;
 wire \user_module.data[22][3] ;
 wire \user_module.data[23][0] ;
 wire \user_module.data[23][1] ;
 wire \user_module.data[23][2] ;
 wire \user_module.data[23][3] ;
 wire \user_module.data[24][0] ;
 wire \user_module.data[24][1] ;
 wire \user_module.data[24][2] ;
 wire \user_module.data[24][3] ;
 wire \user_module.data[25][0] ;
 wire \user_module.data[25][1] ;
 wire \user_module.data[25][2] ;
 wire \user_module.data[25][3] ;
 wire \user_module.data[2][0] ;
 wire \user_module.data[2][1] ;
 wire \user_module.data[2][2] ;
 wire \user_module.data[2][3] ;
 wire \user_module.data[3][0] ;
 wire \user_module.data[3][1] ;
 wire \user_module.data[3][2] ;
 wire \user_module.data[3][3] ;
 wire \user_module.data[4][0] ;
 wire \user_module.data[4][1] ;
 wire \user_module.data[4][2] ;
 wire \user_module.data[4][3] ;
 wire \user_module.data[5][0] ;
 wire \user_module.data[5][1] ;
 wire \user_module.data[5][2] ;
 wire \user_module.data[5][3] ;
 wire \user_module.data[6][0] ;
 wire \user_module.data[6][1] ;
 wire \user_module.data[6][2] ;
 wire \user_module.data[6][3] ;
 wire \user_module.data[7][0] ;
 wire \user_module.data[7][1] ;
 wire \user_module.data[7][2] ;
 wire \user_module.data[7][3] ;
 wire \user_module.data[8][0] ;
 wire \user_module.data[8][1] ;
 wire \user_module.data[8][2] ;
 wire \user_module.data[8][3] ;
 wire \user_module.data[9][0] ;
 wire \user_module.data[9][1] ;
 wire \user_module.data[9][2] ;
 wire \user_module.data[9][3] ;
 wire \user_module.io_in[0] ;
 wire \user_module.io_in[1] ;
 wire \user_module.io_in[2] ;
 wire \user_module.io_in[3] ;
 wire \user_module.io_in[4] ;
 wire \user_module.io_in[5] ;
 wire \user_module.io_in[6] ;
 wire \user_module.io_in[7] ;
 wire \user_module.rd_empty ;
 wire \user_module.rd_ena ;
 wire \user_module.rd_ena_n ;
 wire \user_module.rst_n ;
 wire \user_module.stage[10].l_ce ;
 wire \user_module.stage[10].l_clk ;
 wire \user_module.stage[10].l_data_mux[0] ;
 wire \user_module.stage[10].l_data_mux[1] ;
 wire \user_module.stage[10].l_data_mux[2] ;
 wire \user_module.stage[10].l_data_mux[3] ;
 wire \user_module.stage[10].l_valid_comb ;
 wire \user_module.stage[10].l_valid_n ;
 wire \user_module.stage[10].l_valid_reg ;
 wire \user_module.stage[11].l_ce ;
 wire \user_module.stage[11].l_clk ;
 wire \user_module.stage[11].l_data_mux[0] ;
 wire \user_module.stage[11].l_data_mux[1] ;
 wire \user_module.stage[11].l_data_mux[2] ;
 wire \user_module.stage[11].l_data_mux[3] ;
 wire \user_module.stage[11].l_valid_comb ;
 wire \user_module.stage[11].l_valid_n ;
 wire \user_module.stage[11].l_valid_reg ;
 wire \user_module.stage[12].l_ce ;
 wire \user_module.stage[12].l_clk ;
 wire \user_module.stage[12].l_data_mux[0] ;
 wire \user_module.stage[12].l_data_mux[1] ;
 wire \user_module.stage[12].l_data_mux[2] ;
 wire \user_module.stage[12].l_data_mux[3] ;
 wire \user_module.stage[12].l_valid_comb ;
 wire \user_module.stage[12].l_valid_n ;
 wire \user_module.stage[12].l_valid_reg ;
 wire \user_module.stage[13].l_ce ;
 wire \user_module.stage[13].l_clk ;
 wire \user_module.stage[13].l_data_mux[0] ;
 wire \user_module.stage[13].l_data_mux[1] ;
 wire \user_module.stage[13].l_data_mux[2] ;
 wire \user_module.stage[13].l_data_mux[3] ;
 wire \user_module.stage[13].l_valid_comb ;
 wire \user_module.stage[13].l_valid_n ;
 wire \user_module.stage[13].l_valid_reg ;
 wire \user_module.stage[14].l_ce ;
 wire \user_module.stage[14].l_clk ;
 wire \user_module.stage[14].l_data_mux[0] ;
 wire \user_module.stage[14].l_data_mux[1] ;
 wire \user_module.stage[14].l_data_mux[2] ;
 wire \user_module.stage[14].l_data_mux[3] ;
 wire \user_module.stage[14].l_valid_comb ;
 wire \user_module.stage[14].l_valid_n ;
 wire \user_module.stage[14].l_valid_reg ;
 wire \user_module.stage[15].l_ce ;
 wire \user_module.stage[15].l_clk ;
 wire \user_module.stage[15].l_data_mux[0] ;
 wire \user_module.stage[15].l_data_mux[1] ;
 wire \user_module.stage[15].l_data_mux[2] ;
 wire \user_module.stage[15].l_data_mux[3] ;
 wire \user_module.stage[15].l_valid_comb ;
 wire \user_module.stage[15].l_valid_n ;
 wire \user_module.stage[15].l_valid_reg ;
 wire \user_module.stage[16].l_ce ;
 wire \user_module.stage[16].l_clk ;
 wire \user_module.stage[16].l_data_mux[0] ;
 wire \user_module.stage[16].l_data_mux[1] ;
 wire \user_module.stage[16].l_data_mux[2] ;
 wire \user_module.stage[16].l_data_mux[3] ;
 wire \user_module.stage[16].l_valid_comb ;
 wire \user_module.stage[16].l_valid_n ;
 wire \user_module.stage[16].l_valid_reg ;
 wire \user_module.stage[17].l_ce ;
 wire \user_module.stage[17].l_clk ;
 wire \user_module.stage[17].l_data_mux[0] ;
 wire \user_module.stage[17].l_data_mux[1] ;
 wire \user_module.stage[17].l_data_mux[2] ;
 wire \user_module.stage[17].l_data_mux[3] ;
 wire \user_module.stage[17].l_valid_comb ;
 wire \user_module.stage[17].l_valid_n ;
 wire \user_module.stage[17].l_valid_reg ;
 wire \user_module.stage[18].l_ce ;
 wire \user_module.stage[18].l_clk ;
 wire \user_module.stage[18].l_data_mux[0] ;
 wire \user_module.stage[18].l_data_mux[1] ;
 wire \user_module.stage[18].l_data_mux[2] ;
 wire \user_module.stage[18].l_data_mux[3] ;
 wire \user_module.stage[18].l_valid_comb ;
 wire \user_module.stage[18].l_valid_n ;
 wire \user_module.stage[18].l_valid_reg ;
 wire \user_module.stage[19].l_ce ;
 wire \user_module.stage[19].l_clk ;
 wire \user_module.stage[19].l_data_mux[0] ;
 wire \user_module.stage[19].l_data_mux[1] ;
 wire \user_module.stage[19].l_data_mux[2] ;
 wire \user_module.stage[19].l_data_mux[3] ;
 wire \user_module.stage[19].l_valid_comb ;
 wire \user_module.stage[19].l_valid_n ;
 wire \user_module.stage[19].l_valid_reg ;
 wire \user_module.stage[1].l_ce ;
 wire \user_module.stage[1].l_clk ;
 wire \user_module.stage[1].l_data_mux[0] ;
 wire \user_module.stage[1].l_data_mux[1] ;
 wire \user_module.stage[1].l_data_mux[2] ;
 wire \user_module.stage[1].l_data_mux[3] ;
 wire \user_module.stage[1].l_valid_comb ;
 wire \user_module.stage[1].l_valid_n ;
 wire \user_module.stage[1].l_valid_reg ;
 wire \user_module.stage[20].l_ce ;
 wire \user_module.stage[20].l_clk ;
 wire \user_module.stage[20].l_data_mux[0] ;
 wire \user_module.stage[20].l_data_mux[1] ;
 wire \user_module.stage[20].l_data_mux[2] ;
 wire \user_module.stage[20].l_data_mux[3] ;
 wire \user_module.stage[20].l_valid_comb ;
 wire \user_module.stage[20].l_valid_n ;
 wire \user_module.stage[20].l_valid_reg ;
 wire \user_module.stage[21].l_ce ;
 wire \user_module.stage[21].l_clk ;
 wire \user_module.stage[21].l_data_mux[0] ;
 wire \user_module.stage[21].l_data_mux[1] ;
 wire \user_module.stage[21].l_data_mux[2] ;
 wire \user_module.stage[21].l_data_mux[3] ;
 wire \user_module.stage[21].l_valid_comb ;
 wire \user_module.stage[21].l_valid_n ;
 wire \user_module.stage[21].l_valid_reg ;
 wire \user_module.stage[22].l_ce ;
 wire \user_module.stage[22].l_clk ;
 wire \user_module.stage[22].l_data_mux[0] ;
 wire \user_module.stage[22].l_data_mux[1] ;
 wire \user_module.stage[22].l_data_mux[2] ;
 wire \user_module.stage[22].l_data_mux[3] ;
 wire \user_module.stage[22].l_valid_comb ;
 wire \user_module.stage[22].l_valid_n ;
 wire \user_module.stage[22].l_valid_reg ;
 wire \user_module.stage[23].l_ce ;
 wire \user_module.stage[23].l_clk ;
 wire \user_module.stage[23].l_data_mux[0] ;
 wire \user_module.stage[23].l_data_mux[1] ;
 wire \user_module.stage[23].l_data_mux[2] ;
 wire \user_module.stage[23].l_data_mux[3] ;
 wire \user_module.stage[23].l_valid_comb ;
 wire \user_module.stage[23].l_valid_n ;
 wire \user_module.stage[23].l_valid_reg ;
 wire \user_module.stage[24].l_ce ;
 wire \user_module.stage[24].l_clk ;
 wire \user_module.stage[24].l_valid_comb ;
 wire \user_module.stage[24].l_valid_n ;
 wire \user_module.stage[24].l_valid_reg ;
 wire \user_module.stage[2].l_ce ;
 wire \user_module.stage[2].l_clk ;
 wire \user_module.stage[2].l_data_mux[0] ;
 wire \user_module.stage[2].l_data_mux[1] ;
 wire \user_module.stage[2].l_data_mux[2] ;
 wire \user_module.stage[2].l_data_mux[3] ;
 wire \user_module.stage[2].l_valid_comb ;
 wire \user_module.stage[2].l_valid_n ;
 wire \user_module.stage[2].l_valid_reg ;
 wire \user_module.stage[3].l_ce ;
 wire \user_module.stage[3].l_clk ;
 wire \user_module.stage[3].l_data_mux[0] ;
 wire \user_module.stage[3].l_data_mux[1] ;
 wire \user_module.stage[3].l_data_mux[2] ;
 wire \user_module.stage[3].l_data_mux[3] ;
 wire \user_module.stage[3].l_valid_comb ;
 wire \user_module.stage[3].l_valid_n ;
 wire \user_module.stage[3].l_valid_reg ;
 wire \user_module.stage[4].l_ce ;
 wire \user_module.stage[4].l_clk ;
 wire \user_module.stage[4].l_data_mux[0] ;
 wire \user_module.stage[4].l_data_mux[1] ;
 wire \user_module.stage[4].l_data_mux[2] ;
 wire \user_module.stage[4].l_data_mux[3] ;
 wire \user_module.stage[4].l_valid_comb ;
 wire \user_module.stage[4].l_valid_n ;
 wire \user_module.stage[4].l_valid_reg ;
 wire \user_module.stage[5].l_ce ;
 wire \user_module.stage[5].l_clk ;
 wire \user_module.stage[5].l_data_mux[0] ;
 wire \user_module.stage[5].l_data_mux[1] ;
 wire \user_module.stage[5].l_data_mux[2] ;
 wire \user_module.stage[5].l_data_mux[3] ;
 wire \user_module.stage[5].l_valid_comb ;
 wire \user_module.stage[5].l_valid_n ;
 wire \user_module.stage[5].l_valid_reg ;
 wire \user_module.stage[6].l_ce ;
 wire \user_module.stage[6].l_clk ;
 wire \user_module.stage[6].l_data_mux[0] ;
 wire \user_module.stage[6].l_data_mux[1] ;
 wire \user_module.stage[6].l_data_mux[2] ;
 wire \user_module.stage[6].l_data_mux[3] ;
 wire \user_module.stage[6].l_valid_comb ;
 wire \user_module.stage[6].l_valid_n ;
 wire \user_module.stage[6].l_valid_reg ;
 wire \user_module.stage[7].l_ce ;
 wire \user_module.stage[7].l_clk ;
 wire \user_module.stage[7].l_data_mux[0] ;
 wire \user_module.stage[7].l_data_mux[1] ;
 wire \user_module.stage[7].l_data_mux[2] ;
 wire \user_module.stage[7].l_data_mux[3] ;
 wire \user_module.stage[7].l_valid_comb ;
 wire \user_module.stage[7].l_valid_n ;
 wire \user_module.stage[7].l_valid_reg ;
 wire \user_module.stage[8].l_ce ;
 wire \user_module.stage[8].l_clk ;
 wire \user_module.stage[8].l_data_mux[0] ;
 wire \user_module.stage[8].l_data_mux[1] ;
 wire \user_module.stage[8].l_data_mux[2] ;
 wire \user_module.stage[8].l_data_mux[3] ;
 wire \user_module.stage[8].l_valid_comb ;
 wire \user_module.stage[8].l_valid_n ;
 wire \user_module.stage[8].l_valid_reg ;
 wire \user_module.stage[9].l_ce ;
 wire \user_module.stage[9].l_clk ;
 wire \user_module.stage[9].l_data_mux[0] ;
 wire \user_module.stage[9].l_data_mux[1] ;
 wire \user_module.stage[9].l_data_mux[2] ;
 wire \user_module.stage[9].l_data_mux[3] ;
 wire \user_module.stage[9].l_valid_comb ;
 wire \user_module.stage[9].l_valid_n ;
 wire \user_module.stage[9].l_valid_reg ;
 wire \user_module.wr_ena ;

 sky130_fd_sc_hd__diode_2 ANTENNA_0 (.DIODE(\user_module.data[20][2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\user_module.data[20][3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\user_module.stage[12].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\user_module.stage[8].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_9 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_10_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_12_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_14_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_19_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_1_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_140 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_152 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_1_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_1_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_22_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_22_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_22_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_23_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_24_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_168 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_25_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_26_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_184 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_176 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_188 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_27_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_28_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_168 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_180 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_156 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_29_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_148 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_160 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_172 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_184 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_2_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_148 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_160 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_30_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_30_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_30_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_30_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_140 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_152 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_31_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_31_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_31_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_33_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_33_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_33_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_33_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_33_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_33_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_33_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_3_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_3_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_3_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_3_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_4_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_159 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_171 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_176 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_188 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_5_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_6_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_6_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_6_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_7_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_189 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_7_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_7_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_170 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _5__7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net7));
 sky130_fd_sc_hd__conb_1 _6__8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net8));
 sky130_fd_sc_hd__conb_1 _7__4 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net4));
 sky130_fd_sc_hd__conb_1 _8__5 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net5));
 sky130_fd_sc_hd__conb_1 _9__6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net6));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(data_in),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(latch_enable_in),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(scan_select_in),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input_buf_clk (.A(clk_in),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clk));
 sky130_fd_sc_hd__dlxtp_1 \latch[0]  (.D(\scan_data_in[1] ),
    .GATE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.io_in[0] ));
 sky130_fd_sc_hd__dlxtp_1 \latch[1]  (.D(\scan_data_in[2] ),
    .GATE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.io_in[1] ));
 sky130_fd_sc_hd__dlxtp_1 \latch[2]  (.D(\scan_data_in[3] ),
    .GATE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.io_in[2] ));
 sky130_fd_sc_hd__dlxtp_1 \latch[3]  (.D(\scan_data_in[4] ),
    .GATE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.io_in[3] ));
 sky130_fd_sc_hd__dlxtp_1 \latch[4]  (.D(\scan_data_in[5] ),
    .GATE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.io_in[4] ));
 sky130_fd_sc_hd__dlxtp_1 \latch[5]  (.D(\scan_data_in[6] ),
    .GATE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.io_in[5] ));
 sky130_fd_sc_hd__dlxtp_1 \latch[6]  (.D(\scan_data_in[7] ),
    .GATE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.io_in[6] ));
 sky130_fd_sc_hd__dlxtp_1 \latch[7]  (.D(\scan_data_out[7] ),
    .GATE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.io_in[7] ));
 sky130_fd_sc_hd__dfrtn_1 out_flop (.CLK_N(clk),
    .D(\scan_data_out[7] ),
    .RESET_B(net7),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(data_out_i));
 sky130_fd_sc_hd__buf_4 \output_buffers[0]  (.A(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(latch_enable_out));
 sky130_fd_sc_hd__buf_4 \output_buffers[1]  (.A(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(scan_select_out));
 sky130_fd_sc_hd__buf_4 \output_buffers[2]  (.A(data_out_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(data_out));
 sky130_fd_sc_hd__buf_4 \output_buffers[3]  (.A(clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clk_out));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[0]  (.CLK(clk),
    .D(net1),
    .SCD(net4),
    .SCE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\scan_data_in[1] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[1]  (.CLK(clk),
    .D(\scan_data_in[1] ),
    .SCD(net5),
    .SCE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\scan_data_in[2] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[2]  (.CLK(clk),
    .D(\scan_data_in[2] ),
    .SCD(\user_module.stage[24].l_valid_reg ),
    .SCE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\scan_data_in[3] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[3]  (.CLK(clk),
    .D(\scan_data_in[3] ),
    .SCD(\user_module.rd_empty ),
    .SCE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\scan_data_in[4] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[4]  (.CLK(clk),
    .D(\scan_data_in[4] ),
    .SCD(\user_module.data[1][0] ),
    .SCE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\scan_data_in[5] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[5]  (.CLK(clk),
    .D(\scan_data_in[5] ),
    .SCD(\user_module.data[1][1] ),
    .SCE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\scan_data_in[6] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[6]  (.CLK(clk),
    .D(\scan_data_in[6] ),
    .SCD(\user_module.data[1][2] ),
    .SCE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\scan_data_in[7] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[7]  (.CLK(clk),
    .D(\scan_data_in[7] ),
    .SCD(\user_module.data[1][3] ),
    .SCE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\scan_data_out[7] ));
 sky130_fd_sc_hd__inv_1 \user_module.empty_I  (.A(\user_module.stage[1].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.rd_empty ));
 sky130_fd_sc_hd__clkbuf_4 \user_module.inbuf_clk_I  (.A(\user_module.io_in[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.clk ));
 sky130_fd_sc_hd__buf_6 \user_module.inbuf_rd_ena_I  (.A(\user_module.io_in[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.rd_ena ));
 sky130_fd_sc_hd__inv_6 \user_module.inbuf_rd_ena_n_I  (.A(\user_module.io_in[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.rd_ena_n ));
 sky130_fd_sc_hd__buf_8 \user_module.inbuf_rst_I  (.A(\user_module.io_in[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.rst_n ));
 sky130_fd_sc_hd__buf_4 \user_module.inbuf_wr_data_I[0]  (.A(\user_module.io_in[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.data[25][0] ));
 sky130_fd_sc_hd__buf_4 \user_module.inbuf_wr_data_I[1]  (.A(\user_module.io_in[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.data[25][1] ));
 sky130_fd_sc_hd__buf_4 \user_module.inbuf_wr_data_I[2]  (.A(\user_module.io_in[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.data[25][2] ));
 sky130_fd_sc_hd__buf_4 \user_module.inbuf_wr_data_I[3]  (.A(\user_module.io_in[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.data[25][3] ));
 sky130_fd_sc_hd__buf_12 \user_module.inbuf_wr_ena_I  (.A(\user_module.io_in[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.wr_ena ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[10].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[10].l_valid_n ),
    .A3(\user_module.stage[9].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[10].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[10].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[10].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[10].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[10].data_reg_I[0]  (.CLK(\user_module.stage[10].l_clk ),
    .D(\user_module.stage[10].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[10].data_reg_I[1]  (.CLK(\user_module.stage[10].l_clk ),
    .D(\user_module.stage[10].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[10].data_reg_I[2]  (.CLK(\user_module.stage[10].l_clk ),
    .D(\user_module.stage[10].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[10].data_reg_I[3]  (.CLK(\user_module.stage[10].l_clk ),
    .D(\user_module.stage[10].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[10][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[10].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[11][0] ),
    .S(\user_module.stage[11].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[10].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[10].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[11][1] ),
    .S(\user_module.stage[11].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[10].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[10].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[11][2] ),
    .S(\user_module.stage[11].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[10].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[10].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[11][3] ),
    .S(\user_module.stage[11].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[10].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[10].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[10].l_valid_reg ),
    .B1(\user_module.stage[11].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[10].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[10].valid_n_I  (.A(\user_module.stage[10].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[10].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[10].valid_reg_I  (.CLK(\user_module.stage[10].l_clk ),
    .D(\user_module.stage[10].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[10].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[11].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[11].l_valid_n ),
    .A3(\user_module.stage[10].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[11].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[11].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[11].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[11].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[11].data_reg_I[0]  (.CLK(\user_module.stage[11].l_clk ),
    .D(\user_module.stage[11].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[11].data_reg_I[1]  (.CLK(\user_module.stage[11].l_clk ),
    .D(\user_module.stage[11].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[11].data_reg_I[2]  (.CLK(\user_module.stage[11].l_clk ),
    .D(\user_module.stage[11].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[11].data_reg_I[3]  (.CLK(\user_module.stage[11].l_clk ),
    .D(\user_module.stage[11].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[11][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[11].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[12][0] ),
    .S(\user_module.stage[12].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[11].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[11].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[12][1] ),
    .S(\user_module.stage[12].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[11].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[11].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[12][2] ),
    .S(\user_module.stage[12].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[11].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[11].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[12][3] ),
    .S(\user_module.stage[12].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[11].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[11].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[11].l_valid_reg ),
    .B1(\user_module.stage[12].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[11].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[11].valid_n_I  (.A(\user_module.stage[11].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[11].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[11].valid_reg_I  (.CLK(\user_module.stage[11].l_clk ),
    .D(\user_module.stage[11].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[11].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[12].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[12].l_valid_n ),
    .A3(\user_module.stage[11].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[12].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[12].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[12].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[12].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[12].data_reg_I[0]  (.CLK(\user_module.stage[12].l_clk ),
    .D(\user_module.stage[12].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[12].data_reg_I[1]  (.CLK(\user_module.stage[12].l_clk ),
    .D(\user_module.stage[12].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[12].data_reg_I[2]  (.CLK(\user_module.stage[12].l_clk ),
    .D(\user_module.stage[12].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[12].data_reg_I[3]  (.CLK(\user_module.stage[12].l_clk ),
    .D(\user_module.stage[12].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[12][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[12].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[13][0] ),
    .S(\user_module.stage[13].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[12].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[12].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[13][1] ),
    .S(\user_module.stage[13].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[12].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[12].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[13][2] ),
    .S(\user_module.stage[13].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[12].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[12].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[13][3] ),
    .S(\user_module.stage[13].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[12].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[12].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[12].l_valid_reg ),
    .B1(\user_module.stage[13].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[12].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[12].valid_n_I  (.A(\user_module.stage[12].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[12].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[12].valid_reg_I  (.CLK(\user_module.stage[12].l_clk ),
    .D(\user_module.stage[12].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[12].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[13].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[13].l_valid_n ),
    .A3(\user_module.stage[12].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[13].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[13].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[13].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[13].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[13].data_reg_I[0]  (.CLK(\user_module.stage[13].l_clk ),
    .D(\user_module.stage[13].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[13].data_reg_I[1]  (.CLK(\user_module.stage[13].l_clk ),
    .D(\user_module.stage[13].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[13].data_reg_I[2]  (.CLK(\user_module.stage[13].l_clk ),
    .D(\user_module.stage[13].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[13].data_reg_I[3]  (.CLK(\user_module.stage[13].l_clk ),
    .D(\user_module.stage[13].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[13][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[13].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[14][0] ),
    .S(\user_module.stage[14].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[13].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[13].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[14][1] ),
    .S(\user_module.stage[14].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[13].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[13].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[14][2] ),
    .S(\user_module.stage[14].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[13].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[13].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[14][3] ),
    .S(\user_module.stage[14].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[13].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[13].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[13].l_valid_reg ),
    .B1(\user_module.stage[14].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[13].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[13].valid_n_I  (.A(\user_module.stage[13].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[13].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[13].valid_reg_I  (.CLK(\user_module.stage[13].l_clk ),
    .D(\user_module.stage[13].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[13].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[14].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[14].l_valid_n ),
    .A3(\user_module.stage[13].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[14].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[14].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[14].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[14].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[14].data_reg_I[0]  (.CLK(\user_module.stage[14].l_clk ),
    .D(\user_module.stage[14].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[14].data_reg_I[1]  (.CLK(\user_module.stage[14].l_clk ),
    .D(\user_module.stage[14].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[14].data_reg_I[2]  (.CLK(\user_module.stage[14].l_clk ),
    .D(\user_module.stage[14].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[14].data_reg_I[3]  (.CLK(\user_module.stage[14].l_clk ),
    .D(\user_module.stage[14].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[14][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[14].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[15][0] ),
    .S(\user_module.stage[15].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[14].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[14].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[15][1] ),
    .S(\user_module.stage[15].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[14].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[14].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[15][2] ),
    .S(\user_module.stage[15].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[14].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[14].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[15][3] ),
    .S(\user_module.stage[15].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[14].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[14].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[14].l_valid_reg ),
    .B1(\user_module.stage[15].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[14].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[14].valid_n_I  (.A(\user_module.stage[14].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[14].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[14].valid_reg_I  (.CLK(\user_module.stage[14].l_clk ),
    .D(\user_module.stage[14].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[14].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[15].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[15].l_valid_n ),
    .A3(\user_module.stage[14].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[15].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[15].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[15].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[15].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[15].data_reg_I[0]  (.CLK(\user_module.stage[15].l_clk ),
    .D(\user_module.stage[15].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[15].data_reg_I[1]  (.CLK(\user_module.stage[15].l_clk ),
    .D(\user_module.stage[15].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[15].data_reg_I[2]  (.CLK(\user_module.stage[15].l_clk ),
    .D(\user_module.stage[15].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[15].data_reg_I[3]  (.CLK(\user_module.stage[15].l_clk ),
    .D(\user_module.stage[15].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[15][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[15].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[16][0] ),
    .S(\user_module.stage[16].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[15].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[15].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[16][1] ),
    .S(\user_module.stage[16].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[15].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[15].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[16][2] ),
    .S(\user_module.stage[16].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[15].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[15].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[16][3] ),
    .S(\user_module.stage[16].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[15].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[15].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[15].l_valid_reg ),
    .B1(\user_module.stage[16].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[15].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[15].valid_n_I  (.A(\user_module.stage[15].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[15].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[15].valid_reg_I  (.CLK(\user_module.stage[15].l_clk ),
    .D(\user_module.stage[15].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[15].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[16].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[16].l_valid_n ),
    .A3(\user_module.stage[15].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[16].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[16].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[16].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[16].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[16].data_reg_I[0]  (.CLK(\user_module.stage[16].l_clk ),
    .D(\user_module.stage[16].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[16].data_reg_I[1]  (.CLK(\user_module.stage[16].l_clk ),
    .D(\user_module.stage[16].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[16].data_reg_I[2]  (.CLK(\user_module.stage[16].l_clk ),
    .D(\user_module.stage[16].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[16].data_reg_I[3]  (.CLK(\user_module.stage[16].l_clk ),
    .D(\user_module.stage[16].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[16][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[16].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[17][0] ),
    .S(\user_module.stage[17].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[16].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[16].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[17][1] ),
    .S(\user_module.stage[17].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[16].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[16].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[17][2] ),
    .S(\user_module.stage[17].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[16].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[16].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[17][3] ),
    .S(\user_module.stage[17].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[16].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[16].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[16].l_valid_reg ),
    .B1(\user_module.stage[17].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[16].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[16].valid_n_I  (.A(\user_module.stage[16].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[16].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[16].valid_reg_I  (.CLK(\user_module.stage[16].l_clk ),
    .D(\user_module.stage[16].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[16].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[17].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[17].l_valid_n ),
    .A3(\user_module.stage[16].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[17].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[17].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[17].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[17].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[17].data_reg_I[0]  (.CLK(\user_module.stage[17].l_clk ),
    .D(\user_module.stage[17].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[17].data_reg_I[1]  (.CLK(\user_module.stage[17].l_clk ),
    .D(\user_module.stage[17].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[17].data_reg_I[2]  (.CLK(\user_module.stage[17].l_clk ),
    .D(\user_module.stage[17].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[17].data_reg_I[3]  (.CLK(\user_module.stage[17].l_clk ),
    .D(\user_module.stage[17].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[17][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[17].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[18][0] ),
    .S(\user_module.stage[18].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[17].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[17].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[18][1] ),
    .S(\user_module.stage[18].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[17].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[17].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[18][2] ),
    .S(\user_module.stage[18].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[17].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[17].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[18][3] ),
    .S(\user_module.stage[18].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[17].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[17].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[17].l_valid_reg ),
    .B1(\user_module.stage[18].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[17].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[17].valid_n_I  (.A(\user_module.stage[17].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[17].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[17].valid_reg_I  (.CLK(\user_module.stage[17].l_clk ),
    .D(\user_module.stage[17].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[17].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[18].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[18].l_valid_n ),
    .A3(\user_module.stage[17].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[18].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[18].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[18].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[18].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[18].data_reg_I[0]  (.CLK(\user_module.stage[18].l_clk ),
    .D(\user_module.stage[18].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[18].data_reg_I[1]  (.CLK(\user_module.stage[18].l_clk ),
    .D(\user_module.stage[18].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[18].data_reg_I[2]  (.CLK(\user_module.stage[18].l_clk ),
    .D(\user_module.stage[18].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[18].data_reg_I[3]  (.CLK(\user_module.stage[18].l_clk ),
    .D(\user_module.stage[18].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[18][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[18].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[19][0] ),
    .S(\user_module.stage[19].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[18].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[18].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[19][1] ),
    .S(\user_module.stage[19].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[18].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[18].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[19][2] ),
    .S(\user_module.stage[19].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[18].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[18].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[19][3] ),
    .S(\user_module.stage[19].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[18].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[18].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[18].l_valid_reg ),
    .B1(\user_module.stage[19].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[18].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[18].valid_n_I  (.A(\user_module.stage[18].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[18].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[18].valid_reg_I  (.CLK(\user_module.stage[18].l_clk ),
    .D(\user_module.stage[18].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[18].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[19].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[19].l_valid_n ),
    .A3(\user_module.stage[18].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[19].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[19].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[19].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[19].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[19].data_reg_I[0]  (.CLK(\user_module.stage[19].l_clk ),
    .D(\user_module.stage[19].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[19].data_reg_I[1]  (.CLK(\user_module.stage[19].l_clk ),
    .D(\user_module.stage[19].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[19].data_reg_I[2]  (.CLK(\user_module.stage[19].l_clk ),
    .D(\user_module.stage[19].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[19].data_reg_I[3]  (.CLK(\user_module.stage[19].l_clk ),
    .D(\user_module.stage[19].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[19][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[19].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[20][0] ),
    .S(\user_module.stage[20].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[19].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[19].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[20][1] ),
    .S(\user_module.stage[20].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[19].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[19].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[20][2] ),
    .S(\user_module.stage[20].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[19].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[19].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[20][3] ),
    .S(\user_module.stage[20].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[19].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[19].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[19].l_valid_reg ),
    .B1(\user_module.stage[20].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[19].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[19].valid_n_I  (.A(\user_module.stage[19].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[19].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[19].valid_reg_I  (.CLK(\user_module.stage[19].l_clk ),
    .D(\user_module.stage[19].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[19].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[1].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[1].l_valid_n ),
    .A3(net8),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[1].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[1].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[1].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[1].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[1].data_reg_I[0]  (.CLK(\user_module.stage[1].l_clk ),
    .D(\user_module.stage[1].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[1].data_reg_I[1]  (.CLK(\user_module.stage[1].l_clk ),
    .D(\user_module.stage[1].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[1].data_reg_I[2]  (.CLK(\user_module.stage[1].l_clk ),
    .D(\user_module.stage[1].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[1].data_reg_I[3]  (.CLK(\user_module.stage[1].l_clk ),
    .D(\user_module.stage[1].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[1][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[1].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[2][0] ),
    .S(\user_module.stage[2].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[1].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[1].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[2][1] ),
    .S(\user_module.stage[2].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[1].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[1].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[2][2] ),
    .S(\user_module.stage[2].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[1].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[1].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[2][3] ),
    .S(\user_module.stage[2].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[1].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[1].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[1].l_valid_reg ),
    .B1(\user_module.stage[2].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[1].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[1].valid_n_I  (.A(\user_module.stage[1].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[1].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_1 \user_module.stage[1].valid_reg_I  (.CLK(\user_module.stage[1].l_clk ),
    .D(\user_module.stage[1].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[1].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[20].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[20].l_valid_n ),
    .A3(\user_module.stage[19].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[20].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[20].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[20].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[20].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[20].data_reg_I[0]  (.CLK(\user_module.stage[20].l_clk ),
    .D(\user_module.stage[20].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[20].data_reg_I[1]  (.CLK(\user_module.stage[20].l_clk ),
    .D(\user_module.stage[20].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[20].data_reg_I[2]  (.CLK(\user_module.stage[20].l_clk ),
    .D(\user_module.stage[20].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[20].data_reg_I[3]  (.CLK(\user_module.stage[20].l_clk ),
    .D(\user_module.stage[20].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[20][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[20].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[21][0] ),
    .S(\user_module.stage[21].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[20].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[20].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[21][1] ),
    .S(\user_module.stage[21].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[20].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[20].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[21][2] ),
    .S(\user_module.stage[21].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[20].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[20].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[21][3] ),
    .S(\user_module.stage[21].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[20].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[20].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[20].l_valid_reg ),
    .B1(\user_module.stage[21].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[20].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[20].valid_n_I  (.A(\user_module.stage[20].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[20].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[20].valid_reg_I  (.CLK(\user_module.stage[20].l_clk ),
    .D(\user_module.stage[20].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[20].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[21].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[21].l_valid_n ),
    .A3(\user_module.stage[20].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[21].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[21].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[21].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[21].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[21].data_reg_I[0]  (.CLK(\user_module.stage[21].l_clk ),
    .D(\user_module.stage[21].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[21].data_reg_I[1]  (.CLK(\user_module.stage[21].l_clk ),
    .D(\user_module.stage[21].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[21].data_reg_I[2]  (.CLK(\user_module.stage[21].l_clk ),
    .D(\user_module.stage[21].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[21].data_reg_I[3]  (.CLK(\user_module.stage[21].l_clk ),
    .D(\user_module.stage[21].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[21][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[21].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[22][0] ),
    .S(\user_module.stage[22].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[21].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[21].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[22][1] ),
    .S(\user_module.stage[22].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[21].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[21].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[22][2] ),
    .S(\user_module.stage[22].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[21].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[21].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[22][3] ),
    .S(\user_module.stage[22].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[21].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[21].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[21].l_valid_reg ),
    .B1(\user_module.stage[22].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[21].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[21].valid_n_I  (.A(\user_module.stage[21].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[21].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[21].valid_reg_I  (.CLK(\user_module.stage[21].l_clk ),
    .D(\user_module.stage[21].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[21].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[22].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[22].l_valid_n ),
    .A3(\user_module.stage[21].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[22].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[22].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[22].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[22].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[22].data_reg_I[0]  (.CLK(\user_module.stage[22].l_clk ),
    .D(\user_module.stage[22].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[22].data_reg_I[1]  (.CLK(\user_module.stage[22].l_clk ),
    .D(\user_module.stage[22].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[22].data_reg_I[2]  (.CLK(\user_module.stage[22].l_clk ),
    .D(\user_module.stage[22].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[22].data_reg_I[3]  (.CLK(\user_module.stage[22].l_clk ),
    .D(\user_module.stage[22].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[22][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[22].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[23][0] ),
    .S(\user_module.stage[23].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[22].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[22].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[23][1] ),
    .S(\user_module.stage[23].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[22].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[22].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[23][2] ),
    .S(\user_module.stage[23].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[22].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[22].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[23][3] ),
    .S(\user_module.stage[23].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[22].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[22].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[22].l_valid_reg ),
    .B1(\user_module.stage[23].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[22].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[22].valid_n_I  (.A(\user_module.stage[22].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[22].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[22].valid_reg_I  (.CLK(\user_module.stage[22].l_clk ),
    .D(\user_module.stage[22].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[22].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[23].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[23].l_valid_n ),
    .A3(\user_module.stage[22].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[23].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[23].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[23].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[23].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[23].data_reg_I[0]  (.CLK(\user_module.stage[23].l_clk ),
    .D(\user_module.stage[23].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[23].data_reg_I[1]  (.CLK(\user_module.stage[23].l_clk ),
    .D(\user_module.stage[23].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[23].data_reg_I[2]  (.CLK(\user_module.stage[23].l_clk ),
    .D(\user_module.stage[23].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[23].data_reg_I[3]  (.CLK(\user_module.stage[23].l_clk ),
    .D(\user_module.stage[23].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[23][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[23].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[24][0] ),
    .S(\user_module.stage[24].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[23].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[23].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[24][1] ),
    .S(\user_module.stage[24].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[23].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[23].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[24][2] ),
    .S(\user_module.stage[24].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[23].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[23].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[24][3] ),
    .S(\user_module.stage[24].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[23].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[23].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[23].l_valid_reg ),
    .B1(\user_module.stage[24].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[23].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[23].valid_n_I  (.A(\user_module.stage[23].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[23].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[23].valid_reg_I  (.CLK(\user_module.stage[23].l_clk ),
    .D(\user_module.stage[23].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[23].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[24].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[24].l_valid_n ),
    .A3(\user_module.stage[23].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[24].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[24].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[24].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[24].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[24].data_reg_I[0]  (.CLK(\user_module.stage[24].l_clk ),
    .D(\user_module.data[25][0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[24].data_reg_I[1]  (.CLK(\user_module.stage[24].l_clk ),
    .D(\user_module.data[25][1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[24].data_reg_I[2]  (.CLK(\user_module.stage[24].l_clk ),
    .D(\user_module.data[25][2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[24].data_reg_I[3]  (.CLK(\user_module.stage[24].l_clk ),
    .D(\user_module.data[25][3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[24][3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[24].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[24].l_valid_reg ),
    .B1(net6),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[24].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[24].valid_n_I  (.A(\user_module.stage[24].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[24].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[24].valid_reg_I  (.CLK(\user_module.stage[24].l_clk ),
    .D(\user_module.stage[24].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[24].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[2].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[2].l_valid_n ),
    .A3(\user_module.stage[1].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[2].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[2].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[2].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[2].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[2].data_reg_I[0]  (.CLK(\user_module.stage[2].l_clk ),
    .D(\user_module.stage[2].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[2].data_reg_I[1]  (.CLK(\user_module.stage[2].l_clk ),
    .D(\user_module.stage[2].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[2].data_reg_I[2]  (.CLK(\user_module.stage[2].l_clk ),
    .D(\user_module.stage[2].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[2].data_reg_I[3]  (.CLK(\user_module.stage[2].l_clk ),
    .D(\user_module.stage[2].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[2][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[2].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[3][0] ),
    .S(\user_module.stage[3].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[2].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[2].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[3][1] ),
    .S(\user_module.stage[3].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[2].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[2].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[3][2] ),
    .S(\user_module.stage[3].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[2].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[2].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[3][3] ),
    .S(\user_module.stage[3].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[2].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[2].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[2].l_valid_reg ),
    .B1(\user_module.stage[3].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[2].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[2].valid_n_I  (.A(\user_module.stage[2].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[2].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[2].valid_reg_I  (.CLK(\user_module.stage[2].l_clk ),
    .D(\user_module.stage[2].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[2].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[3].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[3].l_valid_n ),
    .A3(\user_module.stage[2].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[3].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[3].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[3].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[3].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[3].data_reg_I[0]  (.CLK(\user_module.stage[3].l_clk ),
    .D(\user_module.stage[3].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[3].data_reg_I[1]  (.CLK(\user_module.stage[3].l_clk ),
    .D(\user_module.stage[3].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[3].data_reg_I[2]  (.CLK(\user_module.stage[3].l_clk ),
    .D(\user_module.stage[3].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[3].data_reg_I[3]  (.CLK(\user_module.stage[3].l_clk ),
    .D(\user_module.stage[3].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[3][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[3].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[4][0] ),
    .S(\user_module.stage[4].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[3].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[3].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[4][1] ),
    .S(\user_module.stage[4].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[3].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[3].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[4][2] ),
    .S(\user_module.stage[4].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[3].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[3].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[4][3] ),
    .S(\user_module.stage[4].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[3].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[3].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[3].l_valid_reg ),
    .B1(\user_module.stage[4].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[3].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[3].valid_n_I  (.A(\user_module.stage[3].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[3].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[3].valid_reg_I  (.CLK(\user_module.stage[3].l_clk ),
    .D(\user_module.stage[3].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[3].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[4].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[4].l_valid_n ),
    .A3(\user_module.stage[3].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[4].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[4].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[4].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[4].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[4].data_reg_I[0]  (.CLK(\user_module.stage[4].l_clk ),
    .D(\user_module.stage[4].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[4].data_reg_I[1]  (.CLK(\user_module.stage[4].l_clk ),
    .D(\user_module.stage[4].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[4].data_reg_I[2]  (.CLK(\user_module.stage[4].l_clk ),
    .D(\user_module.stage[4].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[4].data_reg_I[3]  (.CLK(\user_module.stage[4].l_clk ),
    .D(\user_module.stage[4].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[4][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[4].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[5][0] ),
    .S(\user_module.stage[5].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[4].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[4].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[5][1] ),
    .S(\user_module.stage[5].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[4].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[4].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[5][2] ),
    .S(\user_module.stage[5].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[4].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[4].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[5][3] ),
    .S(\user_module.stage[5].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[4].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[4].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[4].l_valid_reg ),
    .B1(\user_module.stage[5].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[4].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[4].valid_n_I  (.A(\user_module.stage[4].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[4].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[4].valid_reg_I  (.CLK(\user_module.stage[4].l_clk ),
    .D(\user_module.stage[4].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[4].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[5].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[5].l_valid_n ),
    .A3(\user_module.stage[4].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[5].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[5].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[5].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[5].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[5].data_reg_I[0]  (.CLK(\user_module.stage[5].l_clk ),
    .D(\user_module.stage[5].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[5].data_reg_I[1]  (.CLK(\user_module.stage[5].l_clk ),
    .D(\user_module.stage[5].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[5].data_reg_I[2]  (.CLK(\user_module.stage[5].l_clk ),
    .D(\user_module.stage[5].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[5].data_reg_I[3]  (.CLK(\user_module.stage[5].l_clk ),
    .D(\user_module.stage[5].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[5][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[5].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[6][0] ),
    .S(\user_module.stage[6].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[5].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[5].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[6][1] ),
    .S(\user_module.stage[6].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[5].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[5].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[6][2] ),
    .S(\user_module.stage[6].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[5].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[5].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[6][3] ),
    .S(\user_module.stage[6].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[5].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[5].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[5].l_valid_reg ),
    .B1(\user_module.stage[6].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[5].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[5].valid_n_I  (.A(\user_module.stage[5].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[5].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[5].valid_reg_I  (.CLK(\user_module.stage[5].l_clk ),
    .D(\user_module.stage[5].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[5].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[6].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[6].l_valid_n ),
    .A3(\user_module.stage[5].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[6].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[6].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[6].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[6].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[6].data_reg_I[0]  (.CLK(\user_module.stage[6].l_clk ),
    .D(\user_module.stage[6].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[6].data_reg_I[1]  (.CLK(\user_module.stage[6].l_clk ),
    .D(\user_module.stage[6].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[6].data_reg_I[2]  (.CLK(\user_module.stage[6].l_clk ),
    .D(\user_module.stage[6].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[6].data_reg_I[3]  (.CLK(\user_module.stage[6].l_clk ),
    .D(\user_module.stage[6].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[6][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[6].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[7][0] ),
    .S(\user_module.stage[7].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[6].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[6].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[7][1] ),
    .S(\user_module.stage[7].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[6].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[6].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[7][2] ),
    .S(\user_module.stage[7].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[6].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[6].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[7][3] ),
    .S(\user_module.stage[7].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[6].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[6].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[6].l_valid_reg ),
    .B1(\user_module.stage[7].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[6].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[6].valid_n_I  (.A(\user_module.stage[6].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[6].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[6].valid_reg_I  (.CLK(\user_module.stage[6].l_clk ),
    .D(\user_module.stage[6].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[6].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[7].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[7].l_valid_n ),
    .A3(\user_module.stage[6].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[7].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[7].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[7].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[7].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[7].data_reg_I[0]  (.CLK(\user_module.stage[7].l_clk ),
    .D(\user_module.stage[7].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[7].data_reg_I[1]  (.CLK(\user_module.stage[7].l_clk ),
    .D(\user_module.stage[7].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[7].data_reg_I[2]  (.CLK(\user_module.stage[7].l_clk ),
    .D(\user_module.stage[7].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[7].data_reg_I[3]  (.CLK(\user_module.stage[7].l_clk ),
    .D(\user_module.stage[7].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[7][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[7].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[8][0] ),
    .S(\user_module.stage[8].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[7].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[7].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[8][1] ),
    .S(\user_module.stage[8].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[7].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[7].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[8][2] ),
    .S(\user_module.stage[8].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[7].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[7].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[8][3] ),
    .S(\user_module.stage[8].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[7].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[7].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[7].l_valid_reg ),
    .B1(\user_module.stage[8].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[7].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[7].valid_n_I  (.A(\user_module.stage[7].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[7].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[7].valid_reg_I  (.CLK(\user_module.stage[7].l_clk ),
    .D(\user_module.stage[7].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[7].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[8].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[8].l_valid_n ),
    .A3(\user_module.stage[7].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[8].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[8].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[8].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[8].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[8].data_reg_I[0]  (.CLK(\user_module.stage[8].l_clk ),
    .D(\user_module.stage[8].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[8].data_reg_I[1]  (.CLK(\user_module.stage[8].l_clk ),
    .D(\user_module.stage[8].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[8].data_reg_I[2]  (.CLK(\user_module.stage[8].l_clk ),
    .D(\user_module.stage[8].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[8].data_reg_I[3]  (.CLK(\user_module.stage[8].l_clk ),
    .D(\user_module.stage[8].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[8][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[8].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[9][0] ),
    .S(\user_module.stage[9].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[8].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[8].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[9][1] ),
    .S(\user_module.stage[9].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[8].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[8].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[9][2] ),
    .S(\user_module.stage[9].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[8].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[8].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[9][3] ),
    .S(\user_module.stage[9].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[8].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[8].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[8].l_valid_reg ),
    .B1(\user_module.stage[9].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[8].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[8].valid_n_I  (.A(\user_module.stage[8].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[8].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[8].valid_reg_I  (.CLK(\user_module.stage[8].l_clk ),
    .D(\user_module.stage[8].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[8].l_valid_reg ));
 sky130_fd_sc_hd__a31o_1 \user_module.stage[9].ce_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[9].l_valid_n ),
    .A3(\user_module.stage[8].l_valid_reg ),
    .B1(\user_module.rd_ena ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[9].l_ce ));
 sky130_fd_sc_hd__dlclkp_1 \user_module.stage[9].clk_gate_I  (.CLK(\user_module.clk ),
    .GATE(\user_module.stage[9].l_ce ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .GCLK(\user_module.stage[9].l_clk ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[9].data_reg_I[0]  (.CLK(\user_module.stage[9].l_clk ),
    .D(\user_module.stage[9].l_data_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[9].data_reg_I[1]  (.CLK(\user_module.stage[9].l_clk ),
    .D(\user_module.stage[9].l_data_mux[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[9].data_reg_I[2]  (.CLK(\user_module.stage[9].l_clk ),
    .D(\user_module.stage[9].l_data_mux[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.stage[9].data_reg_I[3]  (.CLK(\user_module.stage[9].l_clk ),
    .D(\user_module.stage[9].l_data_mux[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.data[9][3] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[9].genblk1.data_mux_I[0]  (.A0(\user_module.data[25][0] ),
    .A1(\user_module.data[10][0] ),
    .S(\user_module.stage[10].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[9].l_data_mux[0] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[9].genblk1.data_mux_I[1]  (.A0(\user_module.data[25][1] ),
    .A1(\user_module.data[10][1] ),
    .S(\user_module.stage[10].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[9].l_data_mux[1] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[9].genblk1.data_mux_I[2]  (.A0(\user_module.data[25][2] ),
    .A1(\user_module.data[10][2] ),
    .S(\user_module.stage[10].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[9].l_data_mux[2] ));
 sky130_fd_sc_hd__mux2_1 \user_module.stage[9].genblk1.data_mux_I[3]  (.A0(\user_module.data[25][3] ),
    .A1(\user_module.data[10][3] ),
    .S(\user_module.stage[10].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[9].l_data_mux[3] ));
 sky130_fd_sc_hd__a211o_1 \user_module.stage[9].valid_comb_I  (.A1(\user_module.wr_ena ),
    .A2(\user_module.stage[9].l_valid_reg ),
    .B1(\user_module.stage[10].l_valid_reg ),
    .C1(\user_module.rd_ena_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.stage[9].l_valid_comb ));
 sky130_fd_sc_hd__inv_1 \user_module.stage[9].valid_n_I  (.A(\user_module.stage[9].l_valid_reg ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.stage[9].l_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 \user_module.stage[9].valid_reg_I  (.CLK(\user_module.stage[9].l_clk ),
    .D(\user_module.stage[9].l_valid_comb ),
    .RESET_B(\user_module.rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.stage[9].l_valid_reg ));
endmodule
