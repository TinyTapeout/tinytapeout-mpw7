module user_project_wrapper (user_clock2,
    vccd1,
    vccd2,
    vdda1,
    vdda2,
    vssa1,
    vssa2,
    vssd1,
    vssd2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input vccd1;
 input vccd2;
 input vdda1;
 input vdda2;
 input vssa1;
 input vssa2;
 input vssd1;
 input vssd2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire slow_clk;
 wire ready;
 wire \clk[0] ;
 wire \clk[100] ;
 wire \clk[101] ;
 wire \clk[102] ;
 wire \clk[103] ;
 wire \clk[104] ;
 wire \clk[105] ;
 wire \clk[106] ;
 wire \clk[107] ;
 wire \clk[108] ;
 wire \clk[109] ;
 wire \clk[10] ;
 wire \clk[110] ;
 wire \clk[111] ;
 wire \clk[112] ;
 wire \clk[113] ;
 wire \clk[114] ;
 wire \clk[115] ;
 wire \clk[116] ;
 wire \clk[117] ;
 wire \clk[118] ;
 wire \clk[119] ;
 wire \clk[11] ;
 wire \clk[120] ;
 wire \clk[121] ;
 wire \clk[122] ;
 wire \clk[123] ;
 wire \clk[124] ;
 wire \clk[125] ;
 wire \clk[126] ;
 wire \clk[127] ;
 wire \clk[128] ;
 wire \clk[129] ;
 wire \clk[12] ;
 wire \clk[130] ;
 wire \clk[131] ;
 wire \clk[132] ;
 wire \clk[133] ;
 wire \clk[134] ;
 wire \clk[135] ;
 wire \clk[136] ;
 wire \clk[137] ;
 wire \clk[138] ;
 wire \clk[139] ;
 wire \clk[13] ;
 wire \clk[140] ;
 wire \clk[141] ;
 wire \clk[142] ;
 wire \clk[143] ;
 wire \clk[144] ;
 wire \clk[145] ;
 wire \clk[146] ;
 wire \clk[147] ;
 wire \clk[148] ;
 wire \clk[149] ;
 wire \clk[14] ;
 wire \clk[150] ;
 wire \clk[151] ;
 wire \clk[152] ;
 wire \clk[153] ;
 wire \clk[154] ;
 wire \clk[155] ;
 wire \clk[156] ;
 wire \clk[157] ;
 wire \clk[158] ;
 wire \clk[159] ;
 wire \clk[15] ;
 wire \clk[160] ;
 wire \clk[161] ;
 wire \clk[162] ;
 wire \clk[163] ;
 wire \clk[164] ;
 wire \clk[165] ;
 wire \clk[166] ;
 wire \clk[167] ;
 wire \clk[168] ;
 wire \clk[169] ;
 wire \clk[16] ;
 wire \clk[170] ;
 wire \clk[171] ;
 wire \clk[172] ;
 wire \clk[173] ;
 wire \clk[174] ;
 wire \clk[175] ;
 wire \clk[176] ;
 wire \clk[177] ;
 wire \clk[178] ;
 wire \clk[179] ;
 wire \clk[17] ;
 wire \clk[180] ;
 wire \clk[181] ;
 wire \clk[182] ;
 wire \clk[183] ;
 wire \clk[184] ;
 wire \clk[185] ;
 wire \clk[186] ;
 wire \clk[187] ;
 wire \clk[188] ;
 wire \clk[189] ;
 wire \clk[18] ;
 wire \clk[190] ;
 wire \clk[191] ;
 wire \clk[192] ;
 wire \clk[193] ;
 wire \clk[194] ;
 wire \clk[195] ;
 wire \clk[196] ;
 wire \clk[197] ;
 wire \clk[198] ;
 wire \clk[199] ;
 wire \clk[19] ;
 wire \clk[1] ;
 wire \clk[200] ;
 wire \clk[201] ;
 wire \clk[202] ;
 wire \clk[203] ;
 wire \clk[204] ;
 wire \clk[205] ;
 wire \clk[206] ;
 wire \clk[207] ;
 wire \clk[208] ;
 wire \clk[209] ;
 wire \clk[20] ;
 wire \clk[210] ;
 wire \clk[211] ;
 wire \clk[212] ;
 wire \clk[213] ;
 wire \clk[214] ;
 wire \clk[215] ;
 wire \clk[216] ;
 wire \clk[217] ;
 wire \clk[218] ;
 wire \clk[219] ;
 wire \clk[21] ;
 wire \clk[220] ;
 wire \clk[221] ;
 wire \clk[222] ;
 wire \clk[223] ;
 wire \clk[224] ;
 wire \clk[225] ;
 wire \clk[226] ;
 wire \clk[227] ;
 wire \clk[228] ;
 wire \clk[229] ;
 wire \clk[22] ;
 wire \clk[230] ;
 wire \clk[231] ;
 wire \clk[232] ;
 wire \clk[233] ;
 wire \clk[234] ;
 wire \clk[235] ;
 wire \clk[236] ;
 wire \clk[237] ;
 wire \clk[238] ;
 wire \clk[239] ;
 wire \clk[23] ;
 wire \clk[240] ;
 wire \clk[241] ;
 wire \clk[242] ;
 wire \clk[243] ;
 wire \clk[244] ;
 wire \clk[245] ;
 wire \clk[246] ;
 wire \clk[247] ;
 wire \clk[248] ;
 wire \clk[249] ;
 wire \clk[24] ;
 wire \clk[250] ;
 wire \clk[251] ;
 wire \clk[252] ;
 wire \clk[253] ;
 wire \clk[254] ;
 wire \clk[255] ;
 wire \clk[256] ;
 wire \clk[257] ;
 wire \clk[258] ;
 wire \clk[259] ;
 wire \clk[25] ;
 wire \clk[260] ;
 wire \clk[261] ;
 wire \clk[262] ;
 wire \clk[263] ;
 wire \clk[264] ;
 wire \clk[265] ;
 wire \clk[266] ;
 wire \clk[267] ;
 wire \clk[268] ;
 wire \clk[269] ;
 wire \clk[26] ;
 wire \clk[270] ;
 wire \clk[271] ;
 wire \clk[272] ;
 wire \clk[273] ;
 wire \clk[274] ;
 wire \clk[275] ;
 wire \clk[276] ;
 wire \clk[277] ;
 wire \clk[278] ;
 wire \clk[279] ;
 wire \clk[27] ;
 wire \clk[280] ;
 wire \clk[281] ;
 wire \clk[282] ;
 wire \clk[283] ;
 wire \clk[284] ;
 wire \clk[285] ;
 wire \clk[286] ;
 wire \clk[287] ;
 wire \clk[288] ;
 wire \clk[289] ;
 wire \clk[28] ;
 wire \clk[290] ;
 wire \clk[291] ;
 wire \clk[292] ;
 wire \clk[293] ;
 wire \clk[294] ;
 wire \clk[295] ;
 wire \clk[296] ;
 wire \clk[297] ;
 wire \clk[298] ;
 wire \clk[299] ;
 wire \clk[29] ;
 wire \clk[2] ;
 wire \clk[300] ;
 wire \clk[301] ;
 wire \clk[302] ;
 wire \clk[303] ;
 wire \clk[304] ;
 wire \clk[305] ;
 wire \clk[306] ;
 wire \clk[307] ;
 wire \clk[308] ;
 wire \clk[309] ;
 wire \clk[30] ;
 wire \clk[310] ;
 wire \clk[311] ;
 wire \clk[312] ;
 wire \clk[313] ;
 wire \clk[314] ;
 wire \clk[315] ;
 wire \clk[316] ;
 wire \clk[317] ;
 wire \clk[318] ;
 wire \clk[319] ;
 wire \clk[31] ;
 wire \clk[320] ;
 wire \clk[321] ;
 wire \clk[322] ;
 wire \clk[323] ;
 wire \clk[324] ;
 wire \clk[325] ;
 wire \clk[326] ;
 wire \clk[327] ;
 wire \clk[328] ;
 wire \clk[329] ;
 wire \clk[32] ;
 wire \clk[330] ;
 wire \clk[331] ;
 wire \clk[332] ;
 wire \clk[333] ;
 wire \clk[334] ;
 wire \clk[335] ;
 wire \clk[336] ;
 wire \clk[337] ;
 wire \clk[338] ;
 wire \clk[339] ;
 wire \clk[33] ;
 wire \clk[340] ;
 wire \clk[341] ;
 wire \clk[342] ;
 wire \clk[343] ;
 wire \clk[344] ;
 wire \clk[345] ;
 wire \clk[346] ;
 wire \clk[347] ;
 wire \clk[348] ;
 wire \clk[349] ;
 wire \clk[34] ;
 wire \clk[350] ;
 wire \clk[351] ;
 wire \clk[352] ;
 wire \clk[353] ;
 wire \clk[354] ;
 wire \clk[355] ;
 wire \clk[356] ;
 wire \clk[357] ;
 wire \clk[358] ;
 wire \clk[359] ;
 wire \clk[35] ;
 wire \clk[360] ;
 wire \clk[361] ;
 wire \clk[362] ;
 wire \clk[363] ;
 wire \clk[364] ;
 wire \clk[365] ;
 wire \clk[366] ;
 wire \clk[367] ;
 wire \clk[368] ;
 wire \clk[369] ;
 wire \clk[36] ;
 wire \clk[370] ;
 wire \clk[371] ;
 wire \clk[372] ;
 wire \clk[373] ;
 wire \clk[374] ;
 wire \clk[375] ;
 wire \clk[376] ;
 wire \clk[377] ;
 wire \clk[378] ;
 wire \clk[379] ;
 wire \clk[37] ;
 wire \clk[380] ;
 wire \clk[381] ;
 wire \clk[382] ;
 wire \clk[383] ;
 wire \clk[384] ;
 wire \clk[385] ;
 wire \clk[386] ;
 wire \clk[387] ;
 wire \clk[388] ;
 wire \clk[389] ;
 wire \clk[38] ;
 wire \clk[390] ;
 wire \clk[391] ;
 wire \clk[392] ;
 wire \clk[393] ;
 wire \clk[394] ;
 wire \clk[395] ;
 wire \clk[396] ;
 wire \clk[397] ;
 wire \clk[398] ;
 wire \clk[399] ;
 wire \clk[39] ;
 wire \clk[3] ;
 wire \clk[400] ;
 wire \clk[401] ;
 wire \clk[402] ;
 wire \clk[403] ;
 wire \clk[404] ;
 wire \clk[405] ;
 wire \clk[406] ;
 wire \clk[407] ;
 wire \clk[408] ;
 wire \clk[409] ;
 wire \clk[40] ;
 wire \clk[410] ;
 wire \clk[411] ;
 wire \clk[412] ;
 wire \clk[413] ;
 wire \clk[414] ;
 wire \clk[415] ;
 wire \clk[416] ;
 wire \clk[417] ;
 wire \clk[418] ;
 wire \clk[419] ;
 wire \clk[41] ;
 wire \clk[420] ;
 wire \clk[421] ;
 wire \clk[422] ;
 wire \clk[423] ;
 wire \clk[424] ;
 wire \clk[425] ;
 wire \clk[426] ;
 wire \clk[427] ;
 wire \clk[428] ;
 wire \clk[429] ;
 wire \clk[42] ;
 wire \clk[430] ;
 wire \clk[431] ;
 wire \clk[432] ;
 wire \clk[433] ;
 wire \clk[434] ;
 wire \clk[435] ;
 wire \clk[436] ;
 wire \clk[437] ;
 wire \clk[438] ;
 wire \clk[439] ;
 wire \clk[43] ;
 wire \clk[440] ;
 wire \clk[441] ;
 wire \clk[442] ;
 wire \clk[443] ;
 wire \clk[444] ;
 wire \clk[445] ;
 wire \clk[446] ;
 wire \clk[447] ;
 wire \clk[448] ;
 wire \clk[449] ;
 wire \clk[44] ;
 wire \clk[450] ;
 wire \clk[451] ;
 wire \clk[452] ;
 wire \clk[453] ;
 wire \clk[454] ;
 wire \clk[455] ;
 wire \clk[456] ;
 wire \clk[457] ;
 wire \clk[458] ;
 wire \clk[459] ;
 wire \clk[45] ;
 wire \clk[460] ;
 wire \clk[461] ;
 wire \clk[462] ;
 wire \clk[463] ;
 wire \clk[464] ;
 wire \clk[465] ;
 wire \clk[466] ;
 wire \clk[467] ;
 wire \clk[468] ;
 wire \clk[469] ;
 wire \clk[46] ;
 wire \clk[470] ;
 wire \clk[471] ;
 wire \clk[472] ;
 wire \clk[473] ;
 wire \clk[474] ;
 wire \clk[475] ;
 wire \clk[476] ;
 wire \clk[477] ;
 wire \clk[478] ;
 wire \clk[479] ;
 wire \clk[47] ;
 wire \clk[480] ;
 wire \clk[481] ;
 wire \clk[482] ;
 wire \clk[483] ;
 wire \clk[484] ;
 wire \clk[485] ;
 wire \clk[486] ;
 wire \clk[487] ;
 wire \clk[488] ;
 wire \clk[489] ;
 wire \clk[48] ;
 wire \clk[490] ;
 wire \clk[491] ;
 wire \clk[492] ;
 wire \clk[493] ;
 wire \clk[494] ;
 wire \clk[495] ;
 wire \clk[496] ;
 wire \clk[497] ;
 wire \clk[498] ;
 wire \clk[49] ;
 wire \clk[4] ;
 wire \clk[50] ;
 wire \clk[51] ;
 wire \clk[52] ;
 wire \clk[53] ;
 wire \clk[54] ;
 wire \clk[55] ;
 wire \clk[56] ;
 wire \clk[57] ;
 wire \clk[58] ;
 wire \clk[59] ;
 wire \clk[5] ;
 wire \clk[60] ;
 wire \clk[61] ;
 wire \clk[62] ;
 wire \clk[63] ;
 wire \clk[64] ;
 wire \clk[65] ;
 wire \clk[66] ;
 wire \clk[67] ;
 wire \clk[68] ;
 wire \clk[69] ;
 wire \clk[6] ;
 wire \clk[70] ;
 wire \clk[71] ;
 wire \clk[72] ;
 wire \clk[73] ;
 wire \clk[74] ;
 wire \clk[75] ;
 wire \clk[76] ;
 wire \clk[77] ;
 wire \clk[78] ;
 wire \clk[79] ;
 wire \clk[7] ;
 wire \clk[80] ;
 wire \clk[81] ;
 wire \clk[82] ;
 wire \clk[83] ;
 wire \clk[84] ;
 wire \clk[85] ;
 wire \clk[86] ;
 wire \clk[87] ;
 wire \clk[88] ;
 wire \clk[89] ;
 wire \clk[8] ;
 wire \clk[90] ;
 wire \clk[91] ;
 wire \clk[92] ;
 wire \clk[93] ;
 wire \clk[94] ;
 wire \clk[95] ;
 wire \clk[96] ;
 wire \clk[97] ;
 wire \clk[98] ;
 wire \clk[99] ;
 wire \clk[9] ;
 wire \data[0] ;
 wire \data[100] ;
 wire \data[101] ;
 wire \data[102] ;
 wire \data[103] ;
 wire \data[104] ;
 wire \data[105] ;
 wire \data[106] ;
 wire \data[107] ;
 wire \data[108] ;
 wire \data[109] ;
 wire \data[10] ;
 wire \data[110] ;
 wire \data[111] ;
 wire \data[112] ;
 wire \data[113] ;
 wire \data[114] ;
 wire \data[115] ;
 wire \data[116] ;
 wire \data[117] ;
 wire \data[118] ;
 wire \data[119] ;
 wire \data[11] ;
 wire \data[120] ;
 wire \data[121] ;
 wire \data[122] ;
 wire \data[123] ;
 wire \data[124] ;
 wire \data[125] ;
 wire \data[126] ;
 wire \data[127] ;
 wire \data[128] ;
 wire \data[129] ;
 wire \data[12] ;
 wire \data[130] ;
 wire \data[131] ;
 wire \data[132] ;
 wire \data[133] ;
 wire \data[134] ;
 wire \data[135] ;
 wire \data[136] ;
 wire \data[137] ;
 wire \data[138] ;
 wire \data[139] ;
 wire \data[13] ;
 wire \data[140] ;
 wire \data[141] ;
 wire \data[142] ;
 wire \data[143] ;
 wire \data[144] ;
 wire \data[145] ;
 wire \data[146] ;
 wire \data[147] ;
 wire \data[148] ;
 wire \data[149] ;
 wire \data[14] ;
 wire \data[150] ;
 wire \data[151] ;
 wire \data[152] ;
 wire \data[153] ;
 wire \data[154] ;
 wire \data[155] ;
 wire \data[156] ;
 wire \data[157] ;
 wire \data[158] ;
 wire \data[159] ;
 wire \data[15] ;
 wire \data[160] ;
 wire \data[161] ;
 wire \data[162] ;
 wire \data[163] ;
 wire \data[164] ;
 wire \data[165] ;
 wire \data[166] ;
 wire \data[167] ;
 wire \data[168] ;
 wire \data[169] ;
 wire \data[16] ;
 wire \data[170] ;
 wire \data[171] ;
 wire \data[172] ;
 wire \data[173] ;
 wire \data[174] ;
 wire \data[175] ;
 wire \data[176] ;
 wire \data[177] ;
 wire \data[178] ;
 wire \data[179] ;
 wire \data[17] ;
 wire \data[180] ;
 wire \data[181] ;
 wire \data[182] ;
 wire \data[183] ;
 wire \data[184] ;
 wire \data[185] ;
 wire \data[186] ;
 wire \data[187] ;
 wire \data[188] ;
 wire \data[189] ;
 wire \data[18] ;
 wire \data[190] ;
 wire \data[191] ;
 wire \data[192] ;
 wire \data[193] ;
 wire \data[194] ;
 wire \data[195] ;
 wire \data[196] ;
 wire \data[197] ;
 wire \data[198] ;
 wire \data[199] ;
 wire \data[19] ;
 wire \data[1] ;
 wire \data[200] ;
 wire \data[201] ;
 wire \data[202] ;
 wire \data[203] ;
 wire \data[204] ;
 wire \data[205] ;
 wire \data[206] ;
 wire \data[207] ;
 wire \data[208] ;
 wire \data[209] ;
 wire \data[20] ;
 wire \data[210] ;
 wire \data[211] ;
 wire \data[212] ;
 wire \data[213] ;
 wire \data[214] ;
 wire \data[215] ;
 wire \data[216] ;
 wire \data[217] ;
 wire \data[218] ;
 wire \data[219] ;
 wire \data[21] ;
 wire \data[220] ;
 wire \data[221] ;
 wire \data[222] ;
 wire \data[223] ;
 wire \data[224] ;
 wire \data[225] ;
 wire \data[226] ;
 wire \data[227] ;
 wire \data[228] ;
 wire \data[229] ;
 wire \data[22] ;
 wire \data[230] ;
 wire \data[231] ;
 wire \data[232] ;
 wire \data[233] ;
 wire \data[234] ;
 wire \data[235] ;
 wire \data[236] ;
 wire \data[237] ;
 wire \data[238] ;
 wire \data[239] ;
 wire \data[23] ;
 wire \data[240] ;
 wire \data[241] ;
 wire \data[242] ;
 wire \data[243] ;
 wire \data[244] ;
 wire \data[245] ;
 wire \data[246] ;
 wire \data[247] ;
 wire \data[248] ;
 wire \data[249] ;
 wire \data[24] ;
 wire \data[250] ;
 wire \data[251] ;
 wire \data[252] ;
 wire \data[253] ;
 wire \data[254] ;
 wire \data[255] ;
 wire \data[256] ;
 wire \data[257] ;
 wire \data[258] ;
 wire \data[259] ;
 wire \data[25] ;
 wire \data[260] ;
 wire \data[261] ;
 wire \data[262] ;
 wire \data[263] ;
 wire \data[264] ;
 wire \data[265] ;
 wire \data[266] ;
 wire \data[267] ;
 wire \data[268] ;
 wire \data[269] ;
 wire \data[26] ;
 wire \data[270] ;
 wire \data[271] ;
 wire \data[272] ;
 wire \data[273] ;
 wire \data[274] ;
 wire \data[275] ;
 wire \data[276] ;
 wire \data[277] ;
 wire \data[278] ;
 wire \data[279] ;
 wire \data[27] ;
 wire \data[280] ;
 wire \data[281] ;
 wire \data[282] ;
 wire \data[283] ;
 wire \data[284] ;
 wire \data[285] ;
 wire \data[286] ;
 wire \data[287] ;
 wire \data[288] ;
 wire \data[289] ;
 wire \data[28] ;
 wire \data[290] ;
 wire \data[291] ;
 wire \data[292] ;
 wire \data[293] ;
 wire \data[294] ;
 wire \data[295] ;
 wire \data[296] ;
 wire \data[297] ;
 wire \data[298] ;
 wire \data[299] ;
 wire \data[29] ;
 wire \data[2] ;
 wire \data[300] ;
 wire \data[301] ;
 wire \data[302] ;
 wire \data[303] ;
 wire \data[304] ;
 wire \data[305] ;
 wire \data[306] ;
 wire \data[307] ;
 wire \data[308] ;
 wire \data[309] ;
 wire \data[30] ;
 wire \data[310] ;
 wire \data[311] ;
 wire \data[312] ;
 wire \data[313] ;
 wire \data[314] ;
 wire \data[315] ;
 wire \data[316] ;
 wire \data[317] ;
 wire \data[318] ;
 wire \data[319] ;
 wire \data[31] ;
 wire \data[320] ;
 wire \data[321] ;
 wire \data[322] ;
 wire \data[323] ;
 wire \data[324] ;
 wire \data[325] ;
 wire \data[326] ;
 wire \data[327] ;
 wire \data[328] ;
 wire \data[329] ;
 wire \data[32] ;
 wire \data[330] ;
 wire \data[331] ;
 wire \data[332] ;
 wire \data[333] ;
 wire \data[334] ;
 wire \data[335] ;
 wire \data[336] ;
 wire \data[337] ;
 wire \data[338] ;
 wire \data[339] ;
 wire \data[33] ;
 wire \data[340] ;
 wire \data[341] ;
 wire \data[342] ;
 wire \data[343] ;
 wire \data[344] ;
 wire \data[345] ;
 wire \data[346] ;
 wire \data[347] ;
 wire \data[348] ;
 wire \data[349] ;
 wire \data[34] ;
 wire \data[350] ;
 wire \data[351] ;
 wire \data[352] ;
 wire \data[353] ;
 wire \data[354] ;
 wire \data[355] ;
 wire \data[356] ;
 wire \data[357] ;
 wire \data[358] ;
 wire \data[359] ;
 wire \data[35] ;
 wire \data[360] ;
 wire \data[361] ;
 wire \data[362] ;
 wire \data[363] ;
 wire \data[364] ;
 wire \data[365] ;
 wire \data[366] ;
 wire \data[367] ;
 wire \data[368] ;
 wire \data[369] ;
 wire \data[36] ;
 wire \data[370] ;
 wire \data[371] ;
 wire \data[372] ;
 wire \data[373] ;
 wire \data[374] ;
 wire \data[375] ;
 wire \data[376] ;
 wire \data[377] ;
 wire \data[378] ;
 wire \data[379] ;
 wire \data[37] ;
 wire \data[380] ;
 wire \data[381] ;
 wire \data[382] ;
 wire \data[383] ;
 wire \data[384] ;
 wire \data[385] ;
 wire \data[386] ;
 wire \data[387] ;
 wire \data[388] ;
 wire \data[389] ;
 wire \data[38] ;
 wire \data[390] ;
 wire \data[391] ;
 wire \data[392] ;
 wire \data[393] ;
 wire \data[394] ;
 wire \data[395] ;
 wire \data[396] ;
 wire \data[397] ;
 wire \data[398] ;
 wire \data[399] ;
 wire \data[39] ;
 wire \data[3] ;
 wire \data[400] ;
 wire \data[401] ;
 wire \data[402] ;
 wire \data[403] ;
 wire \data[404] ;
 wire \data[405] ;
 wire \data[406] ;
 wire \data[407] ;
 wire \data[408] ;
 wire \data[409] ;
 wire \data[40] ;
 wire \data[410] ;
 wire \data[411] ;
 wire \data[412] ;
 wire \data[413] ;
 wire \data[414] ;
 wire \data[415] ;
 wire \data[416] ;
 wire \data[417] ;
 wire \data[418] ;
 wire \data[419] ;
 wire \data[41] ;
 wire \data[420] ;
 wire \data[421] ;
 wire \data[422] ;
 wire \data[423] ;
 wire \data[424] ;
 wire \data[425] ;
 wire \data[426] ;
 wire \data[427] ;
 wire \data[428] ;
 wire \data[429] ;
 wire \data[42] ;
 wire \data[430] ;
 wire \data[431] ;
 wire \data[432] ;
 wire \data[433] ;
 wire \data[434] ;
 wire \data[435] ;
 wire \data[436] ;
 wire \data[437] ;
 wire \data[438] ;
 wire \data[439] ;
 wire \data[43] ;
 wire \data[440] ;
 wire \data[441] ;
 wire \data[442] ;
 wire \data[443] ;
 wire \data[444] ;
 wire \data[445] ;
 wire \data[446] ;
 wire \data[447] ;
 wire \data[448] ;
 wire \data[449] ;
 wire \data[44] ;
 wire \data[450] ;
 wire \data[451] ;
 wire \data[452] ;
 wire \data[453] ;
 wire \data[454] ;
 wire \data[455] ;
 wire \data[456] ;
 wire \data[457] ;
 wire \data[458] ;
 wire \data[459] ;
 wire \data[45] ;
 wire \data[460] ;
 wire \data[461] ;
 wire \data[462] ;
 wire \data[463] ;
 wire \data[464] ;
 wire \data[465] ;
 wire \data[466] ;
 wire \data[467] ;
 wire \data[468] ;
 wire \data[469] ;
 wire \data[46] ;
 wire \data[470] ;
 wire \data[471] ;
 wire \data[472] ;
 wire \data[473] ;
 wire \data[474] ;
 wire \data[475] ;
 wire \data[476] ;
 wire \data[477] ;
 wire \data[478] ;
 wire \data[479] ;
 wire \data[47] ;
 wire \data[480] ;
 wire \data[481] ;
 wire \data[482] ;
 wire \data[483] ;
 wire \data[484] ;
 wire \data[485] ;
 wire \data[486] ;
 wire \data[487] ;
 wire \data[488] ;
 wire \data[489] ;
 wire \data[48] ;
 wire \data[490] ;
 wire \data[491] ;
 wire \data[492] ;
 wire \data[493] ;
 wire \data[494] ;
 wire \data[495] ;
 wire \data[496] ;
 wire \data[497] ;
 wire \data[498] ;
 wire \data[49] ;
 wire \data[4] ;
 wire \data[50] ;
 wire \data[51] ;
 wire \data[52] ;
 wire \data[53] ;
 wire \data[54] ;
 wire \data[55] ;
 wire \data[56] ;
 wire \data[57] ;
 wire \data[58] ;
 wire \data[59] ;
 wire \data[5] ;
 wire \data[60] ;
 wire \data[61] ;
 wire \data[62] ;
 wire \data[63] ;
 wire \data[64] ;
 wire \data[65] ;
 wire \data[66] ;
 wire \data[67] ;
 wire \data[68] ;
 wire \data[69] ;
 wire \data[6] ;
 wire \data[70] ;
 wire \data[71] ;
 wire \data[72] ;
 wire \data[73] ;
 wire \data[74] ;
 wire \data[75] ;
 wire \data[76] ;
 wire \data[77] ;
 wire \data[78] ;
 wire \data[79] ;
 wire \data[7] ;
 wire \data[80] ;
 wire \data[81] ;
 wire \data[82] ;
 wire \data[83] ;
 wire \data[84] ;
 wire \data[85] ;
 wire \data[86] ;
 wire \data[87] ;
 wire \data[88] ;
 wire \data[89] ;
 wire \data[8] ;
 wire \data[90] ;
 wire \data[91] ;
 wire \data[92] ;
 wire \data[93] ;
 wire \data[94] ;
 wire \data[95] ;
 wire \data[96] ;
 wire \data[97] ;
 wire \data[98] ;
 wire \data[99] ;
 wire \data[9] ;
 wire \latch[0] ;
 wire \latch[100] ;
 wire \latch[101] ;
 wire \latch[102] ;
 wire \latch[103] ;
 wire \latch[104] ;
 wire \latch[105] ;
 wire \latch[106] ;
 wire \latch[107] ;
 wire \latch[108] ;
 wire \latch[109] ;
 wire \latch[10] ;
 wire \latch[110] ;
 wire \latch[111] ;
 wire \latch[112] ;
 wire \latch[113] ;
 wire \latch[114] ;
 wire \latch[115] ;
 wire \latch[116] ;
 wire \latch[117] ;
 wire \latch[118] ;
 wire \latch[119] ;
 wire \latch[11] ;
 wire \latch[120] ;
 wire \latch[121] ;
 wire \latch[122] ;
 wire \latch[123] ;
 wire \latch[124] ;
 wire \latch[125] ;
 wire \latch[126] ;
 wire \latch[127] ;
 wire \latch[128] ;
 wire \latch[129] ;
 wire \latch[12] ;
 wire \latch[130] ;
 wire \latch[131] ;
 wire \latch[132] ;
 wire \latch[133] ;
 wire \latch[134] ;
 wire \latch[135] ;
 wire \latch[136] ;
 wire \latch[137] ;
 wire \latch[138] ;
 wire \latch[139] ;
 wire \latch[13] ;
 wire \latch[140] ;
 wire \latch[141] ;
 wire \latch[142] ;
 wire \latch[143] ;
 wire \latch[144] ;
 wire \latch[145] ;
 wire \latch[146] ;
 wire \latch[147] ;
 wire \latch[148] ;
 wire \latch[149] ;
 wire \latch[14] ;
 wire \latch[150] ;
 wire \latch[151] ;
 wire \latch[152] ;
 wire \latch[153] ;
 wire \latch[154] ;
 wire \latch[155] ;
 wire \latch[156] ;
 wire \latch[157] ;
 wire \latch[158] ;
 wire \latch[159] ;
 wire \latch[15] ;
 wire \latch[160] ;
 wire \latch[161] ;
 wire \latch[162] ;
 wire \latch[163] ;
 wire \latch[164] ;
 wire \latch[165] ;
 wire \latch[166] ;
 wire \latch[167] ;
 wire \latch[168] ;
 wire \latch[169] ;
 wire \latch[16] ;
 wire \latch[170] ;
 wire \latch[171] ;
 wire \latch[172] ;
 wire \latch[173] ;
 wire \latch[174] ;
 wire \latch[175] ;
 wire \latch[176] ;
 wire \latch[177] ;
 wire \latch[178] ;
 wire \latch[179] ;
 wire \latch[17] ;
 wire \latch[180] ;
 wire \latch[181] ;
 wire \latch[182] ;
 wire \latch[183] ;
 wire \latch[184] ;
 wire \latch[185] ;
 wire \latch[186] ;
 wire \latch[187] ;
 wire \latch[188] ;
 wire \latch[189] ;
 wire \latch[18] ;
 wire \latch[190] ;
 wire \latch[191] ;
 wire \latch[192] ;
 wire \latch[193] ;
 wire \latch[194] ;
 wire \latch[195] ;
 wire \latch[196] ;
 wire \latch[197] ;
 wire \latch[198] ;
 wire \latch[199] ;
 wire \latch[19] ;
 wire \latch[1] ;
 wire \latch[200] ;
 wire \latch[201] ;
 wire \latch[202] ;
 wire \latch[203] ;
 wire \latch[204] ;
 wire \latch[205] ;
 wire \latch[206] ;
 wire \latch[207] ;
 wire \latch[208] ;
 wire \latch[209] ;
 wire \latch[20] ;
 wire \latch[210] ;
 wire \latch[211] ;
 wire \latch[212] ;
 wire \latch[213] ;
 wire \latch[214] ;
 wire \latch[215] ;
 wire \latch[216] ;
 wire \latch[217] ;
 wire \latch[218] ;
 wire \latch[219] ;
 wire \latch[21] ;
 wire \latch[220] ;
 wire \latch[221] ;
 wire \latch[222] ;
 wire \latch[223] ;
 wire \latch[224] ;
 wire \latch[225] ;
 wire \latch[226] ;
 wire \latch[227] ;
 wire \latch[228] ;
 wire \latch[229] ;
 wire \latch[22] ;
 wire \latch[230] ;
 wire \latch[231] ;
 wire \latch[232] ;
 wire \latch[233] ;
 wire \latch[234] ;
 wire \latch[235] ;
 wire \latch[236] ;
 wire \latch[237] ;
 wire \latch[238] ;
 wire \latch[239] ;
 wire \latch[23] ;
 wire \latch[240] ;
 wire \latch[241] ;
 wire \latch[242] ;
 wire \latch[243] ;
 wire \latch[244] ;
 wire \latch[245] ;
 wire \latch[246] ;
 wire \latch[247] ;
 wire \latch[248] ;
 wire \latch[249] ;
 wire \latch[24] ;
 wire \latch[250] ;
 wire \latch[251] ;
 wire \latch[252] ;
 wire \latch[253] ;
 wire \latch[254] ;
 wire \latch[255] ;
 wire \latch[256] ;
 wire \latch[257] ;
 wire \latch[258] ;
 wire \latch[259] ;
 wire \latch[25] ;
 wire \latch[260] ;
 wire \latch[261] ;
 wire \latch[262] ;
 wire \latch[263] ;
 wire \latch[264] ;
 wire \latch[265] ;
 wire \latch[266] ;
 wire \latch[267] ;
 wire \latch[268] ;
 wire \latch[269] ;
 wire \latch[26] ;
 wire \latch[270] ;
 wire \latch[271] ;
 wire \latch[272] ;
 wire \latch[273] ;
 wire \latch[274] ;
 wire \latch[275] ;
 wire \latch[276] ;
 wire \latch[277] ;
 wire \latch[278] ;
 wire \latch[279] ;
 wire \latch[27] ;
 wire \latch[280] ;
 wire \latch[281] ;
 wire \latch[282] ;
 wire \latch[283] ;
 wire \latch[284] ;
 wire \latch[285] ;
 wire \latch[286] ;
 wire \latch[287] ;
 wire \latch[288] ;
 wire \latch[289] ;
 wire \latch[28] ;
 wire \latch[290] ;
 wire \latch[291] ;
 wire \latch[292] ;
 wire \latch[293] ;
 wire \latch[294] ;
 wire \latch[295] ;
 wire \latch[296] ;
 wire \latch[297] ;
 wire \latch[298] ;
 wire \latch[299] ;
 wire \latch[29] ;
 wire \latch[2] ;
 wire \latch[300] ;
 wire \latch[301] ;
 wire \latch[302] ;
 wire \latch[303] ;
 wire \latch[304] ;
 wire \latch[305] ;
 wire \latch[306] ;
 wire \latch[307] ;
 wire \latch[308] ;
 wire \latch[309] ;
 wire \latch[30] ;
 wire \latch[310] ;
 wire \latch[311] ;
 wire \latch[312] ;
 wire \latch[313] ;
 wire \latch[314] ;
 wire \latch[315] ;
 wire \latch[316] ;
 wire \latch[317] ;
 wire \latch[318] ;
 wire \latch[319] ;
 wire \latch[31] ;
 wire \latch[320] ;
 wire \latch[321] ;
 wire \latch[322] ;
 wire \latch[323] ;
 wire \latch[324] ;
 wire \latch[325] ;
 wire \latch[326] ;
 wire \latch[327] ;
 wire \latch[328] ;
 wire \latch[329] ;
 wire \latch[32] ;
 wire \latch[330] ;
 wire \latch[331] ;
 wire \latch[332] ;
 wire \latch[333] ;
 wire \latch[334] ;
 wire \latch[335] ;
 wire \latch[336] ;
 wire \latch[337] ;
 wire \latch[338] ;
 wire \latch[339] ;
 wire \latch[33] ;
 wire \latch[340] ;
 wire \latch[341] ;
 wire \latch[342] ;
 wire \latch[343] ;
 wire \latch[344] ;
 wire \latch[345] ;
 wire \latch[346] ;
 wire \latch[347] ;
 wire \latch[348] ;
 wire \latch[349] ;
 wire \latch[34] ;
 wire \latch[350] ;
 wire \latch[351] ;
 wire \latch[352] ;
 wire \latch[353] ;
 wire \latch[354] ;
 wire \latch[355] ;
 wire \latch[356] ;
 wire \latch[357] ;
 wire \latch[358] ;
 wire \latch[359] ;
 wire \latch[35] ;
 wire \latch[360] ;
 wire \latch[361] ;
 wire \latch[362] ;
 wire \latch[363] ;
 wire \latch[364] ;
 wire \latch[365] ;
 wire \latch[366] ;
 wire \latch[367] ;
 wire \latch[368] ;
 wire \latch[369] ;
 wire \latch[36] ;
 wire \latch[370] ;
 wire \latch[371] ;
 wire \latch[372] ;
 wire \latch[373] ;
 wire \latch[374] ;
 wire \latch[375] ;
 wire \latch[376] ;
 wire \latch[377] ;
 wire \latch[378] ;
 wire \latch[379] ;
 wire \latch[37] ;
 wire \latch[380] ;
 wire \latch[381] ;
 wire \latch[382] ;
 wire \latch[383] ;
 wire \latch[384] ;
 wire \latch[385] ;
 wire \latch[386] ;
 wire \latch[387] ;
 wire \latch[388] ;
 wire \latch[389] ;
 wire \latch[38] ;
 wire \latch[390] ;
 wire \latch[391] ;
 wire \latch[392] ;
 wire \latch[393] ;
 wire \latch[394] ;
 wire \latch[395] ;
 wire \latch[396] ;
 wire \latch[397] ;
 wire \latch[398] ;
 wire \latch[399] ;
 wire \latch[39] ;
 wire \latch[3] ;
 wire \latch[400] ;
 wire \latch[401] ;
 wire \latch[402] ;
 wire \latch[403] ;
 wire \latch[404] ;
 wire \latch[405] ;
 wire \latch[406] ;
 wire \latch[407] ;
 wire \latch[408] ;
 wire \latch[409] ;
 wire \latch[40] ;
 wire \latch[410] ;
 wire \latch[411] ;
 wire \latch[412] ;
 wire \latch[413] ;
 wire \latch[414] ;
 wire \latch[415] ;
 wire \latch[416] ;
 wire \latch[417] ;
 wire \latch[418] ;
 wire \latch[419] ;
 wire \latch[41] ;
 wire \latch[420] ;
 wire \latch[421] ;
 wire \latch[422] ;
 wire \latch[423] ;
 wire \latch[424] ;
 wire \latch[425] ;
 wire \latch[426] ;
 wire \latch[427] ;
 wire \latch[428] ;
 wire \latch[429] ;
 wire \latch[42] ;
 wire \latch[430] ;
 wire \latch[431] ;
 wire \latch[432] ;
 wire \latch[433] ;
 wire \latch[434] ;
 wire \latch[435] ;
 wire \latch[436] ;
 wire \latch[437] ;
 wire \latch[438] ;
 wire \latch[439] ;
 wire \latch[43] ;
 wire \latch[440] ;
 wire \latch[441] ;
 wire \latch[442] ;
 wire \latch[443] ;
 wire \latch[444] ;
 wire \latch[445] ;
 wire \latch[446] ;
 wire \latch[447] ;
 wire \latch[448] ;
 wire \latch[449] ;
 wire \latch[44] ;
 wire \latch[450] ;
 wire \latch[451] ;
 wire \latch[452] ;
 wire \latch[453] ;
 wire \latch[454] ;
 wire \latch[455] ;
 wire \latch[456] ;
 wire \latch[457] ;
 wire \latch[458] ;
 wire \latch[459] ;
 wire \latch[45] ;
 wire \latch[460] ;
 wire \latch[461] ;
 wire \latch[462] ;
 wire \latch[463] ;
 wire \latch[464] ;
 wire \latch[465] ;
 wire \latch[466] ;
 wire \latch[467] ;
 wire \latch[468] ;
 wire \latch[469] ;
 wire \latch[46] ;
 wire \latch[470] ;
 wire \latch[471] ;
 wire \latch[472] ;
 wire \latch[473] ;
 wire \latch[474] ;
 wire \latch[475] ;
 wire \latch[476] ;
 wire \latch[477] ;
 wire \latch[478] ;
 wire \latch[479] ;
 wire \latch[47] ;
 wire \latch[480] ;
 wire \latch[481] ;
 wire \latch[482] ;
 wire \latch[483] ;
 wire \latch[484] ;
 wire \latch[485] ;
 wire \latch[486] ;
 wire \latch[487] ;
 wire \latch[488] ;
 wire \latch[489] ;
 wire \latch[48] ;
 wire \latch[490] ;
 wire \latch[491] ;
 wire \latch[492] ;
 wire \latch[493] ;
 wire \latch[494] ;
 wire \latch[495] ;
 wire \latch[496] ;
 wire \latch[497] ;
 wire \latch[498] ;
 wire \latch[49] ;
 wire \latch[4] ;
 wire \latch[50] ;
 wire \latch[51] ;
 wire \latch[52] ;
 wire \latch[53] ;
 wire \latch[54] ;
 wire \latch[55] ;
 wire \latch[56] ;
 wire \latch[57] ;
 wire \latch[58] ;
 wire \latch[59] ;
 wire \latch[5] ;
 wire \latch[60] ;
 wire \latch[61] ;
 wire \latch[62] ;
 wire \latch[63] ;
 wire \latch[64] ;
 wire \latch[65] ;
 wire \latch[66] ;
 wire \latch[67] ;
 wire \latch[68] ;
 wire \latch[69] ;
 wire \latch[6] ;
 wire \latch[70] ;
 wire \latch[71] ;
 wire \latch[72] ;
 wire \latch[73] ;
 wire \latch[74] ;
 wire \latch[75] ;
 wire \latch[76] ;
 wire \latch[77] ;
 wire \latch[78] ;
 wire \latch[79] ;
 wire \latch[7] ;
 wire \latch[80] ;
 wire \latch[81] ;
 wire \latch[82] ;
 wire \latch[83] ;
 wire \latch[84] ;
 wire \latch[85] ;
 wire \latch[86] ;
 wire \latch[87] ;
 wire \latch[88] ;
 wire \latch[89] ;
 wire \latch[8] ;
 wire \latch[90] ;
 wire \latch[91] ;
 wire \latch[92] ;
 wire \latch[93] ;
 wire \latch[94] ;
 wire \latch[95] ;
 wire \latch[96] ;
 wire \latch[97] ;
 wire \latch[98] ;
 wire \latch[99] ;
 wire \latch[9] ;
 wire \scan[0] ;
 wire \scan[100] ;
 wire \scan[101] ;
 wire \scan[102] ;
 wire \scan[103] ;
 wire \scan[104] ;
 wire \scan[105] ;
 wire \scan[106] ;
 wire \scan[107] ;
 wire \scan[108] ;
 wire \scan[109] ;
 wire \scan[10] ;
 wire \scan[110] ;
 wire \scan[111] ;
 wire \scan[112] ;
 wire \scan[113] ;
 wire \scan[114] ;
 wire \scan[115] ;
 wire \scan[116] ;
 wire \scan[117] ;
 wire \scan[118] ;
 wire \scan[119] ;
 wire \scan[11] ;
 wire \scan[120] ;
 wire \scan[121] ;
 wire \scan[122] ;
 wire \scan[123] ;
 wire \scan[124] ;
 wire \scan[125] ;
 wire \scan[126] ;
 wire \scan[127] ;
 wire \scan[128] ;
 wire \scan[129] ;
 wire \scan[12] ;
 wire \scan[130] ;
 wire \scan[131] ;
 wire \scan[132] ;
 wire \scan[133] ;
 wire \scan[134] ;
 wire \scan[135] ;
 wire \scan[136] ;
 wire \scan[137] ;
 wire \scan[138] ;
 wire \scan[139] ;
 wire \scan[13] ;
 wire \scan[140] ;
 wire \scan[141] ;
 wire \scan[142] ;
 wire \scan[143] ;
 wire \scan[144] ;
 wire \scan[145] ;
 wire \scan[146] ;
 wire \scan[147] ;
 wire \scan[148] ;
 wire \scan[149] ;
 wire \scan[14] ;
 wire \scan[150] ;
 wire \scan[151] ;
 wire \scan[152] ;
 wire \scan[153] ;
 wire \scan[154] ;
 wire \scan[155] ;
 wire \scan[156] ;
 wire \scan[157] ;
 wire \scan[158] ;
 wire \scan[159] ;
 wire \scan[15] ;
 wire \scan[160] ;
 wire \scan[161] ;
 wire \scan[162] ;
 wire \scan[163] ;
 wire \scan[164] ;
 wire \scan[165] ;
 wire \scan[166] ;
 wire \scan[167] ;
 wire \scan[168] ;
 wire \scan[169] ;
 wire \scan[16] ;
 wire \scan[170] ;
 wire \scan[171] ;
 wire \scan[172] ;
 wire \scan[173] ;
 wire \scan[174] ;
 wire \scan[175] ;
 wire \scan[176] ;
 wire \scan[177] ;
 wire \scan[178] ;
 wire \scan[179] ;
 wire \scan[17] ;
 wire \scan[180] ;
 wire \scan[181] ;
 wire \scan[182] ;
 wire \scan[183] ;
 wire \scan[184] ;
 wire \scan[185] ;
 wire \scan[186] ;
 wire \scan[187] ;
 wire \scan[188] ;
 wire \scan[189] ;
 wire \scan[18] ;
 wire \scan[190] ;
 wire \scan[191] ;
 wire \scan[192] ;
 wire \scan[193] ;
 wire \scan[194] ;
 wire \scan[195] ;
 wire \scan[196] ;
 wire \scan[197] ;
 wire \scan[198] ;
 wire \scan[199] ;
 wire \scan[19] ;
 wire \scan[1] ;
 wire \scan[200] ;
 wire \scan[201] ;
 wire \scan[202] ;
 wire \scan[203] ;
 wire \scan[204] ;
 wire \scan[205] ;
 wire \scan[206] ;
 wire \scan[207] ;
 wire \scan[208] ;
 wire \scan[209] ;
 wire \scan[20] ;
 wire \scan[210] ;
 wire \scan[211] ;
 wire \scan[212] ;
 wire \scan[213] ;
 wire \scan[214] ;
 wire \scan[215] ;
 wire \scan[216] ;
 wire \scan[217] ;
 wire \scan[218] ;
 wire \scan[219] ;
 wire \scan[21] ;
 wire \scan[220] ;
 wire \scan[221] ;
 wire \scan[222] ;
 wire \scan[223] ;
 wire \scan[224] ;
 wire \scan[225] ;
 wire \scan[226] ;
 wire \scan[227] ;
 wire \scan[228] ;
 wire \scan[229] ;
 wire \scan[22] ;
 wire \scan[230] ;
 wire \scan[231] ;
 wire \scan[232] ;
 wire \scan[233] ;
 wire \scan[234] ;
 wire \scan[235] ;
 wire \scan[236] ;
 wire \scan[237] ;
 wire \scan[238] ;
 wire \scan[239] ;
 wire \scan[23] ;
 wire \scan[240] ;
 wire \scan[241] ;
 wire \scan[242] ;
 wire \scan[243] ;
 wire \scan[244] ;
 wire \scan[245] ;
 wire \scan[246] ;
 wire \scan[247] ;
 wire \scan[248] ;
 wire \scan[249] ;
 wire \scan[24] ;
 wire \scan[250] ;
 wire \scan[251] ;
 wire \scan[252] ;
 wire \scan[253] ;
 wire \scan[254] ;
 wire \scan[255] ;
 wire \scan[256] ;
 wire \scan[257] ;
 wire \scan[258] ;
 wire \scan[259] ;
 wire \scan[25] ;
 wire \scan[260] ;
 wire \scan[261] ;
 wire \scan[262] ;
 wire \scan[263] ;
 wire \scan[264] ;
 wire \scan[265] ;
 wire \scan[266] ;
 wire \scan[267] ;
 wire \scan[268] ;
 wire \scan[269] ;
 wire \scan[26] ;
 wire \scan[270] ;
 wire \scan[271] ;
 wire \scan[272] ;
 wire \scan[273] ;
 wire \scan[274] ;
 wire \scan[275] ;
 wire \scan[276] ;
 wire \scan[277] ;
 wire \scan[278] ;
 wire \scan[279] ;
 wire \scan[27] ;
 wire \scan[280] ;
 wire \scan[281] ;
 wire \scan[282] ;
 wire \scan[283] ;
 wire \scan[284] ;
 wire \scan[285] ;
 wire \scan[286] ;
 wire \scan[287] ;
 wire \scan[288] ;
 wire \scan[289] ;
 wire \scan[28] ;
 wire \scan[290] ;
 wire \scan[291] ;
 wire \scan[292] ;
 wire \scan[293] ;
 wire \scan[294] ;
 wire \scan[295] ;
 wire \scan[296] ;
 wire \scan[297] ;
 wire \scan[298] ;
 wire \scan[299] ;
 wire \scan[29] ;
 wire \scan[2] ;
 wire \scan[300] ;
 wire \scan[301] ;
 wire \scan[302] ;
 wire \scan[303] ;
 wire \scan[304] ;
 wire \scan[305] ;
 wire \scan[306] ;
 wire \scan[307] ;
 wire \scan[308] ;
 wire \scan[309] ;
 wire \scan[30] ;
 wire \scan[310] ;
 wire \scan[311] ;
 wire \scan[312] ;
 wire \scan[313] ;
 wire \scan[314] ;
 wire \scan[315] ;
 wire \scan[316] ;
 wire \scan[317] ;
 wire \scan[318] ;
 wire \scan[319] ;
 wire \scan[31] ;
 wire \scan[320] ;
 wire \scan[321] ;
 wire \scan[322] ;
 wire \scan[323] ;
 wire \scan[324] ;
 wire \scan[325] ;
 wire \scan[326] ;
 wire \scan[327] ;
 wire \scan[328] ;
 wire \scan[329] ;
 wire \scan[32] ;
 wire \scan[330] ;
 wire \scan[331] ;
 wire \scan[332] ;
 wire \scan[333] ;
 wire \scan[334] ;
 wire \scan[335] ;
 wire \scan[336] ;
 wire \scan[337] ;
 wire \scan[338] ;
 wire \scan[339] ;
 wire \scan[33] ;
 wire \scan[340] ;
 wire \scan[341] ;
 wire \scan[342] ;
 wire \scan[343] ;
 wire \scan[344] ;
 wire \scan[345] ;
 wire \scan[346] ;
 wire \scan[347] ;
 wire \scan[348] ;
 wire \scan[349] ;
 wire \scan[34] ;
 wire \scan[350] ;
 wire \scan[351] ;
 wire \scan[352] ;
 wire \scan[353] ;
 wire \scan[354] ;
 wire \scan[355] ;
 wire \scan[356] ;
 wire \scan[357] ;
 wire \scan[358] ;
 wire \scan[359] ;
 wire \scan[35] ;
 wire \scan[360] ;
 wire \scan[361] ;
 wire \scan[362] ;
 wire \scan[363] ;
 wire \scan[364] ;
 wire \scan[365] ;
 wire \scan[366] ;
 wire \scan[367] ;
 wire \scan[368] ;
 wire \scan[369] ;
 wire \scan[36] ;
 wire \scan[370] ;
 wire \scan[371] ;
 wire \scan[372] ;
 wire \scan[373] ;
 wire \scan[374] ;
 wire \scan[375] ;
 wire \scan[376] ;
 wire \scan[377] ;
 wire \scan[378] ;
 wire \scan[379] ;
 wire \scan[37] ;
 wire \scan[380] ;
 wire \scan[381] ;
 wire \scan[382] ;
 wire \scan[383] ;
 wire \scan[384] ;
 wire \scan[385] ;
 wire \scan[386] ;
 wire \scan[387] ;
 wire \scan[388] ;
 wire \scan[389] ;
 wire \scan[38] ;
 wire \scan[390] ;
 wire \scan[391] ;
 wire \scan[392] ;
 wire \scan[393] ;
 wire \scan[394] ;
 wire \scan[395] ;
 wire \scan[396] ;
 wire \scan[397] ;
 wire \scan[398] ;
 wire \scan[399] ;
 wire \scan[39] ;
 wire \scan[3] ;
 wire \scan[400] ;
 wire \scan[401] ;
 wire \scan[402] ;
 wire \scan[403] ;
 wire \scan[404] ;
 wire \scan[405] ;
 wire \scan[406] ;
 wire \scan[407] ;
 wire \scan[408] ;
 wire \scan[409] ;
 wire \scan[40] ;
 wire \scan[410] ;
 wire \scan[411] ;
 wire \scan[412] ;
 wire \scan[413] ;
 wire \scan[414] ;
 wire \scan[415] ;
 wire \scan[416] ;
 wire \scan[417] ;
 wire \scan[418] ;
 wire \scan[419] ;
 wire \scan[41] ;
 wire \scan[420] ;
 wire \scan[421] ;
 wire \scan[422] ;
 wire \scan[423] ;
 wire \scan[424] ;
 wire \scan[425] ;
 wire \scan[426] ;
 wire \scan[427] ;
 wire \scan[428] ;
 wire \scan[429] ;
 wire \scan[42] ;
 wire \scan[430] ;
 wire \scan[431] ;
 wire \scan[432] ;
 wire \scan[433] ;
 wire \scan[434] ;
 wire \scan[435] ;
 wire \scan[436] ;
 wire \scan[437] ;
 wire \scan[438] ;
 wire \scan[439] ;
 wire \scan[43] ;
 wire \scan[440] ;
 wire \scan[441] ;
 wire \scan[442] ;
 wire \scan[443] ;
 wire \scan[444] ;
 wire \scan[445] ;
 wire \scan[446] ;
 wire \scan[447] ;
 wire \scan[448] ;
 wire \scan[449] ;
 wire \scan[44] ;
 wire \scan[450] ;
 wire \scan[451] ;
 wire \scan[452] ;
 wire \scan[453] ;
 wire \scan[454] ;
 wire \scan[455] ;
 wire \scan[456] ;
 wire \scan[457] ;
 wire \scan[458] ;
 wire \scan[459] ;
 wire \scan[45] ;
 wire \scan[460] ;
 wire \scan[461] ;
 wire \scan[462] ;
 wire \scan[463] ;
 wire \scan[464] ;
 wire \scan[465] ;
 wire \scan[466] ;
 wire \scan[467] ;
 wire \scan[468] ;
 wire \scan[469] ;
 wire \scan[46] ;
 wire \scan[470] ;
 wire \scan[471] ;
 wire \scan[472] ;
 wire \scan[473] ;
 wire \scan[474] ;
 wire \scan[475] ;
 wire \scan[476] ;
 wire \scan[477] ;
 wire \scan[478] ;
 wire \scan[479] ;
 wire \scan[47] ;
 wire \scan[480] ;
 wire \scan[481] ;
 wire \scan[482] ;
 wire \scan[483] ;
 wire \scan[484] ;
 wire \scan[485] ;
 wire \scan[486] ;
 wire \scan[487] ;
 wire \scan[488] ;
 wire \scan[489] ;
 wire \scan[48] ;
 wire \scan[490] ;
 wire \scan[491] ;
 wire \scan[492] ;
 wire \scan[493] ;
 wire \scan[494] ;
 wire \scan[495] ;
 wire \scan[496] ;
 wire \scan[497] ;
 wire \scan[498] ;
 wire \scan[49] ;
 wire \scan[4] ;
 wire \scan[50] ;
 wire \scan[51] ;
 wire \scan[52] ;
 wire \scan[53] ;
 wire \scan[54] ;
 wire \scan[55] ;
 wire \scan[56] ;
 wire \scan[57] ;
 wire \scan[58] ;
 wire \scan[59] ;
 wire \scan[5] ;
 wire \scan[60] ;
 wire \scan[61] ;
 wire \scan[62] ;
 wire \scan[63] ;
 wire \scan[64] ;
 wire \scan[65] ;
 wire \scan[66] ;
 wire \scan[67] ;
 wire \scan[68] ;
 wire \scan[69] ;
 wire \scan[6] ;
 wire \scan[70] ;
 wire \scan[71] ;
 wire \scan[72] ;
 wire \scan[73] ;
 wire \scan[74] ;
 wire \scan[75] ;
 wire \scan[76] ;
 wire \scan[77] ;
 wire \scan[78] ;
 wire \scan[79] ;
 wire \scan[7] ;
 wire \scan[80] ;
 wire \scan[81] ;
 wire \scan[82] ;
 wire \scan[83] ;
 wire \scan[84] ;
 wire \scan[85] ;
 wire \scan[86] ;
 wire \scan[87] ;
 wire \scan[88] ;
 wire \scan[89] ;
 wire \scan[8] ;
 wire \scan[90] ;
 wire \scan[91] ;
 wire \scan[92] ;
 wire \scan[93] ;
 wire \scan[94] ;
 wire \scan[95] ;
 wire \scan[96] ;
 wire \scan[97] ;
 wire \scan[98] ;
 wire \scan[99] ;
 wire \scan[9] ;

 scan_controller scan_controller (.clk(wb_clk_i),
    .ready(ready),
    .reset(wb_rst_i),
    .scan_clk(\clk[0] ),
    .scan_data_in(\data[498] ),
    .scan_data_out(\data[0] ),
    .scan_latch_enable(\latch[0] ),
    .scan_select(\scan[0] ),
    .set_clk_div(io_in[11]),
    .slow_clk(slow_clk),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .active_select({io_in[20],
    io_in[19],
    io_in[18],
    io_in[17],
    io_in[16],
    io_in[15],
    io_in[14],
    io_in[13],
    io_in[12]}),
    .inputs({io_in[28],
    io_in[27],
    io_in[26],
    io_in[25],
    io_in[24],
    io_in[23],
    io_in[22],
    io_in[21]}),
    .oeb({io_oeb[37],
    io_oeb[36],
    io_oeb[35],
    io_oeb[34],
    io_oeb[33],
    io_oeb[32],
    io_oeb[31],
    io_oeb[30],
    io_oeb[29]}),
    .outputs({io_out[36],
    io_out[35],
    io_out[34],
    io_out[33],
    io_out[32],
    io_out[31],
    io_out[30],
    io_out[29]}));
 scan_wrapper_334445762078310996 scan_wrapper_334445762078310996_1 (.clk_in(\clk[1] ),
    .clk_out(\clk[2] ),
    .data_in(\data[1] ),
    .data_out(\data[2] ),
    .latch_enable_in(\latch[1] ),
    .latch_enable_out(\latch[2] ),
    .scan_select_in(\scan[1] ),
    .scan_select_out(\scan[2] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_335404063203000914 scan_wrapper_335404063203000914_2 (.clk_in(\clk[2] ),
    .clk_out(\clk[3] ),
    .data_in(\data[2] ),
    .data_out(\data[3] ),
    .latch_enable_in(\latch[2] ),
    .latch_enable_out(\latch[3] ),
    .scan_select_in(\scan[2] ),
    .scan_select_out(\scan[3] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339439899388150354 scan_wrapper_339439899388150354_3 (.clk_in(\clk[3] ),
    .clk_out(\clk[4] ),
    .data_in(\data[3] ),
    .data_out(\data[4] ),
    .latch_enable_in(\latch[3] ),
    .latch_enable_out(\latch[4] ),
    .scan_select_in(\scan[3] ),
    .scan_select_out(\scan[4] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_0 (.clk_in(\clk[0] ),
    .clk_out(\clk[1] ),
    .data_in(\data[0] ),
    .data_out(\data[1] ),
    .latch_enable_in(\latch[0] ),
    .latch_enable_out(\latch[1] ),
    .scan_select_in(\scan[0] ),
    .scan_select_out(\scan[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_100 (.clk_in(\clk[100] ),
    .clk_out(\clk[101] ),
    .data_in(\data[100] ),
    .data_out(\data[101] ),
    .latch_enable_in(\latch[100] ),
    .latch_enable_out(\latch[101] ),
    .scan_select_in(\scan[100] ),
    .scan_select_out(\scan[101] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_101 (.clk_in(\clk[101] ),
    .clk_out(\clk[102] ),
    .data_in(\data[101] ),
    .data_out(\data[102] ),
    .latch_enable_in(\latch[101] ),
    .latch_enable_out(\latch[102] ),
    .scan_select_in(\scan[101] ),
    .scan_select_out(\scan[102] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_102 (.clk_in(\clk[102] ),
    .clk_out(\clk[103] ),
    .data_in(\data[102] ),
    .data_out(\data[103] ),
    .latch_enable_in(\latch[102] ),
    .latch_enable_out(\latch[103] ),
    .scan_select_in(\scan[102] ),
    .scan_select_out(\scan[103] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_103 (.clk_in(\clk[103] ),
    .clk_out(\clk[104] ),
    .data_in(\data[103] ),
    .data_out(\data[104] ),
    .latch_enable_in(\latch[103] ),
    .latch_enable_out(\latch[104] ),
    .scan_select_in(\scan[103] ),
    .scan_select_out(\scan[104] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_104 (.clk_in(\clk[104] ),
    .clk_out(\clk[105] ),
    .data_in(\data[104] ),
    .data_out(\data[105] ),
    .latch_enable_in(\latch[104] ),
    .latch_enable_out(\latch[105] ),
    .scan_select_in(\scan[104] ),
    .scan_select_out(\scan[105] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_105 (.clk_in(\clk[105] ),
    .clk_out(\clk[106] ),
    .data_in(\data[105] ),
    .data_out(\data[106] ),
    .latch_enable_in(\latch[105] ),
    .latch_enable_out(\latch[106] ),
    .scan_select_in(\scan[105] ),
    .scan_select_out(\scan[106] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_106 (.clk_in(\clk[106] ),
    .clk_out(\clk[107] ),
    .data_in(\data[106] ),
    .data_out(\data[107] ),
    .latch_enable_in(\latch[106] ),
    .latch_enable_out(\latch[107] ),
    .scan_select_in(\scan[106] ),
    .scan_select_out(\scan[107] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_107 (.clk_in(\clk[107] ),
    .clk_out(\clk[108] ),
    .data_in(\data[107] ),
    .data_out(\data[108] ),
    .latch_enable_in(\latch[107] ),
    .latch_enable_out(\latch[108] ),
    .scan_select_in(\scan[107] ),
    .scan_select_out(\scan[108] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_108 (.clk_in(\clk[108] ),
    .clk_out(\clk[109] ),
    .data_in(\data[108] ),
    .data_out(\data[109] ),
    .latch_enable_in(\latch[108] ),
    .latch_enable_out(\latch[109] ),
    .scan_select_in(\scan[108] ),
    .scan_select_out(\scan[109] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_109 (.clk_in(\clk[109] ),
    .clk_out(\clk[110] ),
    .data_in(\data[109] ),
    .data_out(\data[110] ),
    .latch_enable_in(\latch[109] ),
    .latch_enable_out(\latch[110] ),
    .scan_select_in(\scan[109] ),
    .scan_select_out(\scan[110] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_110 (.clk_in(\clk[110] ),
    .clk_out(\clk[111] ),
    .data_in(\data[110] ),
    .data_out(\data[111] ),
    .latch_enable_in(\latch[110] ),
    .latch_enable_out(\latch[111] ),
    .scan_select_in(\scan[110] ),
    .scan_select_out(\scan[111] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_111 (.clk_in(\clk[111] ),
    .clk_out(\clk[112] ),
    .data_in(\data[111] ),
    .data_out(\data[112] ),
    .latch_enable_in(\latch[111] ),
    .latch_enable_out(\latch[112] ),
    .scan_select_in(\scan[111] ),
    .scan_select_out(\scan[112] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_112 (.clk_in(\clk[112] ),
    .clk_out(\clk[113] ),
    .data_in(\data[112] ),
    .data_out(\data[113] ),
    .latch_enable_in(\latch[112] ),
    .latch_enable_out(\latch[113] ),
    .scan_select_in(\scan[112] ),
    .scan_select_out(\scan[113] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_113 (.clk_in(\clk[113] ),
    .clk_out(\clk[114] ),
    .data_in(\data[113] ),
    .data_out(\data[114] ),
    .latch_enable_in(\latch[113] ),
    .latch_enable_out(\latch[114] ),
    .scan_select_in(\scan[113] ),
    .scan_select_out(\scan[114] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_114 (.clk_in(\clk[114] ),
    .clk_out(\clk[115] ),
    .data_in(\data[114] ),
    .data_out(\data[115] ),
    .latch_enable_in(\latch[114] ),
    .latch_enable_out(\latch[115] ),
    .scan_select_in(\scan[114] ),
    .scan_select_out(\scan[115] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_115 (.clk_in(\clk[115] ),
    .clk_out(\clk[116] ),
    .data_in(\data[115] ),
    .data_out(\data[116] ),
    .latch_enable_in(\latch[115] ),
    .latch_enable_out(\latch[116] ),
    .scan_select_in(\scan[115] ),
    .scan_select_out(\scan[116] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_116 (.clk_in(\clk[116] ),
    .clk_out(\clk[117] ),
    .data_in(\data[116] ),
    .data_out(\data[117] ),
    .latch_enable_in(\latch[116] ),
    .latch_enable_out(\latch[117] ),
    .scan_select_in(\scan[116] ),
    .scan_select_out(\scan[117] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_117 (.clk_in(\clk[117] ),
    .clk_out(\clk[118] ),
    .data_in(\data[117] ),
    .data_out(\data[118] ),
    .latch_enable_in(\latch[117] ),
    .latch_enable_out(\latch[118] ),
    .scan_select_in(\scan[117] ),
    .scan_select_out(\scan[118] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_118 (.clk_in(\clk[118] ),
    .clk_out(\clk[119] ),
    .data_in(\data[118] ),
    .data_out(\data[119] ),
    .latch_enable_in(\latch[118] ),
    .latch_enable_out(\latch[119] ),
    .scan_select_in(\scan[118] ),
    .scan_select_out(\scan[119] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_119 (.clk_in(\clk[119] ),
    .clk_out(\clk[120] ),
    .data_in(\data[119] ),
    .data_out(\data[120] ),
    .latch_enable_in(\latch[119] ),
    .latch_enable_out(\latch[120] ),
    .scan_select_in(\scan[119] ),
    .scan_select_out(\scan[120] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_120 (.clk_in(\clk[120] ),
    .clk_out(\clk[121] ),
    .data_in(\data[120] ),
    .data_out(\data[121] ),
    .latch_enable_in(\latch[120] ),
    .latch_enable_out(\latch[121] ),
    .scan_select_in(\scan[120] ),
    .scan_select_out(\scan[121] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_121 (.clk_in(\clk[121] ),
    .clk_out(\clk[122] ),
    .data_in(\data[121] ),
    .data_out(\data[122] ),
    .latch_enable_in(\latch[121] ),
    .latch_enable_out(\latch[122] ),
    .scan_select_in(\scan[121] ),
    .scan_select_out(\scan[122] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_122 (.clk_in(\clk[122] ),
    .clk_out(\clk[123] ),
    .data_in(\data[122] ),
    .data_out(\data[123] ),
    .latch_enable_in(\latch[122] ),
    .latch_enable_out(\latch[123] ),
    .scan_select_in(\scan[122] ),
    .scan_select_out(\scan[123] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_123 (.clk_in(\clk[123] ),
    .clk_out(\clk[124] ),
    .data_in(\data[123] ),
    .data_out(\data[124] ),
    .latch_enable_in(\latch[123] ),
    .latch_enable_out(\latch[124] ),
    .scan_select_in(\scan[123] ),
    .scan_select_out(\scan[124] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_124 (.clk_in(\clk[124] ),
    .clk_out(\clk[125] ),
    .data_in(\data[124] ),
    .data_out(\data[125] ),
    .latch_enable_in(\latch[124] ),
    .latch_enable_out(\latch[125] ),
    .scan_select_in(\scan[124] ),
    .scan_select_out(\scan[125] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_125 (.clk_in(\clk[125] ),
    .clk_out(\clk[126] ),
    .data_in(\data[125] ),
    .data_out(\data[126] ),
    .latch_enable_in(\latch[125] ),
    .latch_enable_out(\latch[126] ),
    .scan_select_in(\scan[125] ),
    .scan_select_out(\scan[126] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_126 (.clk_in(\clk[126] ),
    .clk_out(\clk[127] ),
    .data_in(\data[126] ),
    .data_out(\data[127] ),
    .latch_enable_in(\latch[126] ),
    .latch_enable_out(\latch[127] ),
    .scan_select_in(\scan[126] ),
    .scan_select_out(\scan[127] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_127 (.clk_in(\clk[127] ),
    .clk_out(\clk[128] ),
    .data_in(\data[127] ),
    .data_out(\data[128] ),
    .latch_enable_in(\latch[127] ),
    .latch_enable_out(\latch[128] ),
    .scan_select_in(\scan[127] ),
    .scan_select_out(\scan[128] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_128 (.clk_in(\clk[128] ),
    .clk_out(\clk[129] ),
    .data_in(\data[128] ),
    .data_out(\data[129] ),
    .latch_enable_in(\latch[128] ),
    .latch_enable_out(\latch[129] ),
    .scan_select_in(\scan[128] ),
    .scan_select_out(\scan[129] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_129 (.clk_in(\clk[129] ),
    .clk_out(\clk[130] ),
    .data_in(\data[129] ),
    .data_out(\data[130] ),
    .latch_enable_in(\latch[129] ),
    .latch_enable_out(\latch[130] ),
    .scan_select_in(\scan[129] ),
    .scan_select_out(\scan[130] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_130 (.clk_in(\clk[130] ),
    .clk_out(\clk[131] ),
    .data_in(\data[130] ),
    .data_out(\data[131] ),
    .latch_enable_in(\latch[130] ),
    .latch_enable_out(\latch[131] ),
    .scan_select_in(\scan[130] ),
    .scan_select_out(\scan[131] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_131 (.clk_in(\clk[131] ),
    .clk_out(\clk[132] ),
    .data_in(\data[131] ),
    .data_out(\data[132] ),
    .latch_enable_in(\latch[131] ),
    .latch_enable_out(\latch[132] ),
    .scan_select_in(\scan[131] ),
    .scan_select_out(\scan[132] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_132 (.clk_in(\clk[132] ),
    .clk_out(\clk[133] ),
    .data_in(\data[132] ),
    .data_out(\data[133] ),
    .latch_enable_in(\latch[132] ),
    .latch_enable_out(\latch[133] ),
    .scan_select_in(\scan[132] ),
    .scan_select_out(\scan[133] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_133 (.clk_in(\clk[133] ),
    .clk_out(\clk[134] ),
    .data_in(\data[133] ),
    .data_out(\data[134] ),
    .latch_enable_in(\latch[133] ),
    .latch_enable_out(\latch[134] ),
    .scan_select_in(\scan[133] ),
    .scan_select_out(\scan[134] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_134 (.clk_in(\clk[134] ),
    .clk_out(\clk[135] ),
    .data_in(\data[134] ),
    .data_out(\data[135] ),
    .latch_enable_in(\latch[134] ),
    .latch_enable_out(\latch[135] ),
    .scan_select_in(\scan[134] ),
    .scan_select_out(\scan[135] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_135 (.clk_in(\clk[135] ),
    .clk_out(\clk[136] ),
    .data_in(\data[135] ),
    .data_out(\data[136] ),
    .latch_enable_in(\latch[135] ),
    .latch_enable_out(\latch[136] ),
    .scan_select_in(\scan[135] ),
    .scan_select_out(\scan[136] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_136 (.clk_in(\clk[136] ),
    .clk_out(\clk[137] ),
    .data_in(\data[136] ),
    .data_out(\data[137] ),
    .latch_enable_in(\latch[136] ),
    .latch_enable_out(\latch[137] ),
    .scan_select_in(\scan[136] ),
    .scan_select_out(\scan[137] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_137 (.clk_in(\clk[137] ),
    .clk_out(\clk[138] ),
    .data_in(\data[137] ),
    .data_out(\data[138] ),
    .latch_enable_in(\latch[137] ),
    .latch_enable_out(\latch[138] ),
    .scan_select_in(\scan[137] ),
    .scan_select_out(\scan[138] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_138 (.clk_in(\clk[138] ),
    .clk_out(\clk[139] ),
    .data_in(\data[138] ),
    .data_out(\data[139] ),
    .latch_enable_in(\latch[138] ),
    .latch_enable_out(\latch[139] ),
    .scan_select_in(\scan[138] ),
    .scan_select_out(\scan[139] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_139 (.clk_in(\clk[139] ),
    .clk_out(\clk[140] ),
    .data_in(\data[139] ),
    .data_out(\data[140] ),
    .latch_enable_in(\latch[139] ),
    .latch_enable_out(\latch[140] ),
    .scan_select_in(\scan[139] ),
    .scan_select_out(\scan[140] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_140 (.clk_in(\clk[140] ),
    .clk_out(\clk[141] ),
    .data_in(\data[140] ),
    .data_out(\data[141] ),
    .latch_enable_in(\latch[140] ),
    .latch_enable_out(\latch[141] ),
    .scan_select_in(\scan[140] ),
    .scan_select_out(\scan[141] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_141 (.clk_in(\clk[141] ),
    .clk_out(\clk[142] ),
    .data_in(\data[141] ),
    .data_out(\data[142] ),
    .latch_enable_in(\latch[141] ),
    .latch_enable_out(\latch[142] ),
    .scan_select_in(\scan[141] ),
    .scan_select_out(\scan[142] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_142 (.clk_in(\clk[142] ),
    .clk_out(\clk[143] ),
    .data_in(\data[142] ),
    .data_out(\data[143] ),
    .latch_enable_in(\latch[142] ),
    .latch_enable_out(\latch[143] ),
    .scan_select_in(\scan[142] ),
    .scan_select_out(\scan[143] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_143 (.clk_in(\clk[143] ),
    .clk_out(\clk[144] ),
    .data_in(\data[143] ),
    .data_out(\data[144] ),
    .latch_enable_in(\latch[143] ),
    .latch_enable_out(\latch[144] ),
    .scan_select_in(\scan[143] ),
    .scan_select_out(\scan[144] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_144 (.clk_in(\clk[144] ),
    .clk_out(\clk[145] ),
    .data_in(\data[144] ),
    .data_out(\data[145] ),
    .latch_enable_in(\latch[144] ),
    .latch_enable_out(\latch[145] ),
    .scan_select_in(\scan[144] ),
    .scan_select_out(\scan[145] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_145 (.clk_in(\clk[145] ),
    .clk_out(\clk[146] ),
    .data_in(\data[145] ),
    .data_out(\data[146] ),
    .latch_enable_in(\latch[145] ),
    .latch_enable_out(\latch[146] ),
    .scan_select_in(\scan[145] ),
    .scan_select_out(\scan[146] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_146 (.clk_in(\clk[146] ),
    .clk_out(\clk[147] ),
    .data_in(\data[146] ),
    .data_out(\data[147] ),
    .latch_enable_in(\latch[146] ),
    .latch_enable_out(\latch[147] ),
    .scan_select_in(\scan[146] ),
    .scan_select_out(\scan[147] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_147 (.clk_in(\clk[147] ),
    .clk_out(\clk[148] ),
    .data_in(\data[147] ),
    .data_out(\data[148] ),
    .latch_enable_in(\latch[147] ),
    .latch_enable_out(\latch[148] ),
    .scan_select_in(\scan[147] ),
    .scan_select_out(\scan[148] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_148 (.clk_in(\clk[148] ),
    .clk_out(\clk[149] ),
    .data_in(\data[148] ),
    .data_out(\data[149] ),
    .latch_enable_in(\latch[148] ),
    .latch_enable_out(\latch[149] ),
    .scan_select_in(\scan[148] ),
    .scan_select_out(\scan[149] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_149 (.clk_in(\clk[149] ),
    .clk_out(\clk[150] ),
    .data_in(\data[149] ),
    .data_out(\data[150] ),
    .latch_enable_in(\latch[149] ),
    .latch_enable_out(\latch[150] ),
    .scan_select_in(\scan[149] ),
    .scan_select_out(\scan[150] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_150 (.clk_in(\clk[150] ),
    .clk_out(\clk[151] ),
    .data_in(\data[150] ),
    .data_out(\data[151] ),
    .latch_enable_in(\latch[150] ),
    .latch_enable_out(\latch[151] ),
    .scan_select_in(\scan[150] ),
    .scan_select_out(\scan[151] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_151 (.clk_in(\clk[151] ),
    .clk_out(\clk[152] ),
    .data_in(\data[151] ),
    .data_out(\data[152] ),
    .latch_enable_in(\latch[151] ),
    .latch_enable_out(\latch[152] ),
    .scan_select_in(\scan[151] ),
    .scan_select_out(\scan[152] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_152 (.clk_in(\clk[152] ),
    .clk_out(\clk[153] ),
    .data_in(\data[152] ),
    .data_out(\data[153] ),
    .latch_enable_in(\latch[152] ),
    .latch_enable_out(\latch[153] ),
    .scan_select_in(\scan[152] ),
    .scan_select_out(\scan[153] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_153 (.clk_in(\clk[153] ),
    .clk_out(\clk[154] ),
    .data_in(\data[153] ),
    .data_out(\data[154] ),
    .latch_enable_in(\latch[153] ),
    .latch_enable_out(\latch[154] ),
    .scan_select_in(\scan[153] ),
    .scan_select_out(\scan[154] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_154 (.clk_in(\clk[154] ),
    .clk_out(\clk[155] ),
    .data_in(\data[154] ),
    .data_out(\data[155] ),
    .latch_enable_in(\latch[154] ),
    .latch_enable_out(\latch[155] ),
    .scan_select_in(\scan[154] ),
    .scan_select_out(\scan[155] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_155 (.clk_in(\clk[155] ),
    .clk_out(\clk[156] ),
    .data_in(\data[155] ),
    .data_out(\data[156] ),
    .latch_enable_in(\latch[155] ),
    .latch_enable_out(\latch[156] ),
    .scan_select_in(\scan[155] ),
    .scan_select_out(\scan[156] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_156 (.clk_in(\clk[156] ),
    .clk_out(\clk[157] ),
    .data_in(\data[156] ),
    .data_out(\data[157] ),
    .latch_enable_in(\latch[156] ),
    .latch_enable_out(\latch[157] ),
    .scan_select_in(\scan[156] ),
    .scan_select_out(\scan[157] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_157 (.clk_in(\clk[157] ),
    .clk_out(\clk[158] ),
    .data_in(\data[157] ),
    .data_out(\data[158] ),
    .latch_enable_in(\latch[157] ),
    .latch_enable_out(\latch[158] ),
    .scan_select_in(\scan[157] ),
    .scan_select_out(\scan[158] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_158 (.clk_in(\clk[158] ),
    .clk_out(\clk[159] ),
    .data_in(\data[158] ),
    .data_out(\data[159] ),
    .latch_enable_in(\latch[158] ),
    .latch_enable_out(\latch[159] ),
    .scan_select_in(\scan[158] ),
    .scan_select_out(\scan[159] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_159 (.clk_in(\clk[159] ),
    .clk_out(\clk[160] ),
    .data_in(\data[159] ),
    .data_out(\data[160] ),
    .latch_enable_in(\latch[159] ),
    .latch_enable_out(\latch[160] ),
    .scan_select_in(\scan[159] ),
    .scan_select_out(\scan[160] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_160 (.clk_in(\clk[160] ),
    .clk_out(\clk[161] ),
    .data_in(\data[160] ),
    .data_out(\data[161] ),
    .latch_enable_in(\latch[160] ),
    .latch_enable_out(\latch[161] ),
    .scan_select_in(\scan[160] ),
    .scan_select_out(\scan[161] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_161 (.clk_in(\clk[161] ),
    .clk_out(\clk[162] ),
    .data_in(\data[161] ),
    .data_out(\data[162] ),
    .latch_enable_in(\latch[161] ),
    .latch_enable_out(\latch[162] ),
    .scan_select_in(\scan[161] ),
    .scan_select_out(\scan[162] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_162 (.clk_in(\clk[162] ),
    .clk_out(\clk[163] ),
    .data_in(\data[162] ),
    .data_out(\data[163] ),
    .latch_enable_in(\latch[162] ),
    .latch_enable_out(\latch[163] ),
    .scan_select_in(\scan[162] ),
    .scan_select_out(\scan[163] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_163 (.clk_in(\clk[163] ),
    .clk_out(\clk[164] ),
    .data_in(\data[163] ),
    .data_out(\data[164] ),
    .latch_enable_in(\latch[163] ),
    .latch_enable_out(\latch[164] ),
    .scan_select_in(\scan[163] ),
    .scan_select_out(\scan[164] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_164 (.clk_in(\clk[164] ),
    .clk_out(\clk[165] ),
    .data_in(\data[164] ),
    .data_out(\data[165] ),
    .latch_enable_in(\latch[164] ),
    .latch_enable_out(\latch[165] ),
    .scan_select_in(\scan[164] ),
    .scan_select_out(\scan[165] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_165 (.clk_in(\clk[165] ),
    .clk_out(\clk[166] ),
    .data_in(\data[165] ),
    .data_out(\data[166] ),
    .latch_enable_in(\latch[165] ),
    .latch_enable_out(\latch[166] ),
    .scan_select_in(\scan[165] ),
    .scan_select_out(\scan[166] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_166 (.clk_in(\clk[166] ),
    .clk_out(\clk[167] ),
    .data_in(\data[166] ),
    .data_out(\data[167] ),
    .latch_enable_in(\latch[166] ),
    .latch_enable_out(\latch[167] ),
    .scan_select_in(\scan[166] ),
    .scan_select_out(\scan[167] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_167 (.clk_in(\clk[167] ),
    .clk_out(\clk[168] ),
    .data_in(\data[167] ),
    .data_out(\data[168] ),
    .latch_enable_in(\latch[167] ),
    .latch_enable_out(\latch[168] ),
    .scan_select_in(\scan[167] ),
    .scan_select_out(\scan[168] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_168 (.clk_in(\clk[168] ),
    .clk_out(\clk[169] ),
    .data_in(\data[168] ),
    .data_out(\data[169] ),
    .latch_enable_in(\latch[168] ),
    .latch_enable_out(\latch[169] ),
    .scan_select_in(\scan[168] ),
    .scan_select_out(\scan[169] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_169 (.clk_in(\clk[169] ),
    .clk_out(\clk[170] ),
    .data_in(\data[169] ),
    .data_out(\data[170] ),
    .latch_enable_in(\latch[169] ),
    .latch_enable_out(\latch[170] ),
    .scan_select_in(\scan[169] ),
    .scan_select_out(\scan[170] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_170 (.clk_in(\clk[170] ),
    .clk_out(\clk[171] ),
    .data_in(\data[170] ),
    .data_out(\data[171] ),
    .latch_enable_in(\latch[170] ),
    .latch_enable_out(\latch[171] ),
    .scan_select_in(\scan[170] ),
    .scan_select_out(\scan[171] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_171 (.clk_in(\clk[171] ),
    .clk_out(\clk[172] ),
    .data_in(\data[171] ),
    .data_out(\data[172] ),
    .latch_enable_in(\latch[171] ),
    .latch_enable_out(\latch[172] ),
    .scan_select_in(\scan[171] ),
    .scan_select_out(\scan[172] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_172 (.clk_in(\clk[172] ),
    .clk_out(\clk[173] ),
    .data_in(\data[172] ),
    .data_out(\data[173] ),
    .latch_enable_in(\latch[172] ),
    .latch_enable_out(\latch[173] ),
    .scan_select_in(\scan[172] ),
    .scan_select_out(\scan[173] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_173 (.clk_in(\clk[173] ),
    .clk_out(\clk[174] ),
    .data_in(\data[173] ),
    .data_out(\data[174] ),
    .latch_enable_in(\latch[173] ),
    .latch_enable_out(\latch[174] ),
    .scan_select_in(\scan[173] ),
    .scan_select_out(\scan[174] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_174 (.clk_in(\clk[174] ),
    .clk_out(\clk[175] ),
    .data_in(\data[174] ),
    .data_out(\data[175] ),
    .latch_enable_in(\latch[174] ),
    .latch_enable_out(\latch[175] ),
    .scan_select_in(\scan[174] ),
    .scan_select_out(\scan[175] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_175 (.clk_in(\clk[175] ),
    .clk_out(\clk[176] ),
    .data_in(\data[175] ),
    .data_out(\data[176] ),
    .latch_enable_in(\latch[175] ),
    .latch_enable_out(\latch[176] ),
    .scan_select_in(\scan[175] ),
    .scan_select_out(\scan[176] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_176 (.clk_in(\clk[176] ),
    .clk_out(\clk[177] ),
    .data_in(\data[176] ),
    .data_out(\data[177] ),
    .latch_enable_in(\latch[176] ),
    .latch_enable_out(\latch[177] ),
    .scan_select_in(\scan[176] ),
    .scan_select_out(\scan[177] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_177 (.clk_in(\clk[177] ),
    .clk_out(\clk[178] ),
    .data_in(\data[177] ),
    .data_out(\data[178] ),
    .latch_enable_in(\latch[177] ),
    .latch_enable_out(\latch[178] ),
    .scan_select_in(\scan[177] ),
    .scan_select_out(\scan[178] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_178 (.clk_in(\clk[178] ),
    .clk_out(\clk[179] ),
    .data_in(\data[178] ),
    .data_out(\data[179] ),
    .latch_enable_in(\latch[178] ),
    .latch_enable_out(\latch[179] ),
    .scan_select_in(\scan[178] ),
    .scan_select_out(\scan[179] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_179 (.clk_in(\clk[179] ),
    .clk_out(\clk[180] ),
    .data_in(\data[179] ),
    .data_out(\data[180] ),
    .latch_enable_in(\latch[179] ),
    .latch_enable_out(\latch[180] ),
    .scan_select_in(\scan[179] ),
    .scan_select_out(\scan[180] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_18 (.clk_in(\clk[18] ),
    .clk_out(\clk[19] ),
    .data_in(\data[18] ),
    .data_out(\data[19] ),
    .latch_enable_in(\latch[18] ),
    .latch_enable_out(\latch[19] ),
    .scan_select_in(\scan[18] ),
    .scan_select_out(\scan[19] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_180 (.clk_in(\clk[180] ),
    .clk_out(\clk[181] ),
    .data_in(\data[180] ),
    .data_out(\data[181] ),
    .latch_enable_in(\latch[180] ),
    .latch_enable_out(\latch[181] ),
    .scan_select_in(\scan[180] ),
    .scan_select_out(\scan[181] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_181 (.clk_in(\clk[181] ),
    .clk_out(\clk[182] ),
    .data_in(\data[181] ),
    .data_out(\data[182] ),
    .latch_enable_in(\latch[181] ),
    .latch_enable_out(\latch[182] ),
    .scan_select_in(\scan[181] ),
    .scan_select_out(\scan[182] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_182 (.clk_in(\clk[182] ),
    .clk_out(\clk[183] ),
    .data_in(\data[182] ),
    .data_out(\data[183] ),
    .latch_enable_in(\latch[182] ),
    .latch_enable_out(\latch[183] ),
    .scan_select_in(\scan[182] ),
    .scan_select_out(\scan[183] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_183 (.clk_in(\clk[183] ),
    .clk_out(\clk[184] ),
    .data_in(\data[183] ),
    .data_out(\data[184] ),
    .latch_enable_in(\latch[183] ),
    .latch_enable_out(\latch[184] ),
    .scan_select_in(\scan[183] ),
    .scan_select_out(\scan[184] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_184 (.clk_in(\clk[184] ),
    .clk_out(\clk[185] ),
    .data_in(\data[184] ),
    .data_out(\data[185] ),
    .latch_enable_in(\latch[184] ),
    .latch_enable_out(\latch[185] ),
    .scan_select_in(\scan[184] ),
    .scan_select_out(\scan[185] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_185 (.clk_in(\clk[185] ),
    .clk_out(\clk[186] ),
    .data_in(\data[185] ),
    .data_out(\data[186] ),
    .latch_enable_in(\latch[185] ),
    .latch_enable_out(\latch[186] ),
    .scan_select_in(\scan[185] ),
    .scan_select_out(\scan[186] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_186 (.clk_in(\clk[186] ),
    .clk_out(\clk[187] ),
    .data_in(\data[186] ),
    .data_out(\data[187] ),
    .latch_enable_in(\latch[186] ),
    .latch_enable_out(\latch[187] ),
    .scan_select_in(\scan[186] ),
    .scan_select_out(\scan[187] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_187 (.clk_in(\clk[187] ),
    .clk_out(\clk[188] ),
    .data_in(\data[187] ),
    .data_out(\data[188] ),
    .latch_enable_in(\latch[187] ),
    .latch_enable_out(\latch[188] ),
    .scan_select_in(\scan[187] ),
    .scan_select_out(\scan[188] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_188 (.clk_in(\clk[188] ),
    .clk_out(\clk[189] ),
    .data_in(\data[188] ),
    .data_out(\data[189] ),
    .latch_enable_in(\latch[188] ),
    .latch_enable_out(\latch[189] ),
    .scan_select_in(\scan[188] ),
    .scan_select_out(\scan[189] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_189 (.clk_in(\clk[189] ),
    .clk_out(\clk[190] ),
    .data_in(\data[189] ),
    .data_out(\data[190] ),
    .latch_enable_in(\latch[189] ),
    .latch_enable_out(\latch[190] ),
    .scan_select_in(\scan[189] ),
    .scan_select_out(\scan[190] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_19 (.clk_in(\clk[19] ),
    .clk_out(\clk[20] ),
    .data_in(\data[19] ),
    .data_out(\data[20] ),
    .latch_enable_in(\latch[19] ),
    .latch_enable_out(\latch[20] ),
    .scan_select_in(\scan[19] ),
    .scan_select_out(\scan[20] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_190 (.clk_in(\clk[190] ),
    .clk_out(\clk[191] ),
    .data_in(\data[190] ),
    .data_out(\data[191] ),
    .latch_enable_in(\latch[190] ),
    .latch_enable_out(\latch[191] ),
    .scan_select_in(\scan[190] ),
    .scan_select_out(\scan[191] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_191 (.clk_in(\clk[191] ),
    .clk_out(\clk[192] ),
    .data_in(\data[191] ),
    .data_out(\data[192] ),
    .latch_enable_in(\latch[191] ),
    .latch_enable_out(\latch[192] ),
    .scan_select_in(\scan[191] ),
    .scan_select_out(\scan[192] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_192 (.clk_in(\clk[192] ),
    .clk_out(\clk[193] ),
    .data_in(\data[192] ),
    .data_out(\data[193] ),
    .latch_enable_in(\latch[192] ),
    .latch_enable_out(\latch[193] ),
    .scan_select_in(\scan[192] ),
    .scan_select_out(\scan[193] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_193 (.clk_in(\clk[193] ),
    .clk_out(\clk[194] ),
    .data_in(\data[193] ),
    .data_out(\data[194] ),
    .latch_enable_in(\latch[193] ),
    .latch_enable_out(\latch[194] ),
    .scan_select_in(\scan[193] ),
    .scan_select_out(\scan[194] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_194 (.clk_in(\clk[194] ),
    .clk_out(\clk[195] ),
    .data_in(\data[194] ),
    .data_out(\data[195] ),
    .latch_enable_in(\latch[194] ),
    .latch_enable_out(\latch[195] ),
    .scan_select_in(\scan[194] ),
    .scan_select_out(\scan[195] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_195 (.clk_in(\clk[195] ),
    .clk_out(\clk[196] ),
    .data_in(\data[195] ),
    .data_out(\data[196] ),
    .latch_enable_in(\latch[195] ),
    .latch_enable_out(\latch[196] ),
    .scan_select_in(\scan[195] ),
    .scan_select_out(\scan[196] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_196 (.clk_in(\clk[196] ),
    .clk_out(\clk[197] ),
    .data_in(\data[196] ),
    .data_out(\data[197] ),
    .latch_enable_in(\latch[196] ),
    .latch_enable_out(\latch[197] ),
    .scan_select_in(\scan[196] ),
    .scan_select_out(\scan[197] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_197 (.clk_in(\clk[197] ),
    .clk_out(\clk[198] ),
    .data_in(\data[197] ),
    .data_out(\data[198] ),
    .latch_enable_in(\latch[197] ),
    .latch_enable_out(\latch[198] ),
    .scan_select_in(\scan[197] ),
    .scan_select_out(\scan[198] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_198 (.clk_in(\clk[198] ),
    .clk_out(\clk[199] ),
    .data_in(\data[198] ),
    .data_out(\data[199] ),
    .latch_enable_in(\latch[198] ),
    .latch_enable_out(\latch[199] ),
    .scan_select_in(\scan[198] ),
    .scan_select_out(\scan[199] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_199 (.clk_in(\clk[199] ),
    .clk_out(\clk[200] ),
    .data_in(\data[199] ),
    .data_out(\data[200] ),
    .latch_enable_in(\latch[199] ),
    .latch_enable_out(\latch[200] ),
    .scan_select_in(\scan[199] ),
    .scan_select_out(\scan[200] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_20 (.clk_in(\clk[20] ),
    .clk_out(\clk[21] ),
    .data_in(\data[20] ),
    .data_out(\data[21] ),
    .latch_enable_in(\latch[20] ),
    .latch_enable_out(\latch[21] ),
    .scan_select_in(\scan[20] ),
    .scan_select_out(\scan[21] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_200 (.clk_in(\clk[200] ),
    .clk_out(\clk[201] ),
    .data_in(\data[200] ),
    .data_out(\data[201] ),
    .latch_enable_in(\latch[200] ),
    .latch_enable_out(\latch[201] ),
    .scan_select_in(\scan[200] ),
    .scan_select_out(\scan[201] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_201 (.clk_in(\clk[201] ),
    .clk_out(\clk[202] ),
    .data_in(\data[201] ),
    .data_out(\data[202] ),
    .latch_enable_in(\latch[201] ),
    .latch_enable_out(\latch[202] ),
    .scan_select_in(\scan[201] ),
    .scan_select_out(\scan[202] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_202 (.clk_in(\clk[202] ),
    .clk_out(\clk[203] ),
    .data_in(\data[202] ),
    .data_out(\data[203] ),
    .latch_enable_in(\latch[202] ),
    .latch_enable_out(\latch[203] ),
    .scan_select_in(\scan[202] ),
    .scan_select_out(\scan[203] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_203 (.clk_in(\clk[203] ),
    .clk_out(\clk[204] ),
    .data_in(\data[203] ),
    .data_out(\data[204] ),
    .latch_enable_in(\latch[203] ),
    .latch_enable_out(\latch[204] ),
    .scan_select_in(\scan[203] ),
    .scan_select_out(\scan[204] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_204 (.clk_in(\clk[204] ),
    .clk_out(\clk[205] ),
    .data_in(\data[204] ),
    .data_out(\data[205] ),
    .latch_enable_in(\latch[204] ),
    .latch_enable_out(\latch[205] ),
    .scan_select_in(\scan[204] ),
    .scan_select_out(\scan[205] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_205 (.clk_in(\clk[205] ),
    .clk_out(\clk[206] ),
    .data_in(\data[205] ),
    .data_out(\data[206] ),
    .latch_enable_in(\latch[205] ),
    .latch_enable_out(\latch[206] ),
    .scan_select_in(\scan[205] ),
    .scan_select_out(\scan[206] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_206 (.clk_in(\clk[206] ),
    .clk_out(\clk[207] ),
    .data_in(\data[206] ),
    .data_out(\data[207] ),
    .latch_enable_in(\latch[206] ),
    .latch_enable_out(\latch[207] ),
    .scan_select_in(\scan[206] ),
    .scan_select_out(\scan[207] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_207 (.clk_in(\clk[207] ),
    .clk_out(\clk[208] ),
    .data_in(\data[207] ),
    .data_out(\data[208] ),
    .latch_enable_in(\latch[207] ),
    .latch_enable_out(\latch[208] ),
    .scan_select_in(\scan[207] ),
    .scan_select_out(\scan[208] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_208 (.clk_in(\clk[208] ),
    .clk_out(\clk[209] ),
    .data_in(\data[208] ),
    .data_out(\data[209] ),
    .latch_enable_in(\latch[208] ),
    .latch_enable_out(\latch[209] ),
    .scan_select_in(\scan[208] ),
    .scan_select_out(\scan[209] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_209 (.clk_in(\clk[209] ),
    .clk_out(\clk[210] ),
    .data_in(\data[209] ),
    .data_out(\data[210] ),
    .latch_enable_in(\latch[209] ),
    .latch_enable_out(\latch[210] ),
    .scan_select_in(\scan[209] ),
    .scan_select_out(\scan[210] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_21 (.clk_in(\clk[21] ),
    .clk_out(\clk[22] ),
    .data_in(\data[21] ),
    .data_out(\data[22] ),
    .latch_enable_in(\latch[21] ),
    .latch_enable_out(\latch[22] ),
    .scan_select_in(\scan[21] ),
    .scan_select_out(\scan[22] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_210 (.clk_in(\clk[210] ),
    .clk_out(\clk[211] ),
    .data_in(\data[210] ),
    .data_out(\data[211] ),
    .latch_enable_in(\latch[210] ),
    .latch_enable_out(\latch[211] ),
    .scan_select_in(\scan[210] ),
    .scan_select_out(\scan[211] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_211 (.clk_in(\clk[211] ),
    .clk_out(\clk[212] ),
    .data_in(\data[211] ),
    .data_out(\data[212] ),
    .latch_enable_in(\latch[211] ),
    .latch_enable_out(\latch[212] ),
    .scan_select_in(\scan[211] ),
    .scan_select_out(\scan[212] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_212 (.clk_in(\clk[212] ),
    .clk_out(\clk[213] ),
    .data_in(\data[212] ),
    .data_out(\data[213] ),
    .latch_enable_in(\latch[212] ),
    .latch_enable_out(\latch[213] ),
    .scan_select_in(\scan[212] ),
    .scan_select_out(\scan[213] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_213 (.clk_in(\clk[213] ),
    .clk_out(\clk[214] ),
    .data_in(\data[213] ),
    .data_out(\data[214] ),
    .latch_enable_in(\latch[213] ),
    .latch_enable_out(\latch[214] ),
    .scan_select_in(\scan[213] ),
    .scan_select_out(\scan[214] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_214 (.clk_in(\clk[214] ),
    .clk_out(\clk[215] ),
    .data_in(\data[214] ),
    .data_out(\data[215] ),
    .latch_enable_in(\latch[214] ),
    .latch_enable_out(\latch[215] ),
    .scan_select_in(\scan[214] ),
    .scan_select_out(\scan[215] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_215 (.clk_in(\clk[215] ),
    .clk_out(\clk[216] ),
    .data_in(\data[215] ),
    .data_out(\data[216] ),
    .latch_enable_in(\latch[215] ),
    .latch_enable_out(\latch[216] ),
    .scan_select_in(\scan[215] ),
    .scan_select_out(\scan[216] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_216 (.clk_in(\clk[216] ),
    .clk_out(\clk[217] ),
    .data_in(\data[216] ),
    .data_out(\data[217] ),
    .latch_enable_in(\latch[216] ),
    .latch_enable_out(\latch[217] ),
    .scan_select_in(\scan[216] ),
    .scan_select_out(\scan[217] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_217 (.clk_in(\clk[217] ),
    .clk_out(\clk[218] ),
    .data_in(\data[217] ),
    .data_out(\data[218] ),
    .latch_enable_in(\latch[217] ),
    .latch_enable_out(\latch[218] ),
    .scan_select_in(\scan[217] ),
    .scan_select_out(\scan[218] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_218 (.clk_in(\clk[218] ),
    .clk_out(\clk[219] ),
    .data_in(\data[218] ),
    .data_out(\data[219] ),
    .latch_enable_in(\latch[218] ),
    .latch_enable_out(\latch[219] ),
    .scan_select_in(\scan[218] ),
    .scan_select_out(\scan[219] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_219 (.clk_in(\clk[219] ),
    .clk_out(\clk[220] ),
    .data_in(\data[219] ),
    .data_out(\data[220] ),
    .latch_enable_in(\latch[219] ),
    .latch_enable_out(\latch[220] ),
    .scan_select_in(\scan[219] ),
    .scan_select_out(\scan[220] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_22 (.clk_in(\clk[22] ),
    .clk_out(\clk[23] ),
    .data_in(\data[22] ),
    .data_out(\data[23] ),
    .latch_enable_in(\latch[22] ),
    .latch_enable_out(\latch[23] ),
    .scan_select_in(\scan[22] ),
    .scan_select_out(\scan[23] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_220 (.clk_in(\clk[220] ),
    .clk_out(\clk[221] ),
    .data_in(\data[220] ),
    .data_out(\data[221] ),
    .latch_enable_in(\latch[220] ),
    .latch_enable_out(\latch[221] ),
    .scan_select_in(\scan[220] ),
    .scan_select_out(\scan[221] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_221 (.clk_in(\clk[221] ),
    .clk_out(\clk[222] ),
    .data_in(\data[221] ),
    .data_out(\data[222] ),
    .latch_enable_in(\latch[221] ),
    .latch_enable_out(\latch[222] ),
    .scan_select_in(\scan[221] ),
    .scan_select_out(\scan[222] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_222 (.clk_in(\clk[222] ),
    .clk_out(\clk[223] ),
    .data_in(\data[222] ),
    .data_out(\data[223] ),
    .latch_enable_in(\latch[222] ),
    .latch_enable_out(\latch[223] ),
    .scan_select_in(\scan[222] ),
    .scan_select_out(\scan[223] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_223 (.clk_in(\clk[223] ),
    .clk_out(\clk[224] ),
    .data_in(\data[223] ),
    .data_out(\data[224] ),
    .latch_enable_in(\latch[223] ),
    .latch_enable_out(\latch[224] ),
    .scan_select_in(\scan[223] ),
    .scan_select_out(\scan[224] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_224 (.clk_in(\clk[224] ),
    .clk_out(\clk[225] ),
    .data_in(\data[224] ),
    .data_out(\data[225] ),
    .latch_enable_in(\latch[224] ),
    .latch_enable_out(\latch[225] ),
    .scan_select_in(\scan[224] ),
    .scan_select_out(\scan[225] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_225 (.clk_in(\clk[225] ),
    .clk_out(\clk[226] ),
    .data_in(\data[225] ),
    .data_out(\data[226] ),
    .latch_enable_in(\latch[225] ),
    .latch_enable_out(\latch[226] ),
    .scan_select_in(\scan[225] ),
    .scan_select_out(\scan[226] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_226 (.clk_in(\clk[226] ),
    .clk_out(\clk[227] ),
    .data_in(\data[226] ),
    .data_out(\data[227] ),
    .latch_enable_in(\latch[226] ),
    .latch_enable_out(\latch[227] ),
    .scan_select_in(\scan[226] ),
    .scan_select_out(\scan[227] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_227 (.clk_in(\clk[227] ),
    .clk_out(\clk[228] ),
    .data_in(\data[227] ),
    .data_out(\data[228] ),
    .latch_enable_in(\latch[227] ),
    .latch_enable_out(\latch[228] ),
    .scan_select_in(\scan[227] ),
    .scan_select_out(\scan[228] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_228 (.clk_in(\clk[228] ),
    .clk_out(\clk[229] ),
    .data_in(\data[228] ),
    .data_out(\data[229] ),
    .latch_enable_in(\latch[228] ),
    .latch_enable_out(\latch[229] ),
    .scan_select_in(\scan[228] ),
    .scan_select_out(\scan[229] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_229 (.clk_in(\clk[229] ),
    .clk_out(\clk[230] ),
    .data_in(\data[229] ),
    .data_out(\data[230] ),
    .latch_enable_in(\latch[229] ),
    .latch_enable_out(\latch[230] ),
    .scan_select_in(\scan[229] ),
    .scan_select_out(\scan[230] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_23 (.clk_in(\clk[23] ),
    .clk_out(\clk[24] ),
    .data_in(\data[23] ),
    .data_out(\data[24] ),
    .latch_enable_in(\latch[23] ),
    .latch_enable_out(\latch[24] ),
    .scan_select_in(\scan[23] ),
    .scan_select_out(\scan[24] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_230 (.clk_in(\clk[230] ),
    .clk_out(\clk[231] ),
    .data_in(\data[230] ),
    .data_out(\data[231] ),
    .latch_enable_in(\latch[230] ),
    .latch_enable_out(\latch[231] ),
    .scan_select_in(\scan[230] ),
    .scan_select_out(\scan[231] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_231 (.clk_in(\clk[231] ),
    .clk_out(\clk[232] ),
    .data_in(\data[231] ),
    .data_out(\data[232] ),
    .latch_enable_in(\latch[231] ),
    .latch_enable_out(\latch[232] ),
    .scan_select_in(\scan[231] ),
    .scan_select_out(\scan[232] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_232 (.clk_in(\clk[232] ),
    .clk_out(\clk[233] ),
    .data_in(\data[232] ),
    .data_out(\data[233] ),
    .latch_enable_in(\latch[232] ),
    .latch_enable_out(\latch[233] ),
    .scan_select_in(\scan[232] ),
    .scan_select_out(\scan[233] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_233 (.clk_in(\clk[233] ),
    .clk_out(\clk[234] ),
    .data_in(\data[233] ),
    .data_out(\data[234] ),
    .latch_enable_in(\latch[233] ),
    .latch_enable_out(\latch[234] ),
    .scan_select_in(\scan[233] ),
    .scan_select_out(\scan[234] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_234 (.clk_in(\clk[234] ),
    .clk_out(\clk[235] ),
    .data_in(\data[234] ),
    .data_out(\data[235] ),
    .latch_enable_in(\latch[234] ),
    .latch_enable_out(\latch[235] ),
    .scan_select_in(\scan[234] ),
    .scan_select_out(\scan[235] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_235 (.clk_in(\clk[235] ),
    .clk_out(\clk[236] ),
    .data_in(\data[235] ),
    .data_out(\data[236] ),
    .latch_enable_in(\latch[235] ),
    .latch_enable_out(\latch[236] ),
    .scan_select_in(\scan[235] ),
    .scan_select_out(\scan[236] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_236 (.clk_in(\clk[236] ),
    .clk_out(\clk[237] ),
    .data_in(\data[236] ),
    .data_out(\data[237] ),
    .latch_enable_in(\latch[236] ),
    .latch_enable_out(\latch[237] ),
    .scan_select_in(\scan[236] ),
    .scan_select_out(\scan[237] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_237 (.clk_in(\clk[237] ),
    .clk_out(\clk[238] ),
    .data_in(\data[237] ),
    .data_out(\data[238] ),
    .latch_enable_in(\latch[237] ),
    .latch_enable_out(\latch[238] ),
    .scan_select_in(\scan[237] ),
    .scan_select_out(\scan[238] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_238 (.clk_in(\clk[238] ),
    .clk_out(\clk[239] ),
    .data_in(\data[238] ),
    .data_out(\data[239] ),
    .latch_enable_in(\latch[238] ),
    .latch_enable_out(\latch[239] ),
    .scan_select_in(\scan[238] ),
    .scan_select_out(\scan[239] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_239 (.clk_in(\clk[239] ),
    .clk_out(\clk[240] ),
    .data_in(\data[239] ),
    .data_out(\data[240] ),
    .latch_enable_in(\latch[239] ),
    .latch_enable_out(\latch[240] ),
    .scan_select_in(\scan[239] ),
    .scan_select_out(\scan[240] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_24 (.clk_in(\clk[24] ),
    .clk_out(\clk[25] ),
    .data_in(\data[24] ),
    .data_out(\data[25] ),
    .latch_enable_in(\latch[24] ),
    .latch_enable_out(\latch[25] ),
    .scan_select_in(\scan[24] ),
    .scan_select_out(\scan[25] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_240 (.clk_in(\clk[240] ),
    .clk_out(\clk[241] ),
    .data_in(\data[240] ),
    .data_out(\data[241] ),
    .latch_enable_in(\latch[240] ),
    .latch_enable_out(\latch[241] ),
    .scan_select_in(\scan[240] ),
    .scan_select_out(\scan[241] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_241 (.clk_in(\clk[241] ),
    .clk_out(\clk[242] ),
    .data_in(\data[241] ),
    .data_out(\data[242] ),
    .latch_enable_in(\latch[241] ),
    .latch_enable_out(\latch[242] ),
    .scan_select_in(\scan[241] ),
    .scan_select_out(\scan[242] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_242 (.clk_in(\clk[242] ),
    .clk_out(\clk[243] ),
    .data_in(\data[242] ),
    .data_out(\data[243] ),
    .latch_enable_in(\latch[242] ),
    .latch_enable_out(\latch[243] ),
    .scan_select_in(\scan[242] ),
    .scan_select_out(\scan[243] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_243 (.clk_in(\clk[243] ),
    .clk_out(\clk[244] ),
    .data_in(\data[243] ),
    .data_out(\data[244] ),
    .latch_enable_in(\latch[243] ),
    .latch_enable_out(\latch[244] ),
    .scan_select_in(\scan[243] ),
    .scan_select_out(\scan[244] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_244 (.clk_in(\clk[244] ),
    .clk_out(\clk[245] ),
    .data_in(\data[244] ),
    .data_out(\data[245] ),
    .latch_enable_in(\latch[244] ),
    .latch_enable_out(\latch[245] ),
    .scan_select_in(\scan[244] ),
    .scan_select_out(\scan[245] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_245 (.clk_in(\clk[245] ),
    .clk_out(\clk[246] ),
    .data_in(\data[245] ),
    .data_out(\data[246] ),
    .latch_enable_in(\latch[245] ),
    .latch_enable_out(\latch[246] ),
    .scan_select_in(\scan[245] ),
    .scan_select_out(\scan[246] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_246 (.clk_in(\clk[246] ),
    .clk_out(\clk[247] ),
    .data_in(\data[246] ),
    .data_out(\data[247] ),
    .latch_enable_in(\latch[246] ),
    .latch_enable_out(\latch[247] ),
    .scan_select_in(\scan[246] ),
    .scan_select_out(\scan[247] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_247 (.clk_in(\clk[247] ),
    .clk_out(\clk[248] ),
    .data_in(\data[247] ),
    .data_out(\data[248] ),
    .latch_enable_in(\latch[247] ),
    .latch_enable_out(\latch[248] ),
    .scan_select_in(\scan[247] ),
    .scan_select_out(\scan[248] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_248 (.clk_in(\clk[248] ),
    .clk_out(\clk[249] ),
    .data_in(\data[248] ),
    .data_out(\data[249] ),
    .latch_enable_in(\latch[248] ),
    .latch_enable_out(\latch[249] ),
    .scan_select_in(\scan[248] ),
    .scan_select_out(\scan[249] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_249 (.clk_in(\clk[249] ),
    .clk_out(\clk[250] ),
    .data_in(\data[249] ),
    .data_out(\data[250] ),
    .latch_enable_in(\latch[249] ),
    .latch_enable_out(\latch[250] ),
    .scan_select_in(\scan[249] ),
    .scan_select_out(\scan[250] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_25 (.clk_in(\clk[25] ),
    .clk_out(\clk[26] ),
    .data_in(\data[25] ),
    .data_out(\data[26] ),
    .latch_enable_in(\latch[25] ),
    .latch_enable_out(\latch[26] ),
    .scan_select_in(\scan[25] ),
    .scan_select_out(\scan[26] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_250 (.clk_in(\clk[250] ),
    .clk_out(\clk[251] ),
    .data_in(\data[250] ),
    .data_out(\data[251] ),
    .latch_enable_in(\latch[250] ),
    .latch_enable_out(\latch[251] ),
    .scan_select_in(\scan[250] ),
    .scan_select_out(\scan[251] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_251 (.clk_in(\clk[251] ),
    .clk_out(\clk[252] ),
    .data_in(\data[251] ),
    .data_out(\data[252] ),
    .latch_enable_in(\latch[251] ),
    .latch_enable_out(\latch[252] ),
    .scan_select_in(\scan[251] ),
    .scan_select_out(\scan[252] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_252 (.clk_in(\clk[252] ),
    .clk_out(\clk[253] ),
    .data_in(\data[252] ),
    .data_out(\data[253] ),
    .latch_enable_in(\latch[252] ),
    .latch_enable_out(\latch[253] ),
    .scan_select_in(\scan[252] ),
    .scan_select_out(\scan[253] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_253 (.clk_in(\clk[253] ),
    .clk_out(\clk[254] ),
    .data_in(\data[253] ),
    .data_out(\data[254] ),
    .latch_enable_in(\latch[253] ),
    .latch_enable_out(\latch[254] ),
    .scan_select_in(\scan[253] ),
    .scan_select_out(\scan[254] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_254 (.clk_in(\clk[254] ),
    .clk_out(\clk[255] ),
    .data_in(\data[254] ),
    .data_out(\data[255] ),
    .latch_enable_in(\latch[254] ),
    .latch_enable_out(\latch[255] ),
    .scan_select_in(\scan[254] ),
    .scan_select_out(\scan[255] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_255 (.clk_in(\clk[255] ),
    .clk_out(\clk[256] ),
    .data_in(\data[255] ),
    .data_out(\data[256] ),
    .latch_enable_in(\latch[255] ),
    .latch_enable_out(\latch[256] ),
    .scan_select_in(\scan[255] ),
    .scan_select_out(\scan[256] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_256 (.clk_in(\clk[256] ),
    .clk_out(\clk[257] ),
    .data_in(\data[256] ),
    .data_out(\data[257] ),
    .latch_enable_in(\latch[256] ),
    .latch_enable_out(\latch[257] ),
    .scan_select_in(\scan[256] ),
    .scan_select_out(\scan[257] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_257 (.clk_in(\clk[257] ),
    .clk_out(\clk[258] ),
    .data_in(\data[257] ),
    .data_out(\data[258] ),
    .latch_enable_in(\latch[257] ),
    .latch_enable_out(\latch[258] ),
    .scan_select_in(\scan[257] ),
    .scan_select_out(\scan[258] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_258 (.clk_in(\clk[258] ),
    .clk_out(\clk[259] ),
    .data_in(\data[258] ),
    .data_out(\data[259] ),
    .latch_enable_in(\latch[258] ),
    .latch_enable_out(\latch[259] ),
    .scan_select_in(\scan[258] ),
    .scan_select_out(\scan[259] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_259 (.clk_in(\clk[259] ),
    .clk_out(\clk[260] ),
    .data_in(\data[259] ),
    .data_out(\data[260] ),
    .latch_enable_in(\latch[259] ),
    .latch_enable_out(\latch[260] ),
    .scan_select_in(\scan[259] ),
    .scan_select_out(\scan[260] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_26 (.clk_in(\clk[26] ),
    .clk_out(\clk[27] ),
    .data_in(\data[26] ),
    .data_out(\data[27] ),
    .latch_enable_in(\latch[26] ),
    .latch_enable_out(\latch[27] ),
    .scan_select_in(\scan[26] ),
    .scan_select_out(\scan[27] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_260 (.clk_in(\clk[260] ),
    .clk_out(\clk[261] ),
    .data_in(\data[260] ),
    .data_out(\data[261] ),
    .latch_enable_in(\latch[260] ),
    .latch_enable_out(\latch[261] ),
    .scan_select_in(\scan[260] ),
    .scan_select_out(\scan[261] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_261 (.clk_in(\clk[261] ),
    .clk_out(\clk[262] ),
    .data_in(\data[261] ),
    .data_out(\data[262] ),
    .latch_enable_in(\latch[261] ),
    .latch_enable_out(\latch[262] ),
    .scan_select_in(\scan[261] ),
    .scan_select_out(\scan[262] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_262 (.clk_in(\clk[262] ),
    .clk_out(\clk[263] ),
    .data_in(\data[262] ),
    .data_out(\data[263] ),
    .latch_enable_in(\latch[262] ),
    .latch_enable_out(\latch[263] ),
    .scan_select_in(\scan[262] ),
    .scan_select_out(\scan[263] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_263 (.clk_in(\clk[263] ),
    .clk_out(\clk[264] ),
    .data_in(\data[263] ),
    .data_out(\data[264] ),
    .latch_enable_in(\latch[263] ),
    .latch_enable_out(\latch[264] ),
    .scan_select_in(\scan[263] ),
    .scan_select_out(\scan[264] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_264 (.clk_in(\clk[264] ),
    .clk_out(\clk[265] ),
    .data_in(\data[264] ),
    .data_out(\data[265] ),
    .latch_enable_in(\latch[264] ),
    .latch_enable_out(\latch[265] ),
    .scan_select_in(\scan[264] ),
    .scan_select_out(\scan[265] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_265 (.clk_in(\clk[265] ),
    .clk_out(\clk[266] ),
    .data_in(\data[265] ),
    .data_out(\data[266] ),
    .latch_enable_in(\latch[265] ),
    .latch_enable_out(\latch[266] ),
    .scan_select_in(\scan[265] ),
    .scan_select_out(\scan[266] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_266 (.clk_in(\clk[266] ),
    .clk_out(\clk[267] ),
    .data_in(\data[266] ),
    .data_out(\data[267] ),
    .latch_enable_in(\latch[266] ),
    .latch_enable_out(\latch[267] ),
    .scan_select_in(\scan[266] ),
    .scan_select_out(\scan[267] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_267 (.clk_in(\clk[267] ),
    .clk_out(\clk[268] ),
    .data_in(\data[267] ),
    .data_out(\data[268] ),
    .latch_enable_in(\latch[267] ),
    .latch_enable_out(\latch[268] ),
    .scan_select_in(\scan[267] ),
    .scan_select_out(\scan[268] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_268 (.clk_in(\clk[268] ),
    .clk_out(\clk[269] ),
    .data_in(\data[268] ),
    .data_out(\data[269] ),
    .latch_enable_in(\latch[268] ),
    .latch_enable_out(\latch[269] ),
    .scan_select_in(\scan[268] ),
    .scan_select_out(\scan[269] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_269 (.clk_in(\clk[269] ),
    .clk_out(\clk[270] ),
    .data_in(\data[269] ),
    .data_out(\data[270] ),
    .latch_enable_in(\latch[269] ),
    .latch_enable_out(\latch[270] ),
    .scan_select_in(\scan[269] ),
    .scan_select_out(\scan[270] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_27 (.clk_in(\clk[27] ),
    .clk_out(\clk[28] ),
    .data_in(\data[27] ),
    .data_out(\data[28] ),
    .latch_enable_in(\latch[27] ),
    .latch_enable_out(\latch[28] ),
    .scan_select_in(\scan[27] ),
    .scan_select_out(\scan[28] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_270 (.clk_in(\clk[270] ),
    .clk_out(\clk[271] ),
    .data_in(\data[270] ),
    .data_out(\data[271] ),
    .latch_enable_in(\latch[270] ),
    .latch_enable_out(\latch[271] ),
    .scan_select_in(\scan[270] ),
    .scan_select_out(\scan[271] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_271 (.clk_in(\clk[271] ),
    .clk_out(\clk[272] ),
    .data_in(\data[271] ),
    .data_out(\data[272] ),
    .latch_enable_in(\latch[271] ),
    .latch_enable_out(\latch[272] ),
    .scan_select_in(\scan[271] ),
    .scan_select_out(\scan[272] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_272 (.clk_in(\clk[272] ),
    .clk_out(\clk[273] ),
    .data_in(\data[272] ),
    .data_out(\data[273] ),
    .latch_enable_in(\latch[272] ),
    .latch_enable_out(\latch[273] ),
    .scan_select_in(\scan[272] ),
    .scan_select_out(\scan[273] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_273 (.clk_in(\clk[273] ),
    .clk_out(\clk[274] ),
    .data_in(\data[273] ),
    .data_out(\data[274] ),
    .latch_enable_in(\latch[273] ),
    .latch_enable_out(\latch[274] ),
    .scan_select_in(\scan[273] ),
    .scan_select_out(\scan[274] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_274 (.clk_in(\clk[274] ),
    .clk_out(\clk[275] ),
    .data_in(\data[274] ),
    .data_out(\data[275] ),
    .latch_enable_in(\latch[274] ),
    .latch_enable_out(\latch[275] ),
    .scan_select_in(\scan[274] ),
    .scan_select_out(\scan[275] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_275 (.clk_in(\clk[275] ),
    .clk_out(\clk[276] ),
    .data_in(\data[275] ),
    .data_out(\data[276] ),
    .latch_enable_in(\latch[275] ),
    .latch_enable_out(\latch[276] ),
    .scan_select_in(\scan[275] ),
    .scan_select_out(\scan[276] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_276 (.clk_in(\clk[276] ),
    .clk_out(\clk[277] ),
    .data_in(\data[276] ),
    .data_out(\data[277] ),
    .latch_enable_in(\latch[276] ),
    .latch_enable_out(\latch[277] ),
    .scan_select_in(\scan[276] ),
    .scan_select_out(\scan[277] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_277 (.clk_in(\clk[277] ),
    .clk_out(\clk[278] ),
    .data_in(\data[277] ),
    .data_out(\data[278] ),
    .latch_enable_in(\latch[277] ),
    .latch_enable_out(\latch[278] ),
    .scan_select_in(\scan[277] ),
    .scan_select_out(\scan[278] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_278 (.clk_in(\clk[278] ),
    .clk_out(\clk[279] ),
    .data_in(\data[278] ),
    .data_out(\data[279] ),
    .latch_enable_in(\latch[278] ),
    .latch_enable_out(\latch[279] ),
    .scan_select_in(\scan[278] ),
    .scan_select_out(\scan[279] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_279 (.clk_in(\clk[279] ),
    .clk_out(\clk[280] ),
    .data_in(\data[279] ),
    .data_out(\data[280] ),
    .latch_enable_in(\latch[279] ),
    .latch_enable_out(\latch[280] ),
    .scan_select_in(\scan[279] ),
    .scan_select_out(\scan[280] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_28 (.clk_in(\clk[28] ),
    .clk_out(\clk[29] ),
    .data_in(\data[28] ),
    .data_out(\data[29] ),
    .latch_enable_in(\latch[28] ),
    .latch_enable_out(\latch[29] ),
    .scan_select_in(\scan[28] ),
    .scan_select_out(\scan[29] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_280 (.clk_in(\clk[280] ),
    .clk_out(\clk[281] ),
    .data_in(\data[280] ),
    .data_out(\data[281] ),
    .latch_enable_in(\latch[280] ),
    .latch_enable_out(\latch[281] ),
    .scan_select_in(\scan[280] ),
    .scan_select_out(\scan[281] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_281 (.clk_in(\clk[281] ),
    .clk_out(\clk[282] ),
    .data_in(\data[281] ),
    .data_out(\data[282] ),
    .latch_enable_in(\latch[281] ),
    .latch_enable_out(\latch[282] ),
    .scan_select_in(\scan[281] ),
    .scan_select_out(\scan[282] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_282 (.clk_in(\clk[282] ),
    .clk_out(\clk[283] ),
    .data_in(\data[282] ),
    .data_out(\data[283] ),
    .latch_enable_in(\latch[282] ),
    .latch_enable_out(\latch[283] ),
    .scan_select_in(\scan[282] ),
    .scan_select_out(\scan[283] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_283 (.clk_in(\clk[283] ),
    .clk_out(\clk[284] ),
    .data_in(\data[283] ),
    .data_out(\data[284] ),
    .latch_enable_in(\latch[283] ),
    .latch_enable_out(\latch[284] ),
    .scan_select_in(\scan[283] ),
    .scan_select_out(\scan[284] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_284 (.clk_in(\clk[284] ),
    .clk_out(\clk[285] ),
    .data_in(\data[284] ),
    .data_out(\data[285] ),
    .latch_enable_in(\latch[284] ),
    .latch_enable_out(\latch[285] ),
    .scan_select_in(\scan[284] ),
    .scan_select_out(\scan[285] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_285 (.clk_in(\clk[285] ),
    .clk_out(\clk[286] ),
    .data_in(\data[285] ),
    .data_out(\data[286] ),
    .latch_enable_in(\latch[285] ),
    .latch_enable_out(\latch[286] ),
    .scan_select_in(\scan[285] ),
    .scan_select_out(\scan[286] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_286 (.clk_in(\clk[286] ),
    .clk_out(\clk[287] ),
    .data_in(\data[286] ),
    .data_out(\data[287] ),
    .latch_enable_in(\latch[286] ),
    .latch_enable_out(\latch[287] ),
    .scan_select_in(\scan[286] ),
    .scan_select_out(\scan[287] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_287 (.clk_in(\clk[287] ),
    .clk_out(\clk[288] ),
    .data_in(\data[287] ),
    .data_out(\data[288] ),
    .latch_enable_in(\latch[287] ),
    .latch_enable_out(\latch[288] ),
    .scan_select_in(\scan[287] ),
    .scan_select_out(\scan[288] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_288 (.clk_in(\clk[288] ),
    .clk_out(\clk[289] ),
    .data_in(\data[288] ),
    .data_out(\data[289] ),
    .latch_enable_in(\latch[288] ),
    .latch_enable_out(\latch[289] ),
    .scan_select_in(\scan[288] ),
    .scan_select_out(\scan[289] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_289 (.clk_in(\clk[289] ),
    .clk_out(\clk[290] ),
    .data_in(\data[289] ),
    .data_out(\data[290] ),
    .latch_enable_in(\latch[289] ),
    .latch_enable_out(\latch[290] ),
    .scan_select_in(\scan[289] ),
    .scan_select_out(\scan[290] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_29 (.clk_in(\clk[29] ),
    .clk_out(\clk[30] ),
    .data_in(\data[29] ),
    .data_out(\data[30] ),
    .latch_enable_in(\latch[29] ),
    .latch_enable_out(\latch[30] ),
    .scan_select_in(\scan[29] ),
    .scan_select_out(\scan[30] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_290 (.clk_in(\clk[290] ),
    .clk_out(\clk[291] ),
    .data_in(\data[290] ),
    .data_out(\data[291] ),
    .latch_enable_in(\latch[290] ),
    .latch_enable_out(\latch[291] ),
    .scan_select_in(\scan[290] ),
    .scan_select_out(\scan[291] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_291 (.clk_in(\clk[291] ),
    .clk_out(\clk[292] ),
    .data_in(\data[291] ),
    .data_out(\data[292] ),
    .latch_enable_in(\latch[291] ),
    .latch_enable_out(\latch[292] ),
    .scan_select_in(\scan[291] ),
    .scan_select_out(\scan[292] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_292 (.clk_in(\clk[292] ),
    .clk_out(\clk[293] ),
    .data_in(\data[292] ),
    .data_out(\data[293] ),
    .latch_enable_in(\latch[292] ),
    .latch_enable_out(\latch[293] ),
    .scan_select_in(\scan[292] ),
    .scan_select_out(\scan[293] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_293 (.clk_in(\clk[293] ),
    .clk_out(\clk[294] ),
    .data_in(\data[293] ),
    .data_out(\data[294] ),
    .latch_enable_in(\latch[293] ),
    .latch_enable_out(\latch[294] ),
    .scan_select_in(\scan[293] ),
    .scan_select_out(\scan[294] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_294 (.clk_in(\clk[294] ),
    .clk_out(\clk[295] ),
    .data_in(\data[294] ),
    .data_out(\data[295] ),
    .latch_enable_in(\latch[294] ),
    .latch_enable_out(\latch[295] ),
    .scan_select_in(\scan[294] ),
    .scan_select_out(\scan[295] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_295 (.clk_in(\clk[295] ),
    .clk_out(\clk[296] ),
    .data_in(\data[295] ),
    .data_out(\data[296] ),
    .latch_enable_in(\latch[295] ),
    .latch_enable_out(\latch[296] ),
    .scan_select_in(\scan[295] ),
    .scan_select_out(\scan[296] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_296 (.clk_in(\clk[296] ),
    .clk_out(\clk[297] ),
    .data_in(\data[296] ),
    .data_out(\data[297] ),
    .latch_enable_in(\latch[296] ),
    .latch_enable_out(\latch[297] ),
    .scan_select_in(\scan[296] ),
    .scan_select_out(\scan[297] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_297 (.clk_in(\clk[297] ),
    .clk_out(\clk[298] ),
    .data_in(\data[297] ),
    .data_out(\data[298] ),
    .latch_enable_in(\latch[297] ),
    .latch_enable_out(\latch[298] ),
    .scan_select_in(\scan[297] ),
    .scan_select_out(\scan[298] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_298 (.clk_in(\clk[298] ),
    .clk_out(\clk[299] ),
    .data_in(\data[298] ),
    .data_out(\data[299] ),
    .latch_enable_in(\latch[298] ),
    .latch_enable_out(\latch[299] ),
    .scan_select_in(\scan[298] ),
    .scan_select_out(\scan[299] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_299 (.clk_in(\clk[299] ),
    .clk_out(\clk[300] ),
    .data_in(\data[299] ),
    .data_out(\data[300] ),
    .latch_enable_in(\latch[299] ),
    .latch_enable_out(\latch[300] ),
    .scan_select_in(\scan[299] ),
    .scan_select_out(\scan[300] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_30 (.clk_in(\clk[30] ),
    .clk_out(\clk[31] ),
    .data_in(\data[30] ),
    .data_out(\data[31] ),
    .latch_enable_in(\latch[30] ),
    .latch_enable_out(\latch[31] ),
    .scan_select_in(\scan[30] ),
    .scan_select_out(\scan[31] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_300 (.clk_in(\clk[300] ),
    .clk_out(\clk[301] ),
    .data_in(\data[300] ),
    .data_out(\data[301] ),
    .latch_enable_in(\latch[300] ),
    .latch_enable_out(\latch[301] ),
    .scan_select_in(\scan[300] ),
    .scan_select_out(\scan[301] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_301 (.clk_in(\clk[301] ),
    .clk_out(\clk[302] ),
    .data_in(\data[301] ),
    .data_out(\data[302] ),
    .latch_enable_in(\latch[301] ),
    .latch_enable_out(\latch[302] ),
    .scan_select_in(\scan[301] ),
    .scan_select_out(\scan[302] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_302 (.clk_in(\clk[302] ),
    .clk_out(\clk[303] ),
    .data_in(\data[302] ),
    .data_out(\data[303] ),
    .latch_enable_in(\latch[302] ),
    .latch_enable_out(\latch[303] ),
    .scan_select_in(\scan[302] ),
    .scan_select_out(\scan[303] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_303 (.clk_in(\clk[303] ),
    .clk_out(\clk[304] ),
    .data_in(\data[303] ),
    .data_out(\data[304] ),
    .latch_enable_in(\latch[303] ),
    .latch_enable_out(\latch[304] ),
    .scan_select_in(\scan[303] ),
    .scan_select_out(\scan[304] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_304 (.clk_in(\clk[304] ),
    .clk_out(\clk[305] ),
    .data_in(\data[304] ),
    .data_out(\data[305] ),
    .latch_enable_in(\latch[304] ),
    .latch_enable_out(\latch[305] ),
    .scan_select_in(\scan[304] ),
    .scan_select_out(\scan[305] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_305 (.clk_in(\clk[305] ),
    .clk_out(\clk[306] ),
    .data_in(\data[305] ),
    .data_out(\data[306] ),
    .latch_enable_in(\latch[305] ),
    .latch_enable_out(\latch[306] ),
    .scan_select_in(\scan[305] ),
    .scan_select_out(\scan[306] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_306 (.clk_in(\clk[306] ),
    .clk_out(\clk[307] ),
    .data_in(\data[306] ),
    .data_out(\data[307] ),
    .latch_enable_in(\latch[306] ),
    .latch_enable_out(\latch[307] ),
    .scan_select_in(\scan[306] ),
    .scan_select_out(\scan[307] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_307 (.clk_in(\clk[307] ),
    .clk_out(\clk[308] ),
    .data_in(\data[307] ),
    .data_out(\data[308] ),
    .latch_enable_in(\latch[307] ),
    .latch_enable_out(\latch[308] ),
    .scan_select_in(\scan[307] ),
    .scan_select_out(\scan[308] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_308 (.clk_in(\clk[308] ),
    .clk_out(\clk[309] ),
    .data_in(\data[308] ),
    .data_out(\data[309] ),
    .latch_enable_in(\latch[308] ),
    .latch_enable_out(\latch[309] ),
    .scan_select_in(\scan[308] ),
    .scan_select_out(\scan[309] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_309 (.clk_in(\clk[309] ),
    .clk_out(\clk[310] ),
    .data_in(\data[309] ),
    .data_out(\data[310] ),
    .latch_enable_in(\latch[309] ),
    .latch_enable_out(\latch[310] ),
    .scan_select_in(\scan[309] ),
    .scan_select_out(\scan[310] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_31 (.clk_in(\clk[31] ),
    .clk_out(\clk[32] ),
    .data_in(\data[31] ),
    .data_out(\data[32] ),
    .latch_enable_in(\latch[31] ),
    .latch_enable_out(\latch[32] ),
    .scan_select_in(\scan[31] ),
    .scan_select_out(\scan[32] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_310 (.clk_in(\clk[310] ),
    .clk_out(\clk[311] ),
    .data_in(\data[310] ),
    .data_out(\data[311] ),
    .latch_enable_in(\latch[310] ),
    .latch_enable_out(\latch[311] ),
    .scan_select_in(\scan[310] ),
    .scan_select_out(\scan[311] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_311 (.clk_in(\clk[311] ),
    .clk_out(\clk[312] ),
    .data_in(\data[311] ),
    .data_out(\data[312] ),
    .latch_enable_in(\latch[311] ),
    .latch_enable_out(\latch[312] ),
    .scan_select_in(\scan[311] ),
    .scan_select_out(\scan[312] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_312 (.clk_in(\clk[312] ),
    .clk_out(\clk[313] ),
    .data_in(\data[312] ),
    .data_out(\data[313] ),
    .latch_enable_in(\latch[312] ),
    .latch_enable_out(\latch[313] ),
    .scan_select_in(\scan[312] ),
    .scan_select_out(\scan[313] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_313 (.clk_in(\clk[313] ),
    .clk_out(\clk[314] ),
    .data_in(\data[313] ),
    .data_out(\data[314] ),
    .latch_enable_in(\latch[313] ),
    .latch_enable_out(\latch[314] ),
    .scan_select_in(\scan[313] ),
    .scan_select_out(\scan[314] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_314 (.clk_in(\clk[314] ),
    .clk_out(\clk[315] ),
    .data_in(\data[314] ),
    .data_out(\data[315] ),
    .latch_enable_in(\latch[314] ),
    .latch_enable_out(\latch[315] ),
    .scan_select_in(\scan[314] ),
    .scan_select_out(\scan[315] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_315 (.clk_in(\clk[315] ),
    .clk_out(\clk[316] ),
    .data_in(\data[315] ),
    .data_out(\data[316] ),
    .latch_enable_in(\latch[315] ),
    .latch_enable_out(\latch[316] ),
    .scan_select_in(\scan[315] ),
    .scan_select_out(\scan[316] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_316 (.clk_in(\clk[316] ),
    .clk_out(\clk[317] ),
    .data_in(\data[316] ),
    .data_out(\data[317] ),
    .latch_enable_in(\latch[316] ),
    .latch_enable_out(\latch[317] ),
    .scan_select_in(\scan[316] ),
    .scan_select_out(\scan[317] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_317 (.clk_in(\clk[317] ),
    .clk_out(\clk[318] ),
    .data_in(\data[317] ),
    .data_out(\data[318] ),
    .latch_enable_in(\latch[317] ),
    .latch_enable_out(\latch[318] ),
    .scan_select_in(\scan[317] ),
    .scan_select_out(\scan[318] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_318 (.clk_in(\clk[318] ),
    .clk_out(\clk[319] ),
    .data_in(\data[318] ),
    .data_out(\data[319] ),
    .latch_enable_in(\latch[318] ),
    .latch_enable_out(\latch[319] ),
    .scan_select_in(\scan[318] ),
    .scan_select_out(\scan[319] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_319 (.clk_in(\clk[319] ),
    .clk_out(\clk[320] ),
    .data_in(\data[319] ),
    .data_out(\data[320] ),
    .latch_enable_in(\latch[319] ),
    .latch_enable_out(\latch[320] ),
    .scan_select_in(\scan[319] ),
    .scan_select_out(\scan[320] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_32 (.clk_in(\clk[32] ),
    .clk_out(\clk[33] ),
    .data_in(\data[32] ),
    .data_out(\data[33] ),
    .latch_enable_in(\latch[32] ),
    .latch_enable_out(\latch[33] ),
    .scan_select_in(\scan[32] ),
    .scan_select_out(\scan[33] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_320 (.clk_in(\clk[320] ),
    .clk_out(\clk[321] ),
    .data_in(\data[320] ),
    .data_out(\data[321] ),
    .latch_enable_in(\latch[320] ),
    .latch_enable_out(\latch[321] ),
    .scan_select_in(\scan[320] ),
    .scan_select_out(\scan[321] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_321 (.clk_in(\clk[321] ),
    .clk_out(\clk[322] ),
    .data_in(\data[321] ),
    .data_out(\data[322] ),
    .latch_enable_in(\latch[321] ),
    .latch_enable_out(\latch[322] ),
    .scan_select_in(\scan[321] ),
    .scan_select_out(\scan[322] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_322 (.clk_in(\clk[322] ),
    .clk_out(\clk[323] ),
    .data_in(\data[322] ),
    .data_out(\data[323] ),
    .latch_enable_in(\latch[322] ),
    .latch_enable_out(\latch[323] ),
    .scan_select_in(\scan[322] ),
    .scan_select_out(\scan[323] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_323 (.clk_in(\clk[323] ),
    .clk_out(\clk[324] ),
    .data_in(\data[323] ),
    .data_out(\data[324] ),
    .latch_enable_in(\latch[323] ),
    .latch_enable_out(\latch[324] ),
    .scan_select_in(\scan[323] ),
    .scan_select_out(\scan[324] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_324 (.clk_in(\clk[324] ),
    .clk_out(\clk[325] ),
    .data_in(\data[324] ),
    .data_out(\data[325] ),
    .latch_enable_in(\latch[324] ),
    .latch_enable_out(\latch[325] ),
    .scan_select_in(\scan[324] ),
    .scan_select_out(\scan[325] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_325 (.clk_in(\clk[325] ),
    .clk_out(\clk[326] ),
    .data_in(\data[325] ),
    .data_out(\data[326] ),
    .latch_enable_in(\latch[325] ),
    .latch_enable_out(\latch[326] ),
    .scan_select_in(\scan[325] ),
    .scan_select_out(\scan[326] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_326 (.clk_in(\clk[326] ),
    .clk_out(\clk[327] ),
    .data_in(\data[326] ),
    .data_out(\data[327] ),
    .latch_enable_in(\latch[326] ),
    .latch_enable_out(\latch[327] ),
    .scan_select_in(\scan[326] ),
    .scan_select_out(\scan[327] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_327 (.clk_in(\clk[327] ),
    .clk_out(\clk[328] ),
    .data_in(\data[327] ),
    .data_out(\data[328] ),
    .latch_enable_in(\latch[327] ),
    .latch_enable_out(\latch[328] ),
    .scan_select_in(\scan[327] ),
    .scan_select_out(\scan[328] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_328 (.clk_in(\clk[328] ),
    .clk_out(\clk[329] ),
    .data_in(\data[328] ),
    .data_out(\data[329] ),
    .latch_enable_in(\latch[328] ),
    .latch_enable_out(\latch[329] ),
    .scan_select_in(\scan[328] ),
    .scan_select_out(\scan[329] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_329 (.clk_in(\clk[329] ),
    .clk_out(\clk[330] ),
    .data_in(\data[329] ),
    .data_out(\data[330] ),
    .latch_enable_in(\latch[329] ),
    .latch_enable_out(\latch[330] ),
    .scan_select_in(\scan[329] ),
    .scan_select_out(\scan[330] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_33 (.clk_in(\clk[33] ),
    .clk_out(\clk[34] ),
    .data_in(\data[33] ),
    .data_out(\data[34] ),
    .latch_enable_in(\latch[33] ),
    .latch_enable_out(\latch[34] ),
    .scan_select_in(\scan[33] ),
    .scan_select_out(\scan[34] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_330 (.clk_in(\clk[330] ),
    .clk_out(\clk[331] ),
    .data_in(\data[330] ),
    .data_out(\data[331] ),
    .latch_enable_in(\latch[330] ),
    .latch_enable_out(\latch[331] ),
    .scan_select_in(\scan[330] ),
    .scan_select_out(\scan[331] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_331 (.clk_in(\clk[331] ),
    .clk_out(\clk[332] ),
    .data_in(\data[331] ),
    .data_out(\data[332] ),
    .latch_enable_in(\latch[331] ),
    .latch_enable_out(\latch[332] ),
    .scan_select_in(\scan[331] ),
    .scan_select_out(\scan[332] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_332 (.clk_in(\clk[332] ),
    .clk_out(\clk[333] ),
    .data_in(\data[332] ),
    .data_out(\data[333] ),
    .latch_enable_in(\latch[332] ),
    .latch_enable_out(\latch[333] ),
    .scan_select_in(\scan[332] ),
    .scan_select_out(\scan[333] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_333 (.clk_in(\clk[333] ),
    .clk_out(\clk[334] ),
    .data_in(\data[333] ),
    .data_out(\data[334] ),
    .latch_enable_in(\latch[333] ),
    .latch_enable_out(\latch[334] ),
    .scan_select_in(\scan[333] ),
    .scan_select_out(\scan[334] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_334 (.clk_in(\clk[334] ),
    .clk_out(\clk[335] ),
    .data_in(\data[334] ),
    .data_out(\data[335] ),
    .latch_enable_in(\latch[334] ),
    .latch_enable_out(\latch[335] ),
    .scan_select_in(\scan[334] ),
    .scan_select_out(\scan[335] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_335 (.clk_in(\clk[335] ),
    .clk_out(\clk[336] ),
    .data_in(\data[335] ),
    .data_out(\data[336] ),
    .latch_enable_in(\latch[335] ),
    .latch_enable_out(\latch[336] ),
    .scan_select_in(\scan[335] ),
    .scan_select_out(\scan[336] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_336 (.clk_in(\clk[336] ),
    .clk_out(\clk[337] ),
    .data_in(\data[336] ),
    .data_out(\data[337] ),
    .latch_enable_in(\latch[336] ),
    .latch_enable_out(\latch[337] ),
    .scan_select_in(\scan[336] ),
    .scan_select_out(\scan[337] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_337 (.clk_in(\clk[337] ),
    .clk_out(\clk[338] ),
    .data_in(\data[337] ),
    .data_out(\data[338] ),
    .latch_enable_in(\latch[337] ),
    .latch_enable_out(\latch[338] ),
    .scan_select_in(\scan[337] ),
    .scan_select_out(\scan[338] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_338 (.clk_in(\clk[338] ),
    .clk_out(\clk[339] ),
    .data_in(\data[338] ),
    .data_out(\data[339] ),
    .latch_enable_in(\latch[338] ),
    .latch_enable_out(\latch[339] ),
    .scan_select_in(\scan[338] ),
    .scan_select_out(\scan[339] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_339 (.clk_in(\clk[339] ),
    .clk_out(\clk[340] ),
    .data_in(\data[339] ),
    .data_out(\data[340] ),
    .latch_enable_in(\latch[339] ),
    .latch_enable_out(\latch[340] ),
    .scan_select_in(\scan[339] ),
    .scan_select_out(\scan[340] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_34 (.clk_in(\clk[34] ),
    .clk_out(\clk[35] ),
    .data_in(\data[34] ),
    .data_out(\data[35] ),
    .latch_enable_in(\latch[34] ),
    .latch_enable_out(\latch[35] ),
    .scan_select_in(\scan[34] ),
    .scan_select_out(\scan[35] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_340 (.clk_in(\clk[340] ),
    .clk_out(\clk[341] ),
    .data_in(\data[340] ),
    .data_out(\data[341] ),
    .latch_enable_in(\latch[340] ),
    .latch_enable_out(\latch[341] ),
    .scan_select_in(\scan[340] ),
    .scan_select_out(\scan[341] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_341 (.clk_in(\clk[341] ),
    .clk_out(\clk[342] ),
    .data_in(\data[341] ),
    .data_out(\data[342] ),
    .latch_enable_in(\latch[341] ),
    .latch_enable_out(\latch[342] ),
    .scan_select_in(\scan[341] ),
    .scan_select_out(\scan[342] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_342 (.clk_in(\clk[342] ),
    .clk_out(\clk[343] ),
    .data_in(\data[342] ),
    .data_out(\data[343] ),
    .latch_enable_in(\latch[342] ),
    .latch_enable_out(\latch[343] ),
    .scan_select_in(\scan[342] ),
    .scan_select_out(\scan[343] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_343 (.clk_in(\clk[343] ),
    .clk_out(\clk[344] ),
    .data_in(\data[343] ),
    .data_out(\data[344] ),
    .latch_enable_in(\latch[343] ),
    .latch_enable_out(\latch[344] ),
    .scan_select_in(\scan[343] ),
    .scan_select_out(\scan[344] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_344 (.clk_in(\clk[344] ),
    .clk_out(\clk[345] ),
    .data_in(\data[344] ),
    .data_out(\data[345] ),
    .latch_enable_in(\latch[344] ),
    .latch_enable_out(\latch[345] ),
    .scan_select_in(\scan[344] ),
    .scan_select_out(\scan[345] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_345 (.clk_in(\clk[345] ),
    .clk_out(\clk[346] ),
    .data_in(\data[345] ),
    .data_out(\data[346] ),
    .latch_enable_in(\latch[345] ),
    .latch_enable_out(\latch[346] ),
    .scan_select_in(\scan[345] ),
    .scan_select_out(\scan[346] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_346 (.clk_in(\clk[346] ),
    .clk_out(\clk[347] ),
    .data_in(\data[346] ),
    .data_out(\data[347] ),
    .latch_enable_in(\latch[346] ),
    .latch_enable_out(\latch[347] ),
    .scan_select_in(\scan[346] ),
    .scan_select_out(\scan[347] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_347 (.clk_in(\clk[347] ),
    .clk_out(\clk[348] ),
    .data_in(\data[347] ),
    .data_out(\data[348] ),
    .latch_enable_in(\latch[347] ),
    .latch_enable_out(\latch[348] ),
    .scan_select_in(\scan[347] ),
    .scan_select_out(\scan[348] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_348 (.clk_in(\clk[348] ),
    .clk_out(\clk[349] ),
    .data_in(\data[348] ),
    .data_out(\data[349] ),
    .latch_enable_in(\latch[348] ),
    .latch_enable_out(\latch[349] ),
    .scan_select_in(\scan[348] ),
    .scan_select_out(\scan[349] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_349 (.clk_in(\clk[349] ),
    .clk_out(\clk[350] ),
    .data_in(\data[349] ),
    .data_out(\data[350] ),
    .latch_enable_in(\latch[349] ),
    .latch_enable_out(\latch[350] ),
    .scan_select_in(\scan[349] ),
    .scan_select_out(\scan[350] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_35 (.clk_in(\clk[35] ),
    .clk_out(\clk[36] ),
    .data_in(\data[35] ),
    .data_out(\data[36] ),
    .latch_enable_in(\latch[35] ),
    .latch_enable_out(\latch[36] ),
    .scan_select_in(\scan[35] ),
    .scan_select_out(\scan[36] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_350 (.clk_in(\clk[350] ),
    .clk_out(\clk[351] ),
    .data_in(\data[350] ),
    .data_out(\data[351] ),
    .latch_enable_in(\latch[350] ),
    .latch_enable_out(\latch[351] ),
    .scan_select_in(\scan[350] ),
    .scan_select_out(\scan[351] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_351 (.clk_in(\clk[351] ),
    .clk_out(\clk[352] ),
    .data_in(\data[351] ),
    .data_out(\data[352] ),
    .latch_enable_in(\latch[351] ),
    .latch_enable_out(\latch[352] ),
    .scan_select_in(\scan[351] ),
    .scan_select_out(\scan[352] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_352 (.clk_in(\clk[352] ),
    .clk_out(\clk[353] ),
    .data_in(\data[352] ),
    .data_out(\data[353] ),
    .latch_enable_in(\latch[352] ),
    .latch_enable_out(\latch[353] ),
    .scan_select_in(\scan[352] ),
    .scan_select_out(\scan[353] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_353 (.clk_in(\clk[353] ),
    .clk_out(\clk[354] ),
    .data_in(\data[353] ),
    .data_out(\data[354] ),
    .latch_enable_in(\latch[353] ),
    .latch_enable_out(\latch[354] ),
    .scan_select_in(\scan[353] ),
    .scan_select_out(\scan[354] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_354 (.clk_in(\clk[354] ),
    .clk_out(\clk[355] ),
    .data_in(\data[354] ),
    .data_out(\data[355] ),
    .latch_enable_in(\latch[354] ),
    .latch_enable_out(\latch[355] ),
    .scan_select_in(\scan[354] ),
    .scan_select_out(\scan[355] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_355 (.clk_in(\clk[355] ),
    .clk_out(\clk[356] ),
    .data_in(\data[355] ),
    .data_out(\data[356] ),
    .latch_enable_in(\latch[355] ),
    .latch_enable_out(\latch[356] ),
    .scan_select_in(\scan[355] ),
    .scan_select_out(\scan[356] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_356 (.clk_in(\clk[356] ),
    .clk_out(\clk[357] ),
    .data_in(\data[356] ),
    .data_out(\data[357] ),
    .latch_enable_in(\latch[356] ),
    .latch_enable_out(\latch[357] ),
    .scan_select_in(\scan[356] ),
    .scan_select_out(\scan[357] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_357 (.clk_in(\clk[357] ),
    .clk_out(\clk[358] ),
    .data_in(\data[357] ),
    .data_out(\data[358] ),
    .latch_enable_in(\latch[357] ),
    .latch_enable_out(\latch[358] ),
    .scan_select_in(\scan[357] ),
    .scan_select_out(\scan[358] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_358 (.clk_in(\clk[358] ),
    .clk_out(\clk[359] ),
    .data_in(\data[358] ),
    .data_out(\data[359] ),
    .latch_enable_in(\latch[358] ),
    .latch_enable_out(\latch[359] ),
    .scan_select_in(\scan[358] ),
    .scan_select_out(\scan[359] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_359 (.clk_in(\clk[359] ),
    .clk_out(\clk[360] ),
    .data_in(\data[359] ),
    .data_out(\data[360] ),
    .latch_enable_in(\latch[359] ),
    .latch_enable_out(\latch[360] ),
    .scan_select_in(\scan[359] ),
    .scan_select_out(\scan[360] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_36 (.clk_in(\clk[36] ),
    .clk_out(\clk[37] ),
    .data_in(\data[36] ),
    .data_out(\data[37] ),
    .latch_enable_in(\latch[36] ),
    .latch_enable_out(\latch[37] ),
    .scan_select_in(\scan[36] ),
    .scan_select_out(\scan[37] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_360 (.clk_in(\clk[360] ),
    .clk_out(\clk[361] ),
    .data_in(\data[360] ),
    .data_out(\data[361] ),
    .latch_enable_in(\latch[360] ),
    .latch_enable_out(\latch[361] ),
    .scan_select_in(\scan[360] ),
    .scan_select_out(\scan[361] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_361 (.clk_in(\clk[361] ),
    .clk_out(\clk[362] ),
    .data_in(\data[361] ),
    .data_out(\data[362] ),
    .latch_enable_in(\latch[361] ),
    .latch_enable_out(\latch[362] ),
    .scan_select_in(\scan[361] ),
    .scan_select_out(\scan[362] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_362 (.clk_in(\clk[362] ),
    .clk_out(\clk[363] ),
    .data_in(\data[362] ),
    .data_out(\data[363] ),
    .latch_enable_in(\latch[362] ),
    .latch_enable_out(\latch[363] ),
    .scan_select_in(\scan[362] ),
    .scan_select_out(\scan[363] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_363 (.clk_in(\clk[363] ),
    .clk_out(\clk[364] ),
    .data_in(\data[363] ),
    .data_out(\data[364] ),
    .latch_enable_in(\latch[363] ),
    .latch_enable_out(\latch[364] ),
    .scan_select_in(\scan[363] ),
    .scan_select_out(\scan[364] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_364 (.clk_in(\clk[364] ),
    .clk_out(\clk[365] ),
    .data_in(\data[364] ),
    .data_out(\data[365] ),
    .latch_enable_in(\latch[364] ),
    .latch_enable_out(\latch[365] ),
    .scan_select_in(\scan[364] ),
    .scan_select_out(\scan[365] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_365 (.clk_in(\clk[365] ),
    .clk_out(\clk[366] ),
    .data_in(\data[365] ),
    .data_out(\data[366] ),
    .latch_enable_in(\latch[365] ),
    .latch_enable_out(\latch[366] ),
    .scan_select_in(\scan[365] ),
    .scan_select_out(\scan[366] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_366 (.clk_in(\clk[366] ),
    .clk_out(\clk[367] ),
    .data_in(\data[366] ),
    .data_out(\data[367] ),
    .latch_enable_in(\latch[366] ),
    .latch_enable_out(\latch[367] ),
    .scan_select_in(\scan[366] ),
    .scan_select_out(\scan[367] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_367 (.clk_in(\clk[367] ),
    .clk_out(\clk[368] ),
    .data_in(\data[367] ),
    .data_out(\data[368] ),
    .latch_enable_in(\latch[367] ),
    .latch_enable_out(\latch[368] ),
    .scan_select_in(\scan[367] ),
    .scan_select_out(\scan[368] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_368 (.clk_in(\clk[368] ),
    .clk_out(\clk[369] ),
    .data_in(\data[368] ),
    .data_out(\data[369] ),
    .latch_enable_in(\latch[368] ),
    .latch_enable_out(\latch[369] ),
    .scan_select_in(\scan[368] ),
    .scan_select_out(\scan[369] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_369 (.clk_in(\clk[369] ),
    .clk_out(\clk[370] ),
    .data_in(\data[369] ),
    .data_out(\data[370] ),
    .latch_enable_in(\latch[369] ),
    .latch_enable_out(\latch[370] ),
    .scan_select_in(\scan[369] ),
    .scan_select_out(\scan[370] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_37 (.clk_in(\clk[37] ),
    .clk_out(\clk[38] ),
    .data_in(\data[37] ),
    .data_out(\data[38] ),
    .latch_enable_in(\latch[37] ),
    .latch_enable_out(\latch[38] ),
    .scan_select_in(\scan[37] ),
    .scan_select_out(\scan[38] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_370 (.clk_in(\clk[370] ),
    .clk_out(\clk[371] ),
    .data_in(\data[370] ),
    .data_out(\data[371] ),
    .latch_enable_in(\latch[370] ),
    .latch_enable_out(\latch[371] ),
    .scan_select_in(\scan[370] ),
    .scan_select_out(\scan[371] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_371 (.clk_in(\clk[371] ),
    .clk_out(\clk[372] ),
    .data_in(\data[371] ),
    .data_out(\data[372] ),
    .latch_enable_in(\latch[371] ),
    .latch_enable_out(\latch[372] ),
    .scan_select_in(\scan[371] ),
    .scan_select_out(\scan[372] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_372 (.clk_in(\clk[372] ),
    .clk_out(\clk[373] ),
    .data_in(\data[372] ),
    .data_out(\data[373] ),
    .latch_enable_in(\latch[372] ),
    .latch_enable_out(\latch[373] ),
    .scan_select_in(\scan[372] ),
    .scan_select_out(\scan[373] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_373 (.clk_in(\clk[373] ),
    .clk_out(\clk[374] ),
    .data_in(\data[373] ),
    .data_out(\data[374] ),
    .latch_enable_in(\latch[373] ),
    .latch_enable_out(\latch[374] ),
    .scan_select_in(\scan[373] ),
    .scan_select_out(\scan[374] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_374 (.clk_in(\clk[374] ),
    .clk_out(\clk[375] ),
    .data_in(\data[374] ),
    .data_out(\data[375] ),
    .latch_enable_in(\latch[374] ),
    .latch_enable_out(\latch[375] ),
    .scan_select_in(\scan[374] ),
    .scan_select_out(\scan[375] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_375 (.clk_in(\clk[375] ),
    .clk_out(\clk[376] ),
    .data_in(\data[375] ),
    .data_out(\data[376] ),
    .latch_enable_in(\latch[375] ),
    .latch_enable_out(\latch[376] ),
    .scan_select_in(\scan[375] ),
    .scan_select_out(\scan[376] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_376 (.clk_in(\clk[376] ),
    .clk_out(\clk[377] ),
    .data_in(\data[376] ),
    .data_out(\data[377] ),
    .latch_enable_in(\latch[376] ),
    .latch_enable_out(\latch[377] ),
    .scan_select_in(\scan[376] ),
    .scan_select_out(\scan[377] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_377 (.clk_in(\clk[377] ),
    .clk_out(\clk[378] ),
    .data_in(\data[377] ),
    .data_out(\data[378] ),
    .latch_enable_in(\latch[377] ),
    .latch_enable_out(\latch[378] ),
    .scan_select_in(\scan[377] ),
    .scan_select_out(\scan[378] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_378 (.clk_in(\clk[378] ),
    .clk_out(\clk[379] ),
    .data_in(\data[378] ),
    .data_out(\data[379] ),
    .latch_enable_in(\latch[378] ),
    .latch_enable_out(\latch[379] ),
    .scan_select_in(\scan[378] ),
    .scan_select_out(\scan[379] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_379 (.clk_in(\clk[379] ),
    .clk_out(\clk[380] ),
    .data_in(\data[379] ),
    .data_out(\data[380] ),
    .latch_enable_in(\latch[379] ),
    .latch_enable_out(\latch[380] ),
    .scan_select_in(\scan[379] ),
    .scan_select_out(\scan[380] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_38 (.clk_in(\clk[38] ),
    .clk_out(\clk[39] ),
    .data_in(\data[38] ),
    .data_out(\data[39] ),
    .latch_enable_in(\latch[38] ),
    .latch_enable_out(\latch[39] ),
    .scan_select_in(\scan[38] ),
    .scan_select_out(\scan[39] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_380 (.clk_in(\clk[380] ),
    .clk_out(\clk[381] ),
    .data_in(\data[380] ),
    .data_out(\data[381] ),
    .latch_enable_in(\latch[380] ),
    .latch_enable_out(\latch[381] ),
    .scan_select_in(\scan[380] ),
    .scan_select_out(\scan[381] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_381 (.clk_in(\clk[381] ),
    .clk_out(\clk[382] ),
    .data_in(\data[381] ),
    .data_out(\data[382] ),
    .latch_enable_in(\latch[381] ),
    .latch_enable_out(\latch[382] ),
    .scan_select_in(\scan[381] ),
    .scan_select_out(\scan[382] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_382 (.clk_in(\clk[382] ),
    .clk_out(\clk[383] ),
    .data_in(\data[382] ),
    .data_out(\data[383] ),
    .latch_enable_in(\latch[382] ),
    .latch_enable_out(\latch[383] ),
    .scan_select_in(\scan[382] ),
    .scan_select_out(\scan[383] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_383 (.clk_in(\clk[383] ),
    .clk_out(\clk[384] ),
    .data_in(\data[383] ),
    .data_out(\data[384] ),
    .latch_enable_in(\latch[383] ),
    .latch_enable_out(\latch[384] ),
    .scan_select_in(\scan[383] ),
    .scan_select_out(\scan[384] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_384 (.clk_in(\clk[384] ),
    .clk_out(\clk[385] ),
    .data_in(\data[384] ),
    .data_out(\data[385] ),
    .latch_enable_in(\latch[384] ),
    .latch_enable_out(\latch[385] ),
    .scan_select_in(\scan[384] ),
    .scan_select_out(\scan[385] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_385 (.clk_in(\clk[385] ),
    .clk_out(\clk[386] ),
    .data_in(\data[385] ),
    .data_out(\data[386] ),
    .latch_enable_in(\latch[385] ),
    .latch_enable_out(\latch[386] ),
    .scan_select_in(\scan[385] ),
    .scan_select_out(\scan[386] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_386 (.clk_in(\clk[386] ),
    .clk_out(\clk[387] ),
    .data_in(\data[386] ),
    .data_out(\data[387] ),
    .latch_enable_in(\latch[386] ),
    .latch_enable_out(\latch[387] ),
    .scan_select_in(\scan[386] ),
    .scan_select_out(\scan[387] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_387 (.clk_in(\clk[387] ),
    .clk_out(\clk[388] ),
    .data_in(\data[387] ),
    .data_out(\data[388] ),
    .latch_enable_in(\latch[387] ),
    .latch_enable_out(\latch[388] ),
    .scan_select_in(\scan[387] ),
    .scan_select_out(\scan[388] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_388 (.clk_in(\clk[388] ),
    .clk_out(\clk[389] ),
    .data_in(\data[388] ),
    .data_out(\data[389] ),
    .latch_enable_in(\latch[388] ),
    .latch_enable_out(\latch[389] ),
    .scan_select_in(\scan[388] ),
    .scan_select_out(\scan[389] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_389 (.clk_in(\clk[389] ),
    .clk_out(\clk[390] ),
    .data_in(\data[389] ),
    .data_out(\data[390] ),
    .latch_enable_in(\latch[389] ),
    .latch_enable_out(\latch[390] ),
    .scan_select_in(\scan[389] ),
    .scan_select_out(\scan[390] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_39 (.clk_in(\clk[39] ),
    .clk_out(\clk[40] ),
    .data_in(\data[39] ),
    .data_out(\data[40] ),
    .latch_enable_in(\latch[39] ),
    .latch_enable_out(\latch[40] ),
    .scan_select_in(\scan[39] ),
    .scan_select_out(\scan[40] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_390 (.clk_in(\clk[390] ),
    .clk_out(\clk[391] ),
    .data_in(\data[390] ),
    .data_out(\data[391] ),
    .latch_enable_in(\latch[390] ),
    .latch_enable_out(\latch[391] ),
    .scan_select_in(\scan[390] ),
    .scan_select_out(\scan[391] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_391 (.clk_in(\clk[391] ),
    .clk_out(\clk[392] ),
    .data_in(\data[391] ),
    .data_out(\data[392] ),
    .latch_enable_in(\latch[391] ),
    .latch_enable_out(\latch[392] ),
    .scan_select_in(\scan[391] ),
    .scan_select_out(\scan[392] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_392 (.clk_in(\clk[392] ),
    .clk_out(\clk[393] ),
    .data_in(\data[392] ),
    .data_out(\data[393] ),
    .latch_enable_in(\latch[392] ),
    .latch_enable_out(\latch[393] ),
    .scan_select_in(\scan[392] ),
    .scan_select_out(\scan[393] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_393 (.clk_in(\clk[393] ),
    .clk_out(\clk[394] ),
    .data_in(\data[393] ),
    .data_out(\data[394] ),
    .latch_enable_in(\latch[393] ),
    .latch_enable_out(\latch[394] ),
    .scan_select_in(\scan[393] ),
    .scan_select_out(\scan[394] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_394 (.clk_in(\clk[394] ),
    .clk_out(\clk[395] ),
    .data_in(\data[394] ),
    .data_out(\data[395] ),
    .latch_enable_in(\latch[394] ),
    .latch_enable_out(\latch[395] ),
    .scan_select_in(\scan[394] ),
    .scan_select_out(\scan[395] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_395 (.clk_in(\clk[395] ),
    .clk_out(\clk[396] ),
    .data_in(\data[395] ),
    .data_out(\data[396] ),
    .latch_enable_in(\latch[395] ),
    .latch_enable_out(\latch[396] ),
    .scan_select_in(\scan[395] ),
    .scan_select_out(\scan[396] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_396 (.clk_in(\clk[396] ),
    .clk_out(\clk[397] ),
    .data_in(\data[396] ),
    .data_out(\data[397] ),
    .latch_enable_in(\latch[396] ),
    .latch_enable_out(\latch[397] ),
    .scan_select_in(\scan[396] ),
    .scan_select_out(\scan[397] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_397 (.clk_in(\clk[397] ),
    .clk_out(\clk[398] ),
    .data_in(\data[397] ),
    .data_out(\data[398] ),
    .latch_enable_in(\latch[397] ),
    .latch_enable_out(\latch[398] ),
    .scan_select_in(\scan[397] ),
    .scan_select_out(\scan[398] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_398 (.clk_in(\clk[398] ),
    .clk_out(\clk[399] ),
    .data_in(\data[398] ),
    .data_out(\data[399] ),
    .latch_enable_in(\latch[398] ),
    .latch_enable_out(\latch[399] ),
    .scan_select_in(\scan[398] ),
    .scan_select_out(\scan[399] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_399 (.clk_in(\clk[399] ),
    .clk_out(\clk[400] ),
    .data_in(\data[399] ),
    .data_out(\data[400] ),
    .latch_enable_in(\latch[399] ),
    .latch_enable_out(\latch[400] ),
    .scan_select_in(\scan[399] ),
    .scan_select_out(\scan[400] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_40 (.clk_in(\clk[40] ),
    .clk_out(\clk[41] ),
    .data_in(\data[40] ),
    .data_out(\data[41] ),
    .latch_enable_in(\latch[40] ),
    .latch_enable_out(\latch[41] ),
    .scan_select_in(\scan[40] ),
    .scan_select_out(\scan[41] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_400 (.clk_in(\clk[400] ),
    .clk_out(\clk[401] ),
    .data_in(\data[400] ),
    .data_out(\data[401] ),
    .latch_enable_in(\latch[400] ),
    .latch_enable_out(\latch[401] ),
    .scan_select_in(\scan[400] ),
    .scan_select_out(\scan[401] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_401 (.clk_in(\clk[401] ),
    .clk_out(\clk[402] ),
    .data_in(\data[401] ),
    .data_out(\data[402] ),
    .latch_enable_in(\latch[401] ),
    .latch_enable_out(\latch[402] ),
    .scan_select_in(\scan[401] ),
    .scan_select_out(\scan[402] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_402 (.clk_in(\clk[402] ),
    .clk_out(\clk[403] ),
    .data_in(\data[402] ),
    .data_out(\data[403] ),
    .latch_enable_in(\latch[402] ),
    .latch_enable_out(\latch[403] ),
    .scan_select_in(\scan[402] ),
    .scan_select_out(\scan[403] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_403 (.clk_in(\clk[403] ),
    .clk_out(\clk[404] ),
    .data_in(\data[403] ),
    .data_out(\data[404] ),
    .latch_enable_in(\latch[403] ),
    .latch_enable_out(\latch[404] ),
    .scan_select_in(\scan[403] ),
    .scan_select_out(\scan[404] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_404 (.clk_in(\clk[404] ),
    .clk_out(\clk[405] ),
    .data_in(\data[404] ),
    .data_out(\data[405] ),
    .latch_enable_in(\latch[404] ),
    .latch_enable_out(\latch[405] ),
    .scan_select_in(\scan[404] ),
    .scan_select_out(\scan[405] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_405 (.clk_in(\clk[405] ),
    .clk_out(\clk[406] ),
    .data_in(\data[405] ),
    .data_out(\data[406] ),
    .latch_enable_in(\latch[405] ),
    .latch_enable_out(\latch[406] ),
    .scan_select_in(\scan[405] ),
    .scan_select_out(\scan[406] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_406 (.clk_in(\clk[406] ),
    .clk_out(\clk[407] ),
    .data_in(\data[406] ),
    .data_out(\data[407] ),
    .latch_enable_in(\latch[406] ),
    .latch_enable_out(\latch[407] ),
    .scan_select_in(\scan[406] ),
    .scan_select_out(\scan[407] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_407 (.clk_in(\clk[407] ),
    .clk_out(\clk[408] ),
    .data_in(\data[407] ),
    .data_out(\data[408] ),
    .latch_enable_in(\latch[407] ),
    .latch_enable_out(\latch[408] ),
    .scan_select_in(\scan[407] ),
    .scan_select_out(\scan[408] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_408 (.clk_in(\clk[408] ),
    .clk_out(\clk[409] ),
    .data_in(\data[408] ),
    .data_out(\data[409] ),
    .latch_enable_in(\latch[408] ),
    .latch_enable_out(\latch[409] ),
    .scan_select_in(\scan[408] ),
    .scan_select_out(\scan[409] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_409 (.clk_in(\clk[409] ),
    .clk_out(\clk[410] ),
    .data_in(\data[409] ),
    .data_out(\data[410] ),
    .latch_enable_in(\latch[409] ),
    .latch_enable_out(\latch[410] ),
    .scan_select_in(\scan[409] ),
    .scan_select_out(\scan[410] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_41 (.clk_in(\clk[41] ),
    .clk_out(\clk[42] ),
    .data_in(\data[41] ),
    .data_out(\data[42] ),
    .latch_enable_in(\latch[41] ),
    .latch_enable_out(\latch[42] ),
    .scan_select_in(\scan[41] ),
    .scan_select_out(\scan[42] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_410 (.clk_in(\clk[410] ),
    .clk_out(\clk[411] ),
    .data_in(\data[410] ),
    .data_out(\data[411] ),
    .latch_enable_in(\latch[410] ),
    .latch_enable_out(\latch[411] ),
    .scan_select_in(\scan[410] ),
    .scan_select_out(\scan[411] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_411 (.clk_in(\clk[411] ),
    .clk_out(\clk[412] ),
    .data_in(\data[411] ),
    .data_out(\data[412] ),
    .latch_enable_in(\latch[411] ),
    .latch_enable_out(\latch[412] ),
    .scan_select_in(\scan[411] ),
    .scan_select_out(\scan[412] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_412 (.clk_in(\clk[412] ),
    .clk_out(\clk[413] ),
    .data_in(\data[412] ),
    .data_out(\data[413] ),
    .latch_enable_in(\latch[412] ),
    .latch_enable_out(\latch[413] ),
    .scan_select_in(\scan[412] ),
    .scan_select_out(\scan[413] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_413 (.clk_in(\clk[413] ),
    .clk_out(\clk[414] ),
    .data_in(\data[413] ),
    .data_out(\data[414] ),
    .latch_enable_in(\latch[413] ),
    .latch_enable_out(\latch[414] ),
    .scan_select_in(\scan[413] ),
    .scan_select_out(\scan[414] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_414 (.clk_in(\clk[414] ),
    .clk_out(\clk[415] ),
    .data_in(\data[414] ),
    .data_out(\data[415] ),
    .latch_enable_in(\latch[414] ),
    .latch_enable_out(\latch[415] ),
    .scan_select_in(\scan[414] ),
    .scan_select_out(\scan[415] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_415 (.clk_in(\clk[415] ),
    .clk_out(\clk[416] ),
    .data_in(\data[415] ),
    .data_out(\data[416] ),
    .latch_enable_in(\latch[415] ),
    .latch_enable_out(\latch[416] ),
    .scan_select_in(\scan[415] ),
    .scan_select_out(\scan[416] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_416 (.clk_in(\clk[416] ),
    .clk_out(\clk[417] ),
    .data_in(\data[416] ),
    .data_out(\data[417] ),
    .latch_enable_in(\latch[416] ),
    .latch_enable_out(\latch[417] ),
    .scan_select_in(\scan[416] ),
    .scan_select_out(\scan[417] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_417 (.clk_in(\clk[417] ),
    .clk_out(\clk[418] ),
    .data_in(\data[417] ),
    .data_out(\data[418] ),
    .latch_enable_in(\latch[417] ),
    .latch_enable_out(\latch[418] ),
    .scan_select_in(\scan[417] ),
    .scan_select_out(\scan[418] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_418 (.clk_in(\clk[418] ),
    .clk_out(\clk[419] ),
    .data_in(\data[418] ),
    .data_out(\data[419] ),
    .latch_enable_in(\latch[418] ),
    .latch_enable_out(\latch[419] ),
    .scan_select_in(\scan[418] ),
    .scan_select_out(\scan[419] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_419 (.clk_in(\clk[419] ),
    .clk_out(\clk[420] ),
    .data_in(\data[419] ),
    .data_out(\data[420] ),
    .latch_enable_in(\latch[419] ),
    .latch_enable_out(\latch[420] ),
    .scan_select_in(\scan[419] ),
    .scan_select_out(\scan[420] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_42 (.clk_in(\clk[42] ),
    .clk_out(\clk[43] ),
    .data_in(\data[42] ),
    .data_out(\data[43] ),
    .latch_enable_in(\latch[42] ),
    .latch_enable_out(\latch[43] ),
    .scan_select_in(\scan[42] ),
    .scan_select_out(\scan[43] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_420 (.clk_in(\clk[420] ),
    .clk_out(\clk[421] ),
    .data_in(\data[420] ),
    .data_out(\data[421] ),
    .latch_enable_in(\latch[420] ),
    .latch_enable_out(\latch[421] ),
    .scan_select_in(\scan[420] ),
    .scan_select_out(\scan[421] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_421 (.clk_in(\clk[421] ),
    .clk_out(\clk[422] ),
    .data_in(\data[421] ),
    .data_out(\data[422] ),
    .latch_enable_in(\latch[421] ),
    .latch_enable_out(\latch[422] ),
    .scan_select_in(\scan[421] ),
    .scan_select_out(\scan[422] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_422 (.clk_in(\clk[422] ),
    .clk_out(\clk[423] ),
    .data_in(\data[422] ),
    .data_out(\data[423] ),
    .latch_enable_in(\latch[422] ),
    .latch_enable_out(\latch[423] ),
    .scan_select_in(\scan[422] ),
    .scan_select_out(\scan[423] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_423 (.clk_in(\clk[423] ),
    .clk_out(\clk[424] ),
    .data_in(\data[423] ),
    .data_out(\data[424] ),
    .latch_enable_in(\latch[423] ),
    .latch_enable_out(\latch[424] ),
    .scan_select_in(\scan[423] ),
    .scan_select_out(\scan[424] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_424 (.clk_in(\clk[424] ),
    .clk_out(\clk[425] ),
    .data_in(\data[424] ),
    .data_out(\data[425] ),
    .latch_enable_in(\latch[424] ),
    .latch_enable_out(\latch[425] ),
    .scan_select_in(\scan[424] ),
    .scan_select_out(\scan[425] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_425 (.clk_in(\clk[425] ),
    .clk_out(\clk[426] ),
    .data_in(\data[425] ),
    .data_out(\data[426] ),
    .latch_enable_in(\latch[425] ),
    .latch_enable_out(\latch[426] ),
    .scan_select_in(\scan[425] ),
    .scan_select_out(\scan[426] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_426 (.clk_in(\clk[426] ),
    .clk_out(\clk[427] ),
    .data_in(\data[426] ),
    .data_out(\data[427] ),
    .latch_enable_in(\latch[426] ),
    .latch_enable_out(\latch[427] ),
    .scan_select_in(\scan[426] ),
    .scan_select_out(\scan[427] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_427 (.clk_in(\clk[427] ),
    .clk_out(\clk[428] ),
    .data_in(\data[427] ),
    .data_out(\data[428] ),
    .latch_enable_in(\latch[427] ),
    .latch_enable_out(\latch[428] ),
    .scan_select_in(\scan[427] ),
    .scan_select_out(\scan[428] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_428 (.clk_in(\clk[428] ),
    .clk_out(\clk[429] ),
    .data_in(\data[428] ),
    .data_out(\data[429] ),
    .latch_enable_in(\latch[428] ),
    .latch_enable_out(\latch[429] ),
    .scan_select_in(\scan[428] ),
    .scan_select_out(\scan[429] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_429 (.clk_in(\clk[429] ),
    .clk_out(\clk[430] ),
    .data_in(\data[429] ),
    .data_out(\data[430] ),
    .latch_enable_in(\latch[429] ),
    .latch_enable_out(\latch[430] ),
    .scan_select_in(\scan[429] ),
    .scan_select_out(\scan[430] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_43 (.clk_in(\clk[43] ),
    .clk_out(\clk[44] ),
    .data_in(\data[43] ),
    .data_out(\data[44] ),
    .latch_enable_in(\latch[43] ),
    .latch_enable_out(\latch[44] ),
    .scan_select_in(\scan[43] ),
    .scan_select_out(\scan[44] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_430 (.clk_in(\clk[430] ),
    .clk_out(\clk[431] ),
    .data_in(\data[430] ),
    .data_out(\data[431] ),
    .latch_enable_in(\latch[430] ),
    .latch_enable_out(\latch[431] ),
    .scan_select_in(\scan[430] ),
    .scan_select_out(\scan[431] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_431 (.clk_in(\clk[431] ),
    .clk_out(\clk[432] ),
    .data_in(\data[431] ),
    .data_out(\data[432] ),
    .latch_enable_in(\latch[431] ),
    .latch_enable_out(\latch[432] ),
    .scan_select_in(\scan[431] ),
    .scan_select_out(\scan[432] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_432 (.clk_in(\clk[432] ),
    .clk_out(\clk[433] ),
    .data_in(\data[432] ),
    .data_out(\data[433] ),
    .latch_enable_in(\latch[432] ),
    .latch_enable_out(\latch[433] ),
    .scan_select_in(\scan[432] ),
    .scan_select_out(\scan[433] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_433 (.clk_in(\clk[433] ),
    .clk_out(\clk[434] ),
    .data_in(\data[433] ),
    .data_out(\data[434] ),
    .latch_enable_in(\latch[433] ),
    .latch_enable_out(\latch[434] ),
    .scan_select_in(\scan[433] ),
    .scan_select_out(\scan[434] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_434 (.clk_in(\clk[434] ),
    .clk_out(\clk[435] ),
    .data_in(\data[434] ),
    .data_out(\data[435] ),
    .latch_enable_in(\latch[434] ),
    .latch_enable_out(\latch[435] ),
    .scan_select_in(\scan[434] ),
    .scan_select_out(\scan[435] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_435 (.clk_in(\clk[435] ),
    .clk_out(\clk[436] ),
    .data_in(\data[435] ),
    .data_out(\data[436] ),
    .latch_enable_in(\latch[435] ),
    .latch_enable_out(\latch[436] ),
    .scan_select_in(\scan[435] ),
    .scan_select_out(\scan[436] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_436 (.clk_in(\clk[436] ),
    .clk_out(\clk[437] ),
    .data_in(\data[436] ),
    .data_out(\data[437] ),
    .latch_enable_in(\latch[436] ),
    .latch_enable_out(\latch[437] ),
    .scan_select_in(\scan[436] ),
    .scan_select_out(\scan[437] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_437 (.clk_in(\clk[437] ),
    .clk_out(\clk[438] ),
    .data_in(\data[437] ),
    .data_out(\data[438] ),
    .latch_enable_in(\latch[437] ),
    .latch_enable_out(\latch[438] ),
    .scan_select_in(\scan[437] ),
    .scan_select_out(\scan[438] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_438 (.clk_in(\clk[438] ),
    .clk_out(\clk[439] ),
    .data_in(\data[438] ),
    .data_out(\data[439] ),
    .latch_enable_in(\latch[438] ),
    .latch_enable_out(\latch[439] ),
    .scan_select_in(\scan[438] ),
    .scan_select_out(\scan[439] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_439 (.clk_in(\clk[439] ),
    .clk_out(\clk[440] ),
    .data_in(\data[439] ),
    .data_out(\data[440] ),
    .latch_enable_in(\latch[439] ),
    .latch_enable_out(\latch[440] ),
    .scan_select_in(\scan[439] ),
    .scan_select_out(\scan[440] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_44 (.clk_in(\clk[44] ),
    .clk_out(\clk[45] ),
    .data_in(\data[44] ),
    .data_out(\data[45] ),
    .latch_enable_in(\latch[44] ),
    .latch_enable_out(\latch[45] ),
    .scan_select_in(\scan[44] ),
    .scan_select_out(\scan[45] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_440 (.clk_in(\clk[440] ),
    .clk_out(\clk[441] ),
    .data_in(\data[440] ),
    .data_out(\data[441] ),
    .latch_enable_in(\latch[440] ),
    .latch_enable_out(\latch[441] ),
    .scan_select_in(\scan[440] ),
    .scan_select_out(\scan[441] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_441 (.clk_in(\clk[441] ),
    .clk_out(\clk[442] ),
    .data_in(\data[441] ),
    .data_out(\data[442] ),
    .latch_enable_in(\latch[441] ),
    .latch_enable_out(\latch[442] ),
    .scan_select_in(\scan[441] ),
    .scan_select_out(\scan[442] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_442 (.clk_in(\clk[442] ),
    .clk_out(\clk[443] ),
    .data_in(\data[442] ),
    .data_out(\data[443] ),
    .latch_enable_in(\latch[442] ),
    .latch_enable_out(\latch[443] ),
    .scan_select_in(\scan[442] ),
    .scan_select_out(\scan[443] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_443 (.clk_in(\clk[443] ),
    .clk_out(\clk[444] ),
    .data_in(\data[443] ),
    .data_out(\data[444] ),
    .latch_enable_in(\latch[443] ),
    .latch_enable_out(\latch[444] ),
    .scan_select_in(\scan[443] ),
    .scan_select_out(\scan[444] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_444 (.clk_in(\clk[444] ),
    .clk_out(\clk[445] ),
    .data_in(\data[444] ),
    .data_out(\data[445] ),
    .latch_enable_in(\latch[444] ),
    .latch_enable_out(\latch[445] ),
    .scan_select_in(\scan[444] ),
    .scan_select_out(\scan[445] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_445 (.clk_in(\clk[445] ),
    .clk_out(\clk[446] ),
    .data_in(\data[445] ),
    .data_out(\data[446] ),
    .latch_enable_in(\latch[445] ),
    .latch_enable_out(\latch[446] ),
    .scan_select_in(\scan[445] ),
    .scan_select_out(\scan[446] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_446 (.clk_in(\clk[446] ),
    .clk_out(\clk[447] ),
    .data_in(\data[446] ),
    .data_out(\data[447] ),
    .latch_enable_in(\latch[446] ),
    .latch_enable_out(\latch[447] ),
    .scan_select_in(\scan[446] ),
    .scan_select_out(\scan[447] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_447 (.clk_in(\clk[447] ),
    .clk_out(\clk[448] ),
    .data_in(\data[447] ),
    .data_out(\data[448] ),
    .latch_enable_in(\latch[447] ),
    .latch_enable_out(\latch[448] ),
    .scan_select_in(\scan[447] ),
    .scan_select_out(\scan[448] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_448 (.clk_in(\clk[448] ),
    .clk_out(\clk[449] ),
    .data_in(\data[448] ),
    .data_out(\data[449] ),
    .latch_enable_in(\latch[448] ),
    .latch_enable_out(\latch[449] ),
    .scan_select_in(\scan[448] ),
    .scan_select_out(\scan[449] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_449 (.clk_in(\clk[449] ),
    .clk_out(\clk[450] ),
    .data_in(\data[449] ),
    .data_out(\data[450] ),
    .latch_enable_in(\latch[449] ),
    .latch_enable_out(\latch[450] ),
    .scan_select_in(\scan[449] ),
    .scan_select_out(\scan[450] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_45 (.clk_in(\clk[45] ),
    .clk_out(\clk[46] ),
    .data_in(\data[45] ),
    .data_out(\data[46] ),
    .latch_enable_in(\latch[45] ),
    .latch_enable_out(\latch[46] ),
    .scan_select_in(\scan[45] ),
    .scan_select_out(\scan[46] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_450 (.clk_in(\clk[450] ),
    .clk_out(\clk[451] ),
    .data_in(\data[450] ),
    .data_out(\data[451] ),
    .latch_enable_in(\latch[450] ),
    .latch_enable_out(\latch[451] ),
    .scan_select_in(\scan[450] ),
    .scan_select_out(\scan[451] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_451 (.clk_in(\clk[451] ),
    .clk_out(\clk[452] ),
    .data_in(\data[451] ),
    .data_out(\data[452] ),
    .latch_enable_in(\latch[451] ),
    .latch_enable_out(\latch[452] ),
    .scan_select_in(\scan[451] ),
    .scan_select_out(\scan[452] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_452 (.clk_in(\clk[452] ),
    .clk_out(\clk[453] ),
    .data_in(\data[452] ),
    .data_out(\data[453] ),
    .latch_enable_in(\latch[452] ),
    .latch_enable_out(\latch[453] ),
    .scan_select_in(\scan[452] ),
    .scan_select_out(\scan[453] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_453 (.clk_in(\clk[453] ),
    .clk_out(\clk[454] ),
    .data_in(\data[453] ),
    .data_out(\data[454] ),
    .latch_enable_in(\latch[453] ),
    .latch_enable_out(\latch[454] ),
    .scan_select_in(\scan[453] ),
    .scan_select_out(\scan[454] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_454 (.clk_in(\clk[454] ),
    .clk_out(\clk[455] ),
    .data_in(\data[454] ),
    .data_out(\data[455] ),
    .latch_enable_in(\latch[454] ),
    .latch_enable_out(\latch[455] ),
    .scan_select_in(\scan[454] ),
    .scan_select_out(\scan[455] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_455 (.clk_in(\clk[455] ),
    .clk_out(\clk[456] ),
    .data_in(\data[455] ),
    .data_out(\data[456] ),
    .latch_enable_in(\latch[455] ),
    .latch_enable_out(\latch[456] ),
    .scan_select_in(\scan[455] ),
    .scan_select_out(\scan[456] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_456 (.clk_in(\clk[456] ),
    .clk_out(\clk[457] ),
    .data_in(\data[456] ),
    .data_out(\data[457] ),
    .latch_enable_in(\latch[456] ),
    .latch_enable_out(\latch[457] ),
    .scan_select_in(\scan[456] ),
    .scan_select_out(\scan[457] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_457 (.clk_in(\clk[457] ),
    .clk_out(\clk[458] ),
    .data_in(\data[457] ),
    .data_out(\data[458] ),
    .latch_enable_in(\latch[457] ),
    .latch_enable_out(\latch[458] ),
    .scan_select_in(\scan[457] ),
    .scan_select_out(\scan[458] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_458 (.clk_in(\clk[458] ),
    .clk_out(\clk[459] ),
    .data_in(\data[458] ),
    .data_out(\data[459] ),
    .latch_enable_in(\latch[458] ),
    .latch_enable_out(\latch[459] ),
    .scan_select_in(\scan[458] ),
    .scan_select_out(\scan[459] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_459 (.clk_in(\clk[459] ),
    .clk_out(\clk[460] ),
    .data_in(\data[459] ),
    .data_out(\data[460] ),
    .latch_enable_in(\latch[459] ),
    .latch_enable_out(\latch[460] ),
    .scan_select_in(\scan[459] ),
    .scan_select_out(\scan[460] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_46 (.clk_in(\clk[46] ),
    .clk_out(\clk[47] ),
    .data_in(\data[46] ),
    .data_out(\data[47] ),
    .latch_enable_in(\latch[46] ),
    .latch_enable_out(\latch[47] ),
    .scan_select_in(\scan[46] ),
    .scan_select_out(\scan[47] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_460 (.clk_in(\clk[460] ),
    .clk_out(\clk[461] ),
    .data_in(\data[460] ),
    .data_out(\data[461] ),
    .latch_enable_in(\latch[460] ),
    .latch_enable_out(\latch[461] ),
    .scan_select_in(\scan[460] ),
    .scan_select_out(\scan[461] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_461 (.clk_in(\clk[461] ),
    .clk_out(\clk[462] ),
    .data_in(\data[461] ),
    .data_out(\data[462] ),
    .latch_enable_in(\latch[461] ),
    .latch_enable_out(\latch[462] ),
    .scan_select_in(\scan[461] ),
    .scan_select_out(\scan[462] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_462 (.clk_in(\clk[462] ),
    .clk_out(\clk[463] ),
    .data_in(\data[462] ),
    .data_out(\data[463] ),
    .latch_enable_in(\latch[462] ),
    .latch_enable_out(\latch[463] ),
    .scan_select_in(\scan[462] ),
    .scan_select_out(\scan[463] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_463 (.clk_in(\clk[463] ),
    .clk_out(\clk[464] ),
    .data_in(\data[463] ),
    .data_out(\data[464] ),
    .latch_enable_in(\latch[463] ),
    .latch_enable_out(\latch[464] ),
    .scan_select_in(\scan[463] ),
    .scan_select_out(\scan[464] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_464 (.clk_in(\clk[464] ),
    .clk_out(\clk[465] ),
    .data_in(\data[464] ),
    .data_out(\data[465] ),
    .latch_enable_in(\latch[464] ),
    .latch_enable_out(\latch[465] ),
    .scan_select_in(\scan[464] ),
    .scan_select_out(\scan[465] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_465 (.clk_in(\clk[465] ),
    .clk_out(\clk[466] ),
    .data_in(\data[465] ),
    .data_out(\data[466] ),
    .latch_enable_in(\latch[465] ),
    .latch_enable_out(\latch[466] ),
    .scan_select_in(\scan[465] ),
    .scan_select_out(\scan[466] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_466 (.clk_in(\clk[466] ),
    .clk_out(\clk[467] ),
    .data_in(\data[466] ),
    .data_out(\data[467] ),
    .latch_enable_in(\latch[466] ),
    .latch_enable_out(\latch[467] ),
    .scan_select_in(\scan[466] ),
    .scan_select_out(\scan[467] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_467 (.clk_in(\clk[467] ),
    .clk_out(\clk[468] ),
    .data_in(\data[467] ),
    .data_out(\data[468] ),
    .latch_enable_in(\latch[467] ),
    .latch_enable_out(\latch[468] ),
    .scan_select_in(\scan[467] ),
    .scan_select_out(\scan[468] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_468 (.clk_in(\clk[468] ),
    .clk_out(\clk[469] ),
    .data_in(\data[468] ),
    .data_out(\data[469] ),
    .latch_enable_in(\latch[468] ),
    .latch_enable_out(\latch[469] ),
    .scan_select_in(\scan[468] ),
    .scan_select_out(\scan[469] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_469 (.clk_in(\clk[469] ),
    .clk_out(\clk[470] ),
    .data_in(\data[469] ),
    .data_out(\data[470] ),
    .latch_enable_in(\latch[469] ),
    .latch_enable_out(\latch[470] ),
    .scan_select_in(\scan[469] ),
    .scan_select_out(\scan[470] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_47 (.clk_in(\clk[47] ),
    .clk_out(\clk[48] ),
    .data_in(\data[47] ),
    .data_out(\data[48] ),
    .latch_enable_in(\latch[47] ),
    .latch_enable_out(\latch[48] ),
    .scan_select_in(\scan[47] ),
    .scan_select_out(\scan[48] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_470 (.clk_in(\clk[470] ),
    .clk_out(\clk[471] ),
    .data_in(\data[470] ),
    .data_out(\data[471] ),
    .latch_enable_in(\latch[470] ),
    .latch_enable_out(\latch[471] ),
    .scan_select_in(\scan[470] ),
    .scan_select_out(\scan[471] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_471 (.clk_in(\clk[471] ),
    .clk_out(\clk[472] ),
    .data_in(\data[471] ),
    .data_out(\data[472] ),
    .latch_enable_in(\latch[471] ),
    .latch_enable_out(\latch[472] ),
    .scan_select_in(\scan[471] ),
    .scan_select_out(\scan[472] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_472 (.clk_in(\clk[472] ),
    .clk_out(\clk[473] ),
    .data_in(\data[472] ),
    .data_out(\data[473] ),
    .latch_enable_in(\latch[472] ),
    .latch_enable_out(\latch[473] ),
    .scan_select_in(\scan[472] ),
    .scan_select_out(\scan[473] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_473 (.clk_in(\clk[473] ),
    .clk_out(\clk[474] ),
    .data_in(\data[473] ),
    .data_out(\data[474] ),
    .latch_enable_in(\latch[473] ),
    .latch_enable_out(\latch[474] ),
    .scan_select_in(\scan[473] ),
    .scan_select_out(\scan[474] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_474 (.clk_in(\clk[474] ),
    .clk_out(\clk[475] ),
    .data_in(\data[474] ),
    .data_out(\data[475] ),
    .latch_enable_in(\latch[474] ),
    .latch_enable_out(\latch[475] ),
    .scan_select_in(\scan[474] ),
    .scan_select_out(\scan[475] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_475 (.clk_in(\clk[475] ),
    .clk_out(\clk[476] ),
    .data_in(\data[475] ),
    .data_out(\data[476] ),
    .latch_enable_in(\latch[475] ),
    .latch_enable_out(\latch[476] ),
    .scan_select_in(\scan[475] ),
    .scan_select_out(\scan[476] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_476 (.clk_in(\clk[476] ),
    .clk_out(\clk[477] ),
    .data_in(\data[476] ),
    .data_out(\data[477] ),
    .latch_enable_in(\latch[476] ),
    .latch_enable_out(\latch[477] ),
    .scan_select_in(\scan[476] ),
    .scan_select_out(\scan[477] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_477 (.clk_in(\clk[477] ),
    .clk_out(\clk[478] ),
    .data_in(\data[477] ),
    .data_out(\data[478] ),
    .latch_enable_in(\latch[477] ),
    .latch_enable_out(\latch[478] ),
    .scan_select_in(\scan[477] ),
    .scan_select_out(\scan[478] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_478 (.clk_in(\clk[478] ),
    .clk_out(\clk[479] ),
    .data_in(\data[478] ),
    .data_out(\data[479] ),
    .latch_enable_in(\latch[478] ),
    .latch_enable_out(\latch[479] ),
    .scan_select_in(\scan[478] ),
    .scan_select_out(\scan[479] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_479 (.clk_in(\clk[479] ),
    .clk_out(\clk[480] ),
    .data_in(\data[479] ),
    .data_out(\data[480] ),
    .latch_enable_in(\latch[479] ),
    .latch_enable_out(\latch[480] ),
    .scan_select_in(\scan[479] ),
    .scan_select_out(\scan[480] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_48 (.clk_in(\clk[48] ),
    .clk_out(\clk[49] ),
    .data_in(\data[48] ),
    .data_out(\data[49] ),
    .latch_enable_in(\latch[48] ),
    .latch_enable_out(\latch[49] ),
    .scan_select_in(\scan[48] ),
    .scan_select_out(\scan[49] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_480 (.clk_in(\clk[480] ),
    .clk_out(\clk[481] ),
    .data_in(\data[480] ),
    .data_out(\data[481] ),
    .latch_enable_in(\latch[480] ),
    .latch_enable_out(\latch[481] ),
    .scan_select_in(\scan[480] ),
    .scan_select_out(\scan[481] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_481 (.clk_in(\clk[481] ),
    .clk_out(\clk[482] ),
    .data_in(\data[481] ),
    .data_out(\data[482] ),
    .latch_enable_in(\latch[481] ),
    .latch_enable_out(\latch[482] ),
    .scan_select_in(\scan[481] ),
    .scan_select_out(\scan[482] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_482 (.clk_in(\clk[482] ),
    .clk_out(\clk[483] ),
    .data_in(\data[482] ),
    .data_out(\data[483] ),
    .latch_enable_in(\latch[482] ),
    .latch_enable_out(\latch[483] ),
    .scan_select_in(\scan[482] ),
    .scan_select_out(\scan[483] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_483 (.clk_in(\clk[483] ),
    .clk_out(\clk[484] ),
    .data_in(\data[483] ),
    .data_out(\data[484] ),
    .latch_enable_in(\latch[483] ),
    .latch_enable_out(\latch[484] ),
    .scan_select_in(\scan[483] ),
    .scan_select_out(\scan[484] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_484 (.clk_in(\clk[484] ),
    .clk_out(\clk[485] ),
    .data_in(\data[484] ),
    .data_out(\data[485] ),
    .latch_enable_in(\latch[484] ),
    .latch_enable_out(\latch[485] ),
    .scan_select_in(\scan[484] ),
    .scan_select_out(\scan[485] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_485 (.clk_in(\clk[485] ),
    .clk_out(\clk[486] ),
    .data_in(\data[485] ),
    .data_out(\data[486] ),
    .latch_enable_in(\latch[485] ),
    .latch_enable_out(\latch[486] ),
    .scan_select_in(\scan[485] ),
    .scan_select_out(\scan[486] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_486 (.clk_in(\clk[486] ),
    .clk_out(\clk[487] ),
    .data_in(\data[486] ),
    .data_out(\data[487] ),
    .latch_enable_in(\latch[486] ),
    .latch_enable_out(\latch[487] ),
    .scan_select_in(\scan[486] ),
    .scan_select_out(\scan[487] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_487 (.clk_in(\clk[487] ),
    .clk_out(\clk[488] ),
    .data_in(\data[487] ),
    .data_out(\data[488] ),
    .latch_enable_in(\latch[487] ),
    .latch_enable_out(\latch[488] ),
    .scan_select_in(\scan[487] ),
    .scan_select_out(\scan[488] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_488 (.clk_in(\clk[488] ),
    .clk_out(\clk[489] ),
    .data_in(\data[488] ),
    .data_out(\data[489] ),
    .latch_enable_in(\latch[488] ),
    .latch_enable_out(\latch[489] ),
    .scan_select_in(\scan[488] ),
    .scan_select_out(\scan[489] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_489 (.clk_in(\clk[489] ),
    .clk_out(\clk[490] ),
    .data_in(\data[489] ),
    .data_out(\data[490] ),
    .latch_enable_in(\latch[489] ),
    .latch_enable_out(\latch[490] ),
    .scan_select_in(\scan[489] ),
    .scan_select_out(\scan[490] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_49 (.clk_in(\clk[49] ),
    .clk_out(\clk[50] ),
    .data_in(\data[49] ),
    .data_out(\data[50] ),
    .latch_enable_in(\latch[49] ),
    .latch_enable_out(\latch[50] ),
    .scan_select_in(\scan[49] ),
    .scan_select_out(\scan[50] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_490 (.clk_in(\clk[490] ),
    .clk_out(\clk[491] ),
    .data_in(\data[490] ),
    .data_out(\data[491] ),
    .latch_enable_in(\latch[490] ),
    .latch_enable_out(\latch[491] ),
    .scan_select_in(\scan[490] ),
    .scan_select_out(\scan[491] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_491 (.clk_in(\clk[491] ),
    .clk_out(\clk[492] ),
    .data_in(\data[491] ),
    .data_out(\data[492] ),
    .latch_enable_in(\latch[491] ),
    .latch_enable_out(\latch[492] ),
    .scan_select_in(\scan[491] ),
    .scan_select_out(\scan[492] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_492 (.clk_in(\clk[492] ),
    .clk_out(\clk[493] ),
    .data_in(\data[492] ),
    .data_out(\data[493] ),
    .latch_enable_in(\latch[492] ),
    .latch_enable_out(\latch[493] ),
    .scan_select_in(\scan[492] ),
    .scan_select_out(\scan[493] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_493 (.clk_in(\clk[493] ),
    .clk_out(\clk[494] ),
    .data_in(\data[493] ),
    .data_out(\data[494] ),
    .latch_enable_in(\latch[493] ),
    .latch_enable_out(\latch[494] ),
    .scan_select_in(\scan[493] ),
    .scan_select_out(\scan[494] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_494 (.clk_in(\clk[494] ),
    .clk_out(\clk[495] ),
    .data_in(\data[494] ),
    .data_out(\data[495] ),
    .latch_enable_in(\latch[494] ),
    .latch_enable_out(\latch[495] ),
    .scan_select_in(\scan[494] ),
    .scan_select_out(\scan[495] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_495 (.clk_in(\clk[495] ),
    .clk_out(\clk[496] ),
    .data_in(\data[495] ),
    .data_out(\data[496] ),
    .latch_enable_in(\latch[495] ),
    .latch_enable_out(\latch[496] ),
    .scan_select_in(\scan[495] ),
    .scan_select_out(\scan[496] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_496 (.clk_in(\clk[496] ),
    .clk_out(\clk[497] ),
    .data_in(\data[496] ),
    .data_out(\data[497] ),
    .latch_enable_in(\latch[496] ),
    .latch_enable_out(\latch[497] ),
    .scan_select_in(\scan[496] ),
    .scan_select_out(\scan[497] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_497 (.clk_in(\clk[497] ),
    .clk_out(\clk[498] ),
    .data_in(\data[497] ),
    .data_out(\data[498] ),
    .latch_enable_in(\latch[497] ),
    .latch_enable_out(\latch[498] ),
    .scan_select_in(\scan[497] ),
    .scan_select_out(\scan[498] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_50 (.clk_in(\clk[50] ),
    .clk_out(\clk[51] ),
    .data_in(\data[50] ),
    .data_out(\data[51] ),
    .latch_enable_in(\latch[50] ),
    .latch_enable_out(\latch[51] ),
    .scan_select_in(\scan[50] ),
    .scan_select_out(\scan[51] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_51 (.clk_in(\clk[51] ),
    .clk_out(\clk[52] ),
    .data_in(\data[51] ),
    .data_out(\data[52] ),
    .latch_enable_in(\latch[51] ),
    .latch_enable_out(\latch[52] ),
    .scan_select_in(\scan[51] ),
    .scan_select_out(\scan[52] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_52 (.clk_in(\clk[52] ),
    .clk_out(\clk[53] ),
    .data_in(\data[52] ),
    .data_out(\data[53] ),
    .latch_enable_in(\latch[52] ),
    .latch_enable_out(\latch[53] ),
    .scan_select_in(\scan[52] ),
    .scan_select_out(\scan[53] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_53 (.clk_in(\clk[53] ),
    .clk_out(\clk[54] ),
    .data_in(\data[53] ),
    .data_out(\data[54] ),
    .latch_enable_in(\latch[53] ),
    .latch_enable_out(\latch[54] ),
    .scan_select_in(\scan[53] ),
    .scan_select_out(\scan[54] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_54 (.clk_in(\clk[54] ),
    .clk_out(\clk[55] ),
    .data_in(\data[54] ),
    .data_out(\data[55] ),
    .latch_enable_in(\latch[54] ),
    .latch_enable_out(\latch[55] ),
    .scan_select_in(\scan[54] ),
    .scan_select_out(\scan[55] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_55 (.clk_in(\clk[55] ),
    .clk_out(\clk[56] ),
    .data_in(\data[55] ),
    .data_out(\data[56] ),
    .latch_enable_in(\latch[55] ),
    .latch_enable_out(\latch[56] ),
    .scan_select_in(\scan[55] ),
    .scan_select_out(\scan[56] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_56 (.clk_in(\clk[56] ),
    .clk_out(\clk[57] ),
    .data_in(\data[56] ),
    .data_out(\data[57] ),
    .latch_enable_in(\latch[56] ),
    .latch_enable_out(\latch[57] ),
    .scan_select_in(\scan[56] ),
    .scan_select_out(\scan[57] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_57 (.clk_in(\clk[57] ),
    .clk_out(\clk[58] ),
    .data_in(\data[57] ),
    .data_out(\data[58] ),
    .latch_enable_in(\latch[57] ),
    .latch_enable_out(\latch[58] ),
    .scan_select_in(\scan[57] ),
    .scan_select_out(\scan[58] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_58 (.clk_in(\clk[58] ),
    .clk_out(\clk[59] ),
    .data_in(\data[58] ),
    .data_out(\data[59] ),
    .latch_enable_in(\latch[58] ),
    .latch_enable_out(\latch[59] ),
    .scan_select_in(\scan[58] ),
    .scan_select_out(\scan[59] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_59 (.clk_in(\clk[59] ),
    .clk_out(\clk[60] ),
    .data_in(\data[59] ),
    .data_out(\data[60] ),
    .latch_enable_in(\latch[59] ),
    .latch_enable_out(\latch[60] ),
    .scan_select_in(\scan[59] ),
    .scan_select_out(\scan[60] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_60 (.clk_in(\clk[60] ),
    .clk_out(\clk[61] ),
    .data_in(\data[60] ),
    .data_out(\data[61] ),
    .latch_enable_in(\latch[60] ),
    .latch_enable_out(\latch[61] ),
    .scan_select_in(\scan[60] ),
    .scan_select_out(\scan[61] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_61 (.clk_in(\clk[61] ),
    .clk_out(\clk[62] ),
    .data_in(\data[61] ),
    .data_out(\data[62] ),
    .latch_enable_in(\latch[61] ),
    .latch_enable_out(\latch[62] ),
    .scan_select_in(\scan[61] ),
    .scan_select_out(\scan[62] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_62 (.clk_in(\clk[62] ),
    .clk_out(\clk[63] ),
    .data_in(\data[62] ),
    .data_out(\data[63] ),
    .latch_enable_in(\latch[62] ),
    .latch_enable_out(\latch[63] ),
    .scan_select_in(\scan[62] ),
    .scan_select_out(\scan[63] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_63 (.clk_in(\clk[63] ),
    .clk_out(\clk[64] ),
    .data_in(\data[63] ),
    .data_out(\data[64] ),
    .latch_enable_in(\latch[63] ),
    .latch_enable_out(\latch[64] ),
    .scan_select_in(\scan[63] ),
    .scan_select_out(\scan[64] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_64 (.clk_in(\clk[64] ),
    .clk_out(\clk[65] ),
    .data_in(\data[64] ),
    .data_out(\data[65] ),
    .latch_enable_in(\latch[64] ),
    .latch_enable_out(\latch[65] ),
    .scan_select_in(\scan[64] ),
    .scan_select_out(\scan[65] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_65 (.clk_in(\clk[65] ),
    .clk_out(\clk[66] ),
    .data_in(\data[65] ),
    .data_out(\data[66] ),
    .latch_enable_in(\latch[65] ),
    .latch_enable_out(\latch[66] ),
    .scan_select_in(\scan[65] ),
    .scan_select_out(\scan[66] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_66 (.clk_in(\clk[66] ),
    .clk_out(\clk[67] ),
    .data_in(\data[66] ),
    .data_out(\data[67] ),
    .latch_enable_in(\latch[66] ),
    .latch_enable_out(\latch[67] ),
    .scan_select_in(\scan[66] ),
    .scan_select_out(\scan[67] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_67 (.clk_in(\clk[67] ),
    .clk_out(\clk[68] ),
    .data_in(\data[67] ),
    .data_out(\data[68] ),
    .latch_enable_in(\latch[67] ),
    .latch_enable_out(\latch[68] ),
    .scan_select_in(\scan[67] ),
    .scan_select_out(\scan[68] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_68 (.clk_in(\clk[68] ),
    .clk_out(\clk[69] ),
    .data_in(\data[68] ),
    .data_out(\data[69] ),
    .latch_enable_in(\latch[68] ),
    .latch_enable_out(\latch[69] ),
    .scan_select_in(\scan[68] ),
    .scan_select_out(\scan[69] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_69 (.clk_in(\clk[69] ),
    .clk_out(\clk[70] ),
    .data_in(\data[69] ),
    .data_out(\data[70] ),
    .latch_enable_in(\latch[69] ),
    .latch_enable_out(\latch[70] ),
    .scan_select_in(\scan[69] ),
    .scan_select_out(\scan[70] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_70 (.clk_in(\clk[70] ),
    .clk_out(\clk[71] ),
    .data_in(\data[70] ),
    .data_out(\data[71] ),
    .latch_enable_in(\latch[70] ),
    .latch_enable_out(\latch[71] ),
    .scan_select_in(\scan[70] ),
    .scan_select_out(\scan[71] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_71 (.clk_in(\clk[71] ),
    .clk_out(\clk[72] ),
    .data_in(\data[71] ),
    .data_out(\data[72] ),
    .latch_enable_in(\latch[71] ),
    .latch_enable_out(\latch[72] ),
    .scan_select_in(\scan[71] ),
    .scan_select_out(\scan[72] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_72 (.clk_in(\clk[72] ),
    .clk_out(\clk[73] ),
    .data_in(\data[72] ),
    .data_out(\data[73] ),
    .latch_enable_in(\latch[72] ),
    .latch_enable_out(\latch[73] ),
    .scan_select_in(\scan[72] ),
    .scan_select_out(\scan[73] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_73 (.clk_in(\clk[73] ),
    .clk_out(\clk[74] ),
    .data_in(\data[73] ),
    .data_out(\data[74] ),
    .latch_enable_in(\latch[73] ),
    .latch_enable_out(\latch[74] ),
    .scan_select_in(\scan[73] ),
    .scan_select_out(\scan[74] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_74 (.clk_in(\clk[74] ),
    .clk_out(\clk[75] ),
    .data_in(\data[74] ),
    .data_out(\data[75] ),
    .latch_enable_in(\latch[74] ),
    .latch_enable_out(\latch[75] ),
    .scan_select_in(\scan[74] ),
    .scan_select_out(\scan[75] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_75 (.clk_in(\clk[75] ),
    .clk_out(\clk[76] ),
    .data_in(\data[75] ),
    .data_out(\data[76] ),
    .latch_enable_in(\latch[75] ),
    .latch_enable_out(\latch[76] ),
    .scan_select_in(\scan[75] ),
    .scan_select_out(\scan[76] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_76 (.clk_in(\clk[76] ),
    .clk_out(\clk[77] ),
    .data_in(\data[76] ),
    .data_out(\data[77] ),
    .latch_enable_in(\latch[76] ),
    .latch_enable_out(\latch[77] ),
    .scan_select_in(\scan[76] ),
    .scan_select_out(\scan[77] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_77 (.clk_in(\clk[77] ),
    .clk_out(\clk[78] ),
    .data_in(\data[77] ),
    .data_out(\data[78] ),
    .latch_enable_in(\latch[77] ),
    .latch_enable_out(\latch[78] ),
    .scan_select_in(\scan[77] ),
    .scan_select_out(\scan[78] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_78 (.clk_in(\clk[78] ),
    .clk_out(\clk[79] ),
    .data_in(\data[78] ),
    .data_out(\data[79] ),
    .latch_enable_in(\latch[78] ),
    .latch_enable_out(\latch[79] ),
    .scan_select_in(\scan[78] ),
    .scan_select_out(\scan[79] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_79 (.clk_in(\clk[79] ),
    .clk_out(\clk[80] ),
    .data_in(\data[79] ),
    .data_out(\data[80] ),
    .latch_enable_in(\latch[79] ),
    .latch_enable_out(\latch[80] ),
    .scan_select_in(\scan[79] ),
    .scan_select_out(\scan[80] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_80 (.clk_in(\clk[80] ),
    .clk_out(\clk[81] ),
    .data_in(\data[80] ),
    .data_out(\data[81] ),
    .latch_enable_in(\latch[80] ),
    .latch_enable_out(\latch[81] ),
    .scan_select_in(\scan[80] ),
    .scan_select_out(\scan[81] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_81 (.clk_in(\clk[81] ),
    .clk_out(\clk[82] ),
    .data_in(\data[81] ),
    .data_out(\data[82] ),
    .latch_enable_in(\latch[81] ),
    .latch_enable_out(\latch[82] ),
    .scan_select_in(\scan[81] ),
    .scan_select_out(\scan[82] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_82 (.clk_in(\clk[82] ),
    .clk_out(\clk[83] ),
    .data_in(\data[82] ),
    .data_out(\data[83] ),
    .latch_enable_in(\latch[82] ),
    .latch_enable_out(\latch[83] ),
    .scan_select_in(\scan[82] ),
    .scan_select_out(\scan[83] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_83 (.clk_in(\clk[83] ),
    .clk_out(\clk[84] ),
    .data_in(\data[83] ),
    .data_out(\data[84] ),
    .latch_enable_in(\latch[83] ),
    .latch_enable_out(\latch[84] ),
    .scan_select_in(\scan[83] ),
    .scan_select_out(\scan[84] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_84 (.clk_in(\clk[84] ),
    .clk_out(\clk[85] ),
    .data_in(\data[84] ),
    .data_out(\data[85] ),
    .latch_enable_in(\latch[84] ),
    .latch_enable_out(\latch[85] ),
    .scan_select_in(\scan[84] ),
    .scan_select_out(\scan[85] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_85 (.clk_in(\clk[85] ),
    .clk_out(\clk[86] ),
    .data_in(\data[85] ),
    .data_out(\data[86] ),
    .latch_enable_in(\latch[85] ),
    .latch_enable_out(\latch[86] ),
    .scan_select_in(\scan[85] ),
    .scan_select_out(\scan[86] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_86 (.clk_in(\clk[86] ),
    .clk_out(\clk[87] ),
    .data_in(\data[86] ),
    .data_out(\data[87] ),
    .latch_enable_in(\latch[86] ),
    .latch_enable_out(\latch[87] ),
    .scan_select_in(\scan[86] ),
    .scan_select_out(\scan[87] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_87 (.clk_in(\clk[87] ),
    .clk_out(\clk[88] ),
    .data_in(\data[87] ),
    .data_out(\data[88] ),
    .latch_enable_in(\latch[87] ),
    .latch_enable_out(\latch[88] ),
    .scan_select_in(\scan[87] ),
    .scan_select_out(\scan[88] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_88 (.clk_in(\clk[88] ),
    .clk_out(\clk[89] ),
    .data_in(\data[88] ),
    .data_out(\data[89] ),
    .latch_enable_in(\latch[88] ),
    .latch_enable_out(\latch[89] ),
    .scan_select_in(\scan[88] ),
    .scan_select_out(\scan[89] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_89 (.clk_in(\clk[89] ),
    .clk_out(\clk[90] ),
    .data_in(\data[89] ),
    .data_out(\data[90] ),
    .latch_enable_in(\latch[89] ),
    .latch_enable_out(\latch[90] ),
    .scan_select_in(\scan[89] ),
    .scan_select_out(\scan[90] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_90 (.clk_in(\clk[90] ),
    .clk_out(\clk[91] ),
    .data_in(\data[90] ),
    .data_out(\data[91] ),
    .latch_enable_in(\latch[90] ),
    .latch_enable_out(\latch[91] ),
    .scan_select_in(\scan[90] ),
    .scan_select_out(\scan[91] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_91 (.clk_in(\clk[91] ),
    .clk_out(\clk[92] ),
    .data_in(\data[91] ),
    .data_out(\data[92] ),
    .latch_enable_in(\latch[91] ),
    .latch_enable_out(\latch[92] ),
    .scan_select_in(\scan[91] ),
    .scan_select_out(\scan[92] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_92 (.clk_in(\clk[92] ),
    .clk_out(\clk[93] ),
    .data_in(\data[92] ),
    .data_out(\data[93] ),
    .latch_enable_in(\latch[92] ),
    .latch_enable_out(\latch[93] ),
    .scan_select_in(\scan[92] ),
    .scan_select_out(\scan[93] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_93 (.clk_in(\clk[93] ),
    .clk_out(\clk[94] ),
    .data_in(\data[93] ),
    .data_out(\data[94] ),
    .latch_enable_in(\latch[93] ),
    .latch_enable_out(\latch[94] ),
    .scan_select_in(\scan[93] ),
    .scan_select_out(\scan[94] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_94 (.clk_in(\clk[94] ),
    .clk_out(\clk[95] ),
    .data_in(\data[94] ),
    .data_out(\data[95] ),
    .latch_enable_in(\latch[94] ),
    .latch_enable_out(\latch[95] ),
    .scan_select_in(\scan[94] ),
    .scan_select_out(\scan[95] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_95 (.clk_in(\clk[95] ),
    .clk_out(\clk[96] ),
    .data_in(\data[95] ),
    .data_out(\data[96] ),
    .latch_enable_in(\latch[95] ),
    .latch_enable_out(\latch[96] ),
    .scan_select_in(\scan[95] ),
    .scan_select_out(\scan[96] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_96 (.clk_in(\clk[96] ),
    .clk_out(\clk[97] ),
    .data_in(\data[96] ),
    .data_out(\data[97] ),
    .latch_enable_in(\latch[96] ),
    .latch_enable_out(\latch[97] ),
    .scan_select_in(\scan[96] ),
    .scan_select_out(\scan[97] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_97 (.clk_in(\clk[97] ),
    .clk_out(\clk[98] ),
    .data_in(\data[97] ),
    .data_out(\data[98] ),
    .latch_enable_in(\latch[97] ),
    .latch_enable_out(\latch[98] ),
    .scan_select_in(\scan[97] ),
    .scan_select_out(\scan[98] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_98 (.clk_in(\clk[98] ),
    .clk_out(\clk[99] ),
    .data_in(\data[98] ),
    .data_out(\data[99] ),
    .latch_enable_in(\latch[98] ),
    .latch_enable_out(\latch[99] ),
    .scan_select_in(\scan[98] ),
    .scan_select_out(\scan[99] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339501025136214612 scan_wrapper_339501025136214612_99 (.clk_in(\clk[99] ),
    .clk_out(\clk[100] ),
    .data_in(\data[99] ),
    .data_out(\data[100] ),
    .latch_enable_in(\latch[99] ),
    .latch_enable_out(\latch[100] ),
    .scan_select_in(\scan[99] ),
    .scan_select_out(\scan[100] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339502597164499540 scan_wrapper_339502597164499540_4 (.clk_in(\clk[4] ),
    .clk_out(\clk[5] ),
    .data_in(\data[4] ),
    .data_out(\data[5] ),
    .latch_enable_in(\latch[4] ),
    .latch_enable_out(\latch[5] ),
    .scan_select_in(\scan[4] ),
    .scan_select_out(\scan[5] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339732875283792466 scan_wrapper_339732875283792466_5 (.clk_in(\clk[5] ),
    .clk_out(\clk[6] ),
    .data_in(\data[5] ),
    .data_out(\data[6] ),
    .latch_enable_in(\latch[5] ),
    .latch_enable_out(\latch[6] ),
    .scan_select_in(\scan[5] ),
    .scan_select_out(\scan[6] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339800239192932947 scan_wrapper_339800239192932947_14 (.clk_in(\clk[14] ),
    .clk_out(\clk[15] ),
    .data_in(\data[14] ),
    .data_out(\data[15] ),
    .latch_enable_in(\latch[14] ),
    .latch_enable_out(\latch[15] ),
    .scan_select_in(\scan[14] ),
    .scan_select_out(\scan[15] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339865743461974612 scan_wrapper_339865743461974612_6 (.clk_in(\clk[6] ),
    .clk_out(\clk[7] ),
    .data_in(\data[6] ),
    .data_out(\data[7] ),
    .latch_enable_in(\latch[6] ),
    .latch_enable_out(\latch[7] ),
    .scan_select_in(\scan[6] ),
    .scan_select_out(\scan[7] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_339898704941023827 scan_wrapper_339898704941023827_7 (.clk_in(\clk[7] ),
    .clk_out(\clk[8] ),
    .data_in(\data[7] ),
    .data_out(\data[8] ),
    .latch_enable_in(\latch[7] ),
    .latch_enable_out(\latch[8] ),
    .scan_select_in(\scan[7] ),
    .scan_select_out(\scan[8] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_340218629792465491 scan_wrapper_340218629792465491_8 (.clk_in(\clk[8] ),
    .clk_out(\clk[9] ),
    .data_in(\data[8] ),
    .data_out(\data[9] ),
    .latch_enable_in(\latch[8] ),
    .latch_enable_out(\latch[9] ),
    .scan_select_in(\scan[8] ),
    .scan_select_out(\scan[9] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_340285391309374034 scan_wrapper_340285391309374034_10 (.clk_in(\clk[10] ),
    .clk_out(\clk[11] ),
    .data_in(\data[10] ),
    .data_out(\data[11] ),
    .latch_enable_in(\latch[10] ),
    .latch_enable_out(\latch[11] ),
    .scan_select_in(\scan[10] ),
    .scan_select_out(\scan[11] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_340318610245288530 scan_wrapper_340318610245288530_9 (.clk_in(\clk[9] ),
    .clk_out(\clk[10] ),
    .data_in(\data[9] ),
    .data_out(\data[10] ),
    .latch_enable_in(\latch[9] ),
    .latch_enable_out(\latch[10] ),
    .scan_select_in(\scan[9] ),
    .scan_select_out(\scan[10] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_340661930553246290 scan_wrapper_340661930553246290_11 (.clk_in(\clk[11] ),
    .clk_out(\clk[12] ),
    .data_in(\data[11] ),
    .data_out(\data[12] ),
    .latch_enable_in(\latch[11] ),
    .latch_enable_out(\latch[12] ),
    .scan_select_in(\scan[11] ),
    .scan_select_out(\scan[12] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_340805072482992722 scan_wrapper_340805072482992722_12 (.clk_in(\clk[12] ),
    .clk_out(\clk[13] ),
    .data_in(\data[12] ),
    .data_out(\data[13] ),
    .latch_enable_in(\latch[12] ),
    .latch_enable_out(\latch[13] ),
    .scan_select_in(\scan[12] ),
    .scan_select_out(\scan[13] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_341136771628663380 scan_wrapper_341136771628663380_13 (.clk_in(\clk[13] ),
    .clk_out(\clk[14] ),
    .data_in(\data[13] ),
    .data_out(\data[14] ),
    .latch_enable_in(\latch[13] ),
    .latch_enable_out(\latch[14] ),
    .scan_select_in(\scan[13] ),
    .scan_select_out(\scan[14] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_341154068332282450 scan_wrapper_341154068332282450_17 (.clk_in(\clk[17] ),
    .clk_out(\clk[18] ),
    .data_in(\data[17] ),
    .data_out(\data[18] ),
    .latch_enable_in(\latch[17] ),
    .latch_enable_out(\latch[18] ),
    .scan_select_in(\scan[17] ),
    .scan_select_out(\scan[18] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_341154161238213203 scan_wrapper_341154161238213203_15 (.clk_in(\clk[15] ),
    .clk_out(\clk[16] ),
    .data_in(\data[15] ),
    .data_out(\data[16] ),
    .latch_enable_in(\latch[15] ),
    .latch_enable_out(\latch[16] ),
    .scan_select_in(\scan[15] ),
    .scan_select_out(\scan[16] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 scan_wrapper_341159915403870803 scan_wrapper_341159915403870803_16 (.clk_in(\clk[16] ),
    .clk_out(\clk[17] ),
    .data_in(\data[16] ),
    .data_out(\data[17] ),
    .latch_enable_in(\latch[16] ),
    .latch_enable_out(\latch[17] ),
    .scan_select_in(\scan[16] ),
    .scan_select_out(\scan[17] ),
    .vccd1(vccd1),
    .vssd1(vssd1));
 assign io_out[10] = slow_clk;
 assign io_out[37] = ready;
endmodule
