VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO scan_wrapper_341263346544149074
  CLASS BLOCK ;
  FOREIGN scan_wrapper_341263346544149074 ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN clk_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 96.000 96.970 100.000 ;
    END
  END clk_in
  PIN clk_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END clk_out
  PIN data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 47.640 100.000 48.240 ;
    END
  END data_in
  PIN data_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END data_out
  PIN latch_enable_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END latch_enable_in
  PIN latch_enable_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 96.000 0.370 100.000 ;
    END
  END latch_enable_out
  PIN scan_select_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 96.000 48.670 100.000 ;
    END
  END scan_select_in
  PIN scan_select_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END scan_select_out
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.550 5.200 21.150 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.200 5.200 50.800 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.855 5.200 80.455 92.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.370 5.200 35.970 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.025 5.200 65.625 92.720 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 94.300 92.565 ;
      LAYER met1 ;
        RECT 0.070 3.440 96.990 93.460 ;
      LAYER met2 ;
        RECT 0.650 95.720 48.110 96.000 ;
        RECT 48.950 95.720 96.410 96.000 ;
        RECT 0.100 4.280 96.960 95.720 ;
        RECT 0.650 3.410 48.110 4.280 ;
        RECT 48.950 3.410 96.410 4.280 ;
      LAYER met3 ;
        RECT 4.000 52.040 96.000 92.645 ;
        RECT 4.400 50.640 96.000 52.040 ;
        RECT 4.000 48.640 96.000 50.640 ;
        RECT 4.000 47.240 95.600 48.640 ;
        RECT 4.000 5.275 96.000 47.240 ;
      LAYER met4 ;
        RECT 10.415 5.200 19.150 92.720 ;
        RECT 21.550 5.200 33.970 92.720 ;
        RECT 36.370 5.200 48.800 92.720 ;
        RECT 51.200 5.200 63.625 92.720 ;
        RECT 66.025 5.200 78.455 92.720 ;
        RECT 80.855 5.200 84.345 92.720 ;
  END
END scan_wrapper_341263346544149074
END LIBRARY

