magic
tech sky130B
magscale 1 2
timestamp 1662389564
<< metal1 >>
rect 37918 700748 37924 700800
rect 37976 700788 37982 700800
rect 105446 700788 105452 700800
rect 37976 700760 105452 700788
rect 37976 700748 37982 700760
rect 105446 700748 105452 700760
rect 105504 700748 105510 700800
rect 65610 700680 65616 700732
rect 65668 700720 65674 700732
rect 267642 700720 267648 700732
rect 65668 700692 267648 700720
rect 65668 700680 65674 700692
rect 267642 700680 267648 700692
rect 267700 700680 267706 700732
rect 65702 700612 65708 700664
rect 65760 700652 65766 700664
rect 332502 700652 332508 700664
rect 65760 700624 332508 700652
rect 65760 700612 65766 700624
rect 332502 700612 332508 700624
rect 332560 700612 332566 700664
rect 95878 700544 95884 700596
rect 95936 700584 95942 700596
rect 364978 700584 364984 700596
rect 95936 700556 364984 700584
rect 95936 700544 95942 700556
rect 364978 700544 364984 700556
rect 365036 700544 365042 700596
rect 13446 700476 13452 700528
rect 13504 700516 13510 700528
rect 300118 700516 300124 700528
rect 13504 700488 300124 700516
rect 13504 700476 13510 700488
rect 300118 700476 300124 700488
rect 300176 700476 300182 700528
rect 378778 700476 378784 700528
rect 378836 700516 378842 700528
rect 397454 700516 397460 700528
rect 378836 700488 397460 700516
rect 378836 700476 378842 700488
rect 397454 700476 397460 700488
rect 397512 700476 397518 700528
rect 71038 700408 71044 700460
rect 71096 700448 71102 700460
rect 170306 700448 170312 700460
rect 71096 700420 170312 700448
rect 71096 700408 71102 700420
rect 170306 700408 170312 700420
rect 170364 700408 170370 700460
rect 205082 700408 205088 700460
rect 205140 700448 205146 700460
rect 494790 700448 494796 700460
rect 205140 700420 494796 700448
rect 205140 700408 205146 700420
rect 494790 700408 494796 700420
rect 494848 700408 494854 700460
rect 65518 700340 65524 700392
rect 65576 700380 65582 700392
rect 137830 700380 137836 700392
rect 65576 700352 137836 700380
rect 65576 700340 65582 700352
rect 137830 700340 137836 700352
rect 137888 700340 137894 700392
rect 152458 700340 152464 700392
rect 152516 700380 152522 700392
rect 462314 700380 462320 700392
rect 152516 700352 462320 700380
rect 152516 700340 152522 700352
rect 462314 700340 462320 700352
rect 462372 700340 462378 700392
rect 518158 700340 518164 700392
rect 518216 700380 518222 700392
rect 527174 700380 527180 700392
rect 518216 700352 527180 700380
rect 518216 700340 518222 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 65794 700272 65800 700324
rect 65852 700312 65858 700324
rect 202782 700312 202788 700324
rect 65852 700284 202788 700312
rect 65852 700272 65858 700284
rect 202782 700272 202788 700284
rect 202840 700272 202846 700324
rect 233878 700272 233884 700324
rect 233936 700312 233942 700324
rect 559650 700312 559656 700324
rect 233936 700284 559656 700312
rect 233936 700272 233942 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 68278 699660 68284 699712
rect 68336 699700 68342 699712
rect 72970 699700 72976 699712
rect 68336 699672 72976 699700
rect 68336 699660 68342 699672
rect 72970 699660 72976 699672
rect 73028 699660 73034 699712
rect 100018 687352 100024 687404
rect 100076 687392 100082 687404
rect 121086 687392 121092 687404
rect 100076 687364 121092 687392
rect 100076 687352 100082 687364
rect 121086 687352 121092 687364
rect 121144 687352 121150 687404
rect 268010 687352 268016 687404
rect 268068 687392 268074 687404
rect 289078 687392 289084 687404
rect 268068 687364 289084 687392
rect 268068 687352 268074 687364
rect 289078 687352 289084 687364
rect 289136 687352 289142 687404
rect 380342 687352 380348 687404
rect 380400 687392 380406 687404
rect 401134 687392 401140 687404
rect 380400 687364 401140 687392
rect 380400 687352 380406 687364
rect 401134 687352 401140 687364
rect 401192 687352 401198 687404
rect 464338 687352 464344 687404
rect 464396 687392 464402 687404
rect 485038 687392 485044 687404
rect 464396 687364 485044 687392
rect 464396 687352 464402 687364
rect 485038 687352 485044 687364
rect 485096 687352 485102 687404
rect 36906 687284 36912 687336
rect 36964 687324 36970 687336
rect 54294 687324 54300 687336
rect 36964 687296 54300 687324
rect 36964 687284 36970 687296
rect 54294 687284 54300 687296
rect 54352 687284 54358 687336
rect 65886 687284 65892 687336
rect 65944 687324 65950 687336
rect 81986 687324 81992 687336
rect 65944 687296 81992 687324
rect 65944 687284 65950 687296
rect 81986 687284 81992 687296
rect 82044 687284 82050 687336
rect 92934 687284 92940 687336
rect 92992 687324 92998 687336
rect 110322 687324 110328 687336
rect 92992 687296 110328 687324
rect 92992 687284 92998 687296
rect 110322 687284 110328 687296
rect 110380 687284 110386 687336
rect 176930 687284 176936 687336
rect 176988 687324 176994 687336
rect 194318 687324 194324 687336
rect 176988 687296 194324 687324
rect 176988 687284 176994 687296
rect 194318 687284 194324 687296
rect 194376 687284 194382 687336
rect 261478 687284 261484 687336
rect 261536 687324 261542 687336
rect 278314 687324 278320 687336
rect 261536 687296 278320 687324
rect 261536 687284 261542 687296
rect 278314 687284 278320 687296
rect 278372 687284 278378 687336
rect 317138 687284 317144 687336
rect 317196 687324 317202 687336
rect 334342 687324 334348 687336
rect 317196 687296 334348 687324
rect 317196 687284 317202 687296
rect 334342 687284 334348 687296
rect 334400 687284 334406 687336
rect 372982 687284 372988 687336
rect 373040 687324 373046 687336
rect 390002 687324 390008 687336
rect 373040 687296 390008 687324
rect 373040 687284 373046 687296
rect 390002 687284 390008 687296
rect 390060 687284 390066 687336
rect 457438 687284 457444 687336
rect 457496 687324 457502 687336
rect 473998 687324 474004 687336
rect 457496 687296 474004 687324
rect 457496 687284 457502 687296
rect 473998 687284 474004 687296
rect 474056 687284 474062 687336
rect 15286 687216 15292 687268
rect 15344 687256 15350 687268
rect 26326 687256 26332 687268
rect 15344 687228 26332 687256
rect 15344 687216 15350 687228
rect 26326 687216 26332 687228
rect 26384 687216 26390 687268
rect 39298 687216 39304 687268
rect 39356 687256 39362 687268
rect 64598 687256 64604 687268
rect 39356 687228 64604 687256
rect 39356 687216 39362 687228
rect 64598 687216 64604 687228
rect 64656 687216 64662 687268
rect 72326 687216 72332 687268
rect 72384 687256 72390 687268
rect 93118 687256 93124 687268
rect 72384 687228 93124 687256
rect 72384 687216 72390 687228
rect 93118 687216 93124 687228
rect 93176 687216 93182 687268
rect 120994 687216 121000 687268
rect 121052 687256 121058 687268
rect 138290 687256 138296 687268
rect 121052 687228 138296 687256
rect 121052 687216 121058 687228
rect 138290 687216 138296 687228
rect 138348 687216 138354 687268
rect 156322 687216 156328 687268
rect 156380 687256 156386 687268
rect 177298 687256 177304 687268
rect 156380 687228 177304 687256
rect 156380 687216 156386 687228
rect 177298 687216 177304 687228
rect 177356 687216 177362 687268
rect 184014 687216 184020 687268
rect 184072 687256 184078 687268
rect 204714 687256 204720 687268
rect 184072 687228 204720 687256
rect 184072 687216 184078 687228
rect 204714 687216 204720 687228
rect 204772 687216 204778 687268
rect 209038 687216 209044 687268
rect 209096 687256 209102 687268
rect 222194 687256 222200 687268
rect 209096 687228 222200 687256
rect 209096 687216 209102 687228
rect 222194 687216 222200 687228
rect 222252 687216 222258 687268
rect 232958 687216 232964 687268
rect 233016 687256 233022 687268
rect 250346 687256 250352 687268
rect 233016 687228 250352 687256
rect 233016 687216 233022 687228
rect 250346 687216 250352 687228
rect 250404 687216 250410 687268
rect 288986 687216 288992 687268
rect 289044 687256 289050 687268
rect 306006 687256 306012 687268
rect 289044 687228 306012 687256
rect 289044 687216 289050 687228
rect 306006 687216 306012 687228
rect 306064 687216 306070 687268
rect 317046 687216 317052 687268
rect 317104 687256 317110 687268
rect 344646 687256 344652 687268
rect 317104 687228 344652 687256
rect 317104 687216 317110 687228
rect 344646 687216 344652 687228
rect 344704 687216 344710 687268
rect 352006 687216 352012 687268
rect 352064 687256 352070 687268
rect 373258 687256 373264 687268
rect 352064 687228 373264 687256
rect 352064 687216 352070 687228
rect 373258 687216 373264 687228
rect 373316 687216 373322 687268
rect 401042 687216 401048 687268
rect 401100 687256 401106 687268
rect 418338 687256 418344 687268
rect 401100 687228 418344 687256
rect 401100 687216 401106 687228
rect 418338 687216 418344 687228
rect 418396 687216 418402 687268
rect 429838 687216 429844 687268
rect 429896 687256 429902 687268
rect 456610 687256 456616 687268
rect 429896 687228 456616 687256
rect 429896 687216 429902 687228
rect 456610 687216 456616 687228
rect 456668 687216 456674 687268
rect 484946 687216 484952 687268
rect 485004 687256 485010 687268
rect 502334 687256 502340 687268
rect 485004 687228 502340 687256
rect 485004 687216 485010 687228
rect 502334 687216 502340 687228
rect 502392 687216 502398 687268
rect 512914 687216 512920 687268
rect 512972 687256 512978 687268
rect 530302 687256 530308 687268
rect 512972 687228 530308 687256
rect 512972 687216 512978 687228
rect 530302 687216 530308 687228
rect 530360 687216 530366 687268
rect 92750 684224 92756 684276
rect 92808 684264 92814 684276
rect 92934 684264 92940 684276
rect 92808 684236 92940 684264
rect 92808 684224 92814 684236
rect 92934 684224 92940 684236
rect 92992 684224 92998 684276
rect 120718 684224 120724 684276
rect 120776 684264 120782 684276
rect 120994 684264 121000 684276
rect 120776 684236 121000 684264
rect 120776 684224 120782 684236
rect 120994 684224 121000 684236
rect 121052 684224 121058 684276
rect 204714 684224 204720 684276
rect 204772 684264 204778 684276
rect 204990 684264 204996 684276
rect 204772 684236 204996 684264
rect 204772 684224 204778 684236
rect 204990 684224 204996 684236
rect 205048 684224 205054 684276
rect 232774 684224 232780 684276
rect 232832 684264 232838 684276
rect 232958 684264 232964 684276
rect 232832 684236 232964 684264
rect 232832 684224 232838 684236
rect 232958 684224 232964 684236
rect 233016 684224 233022 684276
rect 316862 684224 316868 684276
rect 316920 684264 316926 684276
rect 317046 684264 317052 684276
rect 316920 684236 317052 684264
rect 316920 684224 316926 684236
rect 317046 684224 317052 684236
rect 317104 684224 317110 684276
rect 372798 684224 372804 684276
rect 372856 684264 372862 684276
rect 372982 684264 372988 684276
rect 372856 684236 372988 684264
rect 372856 684224 372862 684236
rect 372982 684224 372988 684236
rect 373040 684224 373046 684276
rect 400766 684224 400772 684276
rect 400824 684264 400830 684276
rect 401042 684264 401048 684276
rect 400824 684236 401048 684264
rect 400824 684224 400830 684236
rect 401042 684224 401048 684236
rect 401100 684224 401106 684276
rect 120810 684156 120816 684208
rect 120868 684196 120874 684208
rect 121086 684196 121092 684208
rect 120868 684168 121092 684196
rect 120868 684156 120874 684168
rect 121086 684156 121092 684168
rect 121144 684156 121150 684208
rect 316770 684156 316776 684208
rect 316828 684196 316834 684208
rect 317138 684196 317144 684208
rect 316828 684168 317144 684196
rect 316828 684156 316834 684168
rect 317138 684156 317144 684168
rect 317196 684156 317202 684208
rect 400858 684156 400864 684208
rect 400916 684196 400922 684208
rect 401134 684196 401140 684208
rect 400916 684168 401140 684196
rect 400916 684156 400922 684168
rect 401134 684156 401140 684168
rect 401192 684156 401198 684208
rect 176746 683272 176752 683324
rect 176804 683272 176810 683324
rect 176764 683108 176792 683272
rect 288802 683136 288808 683188
rect 288860 683136 288866 683188
rect 484854 683136 484860 683188
rect 484912 683136 484918 683188
rect 512822 683136 512828 683188
rect 512880 683136 512886 683188
rect 176838 683108 176844 683120
rect 176764 683080 176844 683108
rect 176838 683068 176844 683080
rect 176896 683068 176902 683120
rect 288820 682972 288848 683136
rect 484872 682984 484900 683136
rect 512840 682984 512868 683136
rect 288894 682972 288900 682984
rect 288820 682944 288900 682972
rect 288894 682932 288900 682944
rect 288952 682932 288958 682984
rect 484854 682932 484860 682984
rect 484912 682932 484918 682984
rect 512822 682932 512828 682984
rect 512880 682932 512886 682984
rect 512730 682592 512736 682644
rect 512788 682632 512794 682644
rect 512914 682632 512920 682644
rect 512788 682604 512920 682632
rect 512788 682592 512794 682604
rect 512914 682592 512920 682604
rect 512972 682592 512978 682644
rect 204806 681708 204812 681760
rect 204864 681748 204870 681760
rect 209038 681748 209044 681760
rect 204864 681720 209044 681748
rect 204864 681708 204870 681720
rect 209038 681708 209044 681720
rect 209096 681708 209102 681760
rect 288802 681028 288808 681080
rect 288860 681068 288866 681080
rect 288986 681068 288992 681080
rect 288860 681040 288992 681068
rect 288860 681028 288866 681040
rect 288986 681028 288992 681040
rect 289044 681028 289050 681080
rect 176746 679464 176752 679516
rect 176804 679504 176810 679516
rect 176930 679504 176936 679516
rect 176804 679476 176936 679504
rect 176804 679464 176810 679476
rect 176930 679464 176936 679476
rect 176988 679464 176994 679516
rect 484762 677900 484768 677952
rect 484820 677940 484826 677952
rect 484946 677940 484952 677952
rect 484820 677912 484952 677940
rect 484820 677900 484826 677912
rect 484946 677900 484952 677912
rect 485004 677900 485010 677952
rect 64874 669060 64880 669112
rect 64932 669100 64938 669112
rect 65886 669100 65892 669112
rect 64932 669072 65892 669100
rect 64932 669060 64938 669072
rect 65886 669060 65892 669072
rect 65944 669060 65950 669112
rect 36814 668584 36820 668636
rect 36872 668624 36878 668636
rect 36998 668624 37004 668636
rect 36872 668596 37004 668624
rect 36872 668584 36878 668596
rect 36998 668584 37004 668596
rect 37056 668584 37062 668636
rect 204898 667836 204904 667888
rect 204956 667876 204962 667888
rect 211706 667876 211712 667888
rect 204956 667848 211712 667876
rect 204956 667836 204962 667848
rect 211706 667836 211712 667848
rect 211764 667836 211770 667888
rect 485038 667836 485044 667888
rect 485096 667876 485102 667888
rect 491662 667876 491668 667888
rect 485096 667848 491668 667876
rect 485096 667836 485102 667848
rect 491662 667836 491668 667848
rect 491720 667836 491726 667888
rect 289078 667360 289084 667412
rect 289136 667400 289142 667412
rect 295702 667400 295708 667412
rect 289136 667372 295708 667400
rect 289136 667360 289142 667372
rect 295702 667360 295708 667372
rect 295760 667360 295766 667412
rect 93118 667156 93124 667208
rect 93176 667196 93182 667208
rect 99742 667196 99748 667208
rect 93176 667168 99748 667196
rect 93176 667156 93182 667168
rect 99742 667156 99748 667168
rect 99800 667156 99806 667208
rect 120810 667156 120816 667208
rect 120868 667196 120874 667208
rect 127710 667196 127716 667208
rect 120868 667168 127716 667196
rect 120868 667156 120874 667168
rect 127710 667156 127716 667168
rect 127768 667156 127774 667208
rect 177298 667156 177304 667208
rect 177356 667196 177362 667208
rect 183646 667196 183652 667208
rect 177356 667168 183652 667196
rect 177356 667156 177362 667168
rect 183646 667156 183652 667168
rect 183704 667156 183710 667208
rect 373258 667156 373264 667208
rect 373316 667196 373322 667208
rect 379698 667196 379704 667208
rect 373316 667168 379704 667196
rect 373316 667156 373322 667168
rect 379698 667156 379704 667168
rect 379756 667156 379762 667208
rect 400858 667156 400864 667208
rect 400916 667196 400922 667208
rect 407758 667196 407764 667208
rect 400916 667168 407764 667196
rect 400916 667156 400922 667168
rect 407758 667156 407764 667168
rect 407816 667156 407822 667208
rect 42702 665116 42708 665168
rect 42760 665156 42766 665168
rect 95234 665156 95240 665168
rect 42760 665128 95240 665156
rect 42760 665116 42766 665128
rect 95234 665116 95240 665128
rect 95292 665116 95298 665168
rect 97902 665116 97908 665168
rect 97960 665156 97966 665168
rect 150434 665156 150440 665168
rect 97960 665128 150440 665156
rect 97960 665116 97966 665128
rect 150434 665116 150440 665128
rect 150492 665116 150498 665168
rect 154482 665116 154488 665168
rect 154540 665156 154546 665168
rect 207014 665156 207020 665168
rect 154540 665128 207020 665156
rect 154540 665116 154546 665128
rect 207014 665116 207020 665128
rect 207072 665116 207078 665168
rect 209682 665116 209688 665168
rect 209740 665156 209746 665168
rect 262214 665156 262220 665168
rect 209740 665128 262220 665156
rect 209740 665116 209746 665128
rect 262214 665116 262220 665128
rect 262272 665116 262278 665168
rect 266262 665116 266268 665168
rect 266320 665156 266326 665168
rect 318794 665156 318800 665168
rect 266320 665128 318800 665156
rect 266320 665116 266326 665128
rect 318794 665116 318800 665128
rect 318852 665116 318858 665168
rect 322842 665116 322848 665168
rect 322900 665156 322906 665168
rect 375374 665156 375380 665168
rect 322900 665128 375380 665156
rect 322900 665116 322906 665128
rect 375374 665116 375380 665128
rect 375432 665116 375438 665168
rect 378042 665116 378048 665168
rect 378100 665156 378106 665168
rect 430574 665156 430580 665168
rect 378100 665128 430580 665156
rect 378100 665116 378106 665128
rect 430574 665116 430580 665128
rect 430632 665116 430638 665168
rect 434622 665116 434628 665168
rect 434680 665156 434686 665168
rect 487154 665156 487160 665168
rect 434680 665128 487160 665156
rect 434680 665116 434686 665128
rect 487154 665116 487160 665128
rect 487212 665116 487218 665168
rect 489822 665116 489828 665168
rect 489880 665156 489886 665168
rect 542354 665156 542360 665168
rect 489880 665128 542360 665156
rect 489880 665116 489886 665128
rect 542354 665116 542360 665128
rect 542412 665116 542418 665168
rect 15286 664708 15292 664760
rect 15344 664748 15350 664760
rect 16114 664748 16120 664760
rect 15344 664720 16120 664748
rect 15344 664708 15350 664720
rect 16114 664708 16120 664720
rect 16172 664708 16178 664760
rect 36538 664708 36544 664760
rect 36596 664748 36602 664760
rect 36906 664748 36912 664760
rect 36596 664720 36912 664748
rect 36596 664708 36602 664720
rect 36906 664708 36912 664720
rect 36964 664708 36970 664760
rect 15378 662328 15384 662380
rect 15436 662368 15442 662380
rect 43622 662368 43628 662380
rect 15436 662340 43628 662368
rect 15436 662328 15442 662340
rect 43622 662328 43628 662340
rect 43680 662328 43686 662380
rect 138658 662328 138664 662380
rect 138716 662368 138722 662380
rect 176838 662368 176844 662380
rect 138716 662340 176844 662368
rect 138716 662328 138722 662340
rect 176838 662328 176844 662340
rect 176896 662328 176902 662380
rect 194318 662328 194324 662380
rect 194376 662368 194382 662380
rect 232866 662368 232872 662380
rect 194376 662340 232872 662368
rect 194376 662328 194382 662340
rect 232866 662328 232872 662340
rect 232924 662328 232930 662380
rect 238846 662328 238852 662380
rect 238904 662368 238910 662380
rect 238904 662340 248414 662368
rect 238904 662328 238910 662340
rect 26326 662260 26332 662312
rect 26384 662300 26390 662312
rect 39298 662300 39304 662312
rect 26384 662272 39304 662300
rect 26384 662260 26390 662272
rect 39298 662260 39304 662272
rect 39356 662260 39362 662312
rect 42886 662260 42892 662312
rect 42944 662300 42950 662312
rect 71774 662300 71780 662312
rect 42944 662272 71780 662300
rect 42944 662260 42950 662272
rect 71774 662260 71780 662272
rect 71832 662260 71838 662312
rect 82630 662260 82636 662312
rect 82688 662300 82694 662312
rect 120902 662300 120908 662312
rect 82688 662272 120908 662300
rect 82688 662260 82694 662272
rect 120902 662260 120908 662272
rect 120960 662260 120966 662312
rect 127066 662260 127072 662312
rect 127124 662300 127130 662312
rect 155954 662300 155960 662312
rect 127124 662272 155960 662300
rect 127124 662260 127130 662272
rect 155954 662260 155960 662272
rect 156012 662260 156018 662312
rect 166626 662260 166632 662312
rect 166684 662300 166690 662312
rect 204990 662300 204996 662312
rect 166684 662272 204996 662300
rect 166684 662260 166690 662272
rect 204990 662260 204996 662272
rect 205048 662260 205054 662312
rect 211246 662260 211252 662312
rect 211304 662300 211310 662312
rect 239766 662300 239772 662312
rect 211304 662272 239772 662300
rect 211304 662260 211310 662272
rect 239766 662260 239772 662272
rect 239824 662260 239830 662312
rect 248386 662300 248414 662340
rect 295426 662328 295432 662380
rect 295484 662368 295490 662380
rect 323670 662368 323676 662380
rect 295484 662340 323676 662368
rect 295484 662328 295490 662340
rect 323670 662328 323676 662340
rect 323728 662328 323734 662380
rect 334618 662328 334624 662380
rect 334676 662368 334682 662380
rect 372890 662368 372896 662380
rect 334676 662340 372896 662368
rect 334676 662328 334682 662340
rect 372890 662328 372896 662340
rect 372948 662328 372954 662380
rect 390462 662328 390468 662380
rect 390520 662368 390526 662380
rect 428734 662368 428740 662380
rect 390520 662340 428740 662368
rect 390520 662328 390526 662340
rect 428734 662328 428740 662340
rect 428792 662328 428798 662380
rect 434806 662328 434812 662380
rect 434864 662368 434870 662380
rect 434864 662340 441614 662368
rect 434864 662328 434870 662340
rect 268010 662300 268016 662312
rect 248386 662272 268016 662300
rect 268010 662260 268016 662272
rect 268068 662260 268074 662312
rect 278314 662260 278320 662312
rect 278372 662300 278378 662312
rect 316954 662300 316960 662312
rect 278372 662272 316960 662300
rect 278372 662260 278378 662272
rect 316954 662260 316960 662272
rect 317012 662260 317018 662312
rect 323026 662260 323032 662312
rect 323084 662300 323090 662312
rect 352006 662300 352012 662312
rect 323084 662272 352012 662300
rect 323084 662260 323090 662272
rect 352006 662260 352012 662272
rect 352064 662260 352070 662312
rect 362310 662260 362316 662312
rect 362368 662300 362374 662312
rect 400950 662300 400956 662312
rect 362368 662272 400956 662300
rect 362368 662260 362374 662272
rect 400950 662260 400956 662272
rect 401008 662260 401014 662312
rect 407206 662260 407212 662312
rect 407264 662300 407270 662312
rect 436002 662300 436008 662312
rect 407264 662272 436008 662300
rect 407264 662260 407270 662272
rect 436002 662260 436008 662272
rect 436060 662260 436066 662312
rect 441586 662300 441614 662340
rect 491386 662328 491392 662380
rect 491444 662368 491450 662380
rect 519998 662368 520004 662380
rect 491444 662340 520004 662368
rect 491444 662328 491450 662340
rect 519998 662328 520004 662340
rect 520056 662328 520062 662380
rect 530302 662328 530308 662380
rect 530360 662368 530366 662380
rect 568758 662368 568764 662380
rect 530360 662340 568764 662368
rect 530360 662328 530366 662340
rect 568758 662328 568764 662340
rect 568816 662328 568822 662380
rect 463786 662300 463792 662312
rect 441586 662272 463792 662300
rect 463786 662260 463792 662272
rect 463844 662260 463850 662312
rect 474642 662260 474648 662312
rect 474700 662300 474706 662312
rect 512822 662300 512828 662312
rect 474700 662272 512828 662300
rect 474700 662260 474706 662272
rect 512822 662260 512828 662272
rect 512880 662260 512886 662312
rect 518986 662260 518992 662312
rect 519044 662300 519050 662312
rect 547874 662300 547880 662312
rect 519044 662272 547880 662300
rect 519044 662260 519050 662272
rect 547874 662260 547880 662272
rect 547932 662260 547938 662312
rect 54570 662192 54576 662244
rect 54628 662232 54634 662244
rect 92842 662232 92848 662244
rect 54628 662204 92848 662232
rect 54628 662192 54634 662204
rect 92842 662192 92848 662204
rect 92900 662192 92906 662244
rect 110322 662192 110328 662244
rect 110380 662232 110386 662244
rect 148778 662232 148784 662244
rect 110380 662204 148784 662232
rect 110380 662192 110386 662204
rect 148778 662192 148784 662204
rect 148836 662192 148842 662244
rect 250714 662192 250720 662244
rect 250772 662232 250778 662244
rect 288894 662232 288900 662244
rect 250772 662204 288900 662232
rect 250772 662192 250778 662204
rect 288894 662192 288900 662204
rect 288952 662192 288958 662244
rect 306282 662192 306288 662244
rect 306340 662232 306346 662244
rect 316862 662232 316868 662244
rect 306340 662204 316868 662232
rect 306340 662192 306346 662204
rect 316862 662192 316868 662204
rect 316920 662192 316926 662244
rect 418338 662192 418344 662244
rect 418396 662232 418402 662244
rect 429838 662232 429844 662244
rect 418396 662204 429844 662232
rect 418396 662192 418402 662204
rect 429838 662192 429844 662204
rect 429896 662192 429902 662244
rect 446306 662192 446312 662244
rect 446364 662232 446370 662244
rect 484854 662232 484860 662244
rect 446364 662204 484860 662232
rect 446364 662192 446370 662204
rect 484854 662192 484860 662204
rect 484912 662192 484918 662244
rect 502334 662192 502340 662244
rect 502392 662232 502398 662244
rect 540790 662232 540796 662244
rect 502392 662204 540796 662232
rect 502392 662192 502398 662204
rect 540790 662192 540796 662204
rect 540848 662192 540854 662244
rect 13630 661648 13636 661700
rect 13688 661688 13694 661700
rect 557994 661688 558000 661700
rect 13688 661660 558000 661688
rect 13688 661648 13694 661660
rect 557994 661648 558000 661660
rect 558052 661648 558058 661700
rect 26602 660288 26608 660340
rect 26660 660328 26666 660340
rect 36814 660328 36820 660340
rect 26660 660300 36820 660328
rect 26660 660288 26666 660300
rect 36814 660288 36820 660300
rect 36872 660288 36878 660340
rect 38010 659744 38016 659796
rect 38068 659784 38074 659796
rect 44174 659784 44180 659796
rect 38068 659756 44180 659784
rect 38068 659744 38074 659756
rect 44174 659744 44180 659756
rect 44232 659744 44238 659796
rect 71866 659744 71872 659796
rect 71924 659784 71930 659796
rect 110598 659784 110604 659796
rect 71924 659756 110604 659784
rect 71924 659744 71930 659756
rect 110598 659744 110604 659756
rect 110656 659744 110662 659796
rect 211246 659744 211252 659796
rect 211304 659784 211310 659796
rect 250622 659784 250628 659796
rect 211304 659756 250628 659784
rect 211304 659744 211310 659756
rect 250622 659744 250628 659756
rect 250680 659744 250686 659796
rect 295426 659744 295432 659796
rect 295484 659784 295490 659796
rect 334618 659784 334624 659796
rect 295484 659756 334624 659784
rect 295484 659744 295490 659756
rect 334618 659744 334624 659756
rect 334676 659744 334682 659796
rect 407206 659744 407212 659796
rect 407264 659784 407270 659796
rect 446306 659784 446312 659796
rect 407264 659756 446312 659784
rect 407264 659744 407270 659756
rect 446306 659744 446312 659756
rect 446364 659744 446370 659796
rect 491386 659744 491392 659796
rect 491444 659784 491450 659796
rect 530302 659784 530308 659796
rect 491444 659756 530308 659784
rect 491444 659744 491450 659756
rect 530302 659744 530308 659756
rect 530360 659744 530366 659796
rect 15562 659676 15568 659728
rect 15620 659716 15626 659728
rect 54294 659716 54300 659728
rect 15620 659688 54300 659716
rect 15620 659676 15626 659688
rect 54294 659676 54300 659688
rect 54352 659676 54358 659728
rect 99466 659676 99472 659728
rect 99524 659716 99530 659728
rect 138290 659716 138296 659728
rect 99524 659688 138296 659716
rect 99524 659676 99530 659688
rect 138290 659676 138296 659688
rect 138348 659676 138354 659728
rect 149790 659676 149796 659728
rect 149848 659716 149854 659728
rect 166626 659716 166632 659728
rect 149848 659688 166632 659716
rect 149848 659676 149854 659688
rect 166626 659676 166632 659688
rect 166684 659676 166690 659728
rect 183646 659676 183652 659728
rect 183704 659716 183710 659728
rect 222286 659716 222292 659728
rect 183704 659688 222292 659716
rect 183704 659676 183710 659688
rect 222286 659676 222292 659688
rect 222344 659676 222350 659728
rect 233970 659676 233976 659728
rect 234028 659716 234034 659728
rect 240318 659716 240324 659728
rect 234028 659688 240324 659716
rect 234028 659676 234034 659688
rect 240318 659676 240324 659688
rect 240376 659676 240382 659728
rect 267826 659676 267832 659728
rect 267884 659716 267890 659728
rect 306466 659716 306472 659728
rect 267884 659688 306472 659716
rect 267884 659676 267890 659688
rect 306466 659676 306472 659688
rect 306524 659676 306530 659728
rect 318058 659676 318064 659728
rect 318116 659716 318122 659728
rect 324314 659716 324320 659728
rect 318116 659688 324320 659716
rect 318116 659676 318122 659688
rect 324314 659676 324320 659688
rect 324372 659676 324378 659728
rect 345750 659676 345756 659728
rect 345808 659716 345814 659728
rect 362310 659716 362316 659728
rect 345808 659688 362316 659716
rect 345808 659676 345814 659688
rect 362310 659676 362316 659688
rect 362368 659676 362374 659728
rect 379606 659676 379612 659728
rect 379664 659716 379670 659728
rect 418614 659716 418620 659728
rect 379664 659688 418620 659716
rect 379664 659676 379670 659688
rect 418614 659676 418620 659688
rect 418672 659676 418678 659728
rect 429838 659676 429844 659728
rect 429896 659716 429902 659728
rect 436094 659716 436100 659728
rect 429896 659688 436100 659716
rect 429896 659676 429902 659688
rect 436094 659676 436100 659688
rect 436152 659676 436158 659728
rect 463786 659676 463792 659728
rect 463844 659716 463850 659728
rect 502610 659716 502616 659728
rect 463844 659688 502616 659716
rect 463844 659676 463850 659688
rect 502610 659676 502616 659688
rect 502668 659676 502674 659728
rect 541618 659676 541624 659728
rect 541676 659716 541682 659728
rect 558638 659716 558644 659728
rect 541676 659688 558644 659716
rect 541676 659676 541682 659688
rect 558638 659676 558644 659688
rect 558696 659676 558702 659728
rect 205082 657296 205088 657348
rect 205140 657296 205146 657348
rect 205100 657144 205128 657296
rect 205082 657092 205088 657144
rect 205140 657092 205146 657144
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 11698 656928 11704 656940
rect 3568 656900 11704 656928
rect 3568 656888 3574 656900
rect 11698 656888 11704 656900
rect 11756 656888 11762 656940
rect 42702 656888 42708 656940
rect 42760 656928 42766 656940
rect 95234 656928 95240 656940
rect 42760 656900 95240 656928
rect 42760 656888 42766 656900
rect 95234 656888 95240 656900
rect 95292 656888 95298 656940
rect 97902 656888 97908 656940
rect 97960 656928 97966 656940
rect 150434 656928 150440 656940
rect 97960 656900 150440 656928
rect 97960 656888 97966 656900
rect 150434 656888 150440 656900
rect 150492 656888 150498 656940
rect 154482 656888 154488 656940
rect 154540 656928 154546 656940
rect 207014 656928 207020 656940
rect 154540 656900 207020 656928
rect 154540 656888 154546 656900
rect 207014 656888 207020 656900
rect 207072 656888 207078 656940
rect 209682 656888 209688 656940
rect 209740 656928 209746 656940
rect 262214 656928 262220 656940
rect 209740 656900 262220 656928
rect 209740 656888 209746 656900
rect 262214 656888 262220 656900
rect 262272 656888 262278 656940
rect 266262 656888 266268 656940
rect 266320 656928 266326 656940
rect 318794 656928 318800 656940
rect 266320 656900 318800 656928
rect 266320 656888 266326 656900
rect 318794 656888 318800 656900
rect 318852 656888 318858 656940
rect 322842 656888 322848 656940
rect 322900 656928 322906 656940
rect 375374 656928 375380 656940
rect 322900 656900 375380 656928
rect 322900 656888 322906 656900
rect 375374 656888 375380 656900
rect 375432 656888 375438 656940
rect 378042 656888 378048 656940
rect 378100 656928 378106 656940
rect 430574 656928 430580 656940
rect 378100 656900 430580 656928
rect 378100 656888 378106 656900
rect 430574 656888 430580 656900
rect 430632 656888 430638 656940
rect 434622 656888 434628 656940
rect 434680 656928 434686 656940
rect 487154 656928 487160 656940
rect 434680 656900 487160 656928
rect 434680 656888 434686 656900
rect 487154 656888 487160 656900
rect 487212 656888 487218 656940
rect 489822 656888 489828 656940
rect 489880 656928 489886 656940
rect 542354 656928 542360 656940
rect 489880 656900 542360 656928
rect 489880 656888 489886 656900
rect 542354 656888 542360 656900
rect 542412 656888 542418 656940
rect 71774 655664 71780 655716
rect 71832 655704 71838 655716
rect 71958 655704 71964 655716
rect 71832 655676 71964 655704
rect 71832 655664 71838 655676
rect 71958 655664 71964 655676
rect 72016 655664 72022 655716
rect 99374 655664 99380 655716
rect 99432 655704 99438 655716
rect 99926 655704 99932 655716
rect 99432 655676 99932 655704
rect 99432 655664 99438 655676
rect 99926 655664 99932 655676
rect 99984 655664 99990 655716
rect 183554 655664 183560 655716
rect 183612 655704 183618 655716
rect 184014 655704 184020 655716
rect 183612 655676 184020 655704
rect 183612 655664 183618 655676
rect 184014 655664 184020 655676
rect 184072 655664 184078 655716
rect 211154 655664 211160 655716
rect 211212 655704 211218 655716
rect 211982 655704 211988 655716
rect 211212 655676 211988 655704
rect 211212 655664 211218 655676
rect 211982 655664 211988 655676
rect 212040 655664 212046 655716
rect 267734 655664 267740 655716
rect 267792 655704 267798 655716
rect 267918 655704 267924 655716
rect 267792 655676 267924 655704
rect 267792 655664 267798 655676
rect 267918 655664 267924 655676
rect 267976 655664 267982 655716
rect 295334 655664 295340 655716
rect 295392 655704 295398 655716
rect 295978 655704 295984 655716
rect 295392 655676 295984 655704
rect 295392 655664 295398 655676
rect 295978 655664 295984 655676
rect 296036 655664 296042 655716
rect 379514 655664 379520 655716
rect 379572 655704 379578 655716
rect 379974 655704 379980 655716
rect 379572 655676 379980 655704
rect 379572 655664 379578 655676
rect 379974 655664 379980 655676
rect 380032 655664 380038 655716
rect 407114 655664 407120 655716
rect 407172 655704 407178 655716
rect 407942 655704 407948 655716
rect 407172 655676 407948 655704
rect 407172 655664 407178 655676
rect 407942 655664 407948 655676
rect 408000 655664 408006 655716
rect 463694 655664 463700 655716
rect 463752 655704 463758 655716
rect 464062 655704 464068 655716
rect 463752 655676 464068 655704
rect 463752 655664 463758 655676
rect 464062 655664 464068 655676
rect 464120 655664 464126 655716
rect 491294 655664 491300 655716
rect 491352 655704 491358 655716
rect 492030 655704 492036 655716
rect 491352 655676 492036 655704
rect 491352 655664 491358 655676
rect 492030 655664 492036 655676
rect 492088 655664 492094 655716
rect 15194 634720 15200 634772
rect 15252 634760 15258 634772
rect 36906 634760 36912 634772
rect 15252 634732 36912 634760
rect 15252 634720 15258 634732
rect 36906 634720 36912 634732
rect 36964 634720 36970 634772
rect 37090 634720 37096 634772
rect 37148 634760 37154 634772
rect 64874 634760 64880 634772
rect 37148 634732 64880 634760
rect 37148 634720 37154 634732
rect 64874 634720 64880 634732
rect 64932 634720 64938 634772
rect 65058 634720 65064 634772
rect 65116 634760 65122 634772
rect 92934 634760 92940 634772
rect 65116 634732 92940 634760
rect 65116 634720 65122 634732
rect 92934 634720 92940 634732
rect 92992 634720 92998 634772
rect 93026 634720 93032 634772
rect 93084 634760 93090 634772
rect 120902 634760 120908 634772
rect 93084 634732 120908 634760
rect 93084 634720 93090 634732
rect 120902 634720 120908 634732
rect 120960 634720 120966 634772
rect 121086 634720 121092 634772
rect 121144 634760 121150 634772
rect 148594 634760 148600 634772
rect 121144 634732 148600 634760
rect 121144 634720 121150 634732
rect 148594 634720 148600 634732
rect 148652 634720 148658 634772
rect 149698 634720 149704 634772
rect 149756 634760 149762 634772
rect 176930 634760 176936 634772
rect 149756 634732 176936 634760
rect 149756 634720 149762 634732
rect 176930 634720 176936 634732
rect 176988 634720 176994 634772
rect 177022 634720 177028 634772
rect 177080 634760 177086 634772
rect 204898 634760 204904 634772
rect 177080 634732 204904 634760
rect 177080 634720 177086 634732
rect 204898 634720 204904 634732
rect 204956 634720 204962 634772
rect 205174 634720 205180 634772
rect 205232 634760 205238 634772
rect 232590 634760 232596 634772
rect 205232 634732 232596 634760
rect 205232 634720 205238 634732
rect 232590 634720 232596 634732
rect 232648 634720 232654 634772
rect 233050 634720 233056 634772
rect 233108 634760 233114 634772
rect 260926 634760 260932 634772
rect 233108 634732 260932 634760
rect 233108 634720 233114 634732
rect 260926 634720 260932 634732
rect 260984 634720 260990 634772
rect 261018 634720 261024 634772
rect 261076 634760 261082 634772
rect 288894 634760 288900 634772
rect 261076 634732 288900 634760
rect 261076 634720 261082 634732
rect 288894 634720 288900 634732
rect 288952 634720 288958 634772
rect 289078 634720 289084 634772
rect 289136 634760 289142 634772
rect 316586 634760 316592 634772
rect 289136 634732 316592 634760
rect 289136 634720 289142 634732
rect 316586 634720 316592 634732
rect 316644 634720 316650 634772
rect 317046 634720 317052 634772
rect 317104 634760 317110 634772
rect 344922 634760 344928 634772
rect 317104 634732 344928 634760
rect 317104 634720 317110 634732
rect 344922 634720 344928 634732
rect 344980 634720 344986 634772
rect 345658 634720 345664 634772
rect 345716 634760 345722 634772
rect 372614 634760 372620 634772
rect 345716 634732 372620 634760
rect 345716 634720 345722 634732
rect 372614 634720 372620 634732
rect 372672 634720 372678 634772
rect 373074 634720 373080 634772
rect 373132 634760 373138 634772
rect 400950 634760 400956 634772
rect 373132 634732 400956 634760
rect 373132 634720 373138 634732
rect 400950 634720 400956 634732
rect 401008 634720 401014 634772
rect 401042 634720 401048 634772
rect 401100 634760 401106 634772
rect 428918 634760 428924 634772
rect 401100 634732 428924 634760
rect 401100 634720 401106 634732
rect 428918 634720 428924 634732
rect 428976 634720 428982 634772
rect 429102 634720 429108 634772
rect 429160 634760 429166 634772
rect 456794 634760 456800 634772
rect 429160 634732 456800 634760
rect 429160 634720 429166 634732
rect 456794 634720 456800 634732
rect 456852 634720 456858 634772
rect 457070 634720 457076 634772
rect 457128 634760 457134 634772
rect 484946 634760 484952 634772
rect 457128 634732 484952 634760
rect 457128 634720 457134 634732
rect 484946 634720 484952 634732
rect 485004 634720 485010 634772
rect 485038 634720 485044 634772
rect 485096 634760 485102 634772
rect 512914 634760 512920 634772
rect 485096 634732 512920 634760
rect 485096 634720 485102 634732
rect 512914 634720 512920 634732
rect 512972 634720 512978 634772
rect 513098 634720 513104 634772
rect 513156 634760 513162 634772
rect 540606 634760 540612 634772
rect 513156 634732 540612 634760
rect 513156 634720 513162 634732
rect 540606 634720 540612 634732
rect 540664 634720 540670 634772
rect 541066 634720 541072 634772
rect 541124 634760 541130 634772
rect 568942 634760 568948 634772
rect 541124 634732 568948 634760
rect 541124 634720 541130 634732
rect 568942 634720 568948 634732
rect 569000 634720 569006 634772
rect 26602 634652 26608 634704
rect 26660 634692 26666 634704
rect 38010 634692 38016 634704
rect 26660 634664 38016 634692
rect 26660 634652 26666 634664
rect 38010 634652 38016 634664
rect 38068 634652 38074 634704
rect 54938 634652 54944 634704
rect 54996 634692 55002 634704
rect 71774 634692 71780 634704
rect 54996 634664 71780 634692
rect 54996 634652 55002 634664
rect 71774 634652 71780 634664
rect 71832 634652 71838 634704
rect 82630 634652 82636 634704
rect 82688 634692 82694 634704
rect 99374 634692 99380 634704
rect 82688 634664 99380 634692
rect 82688 634652 82694 634664
rect 99374 634652 99380 634664
rect 99432 634652 99438 634704
rect 128630 634652 128636 634704
rect 128688 634692 128694 634704
rect 149790 634692 149796 634704
rect 128688 634664 149796 634692
rect 128688 634652 128694 634664
rect 149790 634652 149796 634664
rect 149848 634652 149854 634704
rect 166626 634652 166632 634704
rect 166684 634692 166690 634704
rect 183554 634692 183560 634704
rect 166684 634664 183560 634692
rect 166684 634652 166690 634664
rect 183554 634652 183560 634664
rect 183612 634652 183618 634704
rect 194594 634652 194600 634704
rect 194652 634692 194658 634704
rect 211154 634692 211160 634704
rect 194652 634664 211160 634692
rect 194652 634652 194658 634664
rect 211154 634652 211160 634664
rect 211212 634652 211218 634704
rect 222930 634652 222936 634704
rect 222988 634692 222994 634704
rect 233970 634692 233976 634704
rect 222988 634664 233976 634692
rect 222988 634652 222994 634664
rect 233970 634652 233976 634664
rect 234028 634652 234034 634704
rect 250622 634652 250628 634704
rect 250680 634692 250686 634704
rect 267734 634692 267740 634704
rect 250680 634664 267740 634692
rect 250680 634652 250686 634664
rect 267734 634652 267740 634664
rect 267792 634652 267798 634704
rect 278590 634652 278596 634704
rect 278648 634692 278654 634704
rect 295334 634692 295340 634704
rect 278648 634664 295340 634692
rect 278648 634652 278654 634664
rect 295334 634652 295340 634664
rect 295392 634652 295398 634704
rect 306926 634652 306932 634704
rect 306984 634692 306990 634704
rect 318058 634692 318064 634704
rect 306984 634664 318064 634692
rect 306984 634652 306990 634664
rect 318058 634652 318064 634664
rect 318116 634652 318122 634704
rect 324314 634652 324320 634704
rect 324372 634692 324378 634704
rect 345750 634692 345756 634704
rect 324372 634664 345756 634692
rect 324372 634652 324378 634664
rect 345750 634652 345756 634664
rect 345808 634652 345814 634704
rect 362862 634652 362868 634704
rect 362920 634692 362926 634704
rect 379514 634692 379520 634704
rect 362920 634664 379520 634692
rect 362920 634652 362926 634664
rect 379514 634652 379520 634664
rect 379572 634652 379578 634704
rect 390646 634652 390652 634704
rect 390704 634692 390710 634704
rect 407114 634692 407120 634704
rect 390704 634664 407120 634692
rect 390704 634652 390710 634664
rect 407114 634652 407120 634664
rect 407172 634652 407178 634704
rect 418614 634652 418620 634704
rect 418672 634692 418678 634704
rect 429838 634692 429844 634704
rect 418672 634664 429844 634692
rect 418672 634652 418678 634664
rect 429838 634652 429844 634664
rect 429896 634652 429902 634704
rect 446950 634652 446956 634704
rect 447008 634692 447014 634704
rect 463694 634692 463700 634704
rect 447008 634664 463700 634692
rect 447008 634652 447014 634664
rect 463694 634652 463700 634664
rect 463752 634652 463758 634704
rect 474642 634652 474648 634704
rect 474700 634692 474706 634704
rect 491294 634692 491300 634704
rect 474700 634664 491300 634692
rect 474700 634652 474706 634664
rect 491294 634652 491300 634664
rect 491352 634652 491358 634704
rect 520642 634652 520648 634704
rect 520700 634692 520706 634704
rect 541618 634692 541624 634704
rect 520700 634664 541624 634692
rect 520700 634652 520706 634664
rect 541618 634652 541624 634664
rect 541676 634652 541682 634704
rect 138934 634584 138940 634636
rect 138992 634624 138998 634636
rect 155954 634624 155960 634636
rect 138992 634596 155960 634624
rect 138992 634584 138998 634596
rect 155954 634584 155960 634596
rect 156012 634584 156018 634636
rect 334618 634584 334624 634636
rect 334676 634624 334682 634636
rect 351914 634624 351920 634636
rect 334676 634596 351920 634624
rect 334676 634584 334682 634596
rect 351914 634584 351920 634596
rect 351972 634584 351978 634636
rect 530946 634584 530952 634636
rect 531004 634624 531010 634636
rect 547966 634624 547972 634636
rect 531004 634596 547972 634624
rect 531004 634584 531010 634596
rect 547966 634584 547972 634596
rect 548024 634584 548030 634636
rect 558638 634040 558644 634092
rect 558696 634080 558702 634092
rect 568942 634080 568948 634092
rect 558696 634052 568948 634080
rect 558696 634040 558702 634052
rect 568942 634040 568948 634052
rect 569000 634040 569006 634092
rect 548334 632680 548340 632732
rect 548392 632720 548398 632732
rect 569034 632720 569040 632732
rect 548392 632692 569040 632720
rect 548392 632680 548398 632692
rect 569034 632680 569040 632692
rect 569092 632680 569098 632732
rect 100018 632204 100024 632256
rect 100076 632244 100082 632256
rect 121086 632244 121092 632256
rect 100076 632216 121092 632244
rect 100076 632204 100082 632216
rect 121086 632204 121092 632216
rect 121144 632204 121150 632256
rect 184014 632204 184020 632256
rect 184072 632244 184078 632256
rect 204898 632244 204904 632256
rect 184072 632216 204904 632244
rect 184072 632204 184078 632216
rect 204898 632204 204904 632216
rect 204956 632204 204962 632256
rect 268010 632204 268016 632256
rect 268068 632244 268074 632256
rect 289078 632244 289084 632256
rect 268068 632216 289084 632244
rect 268068 632204 268074 632216
rect 289078 632204 289084 632216
rect 289136 632204 289142 632256
rect 380342 632204 380348 632256
rect 380400 632244 380406 632256
rect 401134 632244 401140 632256
rect 380400 632216 401140 632244
rect 380400 632204 380406 632216
rect 401134 632204 401140 632216
rect 401192 632204 401198 632256
rect 464338 632204 464344 632256
rect 464396 632244 464402 632256
rect 485038 632244 485044 632256
rect 464396 632216 485044 632244
rect 464396 632204 464402 632216
rect 485038 632204 485044 632216
rect 485096 632204 485102 632256
rect 37090 632136 37096 632188
rect 37148 632176 37154 632188
rect 54294 632176 54300 632188
rect 37148 632148 54300 632176
rect 37148 632136 37154 632148
rect 54294 632136 54300 632148
rect 54352 632136 54358 632188
rect 65886 632136 65892 632188
rect 65944 632176 65950 632188
rect 81986 632176 81992 632188
rect 65944 632148 81992 632176
rect 65944 632136 65950 632148
rect 81986 632136 81992 632148
rect 82044 632136 82050 632188
rect 92842 632136 92848 632188
rect 92900 632176 92906 632188
rect 110322 632176 110328 632188
rect 92900 632148 110328 632176
rect 92900 632136 92906 632148
rect 110322 632136 110328 632148
rect 110380 632136 110386 632188
rect 176838 632136 176844 632188
rect 176896 632176 176902 632188
rect 194318 632176 194324 632188
rect 176896 632148 194324 632176
rect 176896 632136 176902 632148
rect 194318 632136 194324 632148
rect 194376 632136 194382 632188
rect 261478 632136 261484 632188
rect 261536 632176 261542 632188
rect 278314 632176 278320 632188
rect 261536 632148 278320 632176
rect 261536 632136 261542 632148
rect 278314 632136 278320 632148
rect 278372 632136 278378 632188
rect 317138 632136 317144 632188
rect 317196 632176 317202 632188
rect 334342 632176 334348 632188
rect 317196 632148 334348 632176
rect 317196 632136 317202 632148
rect 334342 632136 334348 632148
rect 334400 632136 334406 632188
rect 372982 632136 372988 632188
rect 373040 632176 373046 632188
rect 390002 632176 390008 632188
rect 373040 632148 390008 632176
rect 373040 632136 373046 632148
rect 390002 632136 390008 632148
rect 390060 632136 390066 632188
rect 457438 632136 457444 632188
rect 457496 632176 457502 632188
rect 473998 632176 474004 632188
rect 457496 632148 474004 632176
rect 457496 632136 457502 632148
rect 473998 632136 474004 632148
rect 474056 632136 474062 632188
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4798 632108 4804 632120
rect 2832 632080 4804 632108
rect 2832 632068 2838 632080
rect 4798 632068 4804 632080
rect 4856 632068 4862 632120
rect 15286 632068 15292 632120
rect 15344 632108 15350 632120
rect 26326 632108 26332 632120
rect 15344 632080 26332 632108
rect 15344 632068 15350 632080
rect 26326 632068 26332 632080
rect 26384 632068 26390 632120
rect 39298 632068 39304 632120
rect 39356 632108 39362 632120
rect 64598 632108 64604 632120
rect 39356 632080 64604 632108
rect 39356 632068 39362 632080
rect 64598 632068 64604 632080
rect 64656 632068 64662 632120
rect 72326 632068 72332 632120
rect 72384 632108 72390 632120
rect 93118 632108 93124 632120
rect 72384 632080 93124 632108
rect 72384 632068 72390 632080
rect 93118 632068 93124 632080
rect 93176 632068 93182 632120
rect 120994 632068 121000 632120
rect 121052 632108 121058 632120
rect 138290 632108 138296 632120
rect 121052 632080 138296 632108
rect 121052 632068 121058 632080
rect 138290 632068 138296 632080
rect 138348 632068 138354 632120
rect 156322 632068 156328 632120
rect 156380 632108 156386 632120
rect 177298 632108 177304 632120
rect 156380 632080 177304 632108
rect 156380 632068 156386 632080
rect 177298 632068 177304 632080
rect 177356 632068 177362 632120
rect 204806 632068 204812 632120
rect 204864 632108 204870 632120
rect 222194 632108 222200 632120
rect 204864 632080 222200 632108
rect 204864 632068 204870 632080
rect 222194 632068 222200 632080
rect 222252 632068 222258 632120
rect 232958 632068 232964 632120
rect 233016 632108 233022 632120
rect 250346 632108 250352 632120
rect 233016 632080 250352 632108
rect 233016 632068 233022 632080
rect 250346 632068 250352 632080
rect 250404 632068 250410 632120
rect 288894 632068 288900 632120
rect 288952 632108 288958 632120
rect 306006 632108 306012 632120
rect 288952 632080 306012 632108
rect 288952 632068 288958 632080
rect 306006 632068 306012 632080
rect 306064 632068 306070 632120
rect 317046 632068 317052 632120
rect 317104 632108 317110 632120
rect 344646 632108 344652 632120
rect 317104 632080 344652 632108
rect 317104 632068 317110 632080
rect 344646 632068 344652 632080
rect 344704 632068 344710 632120
rect 352006 632068 352012 632120
rect 352064 632108 352070 632120
rect 373258 632108 373264 632120
rect 352064 632080 373264 632108
rect 352064 632068 352070 632080
rect 373258 632068 373264 632080
rect 373316 632068 373322 632120
rect 401042 632068 401048 632120
rect 401100 632108 401106 632120
rect 418338 632108 418344 632120
rect 401100 632080 418344 632108
rect 401100 632068 401106 632080
rect 418338 632068 418344 632080
rect 418396 632068 418402 632120
rect 429838 632068 429844 632120
rect 429896 632108 429902 632120
rect 456610 632108 456616 632120
rect 429896 632080 456616 632108
rect 429896 632068 429902 632080
rect 456610 632068 456616 632080
rect 456668 632068 456674 632120
rect 484854 632068 484860 632120
rect 484912 632108 484918 632120
rect 502334 632108 502340 632120
rect 484912 632080 502340 632108
rect 484912 632068 484918 632080
rect 502334 632068 502340 632080
rect 502392 632068 502398 632120
rect 514846 632068 514852 632120
rect 514904 632108 514910 632120
rect 530302 632108 530308 632120
rect 514904 632080 530308 632108
rect 514904 632068 514910 632080
rect 530302 632068 530308 632080
rect 530360 632068 530366 632120
rect 36722 630232 36728 630284
rect 36780 630272 36786 630284
rect 37090 630272 37096 630284
rect 36780 630244 37096 630272
rect 36780 630232 36786 630244
rect 37090 630232 37096 630244
rect 37148 630232 37154 630284
rect 120718 630232 120724 630284
rect 120776 630272 120782 630284
rect 120994 630272 121000 630284
rect 120776 630244 121000 630272
rect 120776 630232 120782 630244
rect 120994 630232 121000 630244
rect 121052 630232 121058 630284
rect 204714 630232 204720 630284
rect 204772 630272 204778 630284
rect 204990 630272 204996 630284
rect 204772 630244 204996 630272
rect 204772 630232 204778 630244
rect 204990 630232 204996 630244
rect 205048 630232 205054 630284
rect 120810 630164 120816 630216
rect 120868 630204 120874 630216
rect 121086 630204 121092 630216
rect 120868 630176 121092 630204
rect 120868 630164 120874 630176
rect 121086 630164 121092 630176
rect 121144 630164 121150 630216
rect 400858 630164 400864 630216
rect 400916 630204 400922 630216
rect 401134 630204 401140 630216
rect 400916 630176 401140 630204
rect 400916 630164 400922 630176
rect 401134 630164 401140 630176
rect 401192 630164 401198 630216
rect 316770 628668 316776 628720
rect 316828 628708 316834 628720
rect 317138 628708 317144 628720
rect 316828 628680 317144 628708
rect 316828 628668 316834 628680
rect 317138 628668 317144 628680
rect 317196 628668 317202 628720
rect 232774 628600 232780 628652
rect 232832 628640 232838 628652
rect 232958 628640 232964 628652
rect 232832 628612 232964 628640
rect 232832 628600 232838 628612
rect 232958 628600 232964 628612
rect 233016 628600 233022 628652
rect 316862 628600 316868 628652
rect 316920 628640 316926 628652
rect 317046 628640 317052 628652
rect 316920 628612 317052 628640
rect 316920 628600 316926 628612
rect 317046 628600 317052 628612
rect 317104 628600 317110 628652
rect 372798 628600 372804 628652
rect 372856 628640 372862 628652
rect 372982 628640 372988 628652
rect 372856 628612 372988 628640
rect 372856 628600 372862 628612
rect 372982 628600 372988 628612
rect 373040 628600 373046 628652
rect 400766 628600 400772 628652
rect 400824 628640 400830 628652
rect 401042 628640 401048 628652
rect 400824 628612 401048 628640
rect 400824 628600 400830 628612
rect 401042 628600 401048 628612
rect 401100 628600 401106 628652
rect 512730 628600 512736 628652
rect 512788 628640 512794 628652
rect 514846 628640 514852 628652
rect 512788 628612 514852 628640
rect 512788 628600 512794 628612
rect 514846 628600 514852 628612
rect 514904 628600 514910 628652
rect 568758 625812 568764 625864
rect 568816 625852 568822 625864
rect 568942 625852 568948 625864
rect 568816 625824 568948 625852
rect 568816 625812 568822 625824
rect 568942 625812 568948 625824
rect 569000 625812 569006 625864
rect 92750 613980 92756 614032
rect 92808 614020 92814 614032
rect 92934 614020 92940 614032
rect 92808 613992 92940 614020
rect 92808 613980 92814 613992
rect 92934 613980 92940 613992
rect 92992 613980 92998 614032
rect 93118 613368 93124 613420
rect 93176 613408 93182 613420
rect 99742 613408 99748 613420
rect 93176 613380 99748 613408
rect 93176 613368 93182 613380
rect 99742 613368 99748 613380
rect 99800 613368 99806 613420
rect 120810 613368 120816 613420
rect 120868 613408 120874 613420
rect 127710 613408 127716 613420
rect 120868 613380 127716 613408
rect 120868 613368 120874 613380
rect 127710 613368 127716 613380
rect 127768 613368 127774 613420
rect 177298 613368 177304 613420
rect 177356 613408 177362 613420
rect 183646 613408 183652 613420
rect 177356 613380 183652 613408
rect 177356 613368 177362 613380
rect 183646 613368 183652 613380
rect 183704 613368 183710 613420
rect 373258 613368 373264 613420
rect 373316 613408 373322 613420
rect 379698 613408 379704 613420
rect 373316 613380 379704 613408
rect 373316 613368 373322 613380
rect 379698 613368 379704 613380
rect 379756 613368 379762 613420
rect 400858 613368 400864 613420
rect 400916 613408 400922 613420
rect 407758 613408 407764 613420
rect 400916 613380 407764 613408
rect 400916 613368 400922 613380
rect 407758 613368 407764 613380
rect 407816 613368 407822 613420
rect 64874 613096 64880 613148
rect 64932 613136 64938 613148
rect 65886 613136 65892 613148
rect 64932 613108 65892 613136
rect 64932 613096 64938 613108
rect 65886 613096 65892 613108
rect 65944 613096 65950 613148
rect 204898 613096 204904 613148
rect 204956 613136 204962 613148
rect 211706 613136 211712 613148
rect 204956 613108 211712 613136
rect 204956 613096 204962 613108
rect 211706 613096 211712 613108
rect 211764 613096 211770 613148
rect 485038 613096 485044 613148
rect 485096 613136 485102 613148
rect 491662 613136 491668 613148
rect 485096 613108 491668 613136
rect 485096 613096 485102 613108
rect 491662 613096 491668 613108
rect 491720 613096 491726 613148
rect 289078 612756 289084 612808
rect 289136 612796 289142 612808
rect 295702 612796 295708 612808
rect 289136 612768 295708 612796
rect 289136 612756 289142 612768
rect 295702 612756 295708 612768
rect 295760 612756 295766 612808
rect 42702 611260 42708 611312
rect 42760 611300 42766 611312
rect 95234 611300 95240 611312
rect 42760 611272 95240 611300
rect 42760 611260 42766 611272
rect 95234 611260 95240 611272
rect 95292 611260 95298 611312
rect 97902 611260 97908 611312
rect 97960 611300 97966 611312
rect 150434 611300 150440 611312
rect 97960 611272 150440 611300
rect 97960 611260 97966 611272
rect 150434 611260 150440 611272
rect 150492 611260 150498 611312
rect 154482 611260 154488 611312
rect 154540 611300 154546 611312
rect 207014 611300 207020 611312
rect 154540 611272 207020 611300
rect 154540 611260 154546 611272
rect 207014 611260 207020 611272
rect 207072 611260 207078 611312
rect 209682 611260 209688 611312
rect 209740 611300 209746 611312
rect 262214 611300 262220 611312
rect 209740 611272 262220 611300
rect 209740 611260 209746 611272
rect 262214 611260 262220 611272
rect 262272 611260 262278 611312
rect 266262 611260 266268 611312
rect 266320 611300 266326 611312
rect 318794 611300 318800 611312
rect 266320 611272 318800 611300
rect 266320 611260 266326 611272
rect 318794 611260 318800 611272
rect 318852 611260 318858 611312
rect 322842 611260 322848 611312
rect 322900 611300 322906 611312
rect 375374 611300 375380 611312
rect 322900 611272 375380 611300
rect 322900 611260 322906 611272
rect 375374 611260 375380 611272
rect 375432 611260 375438 611312
rect 378042 611260 378048 611312
rect 378100 611300 378106 611312
rect 430574 611300 430580 611312
rect 378100 611272 430580 611300
rect 378100 611260 378106 611272
rect 430574 611260 430580 611272
rect 430632 611260 430638 611312
rect 434622 611260 434628 611312
rect 434680 611300 434686 611312
rect 487154 611300 487160 611312
rect 434680 611272 487160 611300
rect 434680 611260 434686 611272
rect 487154 611260 487160 611272
rect 487212 611260 487218 611312
rect 489822 611260 489828 611312
rect 489880 611300 489886 611312
rect 542354 611300 542360 611312
rect 489880 611272 542360 611300
rect 489880 611260 489886 611272
rect 542354 611260 542360 611272
rect 542412 611260 542418 611312
rect 176746 610784 176752 610836
rect 176804 610824 176810 610836
rect 176930 610824 176936 610836
rect 176804 610796 176936 610824
rect 176804 610784 176810 610796
rect 176930 610784 176936 610796
rect 176988 610784 176994 610836
rect 288802 610784 288808 610836
rect 288860 610824 288866 610836
rect 288986 610824 288992 610836
rect 288860 610796 288992 610824
rect 288860 610784 288866 610796
rect 288986 610784 288992 610796
rect 289044 610784 289050 610836
rect 484762 610784 484768 610836
rect 484820 610824 484826 610836
rect 484946 610824 484952 610836
rect 484820 610796 484952 610824
rect 484820 610784 484826 610796
rect 484946 610784 484952 610796
rect 485004 610784 485010 610836
rect 547874 610648 547880 610700
rect 547932 610688 547938 610700
rect 548150 610688 548156 610700
rect 547932 610660 548156 610688
rect 547932 610648 547938 610660
rect 548150 610648 548156 610660
rect 548208 610648 548214 610700
rect 15286 610104 15292 610156
rect 15344 610104 15350 610156
rect 15304 609940 15332 610104
rect 15930 609940 15936 609952
rect 15304 609912 15936 609940
rect 15930 609900 15936 609912
rect 15988 609900 15994 609952
rect 15378 608540 15384 608592
rect 15436 608580 15442 608592
rect 43990 608580 43996 608592
rect 15436 608552 43996 608580
rect 15436 608540 15442 608552
rect 43990 608540 43996 608552
rect 44048 608540 44054 608592
rect 138290 608540 138296 608592
rect 138348 608580 138354 608592
rect 176930 608580 176936 608592
rect 138348 608552 176936 608580
rect 138348 608540 138354 608552
rect 176930 608540 176936 608552
rect 176988 608540 176994 608592
rect 194318 608540 194324 608592
rect 194376 608580 194382 608592
rect 232866 608580 232872 608592
rect 194376 608552 232872 608580
rect 194376 608540 194382 608552
rect 232866 608540 232872 608552
rect 232924 608540 232930 608592
rect 238846 608540 238852 608592
rect 238904 608580 238910 608592
rect 238904 608552 248414 608580
rect 238904 608540 238910 608552
rect 26326 608472 26332 608524
rect 26384 608512 26390 608524
rect 39298 608512 39304 608524
rect 26384 608484 39304 608512
rect 26384 608472 26390 608484
rect 39298 608472 39304 608484
rect 39356 608472 39362 608524
rect 42886 608472 42892 608524
rect 42944 608512 42950 608524
rect 71774 608512 71780 608524
rect 42944 608484 71780 608512
rect 42944 608472 42950 608484
rect 71774 608472 71780 608484
rect 71832 608472 71838 608524
rect 110322 608472 110328 608524
rect 110380 608512 110386 608524
rect 148778 608512 148784 608524
rect 110380 608484 148784 608512
rect 110380 608472 110386 608484
rect 148778 608472 148784 608484
rect 148836 608472 148842 608524
rect 166626 608472 166632 608524
rect 166684 608512 166690 608524
rect 204990 608512 204996 608524
rect 166684 608484 204996 608512
rect 166684 608472 166690 608484
rect 204990 608472 204996 608484
rect 205048 608472 205054 608524
rect 211246 608472 211252 608524
rect 211304 608512 211310 608524
rect 240042 608512 240048 608524
rect 211304 608484 240048 608512
rect 211304 608472 211310 608484
rect 240042 608472 240048 608484
rect 240100 608472 240106 608524
rect 248386 608512 248414 608552
rect 295426 608540 295432 608592
rect 295484 608580 295490 608592
rect 324038 608580 324044 608592
rect 295484 608552 324044 608580
rect 295484 608540 295490 608552
rect 324038 608540 324044 608552
rect 324096 608540 324102 608592
rect 334342 608540 334348 608592
rect 334400 608580 334406 608592
rect 372890 608580 372896 608592
rect 334400 608552 372896 608580
rect 334400 608540 334406 608552
rect 372890 608540 372896 608552
rect 372948 608540 372954 608592
rect 390462 608540 390468 608592
rect 390520 608580 390526 608592
rect 428734 608580 428740 608592
rect 390520 608552 428740 608580
rect 390520 608540 390526 608552
rect 428734 608540 428740 608552
rect 428792 608540 428798 608592
rect 434806 608540 434812 608592
rect 434864 608580 434870 608592
rect 434864 608552 441614 608580
rect 434864 608540 434870 608552
rect 268010 608512 268016 608524
rect 248386 608484 268016 608512
rect 268010 608472 268016 608484
rect 268068 608472 268074 608524
rect 278314 608472 278320 608524
rect 278372 608512 278378 608524
rect 316954 608512 316960 608524
rect 278372 608484 316960 608512
rect 278372 608472 278378 608484
rect 316954 608472 316960 608484
rect 317012 608472 317018 608524
rect 323026 608472 323032 608524
rect 323084 608512 323090 608524
rect 352006 608512 352012 608524
rect 323084 608484 352012 608512
rect 323084 608472 323090 608484
rect 352006 608472 352012 608484
rect 352064 608472 352070 608524
rect 362310 608472 362316 608524
rect 362368 608512 362374 608524
rect 400950 608512 400956 608524
rect 362368 608484 400956 608512
rect 362368 608472 362374 608484
rect 400950 608472 400956 608484
rect 401008 608472 401014 608524
rect 407206 608472 407212 608524
rect 407264 608512 407270 608524
rect 436002 608512 436008 608524
rect 407264 608484 436008 608512
rect 407264 608472 407270 608484
rect 436002 608472 436008 608484
rect 436060 608472 436066 608524
rect 441586 608512 441614 608552
rect 491386 608540 491392 608592
rect 491444 608580 491450 608592
rect 519998 608580 520004 608592
rect 491444 608552 520004 608580
rect 491444 608540 491450 608552
rect 519998 608540 520004 608552
rect 520056 608540 520062 608592
rect 530302 608540 530308 608592
rect 530360 608580 530366 608592
rect 568850 608580 568856 608592
rect 530360 608552 568856 608580
rect 530360 608540 530366 608552
rect 568850 608540 568856 608552
rect 568908 608540 568914 608592
rect 463694 608512 463700 608524
rect 441586 608484 463700 608512
rect 463694 608472 463700 608484
rect 463752 608472 463758 608524
rect 474642 608472 474648 608524
rect 474700 608512 474706 608524
rect 512822 608512 512828 608524
rect 474700 608484 512828 608512
rect 474700 608472 474706 608484
rect 512822 608472 512828 608484
rect 512880 608472 512886 608524
rect 548150 608472 548156 608524
rect 548208 608512 548214 608524
rect 557994 608512 558000 608524
rect 548208 608484 558000 608512
rect 548208 608472 548214 608484
rect 557994 608472 558000 608484
rect 558052 608472 558058 608524
rect 82630 608404 82636 608456
rect 82688 608444 82694 608456
rect 120902 608444 120908 608456
rect 82688 608416 120908 608444
rect 82688 608404 82694 608416
rect 120902 608404 120908 608416
rect 120960 608404 120966 608456
rect 127066 608404 127072 608456
rect 127124 608444 127130 608456
rect 156046 608444 156052 608456
rect 127124 608416 156052 608444
rect 127124 608404 127130 608416
rect 156046 608404 156052 608416
rect 156104 608404 156110 608456
rect 250346 608404 250352 608456
rect 250404 608444 250410 608456
rect 288986 608444 288992 608456
rect 250404 608416 288992 608444
rect 250404 608404 250410 608416
rect 288986 608404 288992 608416
rect 289044 608404 289050 608456
rect 306282 608404 306288 608456
rect 306340 608444 306346 608456
rect 316862 608444 316868 608456
rect 306340 608416 316868 608444
rect 306340 608404 306346 608416
rect 316862 608404 316868 608416
rect 316920 608404 316926 608456
rect 418338 608404 418344 608456
rect 418396 608444 418402 608456
rect 429838 608444 429844 608456
rect 418396 608416 429844 608444
rect 418396 608404 418402 608416
rect 429838 608404 429844 608416
rect 429896 608404 429902 608456
rect 446306 608404 446312 608456
rect 446364 608444 446370 608456
rect 484946 608444 484952 608456
rect 446364 608416 484952 608444
rect 446364 608404 446370 608416
rect 484946 608404 484952 608416
rect 485004 608404 485010 608456
rect 502334 608404 502340 608456
rect 502392 608444 502398 608456
rect 540790 608444 540796 608456
rect 502392 608416 540796 608444
rect 502392 608404 502398 608416
rect 540790 608404 540796 608416
rect 540848 608404 540854 608456
rect 54294 608336 54300 608388
rect 54352 608376 54358 608388
rect 92934 608376 92940 608388
rect 54352 608348 92940 608376
rect 54352 608336 54358 608348
rect 92934 608336 92940 608348
rect 92992 608336 92998 608388
rect 518986 608336 518992 608388
rect 519044 608376 519050 608388
rect 547874 608376 547880 608388
rect 519044 608348 547880 608376
rect 519044 608336 519050 608348
rect 547874 608336 547880 608348
rect 547932 608336 547938 608388
rect 26602 606432 26608 606484
rect 26660 606472 26666 606484
rect 36814 606472 36820 606484
rect 26660 606444 36820 606472
rect 26660 606432 26666 606444
rect 36814 606432 36820 606444
rect 36872 606432 36878 606484
rect 15378 605956 15384 606008
rect 15436 605996 15442 606008
rect 54294 605996 54300 606008
rect 15436 605968 54300 605996
rect 15436 605956 15442 605968
rect 54294 605956 54300 605968
rect 54352 605956 54358 606008
rect 2774 605888 2780 605940
rect 2832 605928 2838 605940
rect 4890 605928 4896 605940
rect 2832 605900 4896 605928
rect 2832 605888 2838 605900
rect 4890 605888 4896 605900
rect 4948 605888 4954 605940
rect 71866 605888 71872 605940
rect 71924 605928 71930 605940
rect 110598 605928 110604 605940
rect 71924 605900 110604 605928
rect 71924 605888 71930 605900
rect 110598 605888 110604 605900
rect 110656 605888 110662 605940
rect 149882 605888 149888 605940
rect 149940 605928 149946 605940
rect 156322 605928 156328 605940
rect 149940 605900 156328 605928
rect 149940 605888 149946 605900
rect 156322 605888 156328 605900
rect 156380 605888 156386 605940
rect 211246 605888 211252 605940
rect 211304 605928 211310 605940
rect 250622 605928 250628 605940
rect 211304 605900 250628 605928
rect 211304 605888 211310 605900
rect 250622 605888 250628 605900
rect 250680 605888 250686 605940
rect 267826 605888 267832 605940
rect 267884 605928 267890 605940
rect 306374 605928 306380 605940
rect 267884 605900 306380 605928
rect 267884 605888 267890 605900
rect 306374 605888 306380 605900
rect 306432 605888 306438 605940
rect 318058 605888 318064 605940
rect 318116 605928 318122 605940
rect 324314 605928 324320 605940
rect 318116 605900 324320 605928
rect 318116 605888 318122 605900
rect 324314 605888 324320 605900
rect 324372 605888 324378 605940
rect 345750 605888 345756 605940
rect 345808 605928 345814 605940
rect 362310 605928 362316 605940
rect 345808 605900 362316 605928
rect 345808 605888 345814 605900
rect 362310 605888 362316 605900
rect 362368 605888 362374 605940
rect 407206 605888 407212 605940
rect 407264 605928 407270 605940
rect 446306 605928 446312 605940
rect 407264 605900 446312 605928
rect 407264 605888 407270 605900
rect 446306 605888 446312 605900
rect 446364 605888 446370 605940
rect 463786 605888 463792 605940
rect 463844 605928 463850 605940
rect 502610 605928 502616 605940
rect 463844 605900 502616 605928
rect 463844 605888 463850 605900
rect 502610 605888 502616 605900
rect 502668 605888 502674 605940
rect 514018 605888 514024 605940
rect 514076 605928 514082 605940
rect 520274 605928 520280 605940
rect 514076 605900 520280 605928
rect 514076 605888 514082 605900
rect 520274 605888 520280 605900
rect 520332 605888 520338 605940
rect 38102 605820 38108 605872
rect 38160 605860 38166 605872
rect 44174 605860 44180 605872
rect 38160 605832 44180 605860
rect 38160 605820 38166 605832
rect 44174 605820 44180 605832
rect 44232 605820 44238 605872
rect 65886 605820 65892 605872
rect 65944 605860 65950 605872
rect 82630 605860 82636 605872
rect 65944 605832 82636 605860
rect 65944 605820 65950 605832
rect 82630 605820 82636 605832
rect 82688 605820 82694 605872
rect 99374 605820 99380 605872
rect 99432 605860 99438 605872
rect 138290 605860 138296 605872
rect 99432 605832 138296 605860
rect 99432 605820 99438 605832
rect 138290 605820 138296 605832
rect 138348 605820 138354 605872
rect 149790 605820 149796 605872
rect 149848 605860 149854 605872
rect 166626 605860 166632 605872
rect 149848 605832 166632 605860
rect 149848 605820 149854 605832
rect 166626 605820 166632 605832
rect 166684 605820 166690 605872
rect 183554 605820 183560 605872
rect 183612 605860 183618 605872
rect 222378 605860 222384 605872
rect 183612 605832 222384 605860
rect 183612 605820 183618 605832
rect 222378 605820 222384 605832
rect 222436 605820 222442 605872
rect 234062 605820 234068 605872
rect 234120 605860 234126 605872
rect 240318 605860 240324 605872
rect 234120 605832 240324 605860
rect 234120 605820 234126 605832
rect 240318 605820 240324 605832
rect 240376 605820 240382 605872
rect 261478 605820 261484 605872
rect 261536 605860 261542 605872
rect 278590 605860 278596 605872
rect 261536 605832 278596 605860
rect 261536 605820 261542 605832
rect 278590 605820 278596 605832
rect 278648 605820 278654 605872
rect 295334 605820 295340 605872
rect 295392 605860 295398 605872
rect 334618 605860 334624 605872
rect 295392 605832 334624 605860
rect 295392 605820 295398 605832
rect 334618 605820 334624 605832
rect 334676 605820 334682 605872
rect 345658 605820 345664 605872
rect 345716 605860 345722 605872
rect 352006 605860 352012 605872
rect 345716 605832 352012 605860
rect 345716 605820 345722 605832
rect 352006 605820 352012 605832
rect 352064 605820 352070 605872
rect 379514 605820 379520 605872
rect 379572 605860 379578 605872
rect 418614 605860 418620 605872
rect 379572 605832 418620 605860
rect 379572 605820 379578 605832
rect 418614 605820 418620 605832
rect 418672 605820 418678 605872
rect 429930 605820 429936 605872
rect 429988 605860 429994 605872
rect 436094 605860 436100 605872
rect 429988 605832 436100 605860
rect 429988 605820 429994 605832
rect 436094 605820 436100 605832
rect 436152 605820 436158 605872
rect 457438 605820 457444 605872
rect 457496 605860 457502 605872
rect 474642 605860 474648 605872
rect 457496 605832 474648 605860
rect 457496 605820 457502 605832
rect 474642 605820 474648 605832
rect 474700 605820 474706 605872
rect 491294 605820 491300 605872
rect 491352 605860 491358 605872
rect 530302 605860 530308 605872
rect 491352 605832 530308 605860
rect 491352 605820 491358 605832
rect 530302 605820 530308 605832
rect 530360 605820 530366 605872
rect 541618 605820 541624 605872
rect 541676 605860 541682 605872
rect 558638 605860 558644 605872
rect 541676 605832 558644 605860
rect 541676 605820 541682 605832
rect 558638 605820 558644 605832
rect 558696 605820 558702 605872
rect 205082 603304 205088 603356
rect 205140 603304 205146 603356
rect 205100 603152 205128 603304
rect 345014 603236 345020 603288
rect 345072 603276 345078 603288
rect 345842 603276 345848 603288
rect 345072 603248 345848 603276
rect 345072 603236 345078 603248
rect 345842 603236 345848 603248
rect 345900 603236 345906 603288
rect 205082 603100 205088 603152
rect 205140 603100 205146 603152
rect 429102 603100 429108 603152
rect 429160 603140 429166 603152
rect 429838 603140 429844 603152
rect 429160 603112 429844 603140
rect 429160 603100 429166 603112
rect 429838 603100 429844 603112
rect 429896 603100 429902 603152
rect 37274 599700 37280 599752
rect 37332 599740 37338 599752
rect 38010 599740 38016 599752
rect 37332 599712 38016 599740
rect 37332 599700 37338 599712
rect 38010 599700 38016 599712
rect 38068 599700 38074 599752
rect 71774 599700 71780 599752
rect 71832 599740 71838 599752
rect 71958 599740 71964 599752
rect 71832 599712 71964 599740
rect 71832 599700 71838 599712
rect 71958 599700 71964 599712
rect 72016 599700 72022 599752
rect 211154 599700 211160 599752
rect 211212 599740 211218 599752
rect 211982 599740 211988 599752
rect 211212 599712 211988 599740
rect 211212 599700 211218 599712
rect 211982 599700 211988 599712
rect 212040 599700 212046 599752
rect 233234 599700 233240 599752
rect 233292 599740 233298 599752
rect 233970 599740 233976 599752
rect 233292 599712 233976 599740
rect 233292 599700 233298 599712
rect 233970 599700 233976 599712
rect 234028 599700 234034 599752
rect 267734 599700 267740 599752
rect 267792 599740 267798 599752
rect 267918 599740 267924 599752
rect 267792 599712 267924 599740
rect 267792 599700 267798 599712
rect 267918 599700 267924 599712
rect 267976 599700 267982 599752
rect 407114 599700 407120 599752
rect 407172 599740 407178 599752
rect 407942 599740 407948 599752
rect 407172 599712 407948 599740
rect 407172 599700 407178 599712
rect 407942 599700 407948 599712
rect 408000 599700 408006 599752
rect 463694 599700 463700 599752
rect 463752 599740 463758 599752
rect 464062 599740 464068 599752
rect 463752 599712 464068 599740
rect 463752 599700 463758 599712
rect 464062 599700 464068 599712
rect 464120 599700 464126 599752
rect 93118 585760 93124 585812
rect 93176 585800 93182 585812
rect 99466 585800 99472 585812
rect 93176 585772 99472 585800
rect 93176 585760 93182 585772
rect 99466 585760 99472 585772
rect 99524 585760 99530 585812
rect 177114 585760 177120 585812
rect 177172 585800 177178 585812
rect 183646 585800 183652 585812
rect 177172 585772 183652 585800
rect 177172 585760 177178 585772
rect 183646 585760 183652 585772
rect 183704 585760 183710 585812
rect 373166 585760 373172 585812
rect 373224 585800 373230 585812
rect 379606 585800 379612 585812
rect 373224 585772 379612 585800
rect 373224 585760 373230 585772
rect 379606 585760 379612 585772
rect 379664 585760 379670 585812
rect 289722 585148 289728 585200
rect 289780 585188 289786 585200
rect 295426 585188 295432 585200
rect 289780 585160 295432 585188
rect 289780 585148 289786 585160
rect 295426 585148 295432 585160
rect 295484 585148 295490 585200
rect 485130 585148 485136 585200
rect 485188 585188 485194 585200
rect 491386 585188 491392 585200
rect 485188 585160 491392 585188
rect 485188 585148 485194 585160
rect 491386 585148 491392 585160
rect 491444 585148 491450 585200
rect 15194 580932 15200 580984
rect 15252 580972 15258 580984
rect 36906 580972 36912 580984
rect 15252 580944 36912 580972
rect 15252 580932 15258 580944
rect 36906 580932 36912 580944
rect 36964 580932 36970 580984
rect 38010 580932 38016 580984
rect 38068 580972 38074 580984
rect 64874 580972 64880 580984
rect 38068 580944 64880 580972
rect 38068 580932 38074 580944
rect 64874 580932 64880 580944
rect 64932 580932 64938 580984
rect 65058 580932 65064 580984
rect 65116 580972 65122 580984
rect 92934 580972 92940 580984
rect 65116 580944 92940 580972
rect 65116 580932 65122 580944
rect 92934 580932 92940 580944
rect 92992 580932 92998 580984
rect 93026 580932 93032 580984
rect 93084 580972 93090 580984
rect 120902 580972 120908 580984
rect 93084 580944 120908 580972
rect 93084 580932 93090 580944
rect 120902 580932 120908 580944
rect 120960 580932 120966 580984
rect 121086 580932 121092 580984
rect 121144 580972 121150 580984
rect 148594 580972 148600 580984
rect 121144 580944 148600 580972
rect 121144 580932 121150 580944
rect 148594 580932 148600 580944
rect 148652 580932 148658 580984
rect 149698 580932 149704 580984
rect 149756 580972 149762 580984
rect 176930 580972 176936 580984
rect 149756 580944 176936 580972
rect 149756 580932 149762 580944
rect 176930 580932 176936 580944
rect 176988 580932 176994 580984
rect 177022 580932 177028 580984
rect 177080 580972 177086 580984
rect 204898 580972 204904 580984
rect 177080 580944 204904 580972
rect 177080 580932 177086 580944
rect 204898 580932 204904 580944
rect 204956 580932 204962 580984
rect 205174 580932 205180 580984
rect 205232 580972 205238 580984
rect 232590 580972 232596 580984
rect 205232 580944 232596 580972
rect 205232 580932 205238 580944
rect 232590 580932 232596 580944
rect 232648 580932 232654 580984
rect 233970 580932 233976 580984
rect 234028 580972 234034 580984
rect 260926 580972 260932 580984
rect 234028 580944 260932 580972
rect 234028 580932 234034 580944
rect 260926 580932 260932 580944
rect 260984 580932 260990 580984
rect 261018 580932 261024 580984
rect 261076 580972 261082 580984
rect 288894 580972 288900 580984
rect 261076 580944 288900 580972
rect 261076 580932 261082 580944
rect 288894 580932 288900 580944
rect 288952 580932 288958 580984
rect 289078 580932 289084 580984
rect 289136 580972 289142 580984
rect 316586 580972 316592 580984
rect 289136 580944 316592 580972
rect 289136 580932 289142 580944
rect 316586 580932 316592 580944
rect 316644 580932 316650 580984
rect 317046 580932 317052 580984
rect 317104 580972 317110 580984
rect 344922 580972 344928 580984
rect 317104 580944 344928 580972
rect 317104 580932 317110 580944
rect 344922 580932 344928 580944
rect 344980 580932 344986 580984
rect 345842 580932 345848 580984
rect 345900 580972 345906 580984
rect 372614 580972 372620 580984
rect 345900 580944 372620 580972
rect 345900 580932 345906 580944
rect 372614 580932 372620 580944
rect 372672 580932 372678 580984
rect 373074 580932 373080 580984
rect 373132 580972 373138 580984
rect 400950 580972 400956 580984
rect 373132 580944 400956 580972
rect 373132 580932 373138 580944
rect 400950 580932 400956 580944
rect 401008 580932 401014 580984
rect 401042 580932 401048 580984
rect 401100 580972 401106 580984
rect 428918 580972 428924 580984
rect 401100 580944 428924 580972
rect 401100 580932 401106 580944
rect 428918 580932 428924 580944
rect 428976 580932 428982 580984
rect 429838 580932 429844 580984
rect 429896 580972 429902 580984
rect 456794 580972 456800 580984
rect 429896 580944 456800 580972
rect 429896 580932 429902 580944
rect 456794 580932 456800 580944
rect 456852 580932 456858 580984
rect 457070 580932 457076 580984
rect 457128 580972 457134 580984
rect 484946 580972 484952 580984
rect 457128 580944 484952 580972
rect 457128 580932 457134 580944
rect 484946 580932 484952 580944
rect 485004 580932 485010 580984
rect 485038 580932 485044 580984
rect 485096 580972 485102 580984
rect 512914 580972 512920 580984
rect 485096 580944 512920 580972
rect 485096 580932 485102 580944
rect 512914 580932 512920 580944
rect 512972 580932 512978 580984
rect 513098 580932 513104 580984
rect 513156 580972 513162 580984
rect 540606 580972 540612 580984
rect 513156 580944 540612 580972
rect 513156 580932 513162 580944
rect 540606 580932 540612 580944
rect 540664 580932 540670 580984
rect 541066 580932 541072 580984
rect 541124 580972 541130 580984
rect 568942 580972 568948 580984
rect 541124 580944 568948 580972
rect 541124 580932 541130 580944
rect 568942 580932 568948 580944
rect 569000 580932 569006 580984
rect 26602 580864 26608 580916
rect 26660 580904 26666 580916
rect 38102 580904 38108 580916
rect 26660 580876 38108 580904
rect 26660 580864 26666 580876
rect 38102 580864 38108 580876
rect 38160 580864 38166 580916
rect 44634 580864 44640 580916
rect 44692 580904 44698 580916
rect 65886 580904 65892 580916
rect 44692 580876 65892 580904
rect 44692 580864 44698 580876
rect 65886 580864 65892 580876
rect 65944 580864 65950 580916
rect 82630 580864 82636 580916
rect 82688 580904 82694 580916
rect 93118 580904 93124 580916
rect 82688 580876 93124 580904
rect 82688 580864 82694 580876
rect 93118 580864 93124 580876
rect 93176 580864 93182 580916
rect 128630 580864 128636 580916
rect 128688 580904 128694 580916
rect 149790 580904 149796 580916
rect 128688 580876 149796 580904
rect 128688 580864 128694 580876
rect 149790 580864 149796 580876
rect 149848 580864 149854 580916
rect 166626 580864 166632 580916
rect 166684 580904 166690 580916
rect 177114 580904 177120 580916
rect 166684 580876 177120 580904
rect 166684 580864 166690 580876
rect 177114 580864 177120 580876
rect 177172 580864 177178 580916
rect 194594 580864 194600 580916
rect 194652 580904 194658 580916
rect 211154 580904 211160 580916
rect 194652 580876 211160 580904
rect 194652 580864 194658 580876
rect 211154 580864 211160 580876
rect 211212 580864 211218 580916
rect 222930 580864 222936 580916
rect 222988 580904 222994 580916
rect 234062 580904 234068 580916
rect 222988 580876 234068 580904
rect 222988 580864 222994 580876
rect 234062 580864 234068 580876
rect 234120 580864 234126 580916
rect 240318 580864 240324 580916
rect 240376 580904 240382 580916
rect 261478 580904 261484 580916
rect 240376 580876 261484 580904
rect 240376 580864 240382 580876
rect 261478 580864 261484 580876
rect 261536 580864 261542 580916
rect 278590 580864 278596 580916
rect 278648 580904 278654 580916
rect 289722 580904 289728 580916
rect 278648 580876 289728 580904
rect 278648 580864 278654 580876
rect 289722 580864 289728 580876
rect 289780 580864 289786 580916
rect 306926 580864 306932 580916
rect 306984 580904 306990 580916
rect 318058 580904 318064 580916
rect 306984 580876 318064 580904
rect 306984 580864 306990 580876
rect 318058 580864 318064 580876
rect 318116 580864 318122 580916
rect 324314 580864 324320 580916
rect 324372 580904 324378 580916
rect 345750 580904 345756 580916
rect 324372 580876 345756 580904
rect 324372 580864 324378 580876
rect 345750 580864 345756 580876
rect 345808 580864 345814 580916
rect 362862 580864 362868 580916
rect 362920 580904 362926 580916
rect 373166 580904 373172 580916
rect 362920 580876 373172 580904
rect 362920 580864 362926 580876
rect 373166 580864 373172 580876
rect 373224 580864 373230 580916
rect 390646 580864 390652 580916
rect 390704 580904 390710 580916
rect 407114 580904 407120 580916
rect 390704 580876 407120 580904
rect 390704 580864 390710 580876
rect 407114 580864 407120 580876
rect 407172 580864 407178 580916
rect 418614 580864 418620 580916
rect 418672 580904 418678 580916
rect 429930 580904 429936 580916
rect 418672 580876 429936 580904
rect 418672 580864 418678 580876
rect 429930 580864 429936 580876
rect 429988 580864 429994 580916
rect 436646 580864 436652 580916
rect 436704 580904 436710 580916
rect 457438 580904 457444 580916
rect 436704 580876 457444 580904
rect 436704 580864 436710 580876
rect 457438 580864 457444 580876
rect 457496 580864 457502 580916
rect 474642 580864 474648 580916
rect 474700 580904 474706 580916
rect 485130 580904 485136 580916
rect 474700 580876 485136 580904
rect 474700 580864 474706 580876
rect 485130 580864 485136 580876
rect 485188 580864 485194 580916
rect 502610 580864 502616 580916
rect 502668 580904 502674 580916
rect 514018 580904 514024 580916
rect 502668 580876 514024 580904
rect 502668 580864 502674 580876
rect 514018 580864 514024 580876
rect 514076 580864 514082 580916
rect 520642 580864 520648 580916
rect 520700 580904 520706 580916
rect 541618 580904 541624 580916
rect 520700 580876 541624 580904
rect 520700 580864 520706 580876
rect 541618 580864 541624 580876
rect 541676 580864 541682 580916
rect 54846 580796 54852 580848
rect 54904 580836 54910 580848
rect 71774 580836 71780 580848
rect 54904 580808 71780 580836
rect 54904 580796 54910 580808
rect 71774 580796 71780 580808
rect 71832 580796 71838 580848
rect 138934 580796 138940 580848
rect 138992 580836 138998 580848
rect 149882 580836 149888 580848
rect 138992 580808 149888 580836
rect 138992 580796 138998 580808
rect 149882 580796 149888 580808
rect 149940 580796 149946 580848
rect 250622 580796 250628 580848
rect 250680 580836 250686 580848
rect 267734 580836 267740 580848
rect 250680 580808 267740 580836
rect 250680 580796 250686 580808
rect 267734 580796 267740 580808
rect 267792 580796 267798 580848
rect 334618 580796 334624 580848
rect 334676 580836 334682 580848
rect 345658 580836 345664 580848
rect 334676 580808 345664 580836
rect 334676 580796 334682 580808
rect 345658 580796 345664 580808
rect 345716 580796 345722 580848
rect 446950 580796 446956 580848
rect 447008 580836 447014 580848
rect 463694 580836 463700 580848
rect 447008 580808 463700 580836
rect 447008 580796 447014 580808
rect 463694 580796 463700 580808
rect 463752 580796 463758 580848
rect 530946 580796 530952 580848
rect 531004 580836 531010 580848
rect 547966 580836 547972 580848
rect 531004 580808 547972 580836
rect 531004 580796 531010 580808
rect 547966 580796 547972 580808
rect 548024 580796 548030 580848
rect 558638 580252 558644 580304
rect 558696 580292 558702 580304
rect 568758 580292 568764 580304
rect 558696 580264 568764 580292
rect 558696 580252 558702 580264
rect 568758 580252 568764 580264
rect 568816 580252 568822 580304
rect 548334 578892 548340 578944
rect 548392 578932 548398 578944
rect 569034 578932 569040 578944
rect 548392 578904 569040 578932
rect 548392 578892 548398 578904
rect 569034 578892 569040 578904
rect 569092 578892 569098 578944
rect 100018 578348 100024 578400
rect 100076 578388 100082 578400
rect 120994 578388 121000 578400
rect 100076 578360 121000 578388
rect 100076 578348 100082 578360
rect 120994 578348 121000 578360
rect 121052 578348 121058 578400
rect 184014 578348 184020 578400
rect 184072 578388 184078 578400
rect 204898 578388 204904 578400
rect 184072 578360 204904 578388
rect 184072 578348 184078 578360
rect 204898 578348 204904 578360
rect 204956 578348 204962 578400
rect 36906 578280 36912 578332
rect 36964 578320 36970 578332
rect 53926 578320 53932 578332
rect 36964 578292 53932 578320
rect 36964 578280 36970 578292
rect 53926 578280 53932 578292
rect 53984 578280 53990 578332
rect 65886 578280 65892 578332
rect 65944 578320 65950 578332
rect 81986 578320 81992 578332
rect 65944 578292 81992 578320
rect 65944 578280 65950 578292
rect 81986 578280 81992 578292
rect 82044 578280 82050 578332
rect 92842 578280 92848 578332
rect 92900 578320 92906 578332
rect 110322 578320 110328 578332
rect 92900 578292 110328 578320
rect 92900 578280 92906 578292
rect 110322 578280 110328 578292
rect 110380 578280 110386 578332
rect 176746 578280 176752 578332
rect 176804 578320 176810 578332
rect 194318 578320 194324 578332
rect 176804 578292 194324 578320
rect 176804 578280 176810 578292
rect 194318 578280 194324 578292
rect 194376 578280 194382 578332
rect 261478 578280 261484 578332
rect 261536 578320 261542 578332
rect 278314 578320 278320 578332
rect 261536 578292 278320 578320
rect 261536 578280 261542 578292
rect 278314 578280 278320 578292
rect 278372 578280 278378 578332
rect 288894 578280 288900 578332
rect 288952 578320 288958 578332
rect 306006 578320 306012 578332
rect 288952 578292 306012 578320
rect 288952 578280 288958 578292
rect 306006 578280 306012 578292
rect 306064 578280 306070 578332
rect 316770 578280 316776 578332
rect 316828 578320 316834 578332
rect 333974 578320 333980 578332
rect 316828 578292 333980 578320
rect 316828 578280 316834 578292
rect 333974 578280 333980 578292
rect 334032 578280 334038 578332
rect 372890 578280 372896 578332
rect 372948 578320 372954 578332
rect 390002 578320 390008 578332
rect 372948 578292 390008 578320
rect 372948 578280 372954 578292
rect 390002 578280 390008 578292
rect 390060 578280 390066 578332
rect 400766 578280 400772 578332
rect 400824 578320 400830 578332
rect 418338 578320 418344 578332
rect 400824 578292 418344 578320
rect 400824 578280 400830 578292
rect 418338 578280 418344 578292
rect 418396 578280 418402 578332
rect 457438 578280 457444 578332
rect 457496 578320 457502 578332
rect 473998 578320 474004 578332
rect 457496 578292 474004 578320
rect 457496 578280 457502 578292
rect 473998 578280 474004 578292
rect 474056 578280 474062 578332
rect 484854 578280 484860 578332
rect 484912 578320 484918 578332
rect 502334 578320 502340 578332
rect 484912 578292 502340 578320
rect 484912 578280 484918 578292
rect 502334 578280 502340 578292
rect 502392 578280 502398 578332
rect 15286 578212 15292 578264
rect 15344 578252 15350 578264
rect 26326 578252 26332 578264
rect 15344 578224 26332 578252
rect 15344 578212 15350 578224
rect 26326 578212 26332 578224
rect 26384 578212 26390 578264
rect 39298 578212 39304 578264
rect 39356 578252 39362 578264
rect 64230 578252 64236 578264
rect 39356 578224 64236 578252
rect 39356 578212 39362 578224
rect 64230 578212 64236 578224
rect 64288 578212 64294 578264
rect 72326 578212 72332 578264
rect 72384 578252 72390 578264
rect 93118 578252 93124 578264
rect 72384 578224 93124 578252
rect 72384 578212 72390 578224
rect 93118 578212 93124 578224
rect 93176 578212 93182 578264
rect 121086 578212 121092 578264
rect 121144 578252 121150 578264
rect 138014 578252 138020 578264
rect 121144 578224 138020 578252
rect 121144 578212 121150 578224
rect 138014 578212 138020 578224
rect 138072 578212 138078 578264
rect 156322 578212 156328 578264
rect 156380 578252 156386 578264
rect 177298 578252 177304 578264
rect 156380 578224 177304 578252
rect 156380 578212 156386 578224
rect 177298 578212 177304 578224
rect 177356 578212 177362 578264
rect 204806 578212 204812 578264
rect 204864 578252 204870 578264
rect 222194 578252 222200 578264
rect 204864 578224 222200 578252
rect 204864 578212 204870 578224
rect 222194 578212 222200 578224
rect 222252 578212 222258 578264
rect 232774 578212 232780 578264
rect 232832 578252 232838 578264
rect 250070 578252 250076 578264
rect 232832 578224 250076 578252
rect 232832 578212 232838 578224
rect 250070 578212 250076 578224
rect 250128 578212 250134 578264
rect 268010 578212 268016 578264
rect 268068 578252 268074 578264
rect 289078 578252 289084 578264
rect 268068 578224 289084 578252
rect 268068 578212 268074 578224
rect 289078 578212 289084 578224
rect 289136 578212 289142 578264
rect 316862 578212 316868 578264
rect 316920 578252 316926 578264
rect 344278 578252 344284 578264
rect 316920 578224 344284 578252
rect 316920 578212 316926 578224
rect 344278 578212 344284 578224
rect 344336 578212 344342 578264
rect 352006 578212 352012 578264
rect 352064 578252 352070 578264
rect 373258 578252 373264 578264
rect 352064 578224 373264 578252
rect 352064 578212 352070 578224
rect 373258 578212 373264 578224
rect 373316 578212 373322 578264
rect 380342 578212 380348 578264
rect 380400 578252 380406 578264
rect 400858 578252 400864 578264
rect 380400 578224 400864 578252
rect 380400 578212 380406 578224
rect 400858 578212 400864 578224
rect 400916 578212 400922 578264
rect 429838 578212 429844 578264
rect 429896 578252 429902 578264
rect 456610 578252 456616 578264
rect 429896 578224 456616 578252
rect 429896 578212 429902 578224
rect 456610 578212 456616 578224
rect 456668 578212 456674 578264
rect 464338 578212 464344 578264
rect 464396 578252 464402 578264
rect 485038 578252 485044 578264
rect 464396 578224 485044 578252
rect 464396 578212 464402 578224
rect 485038 578212 485044 578224
rect 485096 578212 485102 578264
rect 512730 578212 512736 578264
rect 512788 578252 512794 578264
rect 530302 578252 530308 578264
rect 512788 578224 530308 578252
rect 512788 578212 512794 578224
rect 530302 578212 530308 578224
rect 530360 578212 530366 578264
rect 176746 576376 176752 576428
rect 176804 576376 176810 576428
rect 232774 576376 232780 576428
rect 232832 576376 232838 576428
rect 316770 576376 316776 576428
rect 316828 576376 316834 576428
rect 316862 576376 316868 576428
rect 316920 576376 316926 576428
rect 400766 576376 400772 576428
rect 400824 576376 400830 576428
rect 400858 576376 400864 576428
rect 400916 576376 400922 576428
rect 512730 576376 512736 576428
rect 512788 576376 512794 576428
rect 568758 576376 568764 576428
rect 568816 576376 568822 576428
rect 120718 576240 120724 576292
rect 120776 576280 120782 576292
rect 121086 576280 121092 576292
rect 120776 576252 121092 576280
rect 120776 576240 120782 576252
rect 121086 576240 121092 576252
rect 121144 576240 121150 576292
rect 176764 576224 176792 576376
rect 204714 576240 204720 576292
rect 204772 576280 204778 576292
rect 204990 576280 204996 576292
rect 204772 576252 204996 576280
rect 204772 576240 204778 576252
rect 204990 576240 204996 576252
rect 205048 576240 205054 576292
rect 232792 576224 232820 576376
rect 316788 576224 316816 576376
rect 316880 576224 316908 576376
rect 400784 576224 400812 576376
rect 400876 576224 400904 576376
rect 512748 576224 512776 576376
rect 568776 576224 568804 576376
rect 176746 576172 176752 576224
rect 176804 576172 176810 576224
rect 232774 576172 232780 576224
rect 232832 576172 232838 576224
rect 316770 576172 316776 576224
rect 316828 576172 316834 576224
rect 316862 576172 316868 576224
rect 316920 576172 316926 576224
rect 400766 576172 400772 576224
rect 400824 576172 400830 576224
rect 400858 576172 400864 576224
rect 400916 576172 400922 576224
rect 512730 576172 512736 576224
rect 512788 576172 512794 576224
rect 568758 576172 568764 576224
rect 568816 576172 568822 576224
rect 36814 571208 36820 571260
rect 36872 571248 36878 571260
rect 36998 571248 37004 571260
rect 36872 571220 37004 571248
rect 36872 571208 36878 571220
rect 36998 571208 37004 571220
rect 37056 571208 37062 571260
rect 120902 567944 120908 567996
rect 120960 567944 120966 567996
rect 120920 567792 120948 567944
rect 120902 567740 120908 567792
rect 120960 567740 120966 567792
rect 120810 565088 120816 565140
rect 120868 565128 120874 565140
rect 120994 565128 121000 565140
rect 120868 565100 121000 565128
rect 120868 565088 120874 565100
rect 120994 565088 121000 565100
rect 121052 565088 121058 565140
rect 64874 562300 64880 562352
rect 64932 562340 64938 562352
rect 65886 562340 65892 562352
rect 64932 562312 65892 562340
rect 64932 562300 64938 562312
rect 65886 562300 65892 562312
rect 65944 562300 65950 562352
rect 289078 560192 289084 560244
rect 289136 560232 289142 560244
rect 295702 560232 295708 560244
rect 289136 560204 295708 560232
rect 289136 560192 289142 560204
rect 295702 560192 295708 560204
rect 295760 560192 295766 560244
rect 93118 559512 93124 559564
rect 93176 559552 93182 559564
rect 99742 559552 99748 559564
rect 93176 559524 99748 559552
rect 93176 559512 93182 559524
rect 99742 559512 99748 559524
rect 99800 559512 99806 559564
rect 120810 559512 120816 559564
rect 120868 559552 120874 559564
rect 127710 559552 127716 559564
rect 120868 559524 127716 559552
rect 120868 559512 120874 559524
rect 127710 559512 127716 559524
rect 127768 559512 127774 559564
rect 177298 559512 177304 559564
rect 177356 559552 177362 559564
rect 183738 559552 183744 559564
rect 177356 559524 183744 559552
rect 177356 559512 177362 559524
rect 183738 559512 183744 559524
rect 183796 559512 183802 559564
rect 373258 559512 373264 559564
rect 373316 559552 373322 559564
rect 379698 559552 379704 559564
rect 373316 559524 379704 559552
rect 373316 559512 373322 559524
rect 379698 559512 379704 559524
rect 379756 559512 379762 559564
rect 400858 559512 400864 559564
rect 400916 559552 400922 559564
rect 407758 559552 407764 559564
rect 400916 559524 407764 559552
rect 400916 559512 400922 559524
rect 407758 559512 407764 559524
rect 407816 559512 407822 559564
rect 204898 558900 204904 558952
rect 204956 558940 204962 558952
rect 211706 558940 211712 558952
rect 204956 558912 211712 558940
rect 204956 558900 204962 558912
rect 211706 558900 211712 558912
rect 211764 558900 211770 558952
rect 485038 558900 485044 558952
rect 485096 558940 485102 558952
rect 491662 558940 491668 558952
rect 485096 558912 491668 558940
rect 485096 558900 485102 558912
rect 491662 558900 491668 558912
rect 491720 558900 491726 558952
rect 42702 557472 42708 557524
rect 42760 557512 42766 557524
rect 95234 557512 95240 557524
rect 42760 557484 95240 557512
rect 42760 557472 42766 557484
rect 95234 557472 95240 557484
rect 95292 557472 95298 557524
rect 97902 557472 97908 557524
rect 97960 557512 97966 557524
rect 150434 557512 150440 557524
rect 97960 557484 150440 557512
rect 97960 557472 97966 557484
rect 150434 557472 150440 557484
rect 150492 557472 150498 557524
rect 154482 557472 154488 557524
rect 154540 557512 154546 557524
rect 207014 557512 207020 557524
rect 154540 557484 207020 557512
rect 154540 557472 154546 557484
rect 207014 557472 207020 557484
rect 207072 557472 207078 557524
rect 209682 557472 209688 557524
rect 209740 557512 209746 557524
rect 262214 557512 262220 557524
rect 209740 557484 262220 557512
rect 209740 557472 209746 557484
rect 262214 557472 262220 557484
rect 262272 557472 262278 557524
rect 266262 557472 266268 557524
rect 266320 557512 266326 557524
rect 318794 557512 318800 557524
rect 266320 557484 318800 557512
rect 266320 557472 266326 557484
rect 318794 557472 318800 557484
rect 318852 557472 318858 557524
rect 322842 557472 322848 557524
rect 322900 557512 322906 557524
rect 375374 557512 375380 557524
rect 322900 557484 375380 557512
rect 322900 557472 322906 557484
rect 375374 557472 375380 557484
rect 375432 557472 375438 557524
rect 378042 557472 378048 557524
rect 378100 557512 378106 557524
rect 430574 557512 430580 557524
rect 378100 557484 430580 557512
rect 378100 557472 378106 557484
rect 430574 557472 430580 557484
rect 430632 557472 430638 557524
rect 434622 557472 434628 557524
rect 434680 557512 434686 557524
rect 487154 557512 487160 557524
rect 434680 557484 487160 557512
rect 434680 557472 434686 557484
rect 487154 557472 487160 557484
rect 487212 557472 487218 557524
rect 489822 557472 489828 557524
rect 489880 557512 489886 557524
rect 542354 557512 542360 557524
rect 489880 557484 542360 557512
rect 489880 557472 489886 557484
rect 542354 557472 542360 557484
rect 542412 557472 542418 557524
rect 288802 556792 288808 556844
rect 288860 556832 288866 556844
rect 288986 556832 288992 556844
rect 288860 556804 288992 556832
rect 288860 556792 288866 556804
rect 288986 556792 288992 556804
rect 289044 556792 289050 556844
rect 372798 556792 372804 556844
rect 372856 556832 372862 556844
rect 372982 556832 372988 556844
rect 372856 556804 372988 556832
rect 372856 556792 372862 556804
rect 372982 556792 372988 556804
rect 373040 556792 373046 556844
rect 484762 556792 484768 556844
rect 484820 556832 484826 556844
rect 484946 556832 484952 556844
rect 484820 556804 484952 556832
rect 484820 556792 484826 556804
rect 484946 556792 484952 556804
rect 485004 556792 485010 556844
rect 87414 556588 87420 556640
rect 87472 556628 87478 556640
rect 92750 556628 92756 556640
rect 87472 556600 92756 556628
rect 87472 556588 87478 556600
rect 92750 556588 92756 556600
rect 92808 556588 92814 556640
rect 547874 556112 547880 556164
rect 547932 556152 547938 556164
rect 548150 556152 548156 556164
rect 547932 556124 548156 556152
rect 547932 556112 547938 556124
rect 548150 556112 548156 556124
rect 548208 556112 548214 556164
rect 15378 554684 15384 554736
rect 15436 554724 15442 554736
rect 43990 554724 43996 554736
rect 15436 554696 43996 554724
rect 15436 554684 15442 554696
rect 43990 554684 43996 554696
rect 44048 554684 44054 554736
rect 138290 554684 138296 554736
rect 138348 554724 138354 554736
rect 176838 554724 176844 554736
rect 138348 554696 176844 554724
rect 138348 554684 138354 554696
rect 176838 554684 176844 554696
rect 176896 554684 176902 554736
rect 194318 554684 194324 554736
rect 194376 554724 194382 554736
rect 232866 554724 232872 554736
rect 194376 554696 232872 554724
rect 194376 554684 194382 554696
rect 232866 554684 232872 554696
rect 232924 554684 232930 554736
rect 238846 554684 238852 554736
rect 238904 554724 238910 554736
rect 238904 554696 248414 554724
rect 238904 554684 238910 554696
rect 26326 554616 26332 554668
rect 26384 554656 26390 554668
rect 39298 554656 39304 554668
rect 26384 554628 39304 554656
rect 26384 554616 26390 554628
rect 39298 554616 39304 554628
rect 39356 554616 39362 554668
rect 42886 554616 42892 554668
rect 42944 554656 42950 554668
rect 71774 554656 71780 554668
rect 42944 554628 71780 554656
rect 42944 554616 42950 554628
rect 71774 554616 71780 554628
rect 71832 554616 71838 554668
rect 110322 554616 110328 554668
rect 110380 554656 110386 554668
rect 148778 554656 148784 554668
rect 110380 554628 148784 554656
rect 110380 554616 110386 554628
rect 148778 554616 148784 554628
rect 148836 554616 148842 554668
rect 166626 554616 166632 554668
rect 166684 554656 166690 554668
rect 204990 554656 204996 554668
rect 166684 554628 204996 554656
rect 166684 554616 166690 554628
rect 204990 554616 204996 554628
rect 205048 554616 205054 554668
rect 211246 554616 211252 554668
rect 211304 554656 211310 554668
rect 240042 554656 240048 554668
rect 211304 554628 240048 554656
rect 211304 554616 211310 554628
rect 240042 554616 240048 554628
rect 240100 554616 240106 554668
rect 248386 554656 248414 554696
rect 295426 554684 295432 554736
rect 295484 554724 295490 554736
rect 324038 554724 324044 554736
rect 295484 554696 324044 554724
rect 295484 554684 295490 554696
rect 324038 554684 324044 554696
rect 324096 554684 324102 554736
rect 334342 554684 334348 554736
rect 334400 554724 334406 554736
rect 372982 554724 372988 554736
rect 334400 554696 372988 554724
rect 334400 554684 334406 554696
rect 372982 554684 372988 554696
rect 373040 554684 373046 554736
rect 390462 554684 390468 554736
rect 390520 554724 390526 554736
rect 428734 554724 428740 554736
rect 390520 554696 428740 554724
rect 390520 554684 390526 554696
rect 428734 554684 428740 554696
rect 428792 554684 428798 554736
rect 434806 554684 434812 554736
rect 434864 554724 434870 554736
rect 434864 554696 441614 554724
rect 434864 554684 434870 554696
rect 268010 554656 268016 554668
rect 248386 554628 268016 554656
rect 268010 554616 268016 554628
rect 268068 554616 268074 554668
rect 278314 554616 278320 554668
rect 278372 554656 278378 554668
rect 316954 554656 316960 554668
rect 278372 554628 316960 554656
rect 278372 554616 278378 554628
rect 316954 554616 316960 554628
rect 317012 554616 317018 554668
rect 323026 554616 323032 554668
rect 323084 554656 323090 554668
rect 352006 554656 352012 554668
rect 323084 554628 352012 554656
rect 323084 554616 323090 554628
rect 352006 554616 352012 554628
rect 352064 554616 352070 554668
rect 362310 554616 362316 554668
rect 362368 554656 362374 554668
rect 400950 554656 400956 554668
rect 362368 554628 400956 554656
rect 362368 554616 362374 554628
rect 400950 554616 400956 554628
rect 401008 554616 401014 554668
rect 407206 554616 407212 554668
rect 407264 554656 407270 554668
rect 436002 554656 436008 554668
rect 407264 554628 436008 554656
rect 407264 554616 407270 554628
rect 436002 554616 436008 554628
rect 436060 554616 436066 554668
rect 441586 554656 441614 554696
rect 491386 554684 491392 554736
rect 491444 554724 491450 554736
rect 519998 554724 520004 554736
rect 491444 554696 520004 554724
rect 491444 554684 491450 554696
rect 519998 554684 520004 554696
rect 520056 554684 520062 554736
rect 530302 554684 530308 554736
rect 530360 554724 530366 554736
rect 568850 554724 568856 554736
rect 530360 554696 568856 554724
rect 530360 554684 530366 554696
rect 568850 554684 568856 554696
rect 568908 554684 568914 554736
rect 463694 554656 463700 554668
rect 441586 554628 463700 554656
rect 463694 554616 463700 554628
rect 463752 554616 463758 554668
rect 474642 554616 474648 554668
rect 474700 554656 474706 554668
rect 512822 554656 512828 554668
rect 474700 554628 512828 554656
rect 474700 554616 474706 554628
rect 512822 554616 512828 554628
rect 512880 554616 512886 554668
rect 548150 554616 548156 554668
rect 548208 554656 548214 554668
rect 557994 554656 558000 554668
rect 548208 554628 558000 554656
rect 548208 554616 548214 554628
rect 557994 554616 558000 554628
rect 558052 554616 558058 554668
rect 82630 554548 82636 554600
rect 82688 554588 82694 554600
rect 120902 554588 120908 554600
rect 82688 554560 120908 554588
rect 82688 554548 82694 554560
rect 120902 554548 120908 554560
rect 120960 554548 120966 554600
rect 127066 554548 127072 554600
rect 127124 554588 127130 554600
rect 156046 554588 156052 554600
rect 127124 554560 156052 554588
rect 127124 554548 127130 554560
rect 156046 554548 156052 554560
rect 156104 554548 156110 554600
rect 250346 554548 250352 554600
rect 250404 554588 250410 554600
rect 288986 554588 288992 554600
rect 250404 554560 288992 554588
rect 250404 554548 250410 554560
rect 288986 554548 288992 554560
rect 289044 554548 289050 554600
rect 306282 554548 306288 554600
rect 306340 554588 306346 554600
rect 316862 554588 316868 554600
rect 306340 554560 316868 554588
rect 306340 554548 306346 554560
rect 316862 554548 316868 554560
rect 316920 554548 316926 554600
rect 418338 554548 418344 554600
rect 418396 554588 418402 554600
rect 429838 554588 429844 554600
rect 418396 554560 429844 554588
rect 418396 554548 418402 554560
rect 429838 554548 429844 554560
rect 429896 554548 429902 554600
rect 446306 554548 446312 554600
rect 446364 554588 446370 554600
rect 484946 554588 484952 554600
rect 446364 554560 484952 554588
rect 446364 554548 446370 554560
rect 484946 554548 484952 554560
rect 485004 554548 485010 554600
rect 502334 554548 502340 554600
rect 502392 554588 502398 554600
rect 540790 554588 540796 554600
rect 502392 554560 540796 554588
rect 502392 554548 502398 554560
rect 540790 554548 540796 554560
rect 540848 554548 540854 554600
rect 54294 554480 54300 554532
rect 54352 554520 54358 554532
rect 87414 554520 87420 554532
rect 54352 554492 87420 554520
rect 54352 554480 54358 554492
rect 87414 554480 87420 554492
rect 87472 554480 87478 554532
rect 518986 554480 518992 554532
rect 519044 554520 519050 554532
rect 547874 554520 547880 554532
rect 519044 554492 547880 554520
rect 519044 554480 519050 554492
rect 547874 554480 547880 554492
rect 547932 554480 547938 554532
rect 3602 553392 3608 553444
rect 3660 553432 3666 553444
rect 10318 553432 10324 553444
rect 3660 553404 10324 553432
rect 3660 553392 3666 553404
rect 10318 553392 10324 553404
rect 10376 553392 10382 553444
rect 15286 553324 15292 553376
rect 15344 553364 15350 553376
rect 16022 553364 16028 553376
rect 15344 553336 16028 553364
rect 15344 553324 15350 553336
rect 16022 553324 16028 553336
rect 16080 553324 16086 553376
rect 26602 552644 26608 552696
rect 26660 552684 26666 552696
rect 36814 552684 36820 552696
rect 26660 552656 36820 552684
rect 26660 552644 26666 552656
rect 36814 552644 36820 552656
rect 36872 552644 36878 552696
rect 15562 552168 15568 552220
rect 15620 552208 15626 552220
rect 54294 552208 54300 552220
rect 15620 552180 54300 552208
rect 15620 552168 15626 552180
rect 54294 552168 54300 552180
rect 54352 552168 54358 552220
rect 429838 552168 429844 552220
rect 429896 552208 429902 552220
rect 436094 552208 436100 552220
rect 429896 552180 436100 552208
rect 429896 552168 429902 552180
rect 436094 552168 436100 552180
rect 436152 552168 436158 552220
rect 71774 552100 71780 552152
rect 71832 552140 71838 552152
rect 110598 552140 110604 552152
rect 71832 552112 110604 552140
rect 71832 552100 71838 552112
rect 110598 552100 110604 552112
rect 110656 552100 110662 552152
rect 149882 552100 149888 552152
rect 149940 552140 149946 552152
rect 156322 552140 156328 552152
rect 149940 552112 156328 552140
rect 149940 552100 149946 552112
rect 156322 552100 156328 552112
rect 156380 552100 156386 552152
rect 211154 552100 211160 552152
rect 211212 552140 211218 552152
rect 250622 552140 250628 552152
rect 211212 552112 250628 552140
rect 211212 552100 211218 552112
rect 250622 552100 250628 552112
rect 250680 552100 250686 552152
rect 261478 552100 261484 552152
rect 261536 552140 261542 552152
rect 278590 552140 278596 552152
rect 261536 552112 278596 552140
rect 261536 552100 261542 552112
rect 278590 552100 278596 552112
rect 278648 552100 278654 552152
rect 295334 552100 295340 552152
rect 295392 552140 295398 552152
rect 334618 552140 334624 552152
rect 295392 552112 334624 552140
rect 295392 552100 295398 552112
rect 334618 552100 334624 552112
rect 334676 552100 334682 552152
rect 345750 552100 345756 552152
rect 345808 552140 345814 552152
rect 362310 552140 362316 552152
rect 345808 552112 362316 552140
rect 345808 552100 345814 552112
rect 362310 552100 362316 552112
rect 362368 552100 362374 552152
rect 407114 552100 407120 552152
rect 407172 552140 407178 552152
rect 446306 552140 446312 552152
rect 407172 552112 446312 552140
rect 407172 552100 407178 552112
rect 446306 552100 446312 552112
rect 446364 552100 446370 552152
rect 457438 552100 457444 552152
rect 457496 552140 457502 552152
rect 474642 552140 474648 552152
rect 457496 552112 474648 552140
rect 457496 552100 457502 552112
rect 474642 552100 474648 552112
rect 474700 552100 474706 552152
rect 491294 552100 491300 552152
rect 491352 552140 491358 552152
rect 530302 552140 530308 552152
rect 491352 552112 530308 552140
rect 491352 552100 491358 552112
rect 530302 552100 530308 552112
rect 530360 552100 530366 552152
rect 38010 552032 38016 552084
rect 38068 552072 38074 552084
rect 44174 552072 44180 552084
rect 38068 552044 44180 552072
rect 38068 552032 38074 552044
rect 44174 552032 44180 552044
rect 44232 552032 44238 552084
rect 65886 552032 65892 552084
rect 65944 552072 65950 552084
rect 82630 552072 82636 552084
rect 65944 552044 82636 552072
rect 65944 552032 65950 552044
rect 82630 552032 82636 552044
rect 82688 552032 82694 552084
rect 99374 552032 99380 552084
rect 99432 552072 99438 552084
rect 138290 552072 138296 552084
rect 99432 552044 138296 552072
rect 99432 552032 99438 552044
rect 138290 552032 138296 552044
rect 138348 552032 138354 552084
rect 149790 552032 149796 552084
rect 149848 552072 149854 552084
rect 166626 552072 166632 552084
rect 149848 552044 166632 552072
rect 149848 552032 149854 552044
rect 166626 552032 166632 552044
rect 166684 552032 166690 552084
rect 183554 552032 183560 552084
rect 183612 552072 183618 552084
rect 222286 552072 222292 552084
rect 183612 552044 222292 552072
rect 183612 552032 183618 552044
rect 222286 552032 222292 552044
rect 222344 552032 222350 552084
rect 267734 552032 267740 552084
rect 267792 552072 267798 552084
rect 306466 552072 306472 552084
rect 267792 552044 306472 552072
rect 267792 552032 267798 552044
rect 306466 552032 306472 552044
rect 306524 552032 306530 552084
rect 318058 552032 318064 552084
rect 318116 552072 318122 552084
rect 324314 552072 324320 552084
rect 318116 552044 324320 552072
rect 318116 552032 318122 552044
rect 324314 552032 324320 552044
rect 324372 552032 324378 552084
rect 345842 552032 345848 552084
rect 345900 552072 345906 552084
rect 352006 552072 352012 552084
rect 345900 552044 352012 552072
rect 345900 552032 345906 552044
rect 352006 552032 352012 552044
rect 352064 552032 352070 552084
rect 379514 552032 379520 552084
rect 379572 552072 379578 552084
rect 418614 552072 418620 552084
rect 379572 552044 418620 552072
rect 379572 552032 379578 552044
rect 418614 552032 418620 552044
rect 418672 552032 418678 552084
rect 463694 552032 463700 552084
rect 463752 552072 463758 552084
rect 502610 552072 502616 552084
rect 463752 552044 502616 552072
rect 463752 552032 463758 552044
rect 502610 552032 502616 552044
rect 502668 552032 502674 552084
rect 541618 552032 541624 552084
rect 541676 552072 541682 552084
rect 558638 552072 558644 552084
rect 541676 552044 558644 552072
rect 541676 552032 541682 552044
rect 558638 552032 558644 552044
rect 558696 552032 558702 552084
rect 233970 550536 233976 550588
rect 234028 550576 234034 550588
rect 240134 550576 240140 550588
rect 234028 550548 240140 550576
rect 234028 550536 234034 550548
rect 240134 550536 240140 550548
rect 240192 550536 240198 550588
rect 514018 550536 514024 550588
rect 514076 550576 514082 550588
rect 520274 550576 520280 550588
rect 514076 550548 520280 550576
rect 514076 550536 514082 550548
rect 520274 550536 520280 550548
rect 520332 550536 520338 550588
rect 205082 549312 205088 549364
rect 205140 549312 205146 549364
rect 205100 549160 205128 549312
rect 429102 549244 429108 549296
rect 429160 549284 429166 549296
rect 429930 549284 429936 549296
rect 429160 549256 429936 549284
rect 429160 549244 429166 549256
rect 429930 549244 429936 549256
rect 429988 549244 429994 549296
rect 205082 549108 205088 549160
rect 205140 549108 205146 549160
rect 37274 548496 37280 548548
rect 37332 548536 37338 548548
rect 38102 548536 38108 548548
rect 37332 548508 38108 548536
rect 37332 548496 37338 548508
rect 38102 548496 38108 548508
rect 38160 548496 38166 548548
rect 233234 548496 233240 548548
rect 233292 548536 233298 548548
rect 234062 548536 234068 548548
rect 233292 548508 234068 548536
rect 233292 548496 233298 548508
rect 234062 548496 234068 548508
rect 234120 548496 234126 548548
rect 71774 533604 71780 533656
rect 71832 533644 71838 533656
rect 72050 533644 72056 533656
rect 71832 533616 72056 533644
rect 71832 533604 71838 533616
rect 72050 533604 72056 533616
rect 72108 533604 72114 533656
rect 99374 533604 99380 533656
rect 99432 533644 99438 533656
rect 99926 533644 99932 533656
rect 99432 533616 99932 533644
rect 99432 533604 99438 533616
rect 99926 533604 99932 533616
rect 99984 533604 99990 533656
rect 183554 533604 183560 533656
rect 183612 533644 183618 533656
rect 184014 533644 184020 533656
rect 183612 533616 184020 533644
rect 183612 533604 183618 533616
rect 184014 533604 184020 533616
rect 184072 533604 184078 533656
rect 211154 533604 211160 533656
rect 211212 533644 211218 533656
rect 211982 533644 211988 533656
rect 211212 533616 211988 533644
rect 211212 533604 211218 533616
rect 211982 533604 211988 533616
rect 212040 533604 212046 533656
rect 267734 533604 267740 533656
rect 267792 533644 267798 533656
rect 268010 533644 268016 533656
rect 267792 533616 268016 533644
rect 267792 533604 267798 533616
rect 268010 533604 268016 533616
rect 268068 533604 268074 533656
rect 295334 533604 295340 533656
rect 295392 533644 295398 533656
rect 295978 533644 295984 533656
rect 295392 533616 295984 533644
rect 295392 533604 295398 533616
rect 295978 533604 295984 533616
rect 296036 533604 296042 533656
rect 379514 533604 379520 533656
rect 379572 533644 379578 533656
rect 379974 533644 379980 533656
rect 379572 533616 379980 533644
rect 379572 533604 379578 533616
rect 379974 533604 379980 533616
rect 380032 533604 380038 533656
rect 407114 533604 407120 533656
rect 407172 533644 407178 533656
rect 407942 533644 407948 533656
rect 407172 533616 407948 533644
rect 407172 533604 407178 533616
rect 407942 533604 407948 533616
rect 408000 533604 408006 533656
rect 463694 533604 463700 533656
rect 463752 533644 463758 533656
rect 464062 533644 464068 533656
rect 463752 533616 464068 533644
rect 463752 533604 463758 533616
rect 464062 533604 464068 533616
rect 464120 533604 464126 533656
rect 491294 531904 491300 531956
rect 491352 531944 491358 531956
rect 492030 531944 492036 531956
rect 491352 531916 492036 531944
rect 491352 531904 491358 531916
rect 492030 531904 492036 531916
rect 492088 531904 492094 531956
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 6178 527184 6184 527196
rect 3016 527156 6184 527184
rect 3016 527144 3022 527156
rect 6178 527144 6184 527156
rect 6236 527144 6242 527196
rect 15194 527076 15200 527128
rect 15252 527116 15258 527128
rect 36906 527116 36912 527128
rect 15252 527088 36912 527116
rect 15252 527076 15258 527088
rect 36906 527076 36912 527088
rect 36964 527076 36970 527128
rect 38102 527076 38108 527128
rect 38160 527116 38166 527128
rect 64874 527116 64880 527128
rect 38160 527088 64880 527116
rect 38160 527076 38166 527088
rect 64874 527076 64880 527088
rect 64932 527076 64938 527128
rect 65058 527076 65064 527128
rect 65116 527116 65122 527128
rect 92934 527116 92940 527128
rect 65116 527088 92940 527116
rect 65116 527076 65122 527088
rect 92934 527076 92940 527088
rect 92992 527076 92998 527128
rect 93026 527076 93032 527128
rect 93084 527116 93090 527128
rect 120902 527116 120908 527128
rect 93084 527088 120908 527116
rect 93084 527076 93090 527088
rect 120902 527076 120908 527088
rect 120960 527076 120966 527128
rect 121086 527076 121092 527128
rect 121144 527116 121150 527128
rect 148594 527116 148600 527128
rect 121144 527088 148600 527116
rect 121144 527076 121150 527088
rect 148594 527076 148600 527088
rect 148652 527076 148658 527128
rect 149698 527076 149704 527128
rect 149756 527116 149762 527128
rect 176930 527116 176936 527128
rect 149756 527088 176936 527116
rect 149756 527076 149762 527088
rect 176930 527076 176936 527088
rect 176988 527076 176994 527128
rect 177022 527076 177028 527128
rect 177080 527116 177086 527128
rect 204898 527116 204904 527128
rect 177080 527088 204904 527116
rect 177080 527076 177086 527088
rect 204898 527076 204904 527088
rect 204956 527076 204962 527128
rect 205174 527076 205180 527128
rect 205232 527116 205238 527128
rect 232590 527116 232596 527128
rect 205232 527088 232596 527116
rect 205232 527076 205238 527088
rect 232590 527076 232596 527088
rect 232648 527076 232654 527128
rect 234062 527076 234068 527128
rect 234120 527116 234126 527128
rect 260926 527116 260932 527128
rect 234120 527088 260932 527116
rect 234120 527076 234126 527088
rect 260926 527076 260932 527088
rect 260984 527076 260990 527128
rect 261018 527076 261024 527128
rect 261076 527116 261082 527128
rect 288894 527116 288900 527128
rect 261076 527088 288900 527116
rect 261076 527076 261082 527088
rect 288894 527076 288900 527088
rect 288952 527076 288958 527128
rect 289078 527076 289084 527128
rect 289136 527116 289142 527128
rect 316586 527116 316592 527128
rect 289136 527088 316592 527116
rect 289136 527076 289142 527088
rect 316586 527076 316592 527088
rect 316644 527076 316650 527128
rect 317046 527076 317052 527128
rect 317104 527116 317110 527128
rect 344922 527116 344928 527128
rect 317104 527088 344928 527116
rect 317104 527076 317110 527088
rect 344922 527076 344928 527088
rect 344980 527076 344986 527128
rect 345658 527076 345664 527128
rect 345716 527116 345722 527128
rect 372614 527116 372620 527128
rect 345716 527088 372620 527116
rect 345716 527076 345722 527088
rect 372614 527076 372620 527088
rect 372672 527076 372678 527128
rect 373074 527076 373080 527128
rect 373132 527116 373138 527128
rect 400950 527116 400956 527128
rect 373132 527088 400956 527116
rect 373132 527076 373138 527088
rect 400950 527076 400956 527088
rect 401008 527076 401014 527128
rect 401042 527076 401048 527128
rect 401100 527116 401106 527128
rect 428918 527116 428924 527128
rect 401100 527088 428924 527116
rect 401100 527076 401106 527088
rect 428918 527076 428924 527088
rect 428976 527076 428982 527128
rect 429930 527076 429936 527128
rect 429988 527116 429994 527128
rect 456794 527116 456800 527128
rect 429988 527088 456800 527116
rect 429988 527076 429994 527088
rect 456794 527076 456800 527088
rect 456852 527076 456858 527128
rect 457070 527076 457076 527128
rect 457128 527116 457134 527128
rect 484946 527116 484952 527128
rect 457128 527088 484952 527116
rect 457128 527076 457134 527088
rect 484946 527076 484952 527088
rect 485004 527076 485010 527128
rect 485038 527076 485044 527128
rect 485096 527116 485102 527128
rect 512914 527116 512920 527128
rect 485096 527088 512920 527116
rect 485096 527076 485102 527088
rect 512914 527076 512920 527088
rect 512972 527076 512978 527128
rect 513098 527076 513104 527128
rect 513156 527116 513162 527128
rect 540606 527116 540612 527128
rect 513156 527088 540612 527116
rect 513156 527076 513162 527088
rect 540606 527076 540612 527088
rect 540664 527076 540670 527128
rect 541066 527076 541072 527128
rect 541124 527116 541130 527128
rect 568942 527116 568948 527128
rect 541124 527088 568948 527116
rect 541124 527076 541130 527088
rect 568942 527076 568948 527088
rect 569000 527076 569006 527128
rect 26602 527008 26608 527060
rect 26660 527048 26666 527060
rect 38010 527048 38016 527060
rect 26660 527020 38016 527048
rect 26660 527008 26666 527020
rect 38010 527008 38016 527020
rect 38068 527008 38074 527060
rect 44634 527008 44640 527060
rect 44692 527048 44698 527060
rect 65886 527048 65892 527060
rect 44692 527020 65892 527048
rect 44692 527008 44698 527020
rect 65886 527008 65892 527020
rect 65944 527008 65950 527060
rect 82630 527008 82636 527060
rect 82688 527048 82694 527060
rect 99466 527048 99472 527060
rect 82688 527020 99472 527048
rect 82688 527008 82694 527020
rect 99466 527008 99472 527020
rect 99524 527008 99530 527060
rect 128630 527008 128636 527060
rect 128688 527048 128694 527060
rect 149790 527048 149796 527060
rect 128688 527020 149796 527048
rect 128688 527008 128694 527020
rect 149790 527008 149796 527020
rect 149848 527008 149854 527060
rect 166626 527008 166632 527060
rect 166684 527048 166690 527060
rect 183646 527048 183652 527060
rect 166684 527020 183652 527048
rect 166684 527008 166690 527020
rect 183646 527008 183652 527020
rect 183704 527008 183710 527060
rect 194594 527008 194600 527060
rect 194652 527048 194658 527060
rect 211246 527048 211252 527060
rect 194652 527020 211252 527048
rect 194652 527008 194658 527020
rect 211246 527008 211252 527020
rect 211304 527008 211310 527060
rect 222930 527008 222936 527060
rect 222988 527048 222994 527060
rect 233970 527048 233976 527060
rect 222988 527020 233976 527048
rect 222988 527008 222994 527020
rect 233970 527008 233976 527020
rect 234028 527008 234034 527060
rect 240318 527008 240324 527060
rect 240376 527048 240382 527060
rect 261478 527048 261484 527060
rect 240376 527020 261484 527048
rect 240376 527008 240382 527020
rect 261478 527008 261484 527020
rect 261536 527008 261542 527060
rect 278590 527008 278596 527060
rect 278648 527048 278654 527060
rect 295426 527048 295432 527060
rect 278648 527020 295432 527048
rect 278648 527008 278654 527020
rect 295426 527008 295432 527020
rect 295484 527008 295490 527060
rect 306926 527008 306932 527060
rect 306984 527048 306990 527060
rect 318058 527048 318064 527060
rect 306984 527020 318064 527048
rect 306984 527008 306990 527020
rect 318058 527008 318064 527020
rect 318116 527008 318122 527060
rect 324314 527008 324320 527060
rect 324372 527048 324378 527060
rect 345750 527048 345756 527060
rect 324372 527020 345756 527048
rect 324372 527008 324378 527020
rect 345750 527008 345756 527020
rect 345808 527008 345814 527060
rect 362862 527008 362868 527060
rect 362920 527048 362926 527060
rect 379606 527048 379612 527060
rect 362920 527020 379612 527048
rect 362920 527008 362926 527020
rect 379606 527008 379612 527020
rect 379664 527008 379670 527060
rect 390646 527008 390652 527060
rect 390704 527048 390710 527060
rect 407206 527048 407212 527060
rect 390704 527020 407212 527048
rect 390704 527008 390710 527020
rect 407206 527008 407212 527020
rect 407264 527008 407270 527060
rect 418614 527008 418620 527060
rect 418672 527048 418678 527060
rect 429838 527048 429844 527060
rect 418672 527020 429844 527048
rect 418672 527008 418678 527020
rect 429838 527008 429844 527020
rect 429896 527008 429902 527060
rect 436646 527008 436652 527060
rect 436704 527048 436710 527060
rect 457438 527048 457444 527060
rect 436704 527020 457444 527048
rect 436704 527008 436710 527020
rect 457438 527008 457444 527020
rect 457496 527008 457502 527060
rect 474642 527008 474648 527060
rect 474700 527048 474706 527060
rect 491386 527048 491392 527060
rect 474700 527020 491392 527048
rect 474700 527008 474706 527020
rect 491386 527008 491392 527020
rect 491444 527008 491450 527060
rect 502610 527008 502616 527060
rect 502668 527048 502674 527060
rect 514018 527048 514024 527060
rect 502668 527020 514024 527048
rect 502668 527008 502674 527020
rect 514018 527008 514024 527020
rect 514076 527008 514082 527060
rect 520642 527008 520648 527060
rect 520700 527048 520706 527060
rect 541618 527048 541624 527060
rect 520700 527020 541624 527048
rect 520700 527008 520706 527020
rect 541618 527008 541624 527020
rect 541676 527008 541682 527060
rect 54938 526940 54944 526992
rect 54996 526980 55002 526992
rect 71866 526980 71872 526992
rect 54996 526952 71872 526980
rect 54996 526940 55002 526952
rect 71866 526940 71872 526952
rect 71924 526940 71930 526992
rect 138934 526940 138940 526992
rect 138992 526980 138998 526992
rect 149882 526980 149888 526992
rect 138992 526952 149888 526980
rect 138992 526940 138998 526952
rect 149882 526940 149888 526952
rect 149940 526940 149946 526992
rect 250622 526940 250628 526992
rect 250680 526980 250686 526992
rect 267826 526980 267832 526992
rect 250680 526952 267832 526980
rect 250680 526940 250686 526952
rect 267826 526940 267832 526952
rect 267884 526940 267890 526992
rect 334618 526940 334624 526992
rect 334676 526980 334682 526992
rect 345842 526980 345848 526992
rect 334676 526952 345848 526980
rect 334676 526940 334682 526952
rect 345842 526940 345848 526952
rect 345900 526940 345906 526992
rect 446950 526940 446956 526992
rect 447008 526980 447014 526992
rect 463786 526980 463792 526992
rect 447008 526952 463792 526980
rect 447008 526940 447014 526952
rect 463786 526940 463792 526952
rect 463844 526940 463850 526992
rect 530946 526940 530952 526992
rect 531004 526980 531010 526992
rect 547966 526980 547972 526992
rect 531004 526952 547972 526980
rect 531004 526940 531010 526952
rect 547966 526940 547972 526952
rect 548024 526940 548030 526992
rect 558638 526396 558644 526448
rect 558696 526436 558702 526448
rect 568942 526436 568948 526448
rect 558696 526408 568948 526436
rect 558696 526396 558702 526408
rect 568942 526396 568948 526408
rect 569000 526396 569006 526448
rect 548334 525036 548340 525088
rect 548392 525076 548398 525088
rect 569034 525076 569040 525088
rect 548392 525048 569040 525076
rect 548392 525036 548398 525048
rect 569034 525036 569040 525048
rect 569092 525036 569098 525088
rect 184014 524560 184020 524612
rect 184072 524600 184078 524612
rect 204898 524600 204904 524612
rect 184072 524572 204904 524600
rect 184072 524560 184078 524572
rect 204898 524560 204904 524572
rect 204956 524560 204962 524612
rect 464338 524560 464344 524612
rect 464396 524600 464402 524612
rect 485038 524600 485044 524612
rect 464396 524572 485044 524600
rect 464396 524560 464402 524572
rect 485038 524560 485044 524572
rect 485096 524560 485102 524612
rect 37090 524492 37096 524544
rect 37148 524532 37154 524544
rect 54294 524532 54300 524544
rect 37148 524504 54300 524532
rect 37148 524492 37154 524504
rect 54294 524492 54300 524504
rect 54352 524492 54358 524544
rect 65886 524492 65892 524544
rect 65944 524532 65950 524544
rect 81986 524532 81992 524544
rect 65944 524504 81992 524532
rect 65944 524492 65950 524504
rect 81986 524492 81992 524504
rect 82044 524492 82050 524544
rect 92842 524492 92848 524544
rect 92900 524532 92906 524544
rect 110322 524532 110328 524544
rect 92900 524504 110328 524532
rect 92900 524492 92906 524504
rect 110322 524492 110328 524504
rect 110380 524492 110386 524544
rect 120994 524492 121000 524544
rect 121052 524532 121058 524544
rect 138290 524532 138296 524544
rect 121052 524504 138296 524532
rect 121052 524492 121058 524504
rect 138290 524492 138296 524504
rect 138348 524492 138354 524544
rect 177022 524492 177028 524544
rect 177080 524532 177086 524544
rect 194318 524532 194324 524544
rect 177080 524504 194324 524532
rect 177080 524492 177086 524504
rect 194318 524492 194324 524504
rect 194376 524492 194382 524544
rect 261478 524492 261484 524544
rect 261536 524532 261542 524544
rect 278314 524532 278320 524544
rect 261536 524504 278320 524532
rect 261536 524492 261542 524504
rect 278314 524492 278320 524504
rect 278372 524492 278378 524544
rect 288986 524492 288992 524544
rect 289044 524532 289050 524544
rect 306006 524532 306012 524544
rect 289044 524504 306012 524532
rect 289044 524492 289050 524504
rect 306006 524492 306012 524504
rect 306064 524492 306070 524544
rect 317138 524492 317144 524544
rect 317196 524532 317202 524544
rect 334342 524532 334348 524544
rect 317196 524504 334348 524532
rect 317196 524492 317202 524504
rect 334342 524492 334348 524504
rect 334400 524492 334406 524544
rect 372982 524492 372988 524544
rect 373040 524532 373046 524544
rect 390002 524532 390008 524544
rect 373040 524504 390008 524532
rect 373040 524492 373046 524504
rect 390002 524492 390008 524504
rect 390060 524492 390066 524544
rect 401042 524492 401048 524544
rect 401100 524532 401106 524544
rect 418338 524532 418344 524544
rect 401100 524504 418344 524532
rect 401100 524492 401106 524504
rect 418338 524492 418344 524504
rect 418396 524492 418402 524544
rect 457438 524492 457444 524544
rect 457496 524532 457502 524544
rect 473998 524532 474004 524544
rect 457496 524504 474004 524532
rect 457496 524492 457502 524504
rect 473998 524492 474004 524504
rect 474056 524492 474062 524544
rect 15286 524424 15292 524476
rect 15344 524464 15350 524476
rect 26326 524464 26332 524476
rect 15344 524436 26332 524464
rect 15344 524424 15350 524436
rect 26326 524424 26332 524436
rect 26384 524424 26390 524476
rect 38010 524424 38016 524476
rect 38068 524464 38074 524476
rect 64598 524464 64604 524476
rect 38068 524436 64604 524464
rect 38068 524424 38074 524436
rect 64598 524424 64604 524436
rect 64656 524424 64662 524476
rect 72326 524424 72332 524476
rect 72384 524464 72390 524476
rect 93118 524464 93124 524476
rect 72384 524436 93124 524464
rect 72384 524424 72390 524436
rect 93118 524424 93124 524436
rect 93176 524424 93182 524476
rect 100018 524424 100024 524476
rect 100076 524464 100082 524476
rect 121086 524464 121092 524476
rect 100076 524436 121092 524464
rect 100076 524424 100082 524436
rect 121086 524424 121092 524436
rect 121144 524424 121150 524476
rect 156322 524424 156328 524476
rect 156380 524464 156386 524476
rect 177298 524464 177304 524476
rect 156380 524436 177304 524464
rect 156380 524424 156386 524436
rect 177298 524424 177304 524436
rect 177356 524424 177362 524476
rect 204806 524424 204812 524476
rect 204864 524464 204870 524476
rect 222194 524464 222200 524476
rect 204864 524436 222200 524464
rect 204864 524424 204870 524436
rect 222194 524424 222200 524436
rect 222252 524424 222258 524476
rect 232958 524424 232964 524476
rect 233016 524464 233022 524476
rect 250346 524464 250352 524476
rect 233016 524436 250352 524464
rect 233016 524424 233022 524436
rect 250346 524424 250352 524436
rect 250404 524424 250410 524476
rect 268010 524424 268016 524476
rect 268068 524464 268074 524476
rect 289078 524464 289084 524476
rect 268068 524436 289084 524464
rect 268068 524424 268074 524436
rect 289078 524424 289084 524436
rect 289136 524424 289142 524476
rect 317046 524424 317052 524476
rect 317104 524464 317110 524476
rect 344646 524464 344652 524476
rect 317104 524436 344652 524464
rect 317104 524424 317110 524436
rect 344646 524424 344652 524436
rect 344704 524424 344710 524476
rect 352006 524424 352012 524476
rect 352064 524464 352070 524476
rect 373258 524464 373264 524476
rect 352064 524436 373264 524464
rect 352064 524424 352070 524436
rect 373258 524424 373264 524436
rect 373316 524424 373322 524476
rect 380342 524424 380348 524476
rect 380400 524464 380406 524476
rect 401134 524464 401140 524476
rect 380400 524436 401140 524464
rect 380400 524424 380406 524436
rect 401134 524424 401140 524436
rect 401192 524424 401198 524476
rect 429838 524424 429844 524476
rect 429896 524464 429902 524476
rect 456610 524464 456616 524476
rect 429896 524436 456616 524464
rect 429896 524424 429902 524436
rect 456610 524424 456616 524436
rect 456668 524424 456674 524476
rect 484854 524424 484860 524476
rect 484912 524464 484918 524476
rect 502334 524464 502340 524476
rect 484912 524436 502340 524464
rect 484912 524424 484918 524436
rect 502334 524424 502340 524436
rect 502392 524424 502398 524476
rect 514478 524424 514484 524476
rect 514536 524464 514542 524476
rect 530302 524464 530308 524476
rect 514536 524436 530308 524464
rect 514536 524424 514542 524436
rect 530302 524424 530308 524436
rect 530360 524424 530366 524476
rect 36722 522248 36728 522300
rect 36780 522288 36786 522300
rect 37090 522288 37096 522300
rect 36780 522260 37096 522288
rect 36780 522248 36786 522260
rect 37090 522248 37096 522260
rect 37148 522248 37154 522300
rect 120718 522248 120724 522300
rect 120776 522288 120782 522300
rect 120994 522288 121000 522300
rect 120776 522260 121000 522288
rect 120776 522248 120782 522260
rect 120994 522248 121000 522260
rect 121052 522248 121058 522300
rect 204714 522248 204720 522300
rect 204772 522288 204778 522300
rect 204990 522288 204996 522300
rect 204772 522260 204996 522288
rect 204772 522248 204778 522260
rect 204990 522248 204996 522260
rect 205048 522248 205054 522300
rect 512730 522248 512736 522300
rect 512788 522288 512794 522300
rect 514478 522288 514484 522300
rect 512788 522260 514484 522288
rect 512788 522248 512794 522260
rect 514478 522248 514484 522260
rect 514536 522248 514542 522300
rect 568850 522248 568856 522300
rect 568908 522248 568914 522300
rect 120810 522180 120816 522232
rect 120868 522220 120874 522232
rect 121086 522220 121092 522232
rect 120868 522192 121092 522220
rect 120868 522180 120874 522192
rect 121086 522180 121092 522192
rect 121144 522180 121150 522232
rect 400858 522180 400864 522232
rect 400916 522220 400922 522232
rect 401134 522220 401140 522232
rect 400916 522192 401140 522220
rect 400916 522180 400922 522192
rect 401134 522180 401140 522192
rect 401192 522180 401198 522232
rect 568868 522096 568896 522248
rect 568850 522044 568856 522096
rect 568908 522044 568914 522096
rect 176838 521976 176844 522028
rect 176896 522016 176902 522028
rect 177022 522016 177028 522028
rect 176896 521988 177028 522016
rect 176896 521976 176902 521988
rect 177022 521976 177028 521988
rect 177080 521976 177086 522028
rect 316770 521704 316776 521756
rect 316828 521744 316834 521756
rect 317138 521744 317144 521756
rect 316828 521716 317144 521744
rect 316828 521704 316834 521716
rect 317138 521704 317144 521716
rect 317196 521704 317202 521756
rect 372798 521704 372804 521756
rect 372856 521744 372862 521756
rect 372982 521744 372988 521756
rect 372856 521716 372988 521744
rect 372856 521704 372862 521716
rect 372982 521704 372988 521716
rect 373040 521704 373046 521756
rect 400766 521704 400772 521756
rect 400824 521744 400830 521756
rect 401042 521744 401048 521756
rect 400824 521716 401048 521744
rect 400824 521704 400830 521716
rect 401042 521704 401048 521716
rect 401100 521704 401106 521756
rect 232774 521636 232780 521688
rect 232832 521676 232838 521688
rect 232958 521676 232964 521688
rect 232832 521648 232964 521676
rect 232832 521636 232838 521648
rect 232958 521636 232964 521648
rect 233016 521636 233022 521688
rect 316862 521636 316868 521688
rect 316920 521676 316926 521688
rect 317046 521676 317052 521688
rect 316920 521648 317052 521676
rect 316920 521636 316926 521648
rect 317046 521636 317052 521648
rect 317104 521636 317110 521688
rect 288894 519664 288900 519716
rect 288952 519664 288958 519716
rect 288912 519512 288940 519664
rect 288894 519460 288900 519512
rect 288952 519460 288958 519512
rect 154482 518848 154488 518900
rect 154540 518888 154546 518900
rect 155862 518888 155868 518900
rect 154540 518860 155868 518888
rect 154540 518848 154546 518860
rect 155862 518848 155868 518860
rect 155920 518848 155926 518900
rect 462222 518848 462228 518900
rect 462280 518888 462286 518900
rect 463878 518888 463884 518900
rect 462280 518860 463884 518888
rect 462280 518848 462286 518860
rect 463878 518848 463884 518860
rect 463936 518848 463942 518900
rect 92750 507152 92756 507204
rect 92808 507192 92814 507204
rect 92934 507192 92940 507204
rect 92808 507164 92940 507192
rect 92808 507152 92814 507164
rect 92934 507152 92940 507164
rect 92992 507152 92998 507204
rect 204898 505928 204904 505980
rect 204956 505968 204962 505980
rect 211706 505968 211712 505980
rect 204956 505940 211712 505968
rect 204956 505928 204962 505940
rect 211706 505928 211712 505940
rect 211764 505928 211770 505980
rect 93118 505724 93124 505776
rect 93176 505764 93182 505776
rect 99742 505764 99748 505776
rect 93176 505736 99748 505764
rect 93176 505724 93182 505736
rect 99742 505724 99748 505736
rect 99800 505724 99806 505776
rect 120810 505724 120816 505776
rect 120868 505764 120874 505776
rect 127710 505764 127716 505776
rect 120868 505736 127716 505764
rect 120868 505724 120874 505736
rect 127710 505724 127716 505736
rect 127768 505724 127774 505776
rect 177298 505724 177304 505776
rect 177356 505764 177362 505776
rect 183646 505764 183652 505776
rect 177356 505736 183652 505764
rect 177356 505724 177362 505736
rect 183646 505724 183652 505736
rect 183704 505724 183710 505776
rect 373258 505724 373264 505776
rect 373316 505764 373322 505776
rect 379698 505764 379704 505776
rect 373316 505736 379704 505764
rect 373316 505724 373322 505736
rect 379698 505724 379704 505736
rect 379756 505724 379762 505776
rect 400858 505724 400864 505776
rect 400916 505764 400922 505776
rect 407758 505764 407764 505776
rect 400916 505736 407764 505764
rect 400916 505724 400922 505736
rect 407758 505724 407764 505736
rect 407816 505724 407822 505776
rect 289078 505588 289084 505640
rect 289136 505628 289142 505640
rect 295702 505628 295708 505640
rect 289136 505600 295708 505628
rect 289136 505588 289142 505600
rect 295702 505588 295708 505600
rect 295760 505588 295766 505640
rect 485038 505520 485044 505572
rect 485096 505560 485102 505572
rect 491662 505560 491668 505572
rect 485096 505532 491668 505560
rect 485096 505520 485102 505532
rect 491662 505520 491668 505532
rect 491720 505520 491726 505572
rect 64874 503208 64880 503260
rect 64932 503248 64938 503260
rect 65886 503248 65892 503260
rect 64932 503220 65892 503248
rect 64932 503208 64938 503220
rect 65886 503208 65892 503220
rect 65944 503208 65950 503260
rect 484762 502800 484768 502852
rect 484820 502840 484826 502852
rect 484946 502840 484952 502852
rect 484820 502812 484952 502840
rect 484820 502800 484826 502812
rect 484946 502800 484952 502812
rect 485004 502800 485010 502852
rect 547874 502664 547880 502716
rect 547932 502704 547938 502716
rect 548150 502704 548156 502716
rect 547932 502676 548156 502704
rect 547932 502664 547938 502676
rect 548150 502664 548156 502676
rect 548208 502664 548214 502716
rect 15378 500896 15384 500948
rect 15436 500936 15442 500948
rect 43990 500936 43996 500948
rect 15436 500908 43996 500936
rect 15436 500896 15442 500908
rect 43990 500896 43996 500908
rect 44048 500896 44054 500948
rect 138290 500896 138296 500948
rect 138348 500936 138354 500948
rect 176838 500936 176844 500948
rect 138348 500908 176844 500936
rect 138348 500896 138354 500908
rect 176838 500896 176844 500908
rect 176896 500896 176902 500948
rect 194318 500896 194324 500948
rect 194376 500936 194382 500948
rect 232866 500936 232872 500948
rect 194376 500908 232872 500936
rect 194376 500896 194382 500908
rect 232866 500896 232872 500908
rect 232924 500896 232930 500948
rect 238846 500896 238852 500948
rect 238904 500936 238910 500948
rect 238904 500908 248414 500936
rect 238904 500896 238910 500908
rect 26326 500828 26332 500880
rect 26384 500868 26390 500880
rect 38010 500868 38016 500880
rect 26384 500840 38016 500868
rect 26384 500828 26390 500840
rect 38010 500828 38016 500840
rect 38068 500828 38074 500880
rect 42886 500828 42892 500880
rect 42944 500868 42950 500880
rect 71774 500868 71780 500880
rect 42944 500840 71780 500868
rect 42944 500828 42950 500840
rect 71774 500828 71780 500840
rect 71832 500828 71838 500880
rect 110322 500828 110328 500880
rect 110380 500868 110386 500880
rect 148778 500868 148784 500880
rect 110380 500840 148784 500868
rect 110380 500828 110386 500840
rect 148778 500828 148784 500840
rect 148836 500828 148842 500880
rect 166626 500828 166632 500880
rect 166684 500868 166690 500880
rect 204990 500868 204996 500880
rect 166684 500840 204996 500868
rect 166684 500828 166690 500840
rect 204990 500828 204996 500840
rect 205048 500828 205054 500880
rect 211246 500828 211252 500880
rect 211304 500868 211310 500880
rect 240042 500868 240048 500880
rect 211304 500840 240048 500868
rect 211304 500828 211310 500840
rect 240042 500828 240048 500840
rect 240100 500828 240106 500880
rect 248386 500868 248414 500908
rect 295426 500896 295432 500948
rect 295484 500936 295490 500948
rect 324038 500936 324044 500948
rect 295484 500908 324044 500936
rect 295484 500896 295490 500908
rect 324038 500896 324044 500908
rect 324096 500896 324102 500948
rect 334342 500896 334348 500948
rect 334400 500936 334406 500948
rect 372890 500936 372896 500948
rect 334400 500908 372896 500936
rect 334400 500896 334406 500908
rect 372890 500896 372896 500908
rect 372948 500896 372954 500948
rect 390462 500896 390468 500948
rect 390520 500936 390526 500948
rect 428734 500936 428740 500948
rect 390520 500908 428740 500936
rect 390520 500896 390526 500908
rect 428734 500896 428740 500908
rect 428792 500896 428798 500948
rect 434806 500896 434812 500948
rect 434864 500936 434870 500948
rect 434864 500908 441614 500936
rect 434864 500896 434870 500908
rect 268010 500868 268016 500880
rect 248386 500840 268016 500868
rect 268010 500828 268016 500840
rect 268068 500828 268074 500880
rect 278314 500828 278320 500880
rect 278372 500868 278378 500880
rect 316954 500868 316960 500880
rect 278372 500840 316960 500868
rect 278372 500828 278378 500840
rect 316954 500828 316960 500840
rect 317012 500828 317018 500880
rect 323026 500828 323032 500880
rect 323084 500868 323090 500880
rect 352006 500868 352012 500880
rect 323084 500840 352012 500868
rect 323084 500828 323090 500840
rect 352006 500828 352012 500840
rect 352064 500828 352070 500880
rect 362310 500828 362316 500880
rect 362368 500868 362374 500880
rect 400950 500868 400956 500880
rect 362368 500840 400956 500868
rect 362368 500828 362374 500840
rect 400950 500828 400956 500840
rect 401008 500828 401014 500880
rect 407206 500828 407212 500880
rect 407264 500868 407270 500880
rect 436002 500868 436008 500880
rect 407264 500840 436008 500868
rect 407264 500828 407270 500840
rect 436002 500828 436008 500840
rect 436060 500828 436066 500880
rect 441586 500868 441614 500908
rect 491386 500896 491392 500948
rect 491444 500936 491450 500948
rect 519998 500936 520004 500948
rect 491444 500908 520004 500936
rect 491444 500896 491450 500908
rect 519998 500896 520004 500908
rect 520056 500896 520062 500948
rect 530302 500896 530308 500948
rect 530360 500936 530366 500948
rect 568850 500936 568856 500948
rect 530360 500908 568856 500936
rect 530360 500896 530366 500908
rect 568850 500896 568856 500908
rect 568908 500896 568914 500948
rect 463694 500868 463700 500880
rect 441586 500840 463700 500868
rect 463694 500828 463700 500840
rect 463752 500828 463758 500880
rect 474642 500828 474648 500880
rect 474700 500868 474706 500880
rect 512822 500868 512828 500880
rect 474700 500840 512828 500868
rect 474700 500828 474706 500840
rect 512822 500828 512828 500840
rect 512880 500828 512886 500880
rect 548150 500828 548156 500880
rect 548208 500868 548214 500880
rect 557994 500868 558000 500880
rect 548208 500840 558000 500868
rect 548208 500828 548214 500840
rect 557994 500828 558000 500840
rect 558052 500828 558058 500880
rect 82630 500760 82636 500812
rect 82688 500800 82694 500812
rect 120902 500800 120908 500812
rect 82688 500772 120908 500800
rect 82688 500760 82694 500772
rect 120902 500760 120908 500772
rect 120960 500760 120966 500812
rect 127066 500760 127072 500812
rect 127124 500800 127130 500812
rect 156046 500800 156052 500812
rect 127124 500772 156052 500800
rect 127124 500760 127130 500772
rect 156046 500760 156052 500772
rect 156104 500760 156110 500812
rect 250346 500760 250352 500812
rect 250404 500800 250410 500812
rect 288894 500800 288900 500812
rect 250404 500772 288900 500800
rect 250404 500760 250410 500772
rect 288894 500760 288900 500772
rect 288952 500760 288958 500812
rect 306282 500760 306288 500812
rect 306340 500800 306346 500812
rect 316862 500800 316868 500812
rect 306340 500772 316868 500800
rect 306340 500760 306346 500772
rect 316862 500760 316868 500772
rect 316920 500760 316926 500812
rect 418338 500760 418344 500812
rect 418396 500800 418402 500812
rect 429838 500800 429844 500812
rect 418396 500772 429844 500800
rect 418396 500760 418402 500772
rect 429838 500760 429844 500772
rect 429896 500760 429902 500812
rect 446306 500760 446312 500812
rect 446364 500800 446370 500812
rect 484946 500800 484952 500812
rect 446364 500772 484952 500800
rect 446364 500760 446370 500772
rect 484946 500760 484952 500772
rect 485004 500760 485010 500812
rect 502334 500760 502340 500812
rect 502392 500800 502398 500812
rect 540790 500800 540796 500812
rect 502392 500772 540796 500800
rect 502392 500760 502398 500772
rect 540790 500760 540796 500772
rect 540848 500760 540854 500812
rect 54294 500692 54300 500744
rect 54352 500732 54358 500744
rect 92934 500732 92940 500744
rect 54352 500704 92940 500732
rect 54352 500692 54358 500704
rect 92934 500692 92940 500704
rect 92992 500692 92998 500744
rect 518986 500692 518992 500744
rect 519044 500732 519050 500744
rect 547874 500732 547880 500744
rect 519044 500704 547880 500732
rect 519044 500692 519050 500704
rect 547874 500692 547880 500704
rect 547932 500692 547938 500744
rect 26602 498788 26608 498840
rect 26660 498828 26666 498840
rect 36814 498828 36820 498840
rect 26660 498800 36820 498828
rect 26660 498788 26666 498800
rect 36814 498788 36820 498800
rect 36872 498788 36878 498840
rect 15930 498312 15936 498364
rect 15988 498352 15994 498364
rect 54294 498352 54300 498364
rect 15988 498324 54300 498352
rect 15988 498312 15994 498324
rect 54294 498312 54300 498324
rect 54352 498312 54358 498364
rect 65886 498244 65892 498296
rect 65944 498284 65950 498296
rect 82630 498284 82636 498296
rect 65944 498256 82636 498284
rect 65944 498244 65950 498256
rect 82630 498244 82636 498256
rect 82688 498244 82694 498296
rect 99374 498244 99380 498296
rect 99432 498284 99438 498296
rect 138290 498284 138296 498296
rect 99432 498256 138296 498284
rect 99432 498244 99438 498256
rect 138290 498244 138296 498256
rect 138348 498244 138354 498296
rect 149698 498244 149704 498296
rect 149756 498284 149762 498296
rect 156322 498284 156328 498296
rect 149756 498256 156328 498284
rect 149756 498244 149762 498256
rect 156322 498244 156328 498256
rect 156380 498244 156386 498296
rect 211154 498244 211160 498296
rect 211212 498284 211218 498296
rect 250622 498284 250628 498296
rect 211212 498256 250628 498284
rect 211212 498244 211218 498256
rect 250622 498244 250628 498256
rect 250680 498244 250686 498296
rect 267734 498244 267740 498296
rect 267792 498284 267798 498296
rect 306466 498284 306472 498296
rect 267792 498256 306472 498284
rect 267792 498244 267798 498256
rect 306466 498244 306472 498256
rect 306524 498244 306530 498296
rect 318058 498244 318064 498296
rect 318116 498284 318122 498296
rect 324314 498284 324320 498296
rect 318116 498256 324320 498284
rect 318116 498244 318122 498256
rect 324314 498244 324320 498256
rect 324372 498244 324378 498296
rect 345842 498244 345848 498296
rect 345900 498284 345906 498296
rect 362310 498284 362316 498296
rect 345900 498256 362316 498284
rect 345900 498244 345906 498256
rect 362310 498244 362316 498256
rect 362368 498244 362374 498296
rect 407114 498244 407120 498296
rect 407172 498284 407178 498296
rect 446306 498284 446312 498296
rect 407172 498256 446312 498284
rect 407172 498244 407178 498256
rect 446306 498244 446312 498256
rect 446364 498244 446370 498296
rect 457438 498244 457444 498296
rect 457496 498284 457502 498296
rect 474642 498284 474648 498296
rect 457496 498256 474648 498284
rect 457496 498244 457502 498256
rect 474642 498244 474648 498256
rect 474700 498244 474706 498296
rect 491294 498244 491300 498296
rect 491352 498284 491358 498296
rect 530302 498284 530308 498296
rect 491352 498256 530308 498284
rect 491352 498244 491358 498256
rect 530302 498244 530308 498256
rect 530360 498244 530366 498296
rect 38102 498176 38108 498228
rect 38160 498216 38166 498228
rect 44174 498216 44180 498228
rect 38160 498188 44180 498216
rect 38160 498176 38166 498188
rect 44174 498176 44180 498188
rect 44232 498176 44238 498228
rect 71774 498176 71780 498228
rect 71832 498216 71838 498228
rect 110598 498216 110604 498228
rect 71832 498188 110604 498216
rect 71832 498176 71838 498188
rect 110598 498176 110604 498188
rect 110656 498176 110662 498228
rect 149882 498176 149888 498228
rect 149940 498216 149946 498228
rect 166626 498216 166632 498228
rect 149940 498188 166632 498216
rect 149940 498176 149946 498188
rect 166626 498176 166632 498188
rect 166684 498176 166690 498228
rect 183554 498176 183560 498228
rect 183612 498216 183618 498228
rect 222286 498216 222292 498228
rect 183612 498188 222292 498216
rect 183612 498176 183618 498188
rect 222286 498176 222292 498188
rect 222344 498176 222350 498228
rect 234062 498176 234068 498228
rect 234120 498216 234126 498228
rect 240318 498216 240324 498228
rect 234120 498188 240324 498216
rect 234120 498176 234126 498188
rect 240318 498176 240324 498188
rect 240376 498176 240382 498228
rect 261478 498176 261484 498228
rect 261536 498216 261542 498228
rect 278590 498216 278596 498228
rect 261536 498188 278596 498216
rect 261536 498176 261542 498188
rect 278590 498176 278596 498188
rect 278648 498176 278654 498228
rect 295334 498176 295340 498228
rect 295392 498216 295398 498228
rect 334618 498216 334624 498228
rect 295392 498188 334624 498216
rect 295392 498176 295398 498188
rect 334618 498176 334624 498188
rect 334676 498176 334682 498228
rect 345750 498176 345756 498228
rect 345808 498216 345814 498228
rect 352006 498216 352012 498228
rect 345808 498188 352012 498216
rect 345808 498176 345814 498188
rect 352006 498176 352012 498188
rect 352064 498176 352070 498228
rect 379514 498176 379520 498228
rect 379572 498216 379578 498228
rect 418614 498216 418620 498228
rect 379572 498188 418620 498216
rect 379572 498176 379578 498188
rect 418614 498176 418620 498188
rect 418672 498176 418678 498228
rect 429930 498176 429936 498228
rect 429988 498216 429994 498228
rect 436094 498216 436100 498228
rect 429988 498188 436100 498216
rect 429988 498176 429994 498188
rect 436094 498176 436100 498188
rect 436152 498176 436158 498228
rect 463694 498176 463700 498228
rect 463752 498216 463758 498228
rect 502610 498216 502616 498228
rect 463752 498188 502616 498216
rect 463752 498176 463758 498188
rect 502610 498176 502616 498188
rect 502668 498176 502674 498228
rect 514018 498176 514024 498228
rect 514076 498216 514082 498228
rect 520274 498216 520280 498228
rect 514076 498188 520280 498216
rect 514076 498176 514082 498188
rect 520274 498176 520280 498188
rect 520332 498176 520338 498228
rect 541618 498176 541624 498228
rect 541676 498216 541682 498228
rect 558638 498216 558644 498228
rect 541676 498188 558644 498216
rect 541676 498176 541682 498188
rect 558638 498176 558644 498188
rect 558696 498176 558702 498228
rect 15286 497360 15292 497412
rect 15344 497400 15350 497412
rect 16022 497400 16028 497412
rect 15344 497372 16028 497400
rect 15344 497360 15350 497372
rect 16022 497360 16028 497372
rect 16080 497360 16086 497412
rect 205082 495320 205088 495372
rect 205140 495320 205146 495372
rect 205100 495168 205128 495320
rect 429102 495184 429108 495236
rect 429160 495224 429166 495236
rect 429838 495224 429844 495236
rect 429160 495196 429844 495224
rect 429160 495184 429166 495196
rect 429838 495184 429844 495196
rect 429896 495184 429902 495236
rect 205082 495116 205088 495168
rect 205140 495116 205146 495168
rect 37274 492532 37280 492584
rect 37332 492572 37338 492584
rect 38010 492572 38016 492584
rect 37332 492544 38016 492572
rect 37332 492532 37338 492544
rect 38010 492532 38016 492544
rect 38068 492532 38074 492584
rect 149238 492532 149244 492584
rect 149296 492572 149302 492584
rect 149790 492572 149796 492584
rect 149296 492544 149796 492572
rect 149296 492532 149302 492544
rect 149790 492532 149796 492544
rect 149848 492532 149854 492584
rect 233234 492532 233240 492584
rect 233292 492572 233298 492584
rect 233970 492572 233976 492584
rect 233292 492544 233976 492572
rect 233292 492532 233298 492544
rect 233970 492532 233976 492544
rect 234028 492532 234034 492584
rect 463694 485052 463700 485104
rect 463752 485092 463758 485104
rect 463970 485092 463976 485104
rect 463752 485064 463976 485092
rect 463752 485052 463758 485064
rect 463970 485052 463976 485064
rect 464028 485052 464034 485104
rect 99374 477640 99380 477692
rect 99432 477680 99438 477692
rect 99926 477680 99932 477692
rect 99432 477652 99932 477680
rect 99432 477640 99438 477652
rect 99926 477640 99932 477652
rect 99984 477640 99990 477692
rect 183554 477640 183560 477692
rect 183612 477680 183618 477692
rect 184014 477680 184020 477692
rect 183612 477652 184020 477680
rect 183612 477640 183618 477652
rect 184014 477640 184020 477652
rect 184072 477640 184078 477692
rect 211154 477640 211160 477692
rect 211212 477680 211218 477692
rect 211982 477680 211988 477692
rect 211212 477652 211988 477680
rect 211212 477640 211218 477652
rect 211982 477640 211988 477652
rect 212040 477640 212046 477692
rect 267734 477640 267740 477692
rect 267792 477680 267798 477692
rect 268010 477680 268016 477692
rect 267792 477652 268016 477680
rect 267792 477640 267798 477652
rect 268010 477640 268016 477652
rect 268068 477640 268074 477692
rect 295334 477640 295340 477692
rect 295392 477680 295398 477692
rect 295978 477680 295984 477692
rect 295392 477652 295984 477680
rect 295392 477640 295398 477652
rect 295978 477640 295984 477652
rect 296036 477640 296042 477692
rect 379514 477640 379520 477692
rect 379572 477680 379578 477692
rect 379974 477680 379980 477692
rect 379572 477652 379980 477680
rect 379572 477640 379578 477652
rect 379974 477640 379980 477652
rect 380032 477640 380038 477692
rect 407114 477640 407120 477692
rect 407172 477680 407178 477692
rect 407942 477680 407948 477692
rect 407172 477652 407948 477680
rect 407172 477640 407178 477652
rect 407942 477640 407948 477652
rect 408000 477640 408006 477692
rect 491294 477640 491300 477692
rect 491352 477680 491358 477692
rect 492030 477680 492036 477692
rect 491352 477652 492036 477680
rect 491352 477640 491358 477652
rect 492030 477640 492036 477652
rect 492088 477640 492094 477692
rect 71774 475668 71780 475720
rect 71832 475708 71838 475720
rect 72050 475708 72056 475720
rect 71832 475680 72056 475708
rect 71832 475668 71838 475680
rect 72050 475668 72056 475680
rect 72108 475668 72114 475720
rect 15194 473288 15200 473340
rect 15252 473328 15258 473340
rect 36906 473328 36912 473340
rect 15252 473300 36912 473328
rect 15252 473288 15258 473300
rect 36906 473288 36912 473300
rect 36964 473288 36970 473340
rect 38010 473288 38016 473340
rect 38068 473328 38074 473340
rect 64874 473328 64880 473340
rect 38068 473300 64880 473328
rect 38068 473288 38074 473300
rect 64874 473288 64880 473300
rect 64932 473288 64938 473340
rect 65058 473288 65064 473340
rect 65116 473328 65122 473340
rect 92934 473328 92940 473340
rect 65116 473300 92940 473328
rect 65116 473288 65122 473300
rect 92934 473288 92940 473300
rect 92992 473288 92998 473340
rect 93026 473288 93032 473340
rect 93084 473328 93090 473340
rect 120902 473328 120908 473340
rect 93084 473300 120908 473328
rect 93084 473288 93090 473300
rect 120902 473288 120908 473300
rect 120960 473288 120966 473340
rect 121086 473288 121092 473340
rect 121144 473328 121150 473340
rect 148594 473328 148600 473340
rect 121144 473300 148600 473328
rect 121144 473288 121150 473300
rect 148594 473288 148600 473300
rect 148652 473288 148658 473340
rect 149790 473288 149796 473340
rect 149848 473328 149854 473340
rect 176930 473328 176936 473340
rect 149848 473300 176936 473328
rect 149848 473288 149854 473300
rect 176930 473288 176936 473300
rect 176988 473288 176994 473340
rect 177022 473288 177028 473340
rect 177080 473328 177086 473340
rect 204898 473328 204904 473340
rect 177080 473300 204904 473328
rect 177080 473288 177086 473300
rect 204898 473288 204904 473300
rect 204956 473288 204962 473340
rect 205174 473288 205180 473340
rect 205232 473328 205238 473340
rect 232590 473328 232596 473340
rect 205232 473300 232596 473328
rect 205232 473288 205238 473300
rect 232590 473288 232596 473300
rect 232648 473288 232654 473340
rect 233970 473288 233976 473340
rect 234028 473328 234034 473340
rect 260926 473328 260932 473340
rect 234028 473300 260932 473328
rect 234028 473288 234034 473300
rect 260926 473288 260932 473300
rect 260984 473288 260990 473340
rect 261018 473288 261024 473340
rect 261076 473328 261082 473340
rect 288894 473328 288900 473340
rect 261076 473300 288900 473328
rect 261076 473288 261082 473300
rect 288894 473288 288900 473300
rect 288952 473288 288958 473340
rect 289078 473288 289084 473340
rect 289136 473328 289142 473340
rect 316586 473328 316592 473340
rect 289136 473300 316592 473328
rect 289136 473288 289142 473300
rect 316586 473288 316592 473300
rect 316644 473288 316650 473340
rect 317046 473288 317052 473340
rect 317104 473328 317110 473340
rect 344922 473328 344928 473340
rect 317104 473300 344928 473328
rect 317104 473288 317110 473300
rect 344922 473288 344928 473300
rect 344980 473288 344986 473340
rect 345658 473288 345664 473340
rect 345716 473328 345722 473340
rect 372614 473328 372620 473340
rect 345716 473300 372620 473328
rect 345716 473288 345722 473300
rect 372614 473288 372620 473300
rect 372672 473288 372678 473340
rect 373074 473288 373080 473340
rect 373132 473328 373138 473340
rect 400950 473328 400956 473340
rect 373132 473300 400956 473328
rect 373132 473288 373138 473300
rect 400950 473288 400956 473300
rect 401008 473288 401014 473340
rect 401042 473288 401048 473340
rect 401100 473328 401106 473340
rect 428918 473328 428924 473340
rect 401100 473300 428924 473328
rect 401100 473288 401106 473300
rect 428918 473288 428924 473300
rect 428976 473288 428982 473340
rect 429838 473288 429844 473340
rect 429896 473328 429902 473340
rect 456794 473328 456800 473340
rect 429896 473300 456800 473328
rect 429896 473288 429902 473300
rect 456794 473288 456800 473300
rect 456852 473288 456858 473340
rect 457070 473288 457076 473340
rect 457128 473328 457134 473340
rect 484946 473328 484952 473340
rect 457128 473300 484952 473328
rect 457128 473288 457134 473300
rect 484946 473288 484952 473300
rect 485004 473288 485010 473340
rect 485038 473288 485044 473340
rect 485096 473328 485102 473340
rect 512914 473328 512920 473340
rect 485096 473300 512920 473328
rect 485096 473288 485102 473300
rect 512914 473288 512920 473300
rect 512972 473288 512978 473340
rect 513098 473288 513104 473340
rect 513156 473328 513162 473340
rect 540606 473328 540612 473340
rect 513156 473300 540612 473328
rect 513156 473288 513162 473300
rect 540606 473288 540612 473300
rect 540664 473288 540670 473340
rect 541066 473288 541072 473340
rect 541124 473328 541130 473340
rect 568942 473328 568948 473340
rect 541124 473300 568948 473328
rect 541124 473288 541130 473300
rect 568942 473288 568948 473300
rect 569000 473288 569006 473340
rect 26602 473220 26608 473272
rect 26660 473260 26666 473272
rect 38102 473260 38108 473272
rect 26660 473232 38108 473260
rect 26660 473220 26666 473232
rect 38102 473220 38108 473232
rect 38160 473220 38166 473272
rect 44634 473220 44640 473272
rect 44692 473260 44698 473272
rect 65886 473260 65892 473272
rect 44692 473232 65892 473260
rect 44692 473220 44698 473232
rect 65886 473220 65892 473232
rect 65944 473220 65950 473272
rect 82630 473220 82636 473272
rect 82688 473260 82694 473272
rect 99466 473260 99472 473272
rect 82688 473232 99472 473260
rect 82688 473220 82694 473232
rect 99466 473220 99472 473232
rect 99524 473220 99530 473272
rect 128630 473220 128636 473272
rect 128688 473260 128694 473272
rect 149882 473260 149888 473272
rect 128688 473232 149888 473260
rect 128688 473220 128694 473232
rect 149882 473220 149888 473232
rect 149940 473220 149946 473272
rect 166626 473220 166632 473272
rect 166684 473260 166690 473272
rect 183646 473260 183652 473272
rect 166684 473232 183652 473260
rect 166684 473220 166690 473232
rect 183646 473220 183652 473232
rect 183704 473220 183710 473272
rect 194594 473220 194600 473272
rect 194652 473260 194658 473272
rect 211246 473260 211252 473272
rect 194652 473232 211252 473260
rect 194652 473220 194658 473232
rect 211246 473220 211252 473232
rect 211304 473220 211310 473272
rect 222930 473220 222936 473272
rect 222988 473260 222994 473272
rect 234062 473260 234068 473272
rect 222988 473232 234068 473260
rect 222988 473220 222994 473232
rect 234062 473220 234068 473232
rect 234120 473220 234126 473272
rect 240318 473220 240324 473272
rect 240376 473260 240382 473272
rect 261478 473260 261484 473272
rect 240376 473232 261484 473260
rect 240376 473220 240382 473232
rect 261478 473220 261484 473232
rect 261536 473220 261542 473272
rect 278590 473220 278596 473272
rect 278648 473260 278654 473272
rect 295426 473260 295432 473272
rect 278648 473232 295432 473260
rect 278648 473220 278654 473232
rect 295426 473220 295432 473232
rect 295484 473220 295490 473272
rect 306926 473220 306932 473272
rect 306984 473260 306990 473272
rect 318058 473260 318064 473272
rect 306984 473232 318064 473260
rect 306984 473220 306990 473232
rect 318058 473220 318064 473232
rect 318116 473220 318122 473272
rect 324314 473220 324320 473272
rect 324372 473260 324378 473272
rect 345842 473260 345848 473272
rect 324372 473232 345848 473260
rect 324372 473220 324378 473232
rect 345842 473220 345848 473232
rect 345900 473220 345906 473272
rect 362862 473220 362868 473272
rect 362920 473260 362926 473272
rect 379606 473260 379612 473272
rect 362920 473232 379612 473260
rect 362920 473220 362926 473232
rect 379606 473220 379612 473232
rect 379664 473220 379670 473272
rect 390646 473220 390652 473272
rect 390704 473260 390710 473272
rect 407206 473260 407212 473272
rect 390704 473232 407212 473260
rect 390704 473220 390710 473232
rect 407206 473220 407212 473232
rect 407264 473220 407270 473272
rect 418614 473220 418620 473272
rect 418672 473260 418678 473272
rect 429930 473260 429936 473272
rect 418672 473232 429936 473260
rect 418672 473220 418678 473232
rect 429930 473220 429936 473232
rect 429988 473220 429994 473272
rect 436646 473220 436652 473272
rect 436704 473260 436710 473272
rect 457438 473260 457444 473272
rect 436704 473232 457444 473260
rect 436704 473220 436710 473232
rect 457438 473220 457444 473232
rect 457496 473220 457502 473272
rect 474642 473220 474648 473272
rect 474700 473260 474706 473272
rect 491386 473260 491392 473272
rect 474700 473232 491392 473260
rect 474700 473220 474706 473232
rect 491386 473220 491392 473232
rect 491444 473220 491450 473272
rect 502610 473220 502616 473272
rect 502668 473260 502674 473272
rect 514018 473260 514024 473272
rect 502668 473232 514024 473260
rect 502668 473220 502674 473232
rect 514018 473220 514024 473232
rect 514076 473220 514082 473272
rect 520642 473220 520648 473272
rect 520700 473260 520706 473272
rect 541618 473260 541624 473272
rect 520700 473232 541624 473260
rect 520700 473220 520706 473232
rect 541618 473220 541624 473232
rect 541676 473220 541682 473272
rect 54938 473152 54944 473204
rect 54996 473192 55002 473204
rect 71866 473192 71872 473204
rect 54996 473164 71872 473192
rect 54996 473152 55002 473164
rect 71866 473152 71872 473164
rect 71924 473152 71930 473204
rect 138934 473152 138940 473204
rect 138992 473192 138998 473204
rect 149698 473192 149704 473204
rect 138992 473164 149704 473192
rect 138992 473152 138998 473164
rect 149698 473152 149704 473164
rect 149756 473152 149762 473204
rect 250622 473152 250628 473204
rect 250680 473192 250686 473204
rect 267918 473192 267924 473204
rect 250680 473164 267924 473192
rect 250680 473152 250686 473164
rect 267918 473152 267924 473164
rect 267976 473152 267982 473204
rect 334618 473152 334624 473204
rect 334676 473192 334682 473204
rect 345750 473192 345756 473204
rect 334676 473164 345756 473192
rect 334676 473152 334682 473164
rect 345750 473152 345756 473164
rect 345808 473152 345814 473204
rect 446950 473152 446956 473204
rect 447008 473192 447014 473204
rect 463786 473192 463792 473204
rect 447008 473164 463792 473192
rect 447008 473152 447014 473164
rect 463786 473152 463792 473164
rect 463844 473152 463850 473204
rect 530946 473152 530952 473204
rect 531004 473192 531010 473204
rect 547966 473192 547972 473204
rect 531004 473164 547972 473192
rect 531004 473152 531010 473164
rect 547966 473152 547972 473164
rect 548024 473152 548030 473204
rect 558638 472608 558644 472660
rect 558696 472648 558702 472660
rect 568758 472648 568764 472660
rect 558696 472620 568764 472648
rect 558696 472608 558702 472620
rect 568758 472608 568764 472620
rect 568816 472608 568822 472660
rect 548334 471248 548340 471300
rect 548392 471288 548398 471300
rect 569034 471288 569040 471300
rect 548392 471260 569040 471288
rect 548392 471248 548398 471260
rect 569034 471248 569040 471260
rect 569092 471248 569098 471300
rect 100018 470772 100024 470824
rect 100076 470812 100082 470824
rect 120810 470812 120816 470824
rect 100076 470784 120816 470812
rect 100076 470772 100082 470784
rect 120810 470772 120816 470784
rect 120868 470772 120874 470824
rect 184014 470772 184020 470824
rect 184072 470812 184078 470824
rect 204898 470812 204904 470824
rect 184072 470784 204904 470812
rect 184072 470772 184078 470784
rect 204898 470772 204904 470784
rect 204956 470772 204962 470824
rect 268010 470772 268016 470824
rect 268068 470812 268074 470824
rect 289078 470812 289084 470824
rect 268068 470784 289084 470812
rect 268068 470772 268074 470784
rect 289078 470772 289084 470784
rect 289136 470772 289142 470824
rect 380342 470772 380348 470824
rect 380400 470812 380406 470824
rect 400858 470812 400864 470824
rect 380400 470784 400864 470812
rect 380400 470772 380406 470784
rect 400858 470772 400864 470784
rect 400916 470772 400922 470824
rect 464338 470772 464344 470824
rect 464396 470812 464402 470824
rect 485038 470812 485044 470824
rect 464396 470784 485044 470812
rect 464396 470772 464402 470784
rect 485038 470772 485044 470784
rect 485096 470772 485102 470824
rect 92842 470704 92848 470756
rect 92900 470744 92906 470756
rect 110322 470744 110328 470756
rect 92900 470716 110328 470744
rect 92900 470704 92906 470716
rect 110322 470704 110328 470716
rect 110380 470704 110386 470756
rect 176838 470704 176844 470756
rect 176896 470744 176902 470756
rect 194318 470744 194324 470756
rect 176896 470716 194324 470744
rect 176896 470704 176902 470716
rect 194318 470704 194324 470716
rect 194376 470704 194382 470756
rect 261570 470704 261576 470756
rect 261628 470744 261634 470756
rect 278314 470744 278320 470756
rect 261628 470716 278320 470744
rect 261628 470704 261634 470716
rect 278314 470704 278320 470716
rect 278372 470704 278378 470756
rect 372890 470704 372896 470756
rect 372948 470744 372954 470756
rect 390002 470744 390008 470756
rect 372948 470716 390008 470744
rect 372948 470704 372954 470716
rect 390002 470704 390008 470716
rect 390060 470704 390066 470756
rect 457530 470704 457536 470756
rect 457588 470744 457594 470756
rect 473998 470744 474004 470756
rect 457588 470716 474004 470744
rect 457588 470704 457594 470716
rect 473998 470704 474004 470716
rect 474056 470704 474062 470756
rect 72326 470636 72332 470688
rect 72384 470676 72390 470688
rect 93118 470676 93124 470688
rect 72384 470648 93124 470676
rect 72384 470636 72390 470648
rect 93118 470636 93124 470648
rect 93176 470636 93182 470688
rect 120718 470636 120724 470688
rect 120776 470676 120782 470688
rect 138290 470676 138296 470688
rect 120776 470648 138296 470676
rect 120776 470636 120782 470648
rect 138290 470636 138296 470648
rect 138348 470636 138354 470688
rect 156322 470636 156328 470688
rect 156380 470676 156386 470688
rect 177298 470676 177304 470688
rect 156380 470648 177304 470676
rect 156380 470636 156386 470648
rect 177298 470636 177304 470648
rect 177356 470636 177362 470688
rect 204806 470636 204812 470688
rect 204864 470676 204870 470688
rect 222286 470676 222292 470688
rect 204864 470648 222292 470676
rect 204864 470636 204870 470648
rect 222286 470636 222292 470648
rect 222344 470636 222350 470688
rect 232774 470636 232780 470688
rect 232832 470676 232838 470688
rect 250346 470676 250352 470688
rect 232832 470648 250352 470676
rect 232832 470636 232838 470648
rect 250346 470636 250352 470648
rect 250404 470636 250410 470688
rect 288894 470636 288900 470688
rect 288952 470676 288958 470688
rect 306006 470676 306012 470688
rect 288952 470648 306012 470676
rect 288952 470636 288958 470648
rect 306006 470636 306012 470648
rect 306064 470636 306070 470688
rect 316770 470636 316776 470688
rect 316828 470676 316834 470688
rect 334342 470676 334348 470688
rect 316828 470648 334348 470676
rect 316828 470636 316834 470648
rect 334342 470636 334348 470648
rect 334400 470636 334406 470688
rect 352006 470636 352012 470688
rect 352064 470676 352070 470688
rect 373258 470676 373264 470688
rect 352064 470648 373264 470676
rect 352064 470636 352070 470648
rect 373258 470636 373264 470648
rect 373316 470636 373322 470688
rect 400766 470636 400772 470688
rect 400824 470676 400830 470688
rect 418338 470676 418344 470688
rect 400824 470648 418344 470676
rect 400824 470636 400830 470648
rect 418338 470636 418344 470648
rect 418396 470636 418402 470688
rect 484854 470636 484860 470688
rect 484912 470676 484918 470688
rect 502334 470676 502340 470688
rect 484912 470648 502340 470676
rect 484912 470636 484918 470648
rect 502334 470636 502340 470648
rect 502392 470636 502398 470688
rect 512730 470636 512736 470688
rect 512788 470676 512794 470688
rect 530302 470676 530308 470688
rect 512788 470648 530308 470676
rect 512788 470636 512794 470648
rect 530302 470636 530308 470648
rect 530360 470636 530366 470688
rect 15286 470568 15292 470620
rect 15344 470608 15350 470620
rect 26326 470608 26332 470620
rect 15344 470580 26332 470608
rect 15344 470568 15350 470580
rect 26326 470568 26332 470580
rect 26384 470568 26390 470620
rect 36722 470568 36728 470620
rect 36780 470608 36786 470620
rect 54294 470608 54300 470620
rect 36780 470580 54300 470608
rect 36780 470568 36786 470580
rect 54294 470568 54300 470580
rect 54352 470568 54358 470620
rect 69658 470568 69664 470620
rect 69716 470608 69722 470620
rect 579982 470608 579988 470620
rect 69716 470580 579988 470608
rect 69716 470568 69722 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 36722 468392 36728 468444
rect 36780 468392 36786 468444
rect 120718 468392 120724 468444
rect 120776 468392 120782 468444
rect 120810 468392 120816 468444
rect 120868 468392 120874 468444
rect 232774 468392 232780 468444
rect 232832 468392 232838 468444
rect 316770 468392 316776 468444
rect 316828 468392 316834 468444
rect 400766 468392 400772 468444
rect 400824 468392 400830 468444
rect 400858 468392 400864 468444
rect 400916 468392 400922 468444
rect 512730 468392 512736 468444
rect 512788 468392 512794 468444
rect 568758 468392 568764 468444
rect 568816 468392 568822 468444
rect 36740 468240 36768 468392
rect 120736 468240 120764 468392
rect 120828 468240 120856 468392
rect 204714 468256 204720 468308
rect 204772 468296 204778 468308
rect 204990 468296 204996 468308
rect 204772 468268 204996 468296
rect 204772 468256 204778 468268
rect 204990 468256 204996 468268
rect 205048 468256 205054 468308
rect 232792 468240 232820 468392
rect 316788 468240 316816 468392
rect 400784 468240 400812 468392
rect 400876 468240 400904 468392
rect 512748 468240 512776 468392
rect 568776 468240 568804 468392
rect 36722 468188 36728 468240
rect 36780 468188 36786 468240
rect 120718 468188 120724 468240
rect 120776 468188 120782 468240
rect 120810 468188 120816 468240
rect 120868 468188 120874 468240
rect 232774 468188 232780 468240
rect 232832 468188 232838 468240
rect 316770 468188 316776 468240
rect 316828 468188 316834 468240
rect 400766 468188 400772 468240
rect 400824 468188 400830 468240
rect 400858 468188 400864 468240
rect 400916 468188 400922 468240
rect 512730 468188 512736 468240
rect 512788 468188 512794 468240
rect 568758 468188 568764 468240
rect 568816 468188 568822 468240
rect 289078 452548 289084 452600
rect 289136 452588 289142 452600
rect 295702 452588 295708 452600
rect 289136 452560 295708 452588
rect 289136 452548 289142 452560
rect 295702 452548 295708 452560
rect 295760 452548 295766 452600
rect 92750 451936 92756 451988
rect 92808 451976 92814 451988
rect 92934 451976 92940 451988
rect 92808 451948 92940 451976
rect 92808 451936 92814 451948
rect 92934 451936 92940 451948
rect 92992 451936 92998 451988
rect 93118 451868 93124 451920
rect 93176 451908 93182 451920
rect 99742 451908 99748 451920
rect 93176 451880 99748 451908
rect 93176 451868 93182 451880
rect 99742 451868 99748 451880
rect 99800 451868 99806 451920
rect 120810 451868 120816 451920
rect 120868 451908 120874 451920
rect 127710 451908 127716 451920
rect 120868 451880 127716 451908
rect 120868 451868 120874 451880
rect 127710 451868 127716 451880
rect 127768 451868 127774 451920
rect 177298 451868 177304 451920
rect 177356 451908 177362 451920
rect 183738 451908 183744 451920
rect 177356 451880 183744 451908
rect 177356 451868 177362 451880
rect 183738 451868 183744 451880
rect 183796 451868 183802 451920
rect 373258 451868 373264 451920
rect 373316 451908 373322 451920
rect 379698 451908 379704 451920
rect 373316 451880 379704 451908
rect 373316 451868 373322 451880
rect 379698 451868 379704 451880
rect 379756 451868 379762 451920
rect 400858 451868 400864 451920
rect 400916 451908 400922 451920
rect 407758 451908 407764 451920
rect 400916 451880 407764 451908
rect 400916 451868 400922 451880
rect 407758 451868 407764 451880
rect 407816 451868 407822 451920
rect 204898 451256 204904 451308
rect 204956 451296 204962 451308
rect 211706 451296 211712 451308
rect 204956 451268 211712 451296
rect 204956 451256 204962 451268
rect 211706 451256 211712 451268
rect 211764 451256 211770 451308
rect 485038 451256 485044 451308
rect 485096 451296 485102 451308
rect 491662 451296 491668 451308
rect 485096 451268 491668 451296
rect 485096 451256 485102 451268
rect 491662 451256 491668 451268
rect 491720 451256 491726 451308
rect 2774 448808 2780 448860
rect 2832 448848 2838 448860
rect 4982 448848 4988 448860
rect 2832 448820 4988 448848
rect 2832 448808 2838 448820
rect 4982 448808 4988 448820
rect 5040 448808 5046 448860
rect 176746 448808 176752 448860
rect 176804 448848 176810 448860
rect 176930 448848 176936 448860
rect 176804 448820 176936 448848
rect 176804 448808 176810 448820
rect 176930 448808 176936 448820
rect 176988 448808 176994 448860
rect 288802 448808 288808 448860
rect 288860 448848 288866 448860
rect 288986 448848 288992 448860
rect 288860 448820 288992 448848
rect 288860 448808 288866 448820
rect 288986 448808 288992 448820
rect 289044 448808 289050 448860
rect 372798 448808 372804 448860
rect 372856 448848 372862 448860
rect 372982 448848 372988 448860
rect 372856 448820 372988 448848
rect 372856 448808 372862 448820
rect 372982 448808 372988 448820
rect 373040 448808 373046 448860
rect 484762 448808 484768 448860
rect 484820 448848 484826 448860
rect 484946 448848 484952 448860
rect 484820 448820 484952 448848
rect 484820 448808 484826 448820
rect 484946 448808 484952 448820
rect 485004 448808 485010 448860
rect 547874 448400 547880 448452
rect 547932 448440 547938 448452
rect 548150 448440 548156 448452
rect 547932 448412 548156 448440
rect 547932 448400 547938 448412
rect 548150 448400 548156 448412
rect 548208 448400 548214 448452
rect 15286 448128 15292 448180
rect 15344 448168 15350 448180
rect 16114 448168 16120 448180
rect 15344 448140 16120 448168
rect 15344 448128 15350 448140
rect 16114 448128 16120 448140
rect 16172 448128 16178 448180
rect 15470 445680 15476 445732
rect 15528 445720 15534 445732
rect 43990 445720 43996 445732
rect 15528 445692 43996 445720
rect 15528 445680 15534 445692
rect 43990 445680 43996 445692
rect 44048 445680 44054 445732
rect 54294 445680 54300 445732
rect 54352 445720 54358 445732
rect 92934 445720 92940 445732
rect 54352 445692 92940 445720
rect 54352 445680 54358 445692
rect 92934 445680 92940 445692
rect 92992 445680 92998 445732
rect 110322 445680 110328 445732
rect 110380 445720 110386 445732
rect 148778 445720 148784 445732
rect 110380 445692 148784 445720
rect 110380 445680 110386 445692
rect 148778 445680 148784 445692
rect 148836 445680 148842 445732
rect 194318 445680 194324 445732
rect 194376 445720 194382 445732
rect 232866 445720 232872 445732
rect 194376 445692 232872 445720
rect 194376 445680 194382 445692
rect 232866 445680 232872 445692
rect 232924 445680 232930 445732
rect 238846 445680 238852 445732
rect 238904 445720 238910 445732
rect 238904 445692 248414 445720
rect 238904 445680 238910 445692
rect 26326 445612 26332 445664
rect 26384 445652 26390 445664
rect 64782 445652 64788 445664
rect 26384 445624 64788 445652
rect 26384 445612 26390 445624
rect 64782 445612 64788 445624
rect 64840 445612 64846 445664
rect 82630 445612 82636 445664
rect 82688 445652 82694 445664
rect 120902 445652 120908 445664
rect 82688 445624 120908 445652
rect 82688 445612 82694 445624
rect 120902 445612 120908 445624
rect 120960 445612 120966 445664
rect 138290 445612 138296 445664
rect 138348 445652 138354 445664
rect 176930 445652 176936 445664
rect 138348 445624 176936 445652
rect 138348 445612 138354 445624
rect 176930 445612 176936 445624
rect 176988 445612 176994 445664
rect 211246 445612 211252 445664
rect 211304 445652 211310 445664
rect 240042 445652 240048 445664
rect 211304 445624 240048 445652
rect 211304 445612 211310 445624
rect 240042 445612 240048 445624
rect 240100 445612 240106 445664
rect 248386 445652 248414 445692
rect 295426 445680 295432 445732
rect 295484 445720 295490 445732
rect 324038 445720 324044 445732
rect 295484 445692 324044 445720
rect 295484 445680 295490 445692
rect 324038 445680 324044 445692
rect 324096 445680 324102 445732
rect 334342 445680 334348 445732
rect 334400 445720 334406 445732
rect 372982 445720 372988 445732
rect 334400 445692 372988 445720
rect 334400 445680 334406 445692
rect 372982 445680 372988 445692
rect 373040 445680 373046 445732
rect 390462 445680 390468 445732
rect 390520 445720 390526 445732
rect 428734 445720 428740 445732
rect 390520 445692 428740 445720
rect 390520 445680 390526 445692
rect 428734 445680 428740 445692
rect 428792 445680 428798 445732
rect 434806 445680 434812 445732
rect 434864 445720 434870 445732
rect 434864 445692 441614 445720
rect 434864 445680 434870 445692
rect 268010 445652 268016 445664
rect 248386 445624 268016 445652
rect 268010 445612 268016 445624
rect 268068 445612 268074 445664
rect 306282 445612 306288 445664
rect 306340 445652 306346 445664
rect 344738 445652 344744 445664
rect 306340 445624 344744 445652
rect 306340 445612 306346 445624
rect 344738 445612 344744 445624
rect 344796 445612 344802 445664
rect 362310 445612 362316 445664
rect 362368 445652 362374 445664
rect 400950 445652 400956 445664
rect 362368 445624 400956 445652
rect 362368 445612 362374 445624
rect 400950 445612 400956 445624
rect 401008 445612 401014 445664
rect 407206 445612 407212 445664
rect 407264 445652 407270 445664
rect 436002 445652 436008 445664
rect 407264 445624 436008 445652
rect 407264 445612 407270 445624
rect 436002 445612 436008 445624
rect 436060 445612 436066 445664
rect 441586 445652 441614 445692
rect 491386 445680 491392 445732
rect 491444 445720 491450 445732
rect 519998 445720 520004 445732
rect 491444 445692 520004 445720
rect 491444 445680 491450 445692
rect 519998 445680 520004 445692
rect 520056 445680 520062 445732
rect 530302 445680 530308 445732
rect 530360 445720 530366 445732
rect 568850 445720 568856 445732
rect 530360 445692 568856 445720
rect 530360 445680 530366 445692
rect 568850 445680 568856 445692
rect 568908 445680 568914 445732
rect 463694 445652 463700 445664
rect 441586 445624 463700 445652
rect 463694 445612 463700 445624
rect 463752 445612 463758 445664
rect 474642 445612 474648 445664
rect 474700 445652 474706 445664
rect 512822 445652 512828 445664
rect 474700 445624 512828 445652
rect 474700 445612 474706 445624
rect 512822 445612 512828 445624
rect 512880 445612 512886 445664
rect 518986 445612 518992 445664
rect 519044 445652 519050 445664
rect 547874 445652 547880 445664
rect 519044 445624 547880 445652
rect 519044 445612 519050 445624
rect 547874 445612 547880 445624
rect 547932 445612 547938 445664
rect 42886 445544 42892 445596
rect 42944 445584 42950 445596
rect 71774 445584 71780 445596
rect 42944 445556 71780 445584
rect 42944 445544 42950 445556
rect 71774 445544 71780 445556
rect 71832 445544 71838 445596
rect 127066 445544 127072 445596
rect 127124 445584 127130 445596
rect 156046 445584 156052 445596
rect 127124 445556 156052 445584
rect 127124 445544 127130 445556
rect 156046 445544 156052 445556
rect 156104 445544 156110 445596
rect 166626 445544 166632 445596
rect 166684 445584 166690 445596
rect 204990 445584 204996 445596
rect 166684 445556 204996 445584
rect 166684 445544 166690 445556
rect 204990 445544 204996 445556
rect 205048 445544 205054 445596
rect 278314 445544 278320 445596
rect 278372 445584 278378 445596
rect 316862 445584 316868 445596
rect 278372 445556 316868 445584
rect 278372 445544 278378 445556
rect 316862 445544 316868 445556
rect 316920 445544 316926 445596
rect 323026 445544 323032 445596
rect 323084 445584 323090 445596
rect 352006 445584 352012 445596
rect 323084 445556 352012 445584
rect 323084 445544 323090 445556
rect 352006 445544 352012 445556
rect 352064 445544 352070 445596
rect 446306 445544 446312 445596
rect 446364 445584 446370 445596
rect 484946 445584 484952 445596
rect 446364 445556 484952 445584
rect 446364 445544 446370 445556
rect 484946 445544 484952 445556
rect 485004 445544 485010 445596
rect 502334 445544 502340 445596
rect 502392 445584 502398 445596
rect 540790 445584 540796 445596
rect 502392 445556 540796 445584
rect 502392 445544 502398 445556
rect 540790 445544 540796 445556
rect 540848 445544 540854 445596
rect 548150 445544 548156 445596
rect 548208 445584 548214 445596
rect 557994 445584 558000 445596
rect 548208 445556 558000 445584
rect 548208 445544 548214 445556
rect 557994 445544 558000 445556
rect 558052 445544 558058 445596
rect 250346 445476 250352 445528
rect 250404 445516 250410 445528
rect 288986 445516 288992 445528
rect 250404 445488 288992 445516
rect 250404 445476 250410 445488
rect 288986 445476 288992 445488
rect 289044 445476 289050 445528
rect 26602 445000 26608 445052
rect 26660 445040 26666 445052
rect 36814 445040 36820 445052
rect 26660 445012 36820 445040
rect 26660 445000 26666 445012
rect 36814 445000 36820 445012
rect 36872 445000 36878 445052
rect 15378 444456 15384 444508
rect 15436 444496 15442 444508
rect 54294 444496 54300 444508
rect 15436 444468 54300 444496
rect 15436 444456 15442 444468
rect 54294 444456 54300 444468
rect 54352 444456 54358 444508
rect 65886 444456 65892 444508
rect 65944 444496 65950 444508
rect 82630 444496 82636 444508
rect 65944 444468 82636 444496
rect 65944 444456 65950 444468
rect 82630 444456 82636 444468
rect 82688 444456 82694 444508
rect 99466 444456 99472 444508
rect 99524 444496 99530 444508
rect 138290 444496 138296 444508
rect 99524 444468 138296 444496
rect 99524 444456 99530 444468
rect 138290 444456 138296 444468
rect 138348 444456 138354 444508
rect 149882 444456 149888 444508
rect 149940 444496 149946 444508
rect 156322 444496 156328 444508
rect 149940 444468 156328 444496
rect 149940 444456 149946 444468
rect 156322 444456 156328 444468
rect 156380 444456 156386 444508
rect 211154 444456 211160 444508
rect 211212 444496 211218 444508
rect 250622 444496 250628 444508
rect 211212 444468 250628 444496
rect 211212 444456 211218 444468
rect 250622 444456 250628 444468
rect 250680 444456 250686 444508
rect 261478 444456 261484 444508
rect 261536 444496 261542 444508
rect 278590 444496 278596 444508
rect 261536 444468 278596 444496
rect 261536 444456 261542 444468
rect 278590 444456 278596 444468
rect 278648 444456 278654 444508
rect 295426 444456 295432 444508
rect 295484 444496 295490 444508
rect 334618 444496 334624 444508
rect 295484 444468 334624 444496
rect 295484 444456 295490 444468
rect 334618 444456 334624 444468
rect 334676 444456 334682 444508
rect 345842 444456 345848 444508
rect 345900 444496 345906 444508
rect 362310 444496 362316 444508
rect 345900 444468 362316 444496
rect 345900 444456 345906 444468
rect 362310 444456 362316 444468
rect 362368 444456 362374 444508
rect 407114 444456 407120 444508
rect 407172 444496 407178 444508
rect 446306 444496 446312 444508
rect 407172 444468 446312 444496
rect 407172 444456 407178 444468
rect 446306 444456 446312 444468
rect 446364 444456 446370 444508
rect 457438 444456 457444 444508
rect 457496 444496 457502 444508
rect 474642 444496 474648 444508
rect 457496 444468 474648 444496
rect 457496 444456 457502 444468
rect 474642 444456 474648 444468
rect 474700 444456 474706 444508
rect 491386 444456 491392 444508
rect 491444 444496 491450 444508
rect 530302 444496 530308 444508
rect 491444 444468 530308 444496
rect 491444 444456 491450 444468
rect 530302 444456 530308 444468
rect 530360 444456 530366 444508
rect 71866 444388 71872 444440
rect 71924 444428 71930 444440
rect 110598 444428 110604 444440
rect 71924 444400 110604 444428
rect 71924 444388 71930 444400
rect 110598 444388 110604 444400
rect 110656 444388 110662 444440
rect 149790 444388 149796 444440
rect 149848 444428 149854 444440
rect 166626 444428 166632 444440
rect 149848 444400 166632 444428
rect 149848 444388 149854 444400
rect 166626 444388 166632 444400
rect 166684 444388 166690 444440
rect 183646 444388 183652 444440
rect 183704 444428 183710 444440
rect 222286 444428 222292 444440
rect 183704 444400 222292 444428
rect 183704 444388 183710 444400
rect 222286 444388 222292 444400
rect 222344 444388 222350 444440
rect 267826 444388 267832 444440
rect 267884 444428 267890 444440
rect 306466 444428 306472 444440
rect 267884 444400 306472 444428
rect 267884 444388 267890 444400
rect 306466 444388 306472 444400
rect 306524 444388 306530 444440
rect 318058 444388 318064 444440
rect 318116 444428 318122 444440
rect 324314 444428 324320 444440
rect 318116 444400 324320 444428
rect 318116 444388 318122 444400
rect 324314 444388 324320 444400
rect 324372 444388 324378 444440
rect 345658 444388 345664 444440
rect 345716 444428 345722 444440
rect 352006 444428 352012 444440
rect 345716 444400 352012 444428
rect 345716 444388 345722 444400
rect 352006 444388 352012 444400
rect 352064 444388 352070 444440
rect 379606 444388 379612 444440
rect 379664 444428 379670 444440
rect 418614 444428 418620 444440
rect 379664 444400 418620 444428
rect 379664 444388 379670 444400
rect 418614 444388 418620 444400
rect 418672 444388 418678 444440
rect 463786 444388 463792 444440
rect 463844 444428 463850 444440
rect 502610 444428 502616 444440
rect 463844 444400 502616 444428
rect 463844 444388 463850 444400
rect 502610 444388 502616 444400
rect 502668 444388 502674 444440
rect 514018 444388 514024 444440
rect 514076 444428 514082 444440
rect 520274 444428 520280 444440
rect 514076 444400 520280 444428
rect 514076 444388 514082 444400
rect 520274 444388 520280 444400
rect 520332 444388 520338 444440
rect 541618 444388 541624 444440
rect 541676 444428 541682 444440
rect 558638 444428 558644 444440
rect 541676 444400 558644 444428
rect 541676 444388 541682 444400
rect 558638 444388 558644 444400
rect 558696 444388 558702 444440
rect 429102 441600 429108 441652
rect 429160 441640 429166 441652
rect 429838 441640 429844 441652
rect 429160 441612 429844 441640
rect 429160 441600 429166 441612
rect 429838 441600 429844 441612
rect 429896 441600 429902 441652
rect 205082 441328 205088 441380
rect 205140 441328 205146 441380
rect 205100 441176 205128 441328
rect 345014 441192 345020 441244
rect 345072 441232 345078 441244
rect 345750 441232 345756 441244
rect 345072 441204 345756 441232
rect 345072 441192 345078 441204
rect 345750 441192 345756 441204
rect 345808 441192 345814 441244
rect 205082 441124 205088 441176
rect 205140 441124 205146 441176
rect 93118 439492 93124 439544
rect 93176 439532 93182 439544
rect 99926 439532 99932 439544
rect 93176 439504 99932 439532
rect 93176 439492 93182 439504
rect 99926 439492 99932 439504
rect 99984 439492 99990 439544
rect 177298 439492 177304 439544
rect 177356 439532 177362 439544
rect 184014 439532 184020 439544
rect 177356 439504 184020 439532
rect 177356 439492 177362 439504
rect 184014 439492 184020 439504
rect 184072 439492 184078 439544
rect 373258 439492 373264 439544
rect 373316 439532 373322 439544
rect 379974 439532 379980 439544
rect 373316 439504 379980 439532
rect 373316 439492 373322 439504
rect 379974 439492 379980 439504
rect 380032 439492 380038 439544
rect 457530 439492 457536 439544
rect 457588 439532 457594 439544
rect 464062 439532 464068 439544
rect 457588 439504 464068 439532
rect 457588 439492 457594 439504
rect 464062 439492 464068 439504
rect 464120 439492 464126 439544
rect 37090 438880 37096 438932
rect 37148 438920 37154 438932
rect 44174 438920 44180 438932
rect 37148 438892 44180 438920
rect 37148 438880 37154 438892
rect 44174 438880 44180 438892
rect 44232 438880 44238 438932
rect 65978 438880 65984 438932
rect 66036 438920 66042 438932
rect 71958 438920 71964 438932
rect 66036 438892 71964 438920
rect 66036 438880 66042 438892
rect 71958 438880 71964 438892
rect 72016 438880 72022 438932
rect 261570 438880 261576 438932
rect 261628 438920 261634 438932
rect 267918 438920 267924 438932
rect 261628 438892 267924 438920
rect 261628 438880 261634 438892
rect 267918 438880 267924 438892
rect 267976 438880 267982 438932
rect 289170 438880 289176 438932
rect 289228 438920 289234 438932
rect 295978 438920 295984 438932
rect 289228 438892 295984 438920
rect 289228 438880 289234 438892
rect 295978 438880 295984 438892
rect 296036 438880 296042 438932
rect 485130 438880 485136 438932
rect 485188 438920 485194 438932
rect 492030 438920 492036 438932
rect 485188 438892 492036 438920
rect 485188 438880 485194 438892
rect 492030 438880 492036 438892
rect 492088 438880 492094 438932
rect 37274 436568 37280 436620
rect 37332 436608 37338 436620
rect 38010 436608 38016 436620
rect 37332 436580 38016 436608
rect 37332 436568 37338 436580
rect 38010 436568 38016 436580
rect 38068 436568 38074 436620
rect 233234 436568 233240 436620
rect 233292 436608 233298 436620
rect 233970 436608 233976 436620
rect 233292 436580 233976 436608
rect 233292 436568 233298 436580
rect 233970 436568 233976 436580
rect 234028 436568 234034 436620
rect 211154 427116 211160 427168
rect 211212 427156 211218 427168
rect 211982 427156 211988 427168
rect 211212 427128 211988 427156
rect 211212 427116 211218 427128
rect 211982 427116 211988 427128
rect 212040 427116 212046 427168
rect 407114 427116 407120 427168
rect 407172 427156 407178 427168
rect 407942 427156 407948 427168
rect 407172 427128 407948 427156
rect 407172 427116 407178 427128
rect 407942 427116 407948 427128
rect 408000 427116 408006 427168
rect 15194 419432 15200 419484
rect 15252 419472 15258 419484
rect 36906 419472 36912 419484
rect 15252 419444 36912 419472
rect 15252 419432 15258 419444
rect 36906 419432 36912 419444
rect 36964 419432 36970 419484
rect 38010 419432 38016 419484
rect 38068 419472 38074 419484
rect 64874 419472 64880 419484
rect 38068 419444 64880 419472
rect 38068 419432 38074 419444
rect 64874 419432 64880 419444
rect 64932 419432 64938 419484
rect 65058 419432 65064 419484
rect 65116 419472 65122 419484
rect 92934 419472 92940 419484
rect 65116 419444 92940 419472
rect 65116 419432 65122 419444
rect 92934 419432 92940 419444
rect 92992 419432 92998 419484
rect 93026 419432 93032 419484
rect 93084 419472 93090 419484
rect 120902 419472 120908 419484
rect 93084 419444 120908 419472
rect 93084 419432 93090 419444
rect 120902 419432 120908 419444
rect 120960 419432 120966 419484
rect 121086 419432 121092 419484
rect 121144 419472 121150 419484
rect 148594 419472 148600 419484
rect 121144 419444 148600 419472
rect 121144 419432 121150 419444
rect 148594 419432 148600 419444
rect 148652 419432 148658 419484
rect 149698 419432 149704 419484
rect 149756 419472 149762 419484
rect 176930 419472 176936 419484
rect 149756 419444 176936 419472
rect 149756 419432 149762 419444
rect 176930 419432 176936 419444
rect 176988 419432 176994 419484
rect 177022 419432 177028 419484
rect 177080 419472 177086 419484
rect 204898 419472 204904 419484
rect 177080 419444 204904 419472
rect 177080 419432 177086 419444
rect 204898 419432 204904 419444
rect 204956 419432 204962 419484
rect 205174 419432 205180 419484
rect 205232 419472 205238 419484
rect 232590 419472 232596 419484
rect 205232 419444 232596 419472
rect 205232 419432 205238 419444
rect 232590 419432 232596 419444
rect 232648 419432 232654 419484
rect 233970 419432 233976 419484
rect 234028 419472 234034 419484
rect 260926 419472 260932 419484
rect 234028 419444 260932 419472
rect 234028 419432 234034 419444
rect 260926 419432 260932 419444
rect 260984 419432 260990 419484
rect 261018 419432 261024 419484
rect 261076 419472 261082 419484
rect 288894 419472 288900 419484
rect 261076 419444 288900 419472
rect 261076 419432 261082 419444
rect 288894 419432 288900 419444
rect 288952 419432 288958 419484
rect 289078 419432 289084 419484
rect 289136 419472 289142 419484
rect 316586 419472 316592 419484
rect 289136 419444 316592 419472
rect 289136 419432 289142 419444
rect 316586 419432 316592 419444
rect 316644 419432 316650 419484
rect 317046 419432 317052 419484
rect 317104 419472 317110 419484
rect 344922 419472 344928 419484
rect 317104 419444 344928 419472
rect 317104 419432 317110 419444
rect 344922 419432 344928 419444
rect 344980 419432 344986 419484
rect 345750 419432 345756 419484
rect 345808 419472 345814 419484
rect 372614 419472 372620 419484
rect 345808 419444 372620 419472
rect 345808 419432 345814 419444
rect 372614 419432 372620 419444
rect 372672 419432 372678 419484
rect 373074 419432 373080 419484
rect 373132 419472 373138 419484
rect 400950 419472 400956 419484
rect 373132 419444 400956 419472
rect 373132 419432 373138 419444
rect 400950 419432 400956 419444
rect 401008 419432 401014 419484
rect 401042 419432 401048 419484
rect 401100 419472 401106 419484
rect 428918 419472 428924 419484
rect 401100 419444 428924 419472
rect 401100 419432 401106 419444
rect 428918 419432 428924 419444
rect 428976 419432 428982 419484
rect 429838 419432 429844 419484
rect 429896 419472 429902 419484
rect 456794 419472 456800 419484
rect 429896 419444 456800 419472
rect 429896 419432 429902 419444
rect 456794 419432 456800 419444
rect 456852 419432 456858 419484
rect 457070 419432 457076 419484
rect 457128 419472 457134 419484
rect 484946 419472 484952 419484
rect 457128 419444 484952 419472
rect 457128 419432 457134 419444
rect 484946 419432 484952 419444
rect 485004 419432 485010 419484
rect 485038 419432 485044 419484
rect 485096 419472 485102 419484
rect 512914 419472 512920 419484
rect 485096 419444 512920 419472
rect 485096 419432 485102 419444
rect 512914 419432 512920 419444
rect 512972 419432 512978 419484
rect 513098 419432 513104 419484
rect 513156 419472 513162 419484
rect 540606 419472 540612 419484
rect 513156 419444 540612 419472
rect 513156 419432 513162 419444
rect 540606 419432 540612 419444
rect 540664 419432 540670 419484
rect 541066 419432 541072 419484
rect 541124 419472 541130 419484
rect 568942 419472 568948 419484
rect 541124 419444 568948 419472
rect 541124 419432 541130 419444
rect 568942 419432 568948 419444
rect 569000 419432 569006 419484
rect 26602 419364 26608 419416
rect 26660 419404 26666 419416
rect 37090 419404 37096 419416
rect 26660 419376 37096 419404
rect 26660 419364 26666 419376
rect 37090 419364 37096 419376
rect 37148 419364 37154 419416
rect 44634 419364 44640 419416
rect 44692 419404 44698 419416
rect 65886 419404 65892 419416
rect 44692 419376 65892 419404
rect 44692 419364 44698 419376
rect 65886 419364 65892 419376
rect 65944 419364 65950 419416
rect 82630 419364 82636 419416
rect 82688 419404 82694 419416
rect 93118 419404 93124 419416
rect 82688 419376 93124 419404
rect 82688 419364 82694 419376
rect 93118 419364 93124 419376
rect 93176 419364 93182 419416
rect 128630 419364 128636 419416
rect 128688 419404 128694 419416
rect 149790 419404 149796 419416
rect 128688 419376 149796 419404
rect 128688 419364 128694 419376
rect 149790 419364 149796 419376
rect 149848 419364 149854 419416
rect 166626 419364 166632 419416
rect 166684 419404 166690 419416
rect 177298 419404 177304 419416
rect 166684 419376 177304 419404
rect 166684 419364 166690 419376
rect 177298 419364 177304 419376
rect 177356 419364 177362 419416
rect 194594 419364 194600 419416
rect 194652 419404 194658 419416
rect 211246 419404 211252 419416
rect 194652 419376 211252 419404
rect 194652 419364 194658 419376
rect 211246 419364 211252 419376
rect 211304 419364 211310 419416
rect 222930 419364 222936 419416
rect 222988 419404 222994 419416
rect 240134 419404 240140 419416
rect 222988 419376 240140 419404
rect 222988 419364 222994 419376
rect 240134 419364 240140 419376
rect 240192 419364 240198 419416
rect 240318 419364 240324 419416
rect 240376 419404 240382 419416
rect 261478 419404 261484 419416
rect 240376 419376 261484 419404
rect 240376 419364 240382 419376
rect 261478 419364 261484 419376
rect 261536 419364 261542 419416
rect 278590 419364 278596 419416
rect 278648 419404 278654 419416
rect 289170 419404 289176 419416
rect 278648 419376 289176 419404
rect 278648 419364 278654 419376
rect 289170 419364 289176 419376
rect 289228 419364 289234 419416
rect 306926 419364 306932 419416
rect 306984 419404 306990 419416
rect 318058 419404 318064 419416
rect 306984 419376 318064 419404
rect 306984 419364 306990 419376
rect 318058 419364 318064 419376
rect 318116 419364 318122 419416
rect 324314 419364 324320 419416
rect 324372 419404 324378 419416
rect 345842 419404 345848 419416
rect 324372 419376 345848 419404
rect 324372 419364 324378 419376
rect 345842 419364 345848 419376
rect 345900 419364 345906 419416
rect 362862 419364 362868 419416
rect 362920 419404 362926 419416
rect 373258 419404 373264 419416
rect 362920 419376 373264 419404
rect 362920 419364 362926 419376
rect 373258 419364 373264 419376
rect 373316 419364 373322 419416
rect 390646 419364 390652 419416
rect 390704 419404 390710 419416
rect 407206 419404 407212 419416
rect 390704 419376 407212 419404
rect 390704 419364 390710 419376
rect 407206 419364 407212 419376
rect 407264 419364 407270 419416
rect 418614 419364 418620 419416
rect 418672 419404 418678 419416
rect 436094 419404 436100 419416
rect 418672 419376 436100 419404
rect 418672 419364 418678 419376
rect 436094 419364 436100 419376
rect 436152 419364 436158 419416
rect 436646 419364 436652 419416
rect 436704 419404 436710 419416
rect 457438 419404 457444 419416
rect 436704 419376 457444 419404
rect 436704 419364 436710 419376
rect 457438 419364 457444 419376
rect 457496 419364 457502 419416
rect 474642 419364 474648 419416
rect 474700 419404 474706 419416
rect 485130 419404 485136 419416
rect 474700 419376 485136 419404
rect 474700 419364 474706 419376
rect 485130 419364 485136 419376
rect 485188 419364 485194 419416
rect 502610 419364 502616 419416
rect 502668 419404 502674 419416
rect 514018 419404 514024 419416
rect 502668 419376 514024 419404
rect 502668 419364 502674 419376
rect 514018 419364 514024 419376
rect 514076 419364 514082 419416
rect 520642 419364 520648 419416
rect 520700 419404 520706 419416
rect 541618 419404 541624 419416
rect 520700 419376 541624 419404
rect 520700 419364 520706 419376
rect 541618 419364 541624 419376
rect 541676 419364 541682 419416
rect 54938 419296 54944 419348
rect 54996 419336 55002 419348
rect 65978 419336 65984 419348
rect 54996 419308 65984 419336
rect 54996 419296 55002 419308
rect 65978 419296 65984 419308
rect 66036 419296 66042 419348
rect 138934 419296 138940 419348
rect 138992 419336 138998 419348
rect 149882 419336 149888 419348
rect 138992 419308 149888 419336
rect 138992 419296 138998 419308
rect 149882 419296 149888 419308
rect 149940 419296 149946 419348
rect 250622 419296 250628 419348
rect 250680 419336 250686 419348
rect 261570 419336 261576 419348
rect 250680 419308 261576 419336
rect 250680 419296 250686 419308
rect 261570 419296 261576 419308
rect 261628 419296 261634 419348
rect 334618 419296 334624 419348
rect 334676 419336 334682 419348
rect 345658 419336 345664 419348
rect 334676 419308 345664 419336
rect 334676 419296 334682 419308
rect 345658 419296 345664 419308
rect 345716 419296 345722 419348
rect 446950 419296 446956 419348
rect 447008 419336 447014 419348
rect 457530 419336 457536 419348
rect 447008 419308 457536 419336
rect 447008 419296 447014 419308
rect 457530 419296 457536 419308
rect 457588 419296 457594 419348
rect 530946 419296 530952 419348
rect 531004 419336 531010 419348
rect 547966 419336 547972 419348
rect 531004 419308 547972 419336
rect 531004 419296 531010 419308
rect 547966 419296 547972 419308
rect 548024 419296 548030 419348
rect 558638 418752 558644 418804
rect 558696 418792 558702 418804
rect 568942 418792 568948 418804
rect 558696 418764 568948 418792
rect 558696 418752 558702 418764
rect 568942 418752 568948 418764
rect 569000 418752 569006 418804
rect 548334 417392 548340 417444
rect 548392 417432 548398 417444
rect 569034 417432 569040 417444
rect 548392 417404 569040 417432
rect 548392 417392 548398 417404
rect 569034 417392 569040 417404
rect 569092 417392 569098 417444
rect 100018 416916 100024 416968
rect 100076 416956 100082 416968
rect 121086 416956 121092 416968
rect 100076 416928 121092 416956
rect 100076 416916 100082 416928
rect 121086 416916 121092 416928
rect 121144 416916 121150 416968
rect 268010 416916 268016 416968
rect 268068 416956 268074 416968
rect 289078 416956 289084 416968
rect 268068 416928 289084 416956
rect 268068 416916 268074 416928
rect 289078 416916 289084 416928
rect 289136 416916 289142 416968
rect 380342 416916 380348 416968
rect 380400 416956 380406 416968
rect 401134 416956 401140 416968
rect 380400 416928 401140 416956
rect 380400 416916 380406 416928
rect 401134 416916 401140 416928
rect 401192 416916 401198 416968
rect 464338 416916 464344 416968
rect 464396 416956 464402 416968
rect 485038 416956 485044 416968
rect 464396 416928 485044 416956
rect 464396 416916 464402 416928
rect 485038 416916 485044 416928
rect 485096 416916 485102 416968
rect 92842 416848 92848 416900
rect 92900 416888 92906 416900
rect 110322 416888 110328 416900
rect 92900 416860 110328 416888
rect 92900 416848 92906 416860
rect 110322 416848 110328 416860
rect 110380 416848 110386 416900
rect 176838 416848 176844 416900
rect 176896 416888 176902 416900
rect 194318 416888 194324 416900
rect 176896 416860 194324 416888
rect 176896 416848 176902 416860
rect 194318 416848 194324 416860
rect 194376 416848 194382 416900
rect 204806 416848 204812 416900
rect 204864 416888 204870 416900
rect 222194 416888 222200 416900
rect 204864 416860 222200 416888
rect 204864 416848 204870 416860
rect 222194 416848 222200 416860
rect 222252 416848 222258 416900
rect 261478 416848 261484 416900
rect 261536 416888 261542 416900
rect 278314 416888 278320 416900
rect 261536 416860 278320 416888
rect 261536 416848 261542 416860
rect 278314 416848 278320 416860
rect 278372 416848 278378 416900
rect 372890 416848 372896 416900
rect 372948 416888 372954 416900
rect 390002 416888 390008 416900
rect 372948 416860 390008 416888
rect 372948 416848 372954 416860
rect 390002 416848 390008 416860
rect 390060 416848 390066 416900
rect 457438 416848 457444 416900
rect 457496 416888 457502 416900
rect 473998 416888 474004 416900
rect 457496 416860 474004 416888
rect 457496 416848 457502 416860
rect 473998 416848 474004 416860
rect 474056 416848 474062 416900
rect 15286 416780 15292 416832
rect 15344 416820 15350 416832
rect 26326 416820 26332 416832
rect 15344 416792 26332 416820
rect 15344 416780 15350 416792
rect 26326 416780 26332 416792
rect 26384 416780 26390 416832
rect 36906 416780 36912 416832
rect 36964 416820 36970 416832
rect 54294 416820 54300 416832
rect 36964 416792 54300 416820
rect 36964 416780 36970 416792
rect 54294 416780 54300 416792
rect 54352 416780 54358 416832
rect 72326 416780 72332 416832
rect 72384 416820 72390 416832
rect 93118 416820 93124 416832
rect 72384 416792 93124 416820
rect 72384 416780 72390 416792
rect 93118 416780 93124 416792
rect 93176 416780 93182 416832
rect 120994 416780 121000 416832
rect 121052 416820 121058 416832
rect 138290 416820 138296 416832
rect 121052 416792 138296 416820
rect 121052 416780 121058 416792
rect 138290 416780 138296 416792
rect 138348 416780 138354 416832
rect 156322 416780 156328 416832
rect 156380 416820 156386 416832
rect 177298 416820 177304 416832
rect 156380 416792 177304 416820
rect 156380 416780 156386 416792
rect 177298 416780 177304 416792
rect 177356 416780 177362 416832
rect 184014 416780 184020 416832
rect 184072 416820 184078 416832
rect 204898 416820 204904 416832
rect 184072 416792 204904 416820
rect 184072 416780 184078 416792
rect 204898 416780 204904 416792
rect 204956 416780 204962 416832
rect 232958 416780 232964 416832
rect 233016 416820 233022 416832
rect 250346 416820 250352 416832
rect 233016 416792 250352 416820
rect 233016 416780 233022 416792
rect 250346 416780 250352 416792
rect 250404 416780 250410 416832
rect 288894 416780 288900 416832
rect 288952 416820 288958 416832
rect 306006 416820 306012 416832
rect 288952 416792 306012 416820
rect 288952 416780 288958 416792
rect 306006 416780 306012 416792
rect 306064 416780 306070 416832
rect 316954 416780 316960 416832
rect 317012 416820 317018 416832
rect 334342 416820 334348 416832
rect 317012 416792 334348 416820
rect 317012 416780 317018 416792
rect 334342 416780 334348 416792
rect 334400 416780 334406 416832
rect 352006 416780 352012 416832
rect 352064 416820 352070 416832
rect 373258 416820 373264 416832
rect 352064 416792 373264 416820
rect 352064 416780 352070 416792
rect 373258 416780 373264 416792
rect 373316 416780 373322 416832
rect 401042 416780 401048 416832
rect 401100 416820 401106 416832
rect 418338 416820 418344 416832
rect 401100 416792 418344 416820
rect 401100 416780 401106 416792
rect 418338 416780 418344 416792
rect 418396 416780 418402 416832
rect 484854 416780 484860 416832
rect 484912 416820 484918 416832
rect 502334 416820 502340 416832
rect 484912 416792 502340 416820
rect 484912 416780 484918 416792
rect 502334 416780 502340 416792
rect 502392 416780 502398 416832
rect 512914 416780 512920 416832
rect 512972 416820 512978 416832
rect 530302 416820 530308 416832
rect 512972 416792 530308 416820
rect 512972 416780 512978 416792
rect 530302 416780 530308 416792
rect 530360 416780 530366 416832
rect 120718 414264 120724 414316
rect 120776 414304 120782 414316
rect 120994 414304 121000 414316
rect 120776 414276 121000 414304
rect 120776 414264 120782 414276
rect 120994 414264 121000 414276
rect 121052 414264 121058 414316
rect 232774 414264 232780 414316
rect 232832 414304 232838 414316
rect 232958 414304 232964 414316
rect 232832 414276 232964 414304
rect 232832 414264 232838 414276
rect 232958 414264 232964 414276
rect 233016 414264 233022 414316
rect 400766 414264 400772 414316
rect 400824 414304 400830 414316
rect 401042 414304 401048 414316
rect 400824 414276 401048 414304
rect 400824 414264 400830 414276
rect 401042 414264 401048 414276
rect 401100 414264 401106 414316
rect 36722 414196 36728 414248
rect 36780 414236 36786 414248
rect 36906 414236 36912 414248
rect 36780 414208 36912 414236
rect 36780 414196 36786 414208
rect 36906 414196 36912 414208
rect 36964 414196 36970 414248
rect 120810 414196 120816 414248
rect 120868 414236 120874 414248
rect 121086 414236 121092 414248
rect 120868 414208 121092 414236
rect 120868 414196 120874 414208
rect 121086 414196 121092 414208
rect 121144 414196 121150 414248
rect 204714 414196 204720 414248
rect 204772 414236 204778 414248
rect 204990 414236 204996 414248
rect 204772 414208 204996 414236
rect 204772 414196 204778 414208
rect 204990 414196 204996 414208
rect 205048 414196 205054 414248
rect 400858 414196 400864 414248
rect 400916 414236 400922 414248
rect 401134 414236 401140 414248
rect 400916 414208 401140 414236
rect 400916 414196 400922 414208
rect 401134 414196 401140 414208
rect 401192 414196 401198 414248
rect 512730 412836 512736 412888
rect 512788 412876 512794 412888
rect 512914 412876 512920 412888
rect 512788 412848 512920 412876
rect 512788 412836 512794 412848
rect 512914 412836 512920 412848
rect 512972 412836 512978 412888
rect 36814 412768 36820 412820
rect 36872 412768 36878 412820
rect 316862 412768 316868 412820
rect 316920 412768 316926 412820
rect 512822 412768 512828 412820
rect 512880 412768 512886 412820
rect 36832 412616 36860 412768
rect 316880 412616 316908 412768
rect 512840 412616 512868 412768
rect 36814 412564 36820 412616
rect 36872 412564 36878 412616
rect 316862 412564 316868 412616
rect 316920 412564 316926 412616
rect 512822 412564 512828 412616
rect 512880 412564 512886 412616
rect 568758 410864 568764 410916
rect 568816 410904 568822 410916
rect 568942 410904 568948 410916
rect 568816 410876 568948 410904
rect 568816 410864 568822 410876
rect 568942 410864 568948 410876
rect 569000 410864 569006 410916
rect 3142 410184 3148 410236
rect 3200 410224 3206 410236
rect 8938 410224 8944 410236
rect 3200 410196 8944 410224
rect 3200 410184 3206 410196
rect 8938 410184 8944 410196
rect 8996 410184 9002 410236
rect 316770 408688 316776 408740
rect 316828 408728 316834 408740
rect 316954 408728 316960 408740
rect 316828 408700 316960 408728
rect 316828 408688 316834 408700
rect 316954 408688 316960 408700
rect 317012 408688 317018 408740
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 11790 397508 11796 397520
rect 3384 397480 11796 397508
rect 3384 397468 3390 397480
rect 11790 397468 11796 397480
rect 11848 397468 11854 397520
rect 204898 397400 204904 397452
rect 204956 397440 204962 397452
rect 211706 397440 211712 397452
rect 204956 397412 211712 397440
rect 204956 397400 204962 397412
rect 211706 397400 211712 397412
rect 211764 397400 211770 397452
rect 485038 397400 485044 397452
rect 485096 397440 485102 397452
rect 491662 397440 491668 397452
rect 485096 397412 491668 397440
rect 485096 397400 485102 397412
rect 491662 397400 491668 397412
rect 491720 397400 491726 397452
rect 93118 396720 93124 396772
rect 93176 396760 93182 396772
rect 99742 396760 99748 396772
rect 93176 396732 99748 396760
rect 93176 396720 93182 396732
rect 99742 396720 99748 396732
rect 99800 396720 99806 396772
rect 120810 396720 120816 396772
rect 120868 396760 120874 396772
rect 127710 396760 127716 396772
rect 120868 396732 127716 396760
rect 120868 396720 120874 396732
rect 127710 396720 127716 396732
rect 127768 396720 127774 396772
rect 177298 396720 177304 396772
rect 177356 396760 177362 396772
rect 183646 396760 183652 396772
rect 177356 396732 183652 396760
rect 177356 396720 177362 396732
rect 183646 396720 183652 396732
rect 183704 396720 183710 396772
rect 373258 396720 373264 396772
rect 373316 396760 373322 396772
rect 379698 396760 379704 396772
rect 373316 396732 379704 396760
rect 373316 396720 373322 396732
rect 379698 396720 379704 396732
rect 379756 396720 379762 396772
rect 400858 396720 400864 396772
rect 400916 396760 400922 396772
rect 407758 396760 407764 396772
rect 400916 396732 407764 396760
rect 400916 396720 400922 396732
rect 407758 396720 407764 396732
rect 407816 396720 407822 396772
rect 289078 396448 289084 396500
rect 289136 396488 289142 396500
rect 295702 396488 295708 396500
rect 289136 396460 295708 396488
rect 289136 396448 289142 396460
rect 295702 396448 295708 396460
rect 295760 396448 295766 396500
rect 92750 394816 92756 394868
rect 92808 394816 92814 394868
rect 176746 394816 176752 394868
rect 176804 394816 176810 394868
rect 288802 394816 288808 394868
rect 288860 394816 288866 394868
rect 372798 394816 372804 394868
rect 372856 394816 372862 394868
rect 484762 394816 484768 394868
rect 484820 394816 484826 394868
rect 15286 394680 15292 394732
rect 15344 394720 15350 394732
rect 16114 394720 16120 394732
rect 15344 394692 16120 394720
rect 15344 394680 15350 394692
rect 16114 394680 16120 394692
rect 16172 394680 16178 394732
rect 92768 394664 92796 394816
rect 176764 394664 176792 394816
rect 288820 394664 288848 394816
rect 372816 394664 372844 394816
rect 484780 394664 484808 394816
rect 547874 394680 547880 394732
rect 547932 394720 547938 394732
rect 548150 394720 548156 394732
rect 547932 394692 548156 394720
rect 547932 394680 547938 394692
rect 548150 394680 548156 394692
rect 548208 394680 548214 394732
rect 92750 394612 92756 394664
rect 92808 394612 92814 394664
rect 176746 394612 176752 394664
rect 176804 394612 176810 394664
rect 288802 394612 288808 394664
rect 288860 394612 288866 394664
rect 372798 394612 372804 394664
rect 372856 394612 372862 394664
rect 484762 394612 484768 394664
rect 484820 394612 484826 394664
rect 15378 391892 15384 391944
rect 15436 391932 15442 391944
rect 43990 391932 43996 391944
rect 15436 391904 43996 391932
rect 15436 391892 15442 391904
rect 43990 391892 43996 391904
rect 44048 391892 44054 391944
rect 54294 391892 54300 391944
rect 54352 391932 54358 391944
rect 92750 391932 92756 391944
rect 54352 391904 92756 391932
rect 54352 391892 54358 391904
rect 92750 391892 92756 391904
rect 92808 391892 92814 391944
rect 138290 391892 138296 391944
rect 138348 391932 138354 391944
rect 176746 391932 176752 391944
rect 138348 391904 176752 391932
rect 138348 391892 138354 391904
rect 176746 391892 176752 391904
rect 176804 391892 176810 391944
rect 194318 391892 194324 391944
rect 194376 391932 194382 391944
rect 232866 391932 232872 391944
rect 194376 391904 232872 391932
rect 194376 391892 194382 391904
rect 232866 391892 232872 391904
rect 232924 391892 232930 391944
rect 238846 391892 238852 391944
rect 238904 391932 238910 391944
rect 238904 391904 248414 391932
rect 238904 391892 238910 391904
rect 26326 391824 26332 391876
rect 26384 391864 26390 391876
rect 64782 391864 64788 391876
rect 26384 391836 64788 391864
rect 26384 391824 26390 391836
rect 64782 391824 64788 391836
rect 64840 391824 64846 391876
rect 82630 391824 82636 391876
rect 82688 391864 82694 391876
rect 120902 391864 120908 391876
rect 82688 391836 120908 391864
rect 82688 391824 82694 391836
rect 120902 391824 120908 391836
rect 120960 391824 120966 391876
rect 127066 391824 127072 391876
rect 127124 391864 127130 391876
rect 155954 391864 155960 391876
rect 127124 391836 155960 391864
rect 127124 391824 127130 391836
rect 155954 391824 155960 391836
rect 156012 391824 156018 391876
rect 166626 391824 166632 391876
rect 166684 391864 166690 391876
rect 204990 391864 204996 391876
rect 166684 391836 204996 391864
rect 166684 391824 166690 391836
rect 204990 391824 204996 391836
rect 205048 391824 205054 391876
rect 211246 391824 211252 391876
rect 211304 391864 211310 391876
rect 240042 391864 240048 391876
rect 211304 391836 240048 391864
rect 211304 391824 211310 391836
rect 240042 391824 240048 391836
rect 240100 391824 240106 391876
rect 248386 391864 248414 391904
rect 295426 391892 295432 391944
rect 295484 391932 295490 391944
rect 324038 391932 324044 391944
rect 295484 391904 324044 391932
rect 295484 391892 295490 391904
rect 324038 391892 324044 391904
rect 324096 391892 324102 391944
rect 334342 391892 334348 391944
rect 334400 391932 334406 391944
rect 372798 391932 372804 391944
rect 334400 391904 372804 391932
rect 334400 391892 334406 391904
rect 372798 391892 372804 391904
rect 372856 391892 372862 391944
rect 390462 391892 390468 391944
rect 390520 391932 390526 391944
rect 428734 391932 428740 391944
rect 390520 391904 428740 391932
rect 390520 391892 390526 391904
rect 428734 391892 428740 391904
rect 428792 391892 428798 391944
rect 434806 391892 434812 391944
rect 434864 391932 434870 391944
rect 434864 391904 441614 391932
rect 434864 391892 434870 391904
rect 268010 391864 268016 391876
rect 248386 391836 268016 391864
rect 268010 391824 268016 391836
rect 268068 391824 268074 391876
rect 306282 391824 306288 391876
rect 306340 391864 306346 391876
rect 344738 391864 344744 391876
rect 306340 391836 344744 391864
rect 306340 391824 306346 391836
rect 344738 391824 344744 391836
rect 344796 391824 344802 391876
rect 362310 391824 362316 391876
rect 362368 391864 362374 391876
rect 400950 391864 400956 391876
rect 362368 391836 400956 391864
rect 362368 391824 362374 391836
rect 400950 391824 400956 391836
rect 401008 391824 401014 391876
rect 407206 391824 407212 391876
rect 407264 391864 407270 391876
rect 436002 391864 436008 391876
rect 407264 391836 436008 391864
rect 407264 391824 407270 391836
rect 436002 391824 436008 391836
rect 436060 391824 436066 391876
rect 441586 391864 441614 391904
rect 491386 391892 491392 391944
rect 491444 391932 491450 391944
rect 519998 391932 520004 391944
rect 491444 391904 520004 391932
rect 491444 391892 491450 391904
rect 519998 391892 520004 391904
rect 520056 391892 520062 391944
rect 530302 391892 530308 391944
rect 530360 391932 530366 391944
rect 568850 391932 568856 391944
rect 530360 391904 568856 391932
rect 530360 391892 530366 391904
rect 568850 391892 568856 391904
rect 568908 391892 568914 391944
rect 463786 391864 463792 391876
rect 441586 391836 463792 391864
rect 463786 391824 463792 391836
rect 463844 391824 463850 391876
rect 474642 391824 474648 391876
rect 474700 391864 474706 391876
rect 512822 391864 512828 391876
rect 474700 391836 512828 391864
rect 474700 391824 474706 391836
rect 512822 391824 512828 391836
rect 512880 391824 512886 391876
rect 548150 391824 548156 391876
rect 548208 391864 548214 391876
rect 557994 391864 558000 391876
rect 548208 391836 558000 391864
rect 548208 391824 548214 391836
rect 557994 391824 558000 391836
rect 558052 391824 558058 391876
rect 42886 391756 42892 391808
rect 42944 391796 42950 391808
rect 71774 391796 71780 391808
rect 42944 391768 71780 391796
rect 42944 391756 42950 391768
rect 71774 391756 71780 391768
rect 71832 391756 71838 391808
rect 110322 391756 110328 391808
rect 110380 391796 110386 391808
rect 148778 391796 148784 391808
rect 110380 391768 148784 391796
rect 110380 391756 110386 391768
rect 148778 391756 148784 391768
rect 148836 391756 148842 391808
rect 278314 391756 278320 391808
rect 278372 391796 278378 391808
rect 316862 391796 316868 391808
rect 278372 391768 316868 391796
rect 278372 391756 278378 391768
rect 316862 391756 316868 391768
rect 316920 391756 316926 391808
rect 323026 391756 323032 391808
rect 323084 391796 323090 391808
rect 352006 391796 352012 391808
rect 323084 391768 352012 391796
rect 323084 391756 323090 391768
rect 352006 391756 352012 391768
rect 352064 391756 352070 391808
rect 446306 391756 446312 391808
rect 446364 391796 446370 391808
rect 484762 391796 484768 391808
rect 446364 391768 484768 391796
rect 446364 391756 446370 391768
rect 484762 391756 484768 391768
rect 484820 391756 484826 391808
rect 502334 391756 502340 391808
rect 502392 391796 502398 391808
rect 540790 391796 540796 391808
rect 502392 391768 540796 391796
rect 502392 391756 502398 391768
rect 540790 391756 540796 391768
rect 540848 391756 540854 391808
rect 250346 391688 250352 391740
rect 250404 391728 250410 391740
rect 288802 391728 288808 391740
rect 250404 391700 288808 391728
rect 250404 391688 250410 391700
rect 288802 391688 288808 391700
rect 288860 391688 288866 391740
rect 518986 391688 518992 391740
rect 519044 391728 519050 391740
rect 547874 391728 547880 391740
rect 519044 391700 547880 391728
rect 519044 391688 519050 391700
rect 547874 391688 547880 391700
rect 547932 391688 547938 391740
rect 26602 389784 26608 389836
rect 26660 389824 26666 389836
rect 36814 389824 36820 389836
rect 26660 389796 36820 389824
rect 26660 389784 26666 389796
rect 36814 389784 36820 389796
rect 36872 389784 36878 389836
rect 15378 389308 15384 389360
rect 15436 389348 15442 389360
rect 54294 389348 54300 389360
rect 15436 389320 54300 389348
rect 15436 389308 15442 389320
rect 54294 389308 54300 389320
rect 54352 389308 54358 389360
rect 65886 389240 65892 389292
rect 65944 389280 65950 389292
rect 82630 389280 82636 389292
rect 65944 389252 82636 389280
rect 65944 389240 65950 389252
rect 82630 389240 82636 389252
rect 82688 389240 82694 389292
rect 99466 389240 99472 389292
rect 99524 389280 99530 389292
rect 138290 389280 138296 389292
rect 99524 389252 138296 389280
rect 99524 389240 99530 389252
rect 138290 389240 138296 389252
rect 138348 389240 138354 389292
rect 149698 389240 149704 389292
rect 149756 389280 149762 389292
rect 156322 389280 156328 389292
rect 149756 389252 156328 389280
rect 149756 389240 149762 389252
rect 156322 389240 156328 389252
rect 156380 389240 156386 389292
rect 211246 389240 211252 389292
rect 211304 389280 211310 389292
rect 250622 389280 250628 389292
rect 211304 389252 250628 389280
rect 211304 389240 211310 389252
rect 250622 389240 250628 389252
rect 250680 389240 250686 389292
rect 261478 389240 261484 389292
rect 261536 389280 261542 389292
rect 278590 389280 278596 389292
rect 261536 389252 278596 389280
rect 261536 389240 261542 389252
rect 278590 389240 278596 389252
rect 278648 389240 278654 389292
rect 295426 389240 295432 389292
rect 295484 389280 295490 389292
rect 334618 389280 334624 389292
rect 295484 389252 334624 389280
rect 295484 389240 295490 389252
rect 334618 389240 334624 389252
rect 334676 389240 334682 389292
rect 345750 389240 345756 389292
rect 345808 389280 345814 389292
rect 362310 389280 362316 389292
rect 345808 389252 362316 389280
rect 345808 389240 345814 389252
rect 362310 389240 362316 389252
rect 362368 389240 362374 389292
rect 407206 389240 407212 389292
rect 407264 389280 407270 389292
rect 446306 389280 446312 389292
rect 407264 389252 446312 389280
rect 407264 389240 407270 389252
rect 446306 389240 446312 389252
rect 446364 389240 446370 389292
rect 457438 389240 457444 389292
rect 457496 389280 457502 389292
rect 474642 389280 474648 389292
rect 457496 389252 474648 389280
rect 457496 389240 457502 389252
rect 474642 389240 474648 389252
rect 474700 389240 474706 389292
rect 491386 389240 491392 389292
rect 491444 389280 491450 389292
rect 530302 389280 530308 389292
rect 491444 389252 530308 389280
rect 491444 389240 491450 389252
rect 530302 389240 530308 389252
rect 530360 389240 530366 389292
rect 38010 389172 38016 389224
rect 38068 389212 38074 389224
rect 44174 389212 44180 389224
rect 38068 389184 44180 389212
rect 38068 389172 38074 389184
rect 44174 389172 44180 389184
rect 44232 389172 44238 389224
rect 71774 389172 71780 389224
rect 71832 389212 71838 389224
rect 110598 389212 110604 389224
rect 71832 389184 110604 389212
rect 71832 389172 71838 389184
rect 110598 389172 110604 389184
rect 110656 389172 110662 389224
rect 149790 389172 149796 389224
rect 149848 389212 149854 389224
rect 166626 389212 166632 389224
rect 149848 389184 166632 389212
rect 149848 389172 149854 389184
rect 166626 389172 166632 389184
rect 166684 389172 166690 389224
rect 183554 389172 183560 389224
rect 183612 389212 183618 389224
rect 222286 389212 222292 389224
rect 183612 389184 222292 389212
rect 183612 389172 183618 389184
rect 222286 389172 222292 389184
rect 222344 389172 222350 389224
rect 233970 389172 233976 389224
rect 234028 389212 234034 389224
rect 240318 389212 240324 389224
rect 234028 389184 240324 389212
rect 234028 389172 234034 389184
rect 240318 389172 240324 389184
rect 240376 389172 240382 389224
rect 267826 389172 267832 389224
rect 267884 389212 267890 389224
rect 306466 389212 306472 389224
rect 267884 389184 306472 389212
rect 267884 389172 267890 389184
rect 306466 389172 306472 389184
rect 306524 389172 306530 389224
rect 318058 389172 318064 389224
rect 318116 389212 318122 389224
rect 324314 389212 324320 389224
rect 318116 389184 324320 389212
rect 318116 389172 318122 389184
rect 324314 389172 324320 389184
rect 324372 389172 324378 389224
rect 345658 389172 345664 389224
rect 345716 389212 345722 389224
rect 352006 389212 352012 389224
rect 345716 389184 352012 389212
rect 345716 389172 345722 389184
rect 352006 389172 352012 389184
rect 352064 389172 352070 389224
rect 379606 389172 379612 389224
rect 379664 389212 379670 389224
rect 418614 389212 418620 389224
rect 379664 389184 418620 389212
rect 379664 389172 379670 389184
rect 418614 389172 418620 389184
rect 418672 389172 418678 389224
rect 429838 389172 429844 389224
rect 429896 389212 429902 389224
rect 436094 389212 436100 389224
rect 429896 389184 436100 389212
rect 429896 389172 429902 389184
rect 436094 389172 436100 389184
rect 436152 389172 436158 389224
rect 463694 389172 463700 389224
rect 463752 389212 463758 389224
rect 502610 389212 502616 389224
rect 463752 389184 502616 389212
rect 463752 389172 463758 389184
rect 502610 389172 502616 389184
rect 502668 389172 502674 389224
rect 514018 389172 514024 389224
rect 514076 389212 514082 389224
rect 520274 389212 520280 389224
rect 514076 389184 520280 389212
rect 514076 389172 514082 389184
rect 520274 389172 520280 389184
rect 520332 389172 520338 389224
rect 541618 389172 541624 389224
rect 541676 389212 541682 389224
rect 558638 389212 558644 389224
rect 541676 389184 558644 389212
rect 541676 389172 541682 389184
rect 558638 389172 558644 389184
rect 558696 389172 558702 389224
rect 205082 387336 205088 387388
rect 205140 387336 205146 387388
rect 205100 387184 205128 387336
rect 345014 387200 345020 387252
rect 345072 387240 345078 387252
rect 345842 387240 345848 387252
rect 345072 387212 345848 387240
rect 345072 387200 345078 387212
rect 345842 387200 345848 387212
rect 345900 387200 345906 387252
rect 205082 387132 205088 387184
rect 205140 387132 205146 387184
rect 429102 386384 429108 386436
rect 429160 386424 429166 386436
rect 429930 386424 429936 386436
rect 429160 386396 429936 386424
rect 429160 386384 429166 386396
rect 429930 386384 429936 386396
rect 429988 386384 429994 386436
rect 37274 385432 37280 385484
rect 37332 385472 37338 385484
rect 38102 385472 38108 385484
rect 37332 385444 38108 385472
rect 37332 385432 37338 385444
rect 38102 385432 38108 385444
rect 38160 385432 38166 385484
rect 99374 385432 99380 385484
rect 99432 385472 99438 385484
rect 99926 385472 99932 385484
rect 99432 385444 99932 385472
rect 99432 385432 99438 385444
rect 99926 385432 99932 385444
rect 99984 385432 99990 385484
rect 149238 385432 149244 385484
rect 149296 385472 149302 385484
rect 149882 385472 149888 385484
rect 149296 385444 149888 385472
rect 149296 385432 149302 385444
rect 149882 385432 149888 385444
rect 149940 385432 149946 385484
rect 211154 385432 211160 385484
rect 211212 385472 211218 385484
rect 211982 385472 211988 385484
rect 211212 385444 211988 385472
rect 211212 385432 211218 385444
rect 211982 385432 211988 385444
rect 212040 385432 212046 385484
rect 233234 385432 233240 385484
rect 233292 385472 233298 385484
rect 234062 385472 234068 385484
rect 233292 385444 234068 385472
rect 233292 385432 233298 385444
rect 234062 385432 234068 385444
rect 234120 385432 234126 385484
rect 295334 385432 295340 385484
rect 295392 385472 295398 385484
rect 295978 385472 295984 385484
rect 295392 385444 295984 385472
rect 295392 385432 295398 385444
rect 295978 385432 295984 385444
rect 296036 385432 296042 385484
rect 379514 385432 379520 385484
rect 379572 385472 379578 385484
rect 379974 385472 379980 385484
rect 379572 385444 379980 385472
rect 379572 385432 379578 385444
rect 379974 385432 379980 385444
rect 380032 385432 380038 385484
rect 407114 385432 407120 385484
rect 407172 385472 407178 385484
rect 407942 385472 407948 385484
rect 407172 385444 407948 385472
rect 407172 385432 407178 385444
rect 407942 385432 407948 385444
rect 408000 385432 408006 385484
rect 491294 385432 491300 385484
rect 491352 385472 491358 385484
rect 492030 385472 492036 385484
rect 491352 385444 492036 385472
rect 491352 385432 491358 385444
rect 492030 385432 492036 385444
rect 492088 385432 492094 385484
rect 267734 384752 267740 384804
rect 267792 384792 267798 384804
rect 267918 384792 267924 384804
rect 267792 384764 267924 384792
rect 267792 384752 267798 384764
rect 267918 384752 267924 384764
rect 267976 384752 267982 384804
rect 463694 378768 463700 378820
rect 463752 378808 463758 378820
rect 463970 378808 463976 378820
rect 463752 378780 463976 378808
rect 463752 378768 463758 378780
rect 463970 378768 463976 378780
rect 464028 378768 464034 378820
rect 569218 378156 569224 378208
rect 569276 378196 569282 378208
rect 579798 378196 579804 378208
rect 569276 378168 579804 378196
rect 569276 378156 569282 378168
rect 579798 378156 579804 378168
rect 579856 378156 579862 378208
rect 183554 370540 183560 370592
rect 183612 370580 183618 370592
rect 184014 370580 184020 370592
rect 183612 370552 184020 370580
rect 183612 370540 183618 370552
rect 184014 370540 184020 370552
rect 184072 370540 184078 370592
rect 42702 368432 42708 368484
rect 42760 368472 42766 368484
rect 95234 368472 95240 368484
rect 42760 368444 95240 368472
rect 42760 368432 42766 368444
rect 95234 368432 95240 368444
rect 95292 368432 95298 368484
rect 97902 368432 97908 368484
rect 97960 368472 97966 368484
rect 150434 368472 150440 368484
rect 97960 368444 150440 368472
rect 97960 368432 97966 368444
rect 150434 368432 150440 368444
rect 150492 368432 150498 368484
rect 154482 368432 154488 368484
rect 154540 368472 154546 368484
rect 207014 368472 207020 368484
rect 154540 368444 207020 368472
rect 154540 368432 154546 368444
rect 207014 368432 207020 368444
rect 207072 368432 207078 368484
rect 209682 368432 209688 368484
rect 209740 368472 209746 368484
rect 262214 368472 262220 368484
rect 209740 368444 262220 368472
rect 209740 368432 209746 368444
rect 262214 368432 262220 368444
rect 262272 368432 262278 368484
rect 266262 368432 266268 368484
rect 266320 368472 266326 368484
rect 318794 368472 318800 368484
rect 266320 368444 318800 368472
rect 266320 368432 266326 368444
rect 318794 368432 318800 368444
rect 318852 368432 318858 368484
rect 322842 368432 322848 368484
rect 322900 368472 322906 368484
rect 375374 368472 375380 368484
rect 322900 368444 375380 368472
rect 322900 368432 322906 368444
rect 375374 368432 375380 368444
rect 375432 368432 375438 368484
rect 378042 368432 378048 368484
rect 378100 368472 378106 368484
rect 430574 368472 430580 368484
rect 378100 368444 430580 368472
rect 378100 368432 378106 368444
rect 430574 368432 430580 368444
rect 430632 368432 430638 368484
rect 434622 368432 434628 368484
rect 434680 368472 434686 368484
rect 487154 368472 487160 368484
rect 434680 368444 487160 368472
rect 434680 368432 434686 368444
rect 487154 368432 487160 368444
rect 487212 368432 487218 368484
rect 489822 368432 489828 368484
rect 489880 368472 489886 368484
rect 542354 368472 542360 368484
rect 489880 368444 542360 368472
rect 489880 368432 489886 368444
rect 542354 368432 542360 368444
rect 542412 368432 542418 368484
rect 71774 367684 71780 367736
rect 71832 367724 71838 367736
rect 72050 367724 72056 367736
rect 71832 367696 72056 367724
rect 71832 367684 71838 367696
rect 72050 367684 72056 367696
rect 72108 367684 72114 367736
rect 15194 365644 15200 365696
rect 15252 365684 15258 365696
rect 36906 365684 36912 365696
rect 15252 365656 36912 365684
rect 15252 365644 15258 365656
rect 36906 365644 36912 365656
rect 36964 365644 36970 365696
rect 38102 365644 38108 365696
rect 38160 365684 38166 365696
rect 64874 365684 64880 365696
rect 38160 365656 64880 365684
rect 38160 365644 38166 365656
rect 64874 365644 64880 365656
rect 64932 365644 64938 365696
rect 65058 365644 65064 365696
rect 65116 365684 65122 365696
rect 92934 365684 92940 365696
rect 65116 365656 92940 365684
rect 65116 365644 65122 365656
rect 92934 365644 92940 365656
rect 92992 365644 92998 365696
rect 93026 365644 93032 365696
rect 93084 365684 93090 365696
rect 120902 365684 120908 365696
rect 93084 365656 120908 365684
rect 93084 365644 93090 365656
rect 120902 365644 120908 365656
rect 120960 365644 120966 365696
rect 121086 365644 121092 365696
rect 121144 365684 121150 365696
rect 148594 365684 148600 365696
rect 121144 365656 148600 365684
rect 121144 365644 121150 365656
rect 148594 365644 148600 365656
rect 148652 365644 148658 365696
rect 149882 365644 149888 365696
rect 149940 365684 149946 365696
rect 176930 365684 176936 365696
rect 149940 365656 176936 365684
rect 149940 365644 149946 365656
rect 176930 365644 176936 365656
rect 176988 365644 176994 365696
rect 177022 365644 177028 365696
rect 177080 365684 177086 365696
rect 204898 365684 204904 365696
rect 177080 365656 204904 365684
rect 177080 365644 177086 365656
rect 204898 365644 204904 365656
rect 204956 365644 204962 365696
rect 205174 365644 205180 365696
rect 205232 365684 205238 365696
rect 232590 365684 232596 365696
rect 205232 365656 232596 365684
rect 205232 365644 205238 365656
rect 232590 365644 232596 365656
rect 232648 365644 232654 365696
rect 234062 365644 234068 365696
rect 234120 365684 234126 365696
rect 260926 365684 260932 365696
rect 234120 365656 260932 365684
rect 234120 365644 234126 365656
rect 260926 365644 260932 365656
rect 260984 365644 260990 365696
rect 261018 365644 261024 365696
rect 261076 365684 261082 365696
rect 288894 365684 288900 365696
rect 261076 365656 288900 365684
rect 261076 365644 261082 365656
rect 288894 365644 288900 365656
rect 288952 365644 288958 365696
rect 289078 365644 289084 365696
rect 289136 365684 289142 365696
rect 316586 365684 316592 365696
rect 289136 365656 316592 365684
rect 289136 365644 289142 365656
rect 316586 365644 316592 365656
rect 316644 365644 316650 365696
rect 317046 365644 317052 365696
rect 317104 365684 317110 365696
rect 344922 365684 344928 365696
rect 317104 365656 344928 365684
rect 317104 365644 317110 365656
rect 344922 365644 344928 365656
rect 344980 365644 344986 365696
rect 345842 365644 345848 365696
rect 345900 365684 345906 365696
rect 372614 365684 372620 365696
rect 345900 365656 372620 365684
rect 345900 365644 345906 365656
rect 372614 365644 372620 365656
rect 372672 365644 372678 365696
rect 373074 365644 373080 365696
rect 373132 365684 373138 365696
rect 400950 365684 400956 365696
rect 373132 365656 400956 365684
rect 373132 365644 373138 365656
rect 400950 365644 400956 365656
rect 401008 365644 401014 365696
rect 401042 365644 401048 365696
rect 401100 365684 401106 365696
rect 428918 365684 428924 365696
rect 401100 365656 428924 365684
rect 401100 365644 401106 365656
rect 428918 365644 428924 365656
rect 428976 365644 428982 365696
rect 429930 365644 429936 365696
rect 429988 365684 429994 365696
rect 456794 365684 456800 365696
rect 429988 365656 456800 365684
rect 429988 365644 429994 365656
rect 456794 365644 456800 365656
rect 456852 365644 456858 365696
rect 457070 365644 457076 365696
rect 457128 365684 457134 365696
rect 484946 365684 484952 365696
rect 457128 365656 484952 365684
rect 457128 365644 457134 365656
rect 484946 365644 484952 365656
rect 485004 365644 485010 365696
rect 485038 365644 485044 365696
rect 485096 365684 485102 365696
rect 512914 365684 512920 365696
rect 485096 365656 512920 365684
rect 485096 365644 485102 365656
rect 512914 365644 512920 365656
rect 512972 365644 512978 365696
rect 513098 365644 513104 365696
rect 513156 365684 513162 365696
rect 540606 365684 540612 365696
rect 513156 365656 540612 365684
rect 513156 365644 513162 365656
rect 540606 365644 540612 365656
rect 540664 365644 540670 365696
rect 541066 365644 541072 365696
rect 541124 365684 541130 365696
rect 568942 365684 568948 365696
rect 541124 365656 568948 365684
rect 541124 365644 541130 365656
rect 568942 365644 568948 365656
rect 569000 365644 569006 365696
rect 26602 365576 26608 365628
rect 26660 365616 26666 365628
rect 38010 365616 38016 365628
rect 26660 365588 38016 365616
rect 26660 365576 26666 365588
rect 38010 365576 38016 365588
rect 38068 365576 38074 365628
rect 44634 365576 44640 365628
rect 44692 365616 44698 365628
rect 65886 365616 65892 365628
rect 44692 365588 65892 365616
rect 44692 365576 44698 365588
rect 65886 365576 65892 365588
rect 65944 365576 65950 365628
rect 82630 365576 82636 365628
rect 82688 365616 82694 365628
rect 99374 365616 99380 365628
rect 82688 365588 99380 365616
rect 82688 365576 82694 365588
rect 99374 365576 99380 365588
rect 99432 365576 99438 365628
rect 128630 365576 128636 365628
rect 128688 365616 128694 365628
rect 149790 365616 149796 365628
rect 128688 365588 149796 365616
rect 128688 365576 128694 365588
rect 149790 365576 149796 365588
rect 149848 365576 149854 365628
rect 166626 365576 166632 365628
rect 166684 365616 166690 365628
rect 183646 365616 183652 365628
rect 166684 365588 183652 365616
rect 166684 365576 166690 365588
rect 183646 365576 183652 365588
rect 183704 365576 183710 365628
rect 194594 365576 194600 365628
rect 194652 365616 194658 365628
rect 211154 365616 211160 365628
rect 194652 365588 211160 365616
rect 194652 365576 194658 365588
rect 211154 365576 211160 365588
rect 211212 365576 211218 365628
rect 222930 365576 222936 365628
rect 222988 365616 222994 365628
rect 233970 365616 233976 365628
rect 222988 365588 233976 365616
rect 222988 365576 222994 365588
rect 233970 365576 233976 365588
rect 234028 365576 234034 365628
rect 240318 365576 240324 365628
rect 240376 365616 240382 365628
rect 261478 365616 261484 365628
rect 240376 365588 261484 365616
rect 240376 365576 240382 365588
rect 261478 365576 261484 365588
rect 261536 365576 261542 365628
rect 278590 365576 278596 365628
rect 278648 365616 278654 365628
rect 295334 365616 295340 365628
rect 278648 365588 295340 365616
rect 278648 365576 278654 365588
rect 295334 365576 295340 365588
rect 295392 365576 295398 365628
rect 306926 365576 306932 365628
rect 306984 365616 306990 365628
rect 318058 365616 318064 365628
rect 306984 365588 318064 365616
rect 306984 365576 306990 365588
rect 318058 365576 318064 365588
rect 318116 365576 318122 365628
rect 324314 365576 324320 365628
rect 324372 365616 324378 365628
rect 345750 365616 345756 365628
rect 324372 365588 345756 365616
rect 324372 365576 324378 365588
rect 345750 365576 345756 365588
rect 345808 365576 345814 365628
rect 362862 365576 362868 365628
rect 362920 365616 362926 365628
rect 379514 365616 379520 365628
rect 362920 365588 379520 365616
rect 362920 365576 362926 365588
rect 379514 365576 379520 365588
rect 379572 365576 379578 365628
rect 390646 365576 390652 365628
rect 390704 365616 390710 365628
rect 407114 365616 407120 365628
rect 390704 365588 407120 365616
rect 390704 365576 390710 365588
rect 407114 365576 407120 365588
rect 407172 365576 407178 365628
rect 418614 365576 418620 365628
rect 418672 365616 418678 365628
rect 429838 365616 429844 365628
rect 418672 365588 429844 365616
rect 418672 365576 418678 365588
rect 429838 365576 429844 365588
rect 429896 365576 429902 365628
rect 436646 365576 436652 365628
rect 436704 365616 436710 365628
rect 457438 365616 457444 365628
rect 436704 365588 457444 365616
rect 436704 365576 436710 365588
rect 457438 365576 457444 365588
rect 457496 365576 457502 365628
rect 474642 365576 474648 365628
rect 474700 365616 474706 365628
rect 491294 365616 491300 365628
rect 474700 365588 491300 365616
rect 474700 365576 474706 365588
rect 491294 365576 491300 365588
rect 491352 365576 491358 365628
rect 502610 365576 502616 365628
rect 502668 365616 502674 365628
rect 514018 365616 514024 365628
rect 502668 365588 514024 365616
rect 502668 365576 502674 365588
rect 514018 365576 514024 365588
rect 514076 365576 514082 365628
rect 520642 365576 520648 365628
rect 520700 365616 520706 365628
rect 541618 365616 541624 365628
rect 520700 365588 541624 365616
rect 520700 365576 520706 365588
rect 541618 365576 541624 365588
rect 541676 365576 541682 365628
rect 54938 365508 54944 365560
rect 54996 365548 55002 365560
rect 71866 365548 71872 365560
rect 54996 365520 71872 365548
rect 54996 365508 55002 365520
rect 71866 365508 71872 365520
rect 71924 365508 71930 365560
rect 138934 365508 138940 365560
rect 138992 365548 138998 365560
rect 149698 365548 149704 365560
rect 138992 365520 149704 365548
rect 138992 365508 138998 365520
rect 149698 365508 149704 365520
rect 149756 365508 149762 365560
rect 250622 365508 250628 365560
rect 250680 365548 250686 365560
rect 267734 365548 267740 365560
rect 250680 365520 267740 365548
rect 250680 365508 250686 365520
rect 267734 365508 267740 365520
rect 267792 365508 267798 365560
rect 334618 365508 334624 365560
rect 334676 365548 334682 365560
rect 345658 365548 345664 365560
rect 334676 365520 345664 365548
rect 334676 365508 334682 365520
rect 345658 365508 345664 365520
rect 345716 365508 345722 365560
rect 446950 365508 446956 365560
rect 447008 365548 447014 365560
rect 463786 365548 463792 365560
rect 447008 365520 463792 365548
rect 447008 365508 447014 365520
rect 463786 365508 463792 365520
rect 463844 365508 463850 365560
rect 530946 365508 530952 365560
rect 531004 365548 531010 365560
rect 547966 365548 547972 365560
rect 531004 365520 547972 365548
rect 531004 365508 531010 365520
rect 547966 365508 547972 365520
rect 548024 365508 548030 365560
rect 558638 364964 558644 365016
rect 558696 365004 558702 365016
rect 568758 365004 568764 365016
rect 558696 364976 568764 365004
rect 558696 364964 558702 364976
rect 568758 364964 568764 364976
rect 568816 364964 568822 365016
rect 548334 363604 548340 363656
rect 548392 363644 548398 363656
rect 569034 363644 569040 363656
rect 548392 363616 569040 363644
rect 548392 363604 548398 363616
rect 569034 363604 569040 363616
rect 569092 363604 569098 363656
rect 100018 363060 100024 363112
rect 100076 363100 100082 363112
rect 121086 363100 121092 363112
rect 100076 363072 121092 363100
rect 100076 363060 100082 363072
rect 121086 363060 121092 363072
rect 121144 363060 121150 363112
rect 184014 363060 184020 363112
rect 184072 363100 184078 363112
rect 204898 363100 204904 363112
rect 184072 363072 204904 363100
rect 184072 363060 184078 363072
rect 204898 363060 204904 363072
rect 204956 363060 204962 363112
rect 464338 363060 464344 363112
rect 464396 363100 464402 363112
rect 485038 363100 485044 363112
rect 464396 363072 485044 363100
rect 464396 363060 464402 363072
rect 485038 363060 485044 363072
rect 485096 363060 485102 363112
rect 36906 362992 36912 363044
rect 36964 363032 36970 363044
rect 54294 363032 54300 363044
rect 36964 363004 54300 363032
rect 36964 362992 36970 363004
rect 54294 362992 54300 363004
rect 54352 362992 54358 363044
rect 65886 362992 65892 363044
rect 65944 363032 65950 363044
rect 81986 363032 81992 363044
rect 65944 363004 81992 363032
rect 65944 362992 65950 363004
rect 81986 362992 81992 363004
rect 82044 362992 82050 363044
rect 92842 362992 92848 363044
rect 92900 363032 92906 363044
rect 110322 363032 110328 363044
rect 92900 363004 110328 363032
rect 92900 362992 92906 363004
rect 110322 362992 110328 363004
rect 110380 362992 110386 363044
rect 176838 362992 176844 363044
rect 176896 363032 176902 363044
rect 194318 363032 194324 363044
rect 176896 363004 194324 363032
rect 176896 362992 176902 363004
rect 194318 362992 194324 363004
rect 194376 362992 194382 363044
rect 261478 362992 261484 363044
rect 261536 363032 261542 363044
rect 278314 363032 278320 363044
rect 261536 363004 278320 363032
rect 261536 362992 261542 363004
rect 278314 362992 278320 363004
rect 278372 362992 278378 363044
rect 288894 362992 288900 363044
rect 288952 363032 288958 363044
rect 306006 363032 306012 363044
rect 288952 363004 306012 363032
rect 288952 362992 288958 363004
rect 306006 362992 306012 363004
rect 306064 362992 306070 363044
rect 317138 362992 317144 363044
rect 317196 363032 317202 363044
rect 334342 363032 334348 363044
rect 317196 363004 334348 363032
rect 317196 362992 317202 363004
rect 334342 362992 334348 363004
rect 334400 362992 334406 363044
rect 372890 362992 372896 363044
rect 372948 363032 372954 363044
rect 390002 363032 390008 363044
rect 372948 363004 390008 363032
rect 372948 362992 372954 363004
rect 390002 362992 390008 363004
rect 390060 362992 390066 363044
rect 401042 362992 401048 363044
rect 401100 363032 401106 363044
rect 418338 363032 418344 363044
rect 401100 363004 418344 363032
rect 401100 362992 401106 363004
rect 418338 362992 418344 363004
rect 418396 362992 418402 363044
rect 457438 362992 457444 363044
rect 457496 363032 457502 363044
rect 473998 363032 474004 363044
rect 457496 363004 474004 363032
rect 457496 362992 457502 363004
rect 473998 362992 474004 363004
rect 474056 362992 474062 363044
rect 15286 362924 15292 362976
rect 15344 362964 15350 362976
rect 26326 362964 26332 362976
rect 15344 362936 26332 362964
rect 15344 362924 15350 362936
rect 26326 362924 26332 362936
rect 26384 362924 26390 362976
rect 38010 362924 38016 362976
rect 38068 362964 38074 362976
rect 64598 362964 64604 362976
rect 38068 362936 64604 362964
rect 38068 362924 38074 362936
rect 64598 362924 64604 362936
rect 64656 362924 64662 362976
rect 72326 362924 72332 362976
rect 72384 362964 72390 362976
rect 93118 362964 93124 362976
rect 72384 362936 93124 362964
rect 72384 362924 72390 362936
rect 93118 362924 93124 362936
rect 93176 362924 93182 362976
rect 120994 362924 121000 362976
rect 121052 362964 121058 362976
rect 138290 362964 138296 362976
rect 121052 362936 138296 362964
rect 121052 362924 121058 362936
rect 138290 362924 138296 362936
rect 138348 362924 138354 362976
rect 156322 362924 156328 362976
rect 156380 362964 156386 362976
rect 177298 362964 177304 362976
rect 156380 362936 177304 362964
rect 156380 362924 156386 362936
rect 177298 362924 177304 362936
rect 177356 362924 177362 362976
rect 204806 362924 204812 362976
rect 204864 362964 204870 362976
rect 222194 362964 222200 362976
rect 204864 362936 222200 362964
rect 204864 362924 204870 362936
rect 222194 362924 222200 362936
rect 222252 362924 222258 362976
rect 232958 362924 232964 362976
rect 233016 362964 233022 362976
rect 250346 362964 250352 362976
rect 233016 362936 250352 362964
rect 233016 362924 233022 362936
rect 250346 362924 250352 362936
rect 250404 362924 250410 362976
rect 268010 362924 268016 362976
rect 268068 362964 268074 362976
rect 289078 362964 289084 362976
rect 268068 362936 289084 362964
rect 268068 362924 268074 362936
rect 289078 362924 289084 362936
rect 289136 362924 289142 362976
rect 317046 362924 317052 362976
rect 317104 362964 317110 362976
rect 344646 362964 344652 362976
rect 317104 362936 344652 362964
rect 317104 362924 317110 362936
rect 344646 362924 344652 362936
rect 344704 362924 344710 362976
rect 352006 362924 352012 362976
rect 352064 362964 352070 362976
rect 373258 362964 373264 362976
rect 352064 362936 373264 362964
rect 352064 362924 352070 362936
rect 373258 362924 373264 362936
rect 373316 362924 373322 362976
rect 380342 362924 380348 362976
rect 380400 362964 380406 362976
rect 401134 362964 401140 362976
rect 380400 362936 401140 362964
rect 380400 362924 380406 362936
rect 401134 362924 401140 362936
rect 401192 362924 401198 362976
rect 429838 362924 429844 362976
rect 429896 362964 429902 362976
rect 456610 362964 456616 362976
rect 429896 362936 456616 362964
rect 429896 362924 429902 362936
rect 456610 362924 456616 362936
rect 456668 362924 456674 362976
rect 484946 362924 484952 362976
rect 485004 362964 485010 362976
rect 502334 362964 502340 362976
rect 485004 362936 502340 362964
rect 485004 362924 485010 362936
rect 502334 362924 502340 362936
rect 502392 362924 502398 362976
rect 512914 362924 512920 362976
rect 512972 362964 512978 362976
rect 530302 362964 530308 362976
rect 512972 362936 530308 362964
rect 512972 362924 512978 362936
rect 530302 362924 530308 362936
rect 530360 362924 530366 362976
rect 568758 360408 568764 360460
rect 568816 360408 568822 360460
rect 568776 360256 568804 360408
rect 120718 360204 120724 360256
rect 120776 360244 120782 360256
rect 120994 360244 121000 360256
rect 120776 360216 121000 360244
rect 120776 360204 120782 360216
rect 120994 360204 121000 360216
rect 121052 360204 121058 360256
rect 204714 360204 204720 360256
rect 204772 360244 204778 360256
rect 204990 360244 204996 360256
rect 204772 360216 204996 360244
rect 204772 360204 204778 360216
rect 204990 360204 204996 360216
rect 205048 360204 205054 360256
rect 400858 360204 400864 360256
rect 400916 360244 400922 360256
rect 401134 360244 401140 360256
rect 400916 360216 401140 360244
rect 400916 360204 400922 360216
rect 401134 360204 401140 360216
rect 401192 360204 401198 360256
rect 568758 360204 568764 360256
rect 568816 360204 568822 360256
rect 120810 360136 120816 360188
rect 120868 360176 120874 360188
rect 121086 360176 121092 360188
rect 120868 360148 121092 360176
rect 120868 360136 120874 360148
rect 121086 360136 121092 360148
rect 121144 360136 121150 360188
rect 316770 358844 316776 358896
rect 316828 358884 316834 358896
rect 317138 358884 317144 358896
rect 316828 358856 317144 358884
rect 316828 358844 316834 358856
rect 317138 358844 317144 358856
rect 317196 358844 317202 358896
rect 400766 358844 400772 358896
rect 400824 358884 400830 358896
rect 401042 358884 401048 358896
rect 400824 358856 401048 358884
rect 400824 358844 400830 358856
rect 401042 358844 401048 358856
rect 401100 358844 401106 358896
rect 232774 358776 232780 358828
rect 232832 358816 232838 358828
rect 232958 358816 232964 358828
rect 232832 358788 232964 358816
rect 232832 358776 232838 358788
rect 232958 358776 232964 358788
rect 233016 358776 233022 358828
rect 316862 358776 316868 358828
rect 316920 358816 316926 358828
rect 317046 358816 317052 358828
rect 316920 358788 317052 358816
rect 316920 358776 316926 358788
rect 317046 358776 317052 358788
rect 317104 358776 317110 358828
rect 36814 355376 36820 355428
rect 36872 355416 36878 355428
rect 36998 355416 37004 355428
rect 36872 355388 37004 355416
rect 36872 355376 36878 355388
rect 36998 355376 37004 355388
rect 37056 355376 37062 355428
rect 484854 355376 484860 355428
rect 484912 355376 484918 355428
rect 512822 355376 512828 355428
rect 512880 355416 512886 355428
rect 513006 355416 513012 355428
rect 512880 355388 513012 355416
rect 512880 355376 512886 355388
rect 513006 355376 513012 355388
rect 513064 355376 513070 355428
rect 484872 355224 484900 355376
rect 484854 355172 484860 355224
rect 484912 355172 484918 355224
rect 484762 352248 484768 352300
rect 484820 352288 484826 352300
rect 484946 352288 484952 352300
rect 484820 352260 484952 352288
rect 484820 352248 484826 352260
rect 484946 352248 484952 352260
rect 485004 352248 485010 352300
rect 36814 347760 36820 347812
rect 36872 347800 36878 347812
rect 36998 347800 37004 347812
rect 36872 347772 37004 347800
rect 36872 347760 36878 347772
rect 36998 347760 37004 347772
rect 37056 347760 37062 347812
rect 512822 347760 512828 347812
rect 512880 347800 512886 347812
rect 513006 347800 513012 347812
rect 512880 347772 513012 347800
rect 512880 347760 512886 347772
rect 513006 347760 513012 347772
rect 513064 347760 513070 347812
rect 92750 345652 92756 345704
rect 92808 345692 92814 345704
rect 92934 345692 92940 345704
rect 92808 345664 92940 345692
rect 92808 345652 92814 345664
rect 92934 345652 92940 345664
rect 92992 345652 92998 345704
rect 372798 345652 372804 345704
rect 372856 345692 372862 345704
rect 372982 345692 372988 345704
rect 372856 345664 372988 345692
rect 372856 345652 372862 345664
rect 372982 345652 372988 345664
rect 373040 345652 373046 345704
rect 2774 345176 2780 345228
rect 2832 345216 2838 345228
rect 5074 345216 5080 345228
rect 2832 345188 5080 345216
rect 2832 345176 2838 345188
rect 5074 345176 5080 345188
rect 5132 345176 5138 345228
rect 64874 342864 64880 342916
rect 64932 342904 64938 342916
rect 65886 342904 65892 342916
rect 64932 342876 65892 342904
rect 64932 342864 64938 342876
rect 65886 342864 65892 342876
rect 65944 342864 65950 342916
rect 93118 342864 93124 342916
rect 93176 342904 93182 342916
rect 99742 342904 99748 342916
rect 93176 342876 99748 342904
rect 93176 342864 93182 342876
rect 99742 342864 99748 342876
rect 99800 342864 99806 342916
rect 120810 342864 120816 342916
rect 120868 342904 120874 342916
rect 127710 342904 127716 342916
rect 120868 342876 127716 342904
rect 120868 342864 120874 342876
rect 127710 342864 127716 342876
rect 127768 342864 127774 342916
rect 177298 342864 177304 342916
rect 177356 342904 177362 342916
rect 183646 342904 183652 342916
rect 177356 342876 183652 342904
rect 177356 342864 177362 342876
rect 183646 342864 183652 342876
rect 183704 342864 183710 342916
rect 373258 342864 373264 342916
rect 373316 342904 373322 342916
rect 379698 342904 379704 342916
rect 373316 342876 379704 342904
rect 373316 342864 373322 342876
rect 379698 342864 379704 342876
rect 379756 342864 379762 342916
rect 400858 342864 400864 342916
rect 400916 342904 400922 342916
rect 407758 342904 407764 342916
rect 400916 342876 407764 342904
rect 400916 342864 400922 342876
rect 407758 342864 407764 342876
rect 407816 342864 407822 342916
rect 204898 342592 204904 342644
rect 204956 342632 204962 342644
rect 211706 342632 211712 342644
rect 204956 342604 211712 342632
rect 204956 342592 204962 342604
rect 211706 342592 211712 342604
rect 211764 342592 211770 342644
rect 485038 342592 485044 342644
rect 485096 342632 485102 342644
rect 491662 342632 491668 342644
rect 485096 342604 491668 342632
rect 485096 342592 485102 342604
rect 491662 342592 491668 342604
rect 491720 342592 491726 342644
rect 289078 342524 289084 342576
rect 289136 342564 289142 342576
rect 295702 342564 295708 342576
rect 289136 342536 295708 342564
rect 289136 342524 289142 342536
rect 295702 342524 295708 342536
rect 295760 342524 295766 342576
rect 288802 340892 288808 340944
rect 288860 340932 288866 340944
rect 288986 340932 288992 340944
rect 288860 340904 288992 340932
rect 288860 340892 288866 340904
rect 288986 340892 288992 340904
rect 289044 340892 289050 340944
rect 176746 340824 176752 340876
rect 176804 340864 176810 340876
rect 176930 340864 176936 340876
rect 176804 340836 176936 340864
rect 176804 340824 176810 340836
rect 176930 340824 176936 340836
rect 176988 340824 176994 340876
rect 547874 340688 547880 340740
rect 547932 340728 547938 340740
rect 548150 340728 548156 340740
rect 547932 340700 548156 340728
rect 547932 340688 547938 340700
rect 548150 340688 548156 340700
rect 548208 340688 548214 340740
rect 15286 340144 15292 340196
rect 15344 340144 15350 340196
rect 15304 339980 15332 340144
rect 15930 339980 15936 339992
rect 15304 339952 15936 339980
rect 15930 339940 15936 339952
rect 15988 339940 15994 339992
rect 15378 338036 15384 338088
rect 15436 338076 15442 338088
rect 43990 338076 43996 338088
rect 15436 338048 43996 338076
rect 15436 338036 15442 338048
rect 43990 338036 43996 338048
rect 44048 338036 44054 338088
rect 138290 338036 138296 338088
rect 138348 338076 138354 338088
rect 176930 338076 176936 338088
rect 138348 338048 176936 338076
rect 138348 338036 138354 338048
rect 176930 338036 176936 338048
rect 176988 338036 176994 338088
rect 194318 338036 194324 338088
rect 194376 338076 194382 338088
rect 232866 338076 232872 338088
rect 194376 338048 232872 338076
rect 194376 338036 194382 338048
rect 232866 338036 232872 338048
rect 232924 338036 232930 338088
rect 238846 338036 238852 338088
rect 238904 338076 238910 338088
rect 238904 338048 248414 338076
rect 238904 338036 238910 338048
rect 26326 337968 26332 338020
rect 26384 338008 26390 338020
rect 38010 338008 38016 338020
rect 26384 337980 38016 338008
rect 26384 337968 26390 337980
rect 38010 337968 38016 337980
rect 38068 337968 38074 338020
rect 42886 337968 42892 338020
rect 42944 338008 42950 338020
rect 71774 338008 71780 338020
rect 42944 337980 71780 338008
rect 42944 337968 42950 337980
rect 71774 337968 71780 337980
rect 71832 337968 71838 338020
rect 110322 337968 110328 338020
rect 110380 338008 110386 338020
rect 148778 338008 148784 338020
rect 110380 337980 148784 338008
rect 110380 337968 110386 337980
rect 148778 337968 148784 337980
rect 148836 337968 148842 338020
rect 166626 337968 166632 338020
rect 166684 338008 166690 338020
rect 204990 338008 204996 338020
rect 166684 337980 204996 338008
rect 166684 337968 166690 337980
rect 204990 337968 204996 337980
rect 205048 337968 205054 338020
rect 211246 337968 211252 338020
rect 211304 338008 211310 338020
rect 240042 338008 240048 338020
rect 211304 337980 240048 338008
rect 211304 337968 211310 337980
rect 240042 337968 240048 337980
rect 240100 337968 240106 338020
rect 248386 338008 248414 338048
rect 295426 338036 295432 338088
rect 295484 338076 295490 338088
rect 324038 338076 324044 338088
rect 295484 338048 324044 338076
rect 295484 338036 295490 338048
rect 324038 338036 324044 338048
rect 324096 338036 324102 338088
rect 334342 338036 334348 338088
rect 334400 338076 334406 338088
rect 372982 338076 372988 338088
rect 334400 338048 372988 338076
rect 334400 338036 334406 338048
rect 372982 338036 372988 338048
rect 373040 338036 373046 338088
rect 390462 338036 390468 338088
rect 390520 338076 390526 338088
rect 428734 338076 428740 338088
rect 390520 338048 428740 338076
rect 390520 338036 390526 338048
rect 428734 338036 428740 338048
rect 428792 338036 428798 338088
rect 434806 338036 434812 338088
rect 434864 338076 434870 338088
rect 434864 338048 441614 338076
rect 434864 338036 434870 338048
rect 268010 338008 268016 338020
rect 248386 337980 268016 338008
rect 268010 337968 268016 337980
rect 268068 337968 268074 338020
rect 278314 337968 278320 338020
rect 278372 338008 278378 338020
rect 316954 338008 316960 338020
rect 278372 337980 316960 338008
rect 278372 337968 278378 337980
rect 316954 337968 316960 337980
rect 317012 337968 317018 338020
rect 323026 337968 323032 338020
rect 323084 338008 323090 338020
rect 352006 338008 352012 338020
rect 323084 337980 352012 338008
rect 323084 337968 323090 337980
rect 352006 337968 352012 337980
rect 352064 337968 352070 338020
rect 362310 337968 362316 338020
rect 362368 338008 362374 338020
rect 400950 338008 400956 338020
rect 362368 337980 400956 338008
rect 362368 337968 362374 337980
rect 400950 337968 400956 337980
rect 401008 337968 401014 338020
rect 407206 337968 407212 338020
rect 407264 338008 407270 338020
rect 436002 338008 436008 338020
rect 407264 337980 436008 338008
rect 407264 337968 407270 337980
rect 436002 337968 436008 337980
rect 436060 337968 436066 338020
rect 441586 338008 441614 338048
rect 491386 338036 491392 338088
rect 491444 338076 491450 338088
rect 519998 338076 520004 338088
rect 491444 338048 520004 338076
rect 491444 338036 491450 338048
rect 519998 338036 520004 338048
rect 520056 338036 520062 338088
rect 530302 338036 530308 338088
rect 530360 338076 530366 338088
rect 568850 338076 568856 338088
rect 530360 338048 568856 338076
rect 530360 338036 530366 338048
rect 568850 338036 568856 338048
rect 568908 338036 568914 338088
rect 463694 338008 463700 338020
rect 441586 337980 463700 338008
rect 463694 337968 463700 337980
rect 463752 337968 463758 338020
rect 474642 337968 474648 338020
rect 474700 338008 474706 338020
rect 512822 338008 512828 338020
rect 474700 337980 512828 338008
rect 474700 337968 474706 337980
rect 512822 337968 512828 337980
rect 512880 337968 512886 338020
rect 548150 337968 548156 338020
rect 548208 338008 548214 338020
rect 557994 338008 558000 338020
rect 548208 337980 558000 338008
rect 548208 337968 548214 337980
rect 557994 337968 558000 337980
rect 558052 337968 558058 338020
rect 82630 337900 82636 337952
rect 82688 337940 82694 337952
rect 120902 337940 120908 337952
rect 82688 337912 120908 337940
rect 82688 337900 82694 337912
rect 120902 337900 120908 337912
rect 120960 337900 120966 337952
rect 127066 337900 127072 337952
rect 127124 337940 127130 337952
rect 156046 337940 156052 337952
rect 127124 337912 156052 337940
rect 127124 337900 127130 337912
rect 156046 337900 156052 337912
rect 156104 337900 156110 337952
rect 250346 337900 250352 337952
rect 250404 337940 250410 337952
rect 288986 337940 288992 337952
rect 250404 337912 288992 337940
rect 250404 337900 250410 337912
rect 288986 337900 288992 337912
rect 289044 337900 289050 337952
rect 306282 337900 306288 337952
rect 306340 337940 306346 337952
rect 316862 337940 316868 337952
rect 306340 337912 316868 337940
rect 306340 337900 306346 337912
rect 316862 337900 316868 337912
rect 316920 337900 316926 337952
rect 418338 337900 418344 337952
rect 418396 337940 418402 337952
rect 429838 337940 429844 337952
rect 418396 337912 429844 337940
rect 418396 337900 418402 337912
rect 429838 337900 429844 337912
rect 429896 337900 429902 337952
rect 446306 337900 446312 337952
rect 446364 337940 446370 337952
rect 484854 337940 484860 337952
rect 446364 337912 484860 337940
rect 446364 337900 446370 337912
rect 484854 337900 484860 337912
rect 484912 337900 484918 337952
rect 502334 337900 502340 337952
rect 502392 337940 502398 337952
rect 540790 337940 540796 337952
rect 502392 337912 540796 337940
rect 502392 337900 502398 337912
rect 540790 337900 540796 337912
rect 540848 337900 540854 337952
rect 54294 337832 54300 337884
rect 54352 337872 54358 337884
rect 92934 337872 92940 337884
rect 54352 337844 92940 337872
rect 54352 337832 54358 337844
rect 92934 337832 92940 337844
rect 92992 337832 92998 337884
rect 518986 337832 518992 337884
rect 519044 337872 519050 337884
rect 547874 337872 547880 337884
rect 519044 337844 547880 337872
rect 519044 337832 519050 337844
rect 547874 337832 547880 337844
rect 547932 337832 547938 337884
rect 26602 335996 26608 336048
rect 26660 336036 26666 336048
rect 36814 336036 36820 336048
rect 26660 336008 36820 336036
rect 26660 335996 26666 336008
rect 36814 335996 36820 336008
rect 36872 335996 36878 336048
rect 15378 335452 15384 335504
rect 15436 335492 15442 335504
rect 54294 335492 54300 335504
rect 15436 335464 54300 335492
rect 15436 335452 15442 335464
rect 54294 335452 54300 335464
rect 54352 335452 54358 335504
rect 429838 335452 429844 335504
rect 429896 335492 429902 335504
rect 436094 335492 436100 335504
rect 429896 335464 436100 335492
rect 429896 335452 429902 335464
rect 436094 335452 436100 335464
rect 436152 335452 436158 335504
rect 71774 335384 71780 335436
rect 71832 335424 71838 335436
rect 110598 335424 110604 335436
rect 71832 335396 110604 335424
rect 71832 335384 71838 335396
rect 110598 335384 110604 335396
rect 110656 335384 110662 335436
rect 149698 335384 149704 335436
rect 149756 335424 149762 335436
rect 156322 335424 156328 335436
rect 149756 335396 156328 335424
rect 149756 335384 149762 335396
rect 156322 335384 156328 335396
rect 156380 335384 156386 335436
rect 211154 335384 211160 335436
rect 211212 335424 211218 335436
rect 250622 335424 250628 335436
rect 211212 335396 250628 335424
rect 211212 335384 211218 335396
rect 250622 335384 250628 335396
rect 250680 335384 250686 335436
rect 267826 335384 267832 335436
rect 267884 335424 267890 335436
rect 306374 335424 306380 335436
rect 267884 335396 306380 335424
rect 267884 335384 267890 335396
rect 306374 335384 306380 335396
rect 306432 335384 306438 335436
rect 318058 335384 318064 335436
rect 318116 335424 318122 335436
rect 324314 335424 324320 335436
rect 318116 335396 324320 335424
rect 318116 335384 318122 335396
rect 324314 335384 324320 335396
rect 324372 335384 324378 335436
rect 345750 335384 345756 335436
rect 345808 335424 345814 335436
rect 362310 335424 362316 335436
rect 345808 335396 362316 335424
rect 345808 335384 345814 335396
rect 362310 335384 362316 335396
rect 362368 335384 362374 335436
rect 407206 335384 407212 335436
rect 407264 335424 407270 335436
rect 446306 335424 446312 335436
rect 407264 335396 446312 335424
rect 407264 335384 407270 335396
rect 446306 335384 446312 335396
rect 446364 335384 446370 335436
rect 457438 335384 457444 335436
rect 457496 335424 457502 335436
rect 474642 335424 474648 335436
rect 457496 335396 474648 335424
rect 457496 335384 457502 335396
rect 474642 335384 474648 335396
rect 474700 335384 474706 335436
rect 491386 335384 491392 335436
rect 491444 335424 491450 335436
rect 530302 335424 530308 335436
rect 491444 335396 530308 335424
rect 491444 335384 491450 335396
rect 530302 335384 530308 335396
rect 530360 335384 530366 335436
rect 38010 335316 38016 335368
rect 38068 335356 38074 335368
rect 44174 335356 44180 335368
rect 38068 335328 44180 335356
rect 38068 335316 38074 335328
rect 44174 335316 44180 335328
rect 44232 335316 44238 335368
rect 65886 335316 65892 335368
rect 65944 335356 65950 335368
rect 82630 335356 82636 335368
rect 65944 335328 82636 335356
rect 65944 335316 65950 335328
rect 82630 335316 82636 335328
rect 82688 335316 82694 335368
rect 99374 335316 99380 335368
rect 99432 335356 99438 335368
rect 138290 335356 138296 335368
rect 99432 335328 138296 335356
rect 99432 335316 99438 335328
rect 138290 335316 138296 335328
rect 138348 335316 138354 335368
rect 149882 335316 149888 335368
rect 149940 335356 149946 335368
rect 166626 335356 166632 335368
rect 149940 335328 166632 335356
rect 149940 335316 149946 335328
rect 166626 335316 166632 335328
rect 166684 335316 166690 335368
rect 183554 335316 183560 335368
rect 183612 335356 183618 335368
rect 222378 335356 222384 335368
rect 183612 335328 222384 335356
rect 183612 335316 183618 335328
rect 222378 335316 222384 335328
rect 222436 335316 222442 335368
rect 233970 335316 233976 335368
rect 234028 335356 234034 335368
rect 240318 335356 240324 335368
rect 234028 335328 240324 335356
rect 234028 335316 234034 335328
rect 240318 335316 240324 335328
rect 240376 335316 240382 335368
rect 261478 335316 261484 335368
rect 261536 335356 261542 335368
rect 278590 335356 278596 335368
rect 261536 335328 278596 335356
rect 261536 335316 261542 335328
rect 278590 335316 278596 335328
rect 278648 335316 278654 335368
rect 295426 335316 295432 335368
rect 295484 335356 295490 335368
rect 334618 335356 334624 335368
rect 295484 335328 334624 335356
rect 295484 335316 295490 335328
rect 334618 335316 334624 335328
rect 334676 335316 334682 335368
rect 345658 335316 345664 335368
rect 345716 335356 345722 335368
rect 352006 335356 352012 335368
rect 345716 335328 352012 335356
rect 345716 335316 345722 335328
rect 352006 335316 352012 335328
rect 352064 335316 352070 335368
rect 379606 335316 379612 335368
rect 379664 335356 379670 335368
rect 418614 335356 418620 335368
rect 379664 335328 418620 335356
rect 379664 335316 379670 335328
rect 418614 335316 418620 335328
rect 418672 335316 418678 335368
rect 463786 335316 463792 335368
rect 463844 335356 463850 335368
rect 502610 335356 502616 335368
rect 463844 335328 502616 335356
rect 463844 335316 463850 335328
rect 502610 335316 502616 335328
rect 502668 335316 502674 335368
rect 514018 335316 514024 335368
rect 514076 335356 514082 335368
rect 520274 335356 520280 335368
rect 514076 335328 520280 335356
rect 514076 335316 514082 335328
rect 520274 335316 520280 335328
rect 520332 335316 520338 335368
rect 541618 335316 541624 335368
rect 541676 335356 541682 335368
rect 558638 335356 558644 335368
rect 541676 335328 558644 335356
rect 541676 335316 541682 335328
rect 558638 335316 558644 335328
rect 558696 335316 558702 335368
rect 205082 333344 205088 333396
rect 205140 333344 205146 333396
rect 205100 333192 205128 333344
rect 345014 333208 345020 333260
rect 345072 333248 345078 333260
rect 345842 333248 345848 333260
rect 345072 333220 345848 333248
rect 345072 333208 345078 333220
rect 345842 333208 345848 333220
rect 345900 333208 345906 333260
rect 205082 333140 205088 333192
rect 205140 333140 205146 333192
rect 430574 332704 430580 332716
rect 412606 332676 430580 332704
rect 42702 332596 42708 332648
rect 42760 332636 42766 332648
rect 95234 332636 95240 332648
rect 42760 332608 95240 332636
rect 42760 332596 42766 332608
rect 95234 332596 95240 332608
rect 95292 332596 95298 332648
rect 97902 332596 97908 332648
rect 97960 332636 97966 332648
rect 150434 332636 150440 332648
rect 97960 332608 150440 332636
rect 97960 332596 97966 332608
rect 150434 332596 150440 332608
rect 150492 332596 150498 332648
rect 154482 332596 154488 332648
rect 154540 332636 154546 332648
rect 207014 332636 207020 332648
rect 154540 332608 207020 332636
rect 154540 332596 154546 332608
rect 207014 332596 207020 332608
rect 207072 332596 207078 332648
rect 209682 332596 209688 332648
rect 209740 332636 209746 332648
rect 262214 332636 262220 332648
rect 209740 332608 262220 332636
rect 209740 332596 209746 332608
rect 262214 332596 262220 332608
rect 262272 332596 262278 332648
rect 266262 332596 266268 332648
rect 266320 332636 266326 332648
rect 318794 332636 318800 332648
rect 266320 332608 318800 332636
rect 266320 332596 266326 332608
rect 318794 332596 318800 332608
rect 318852 332596 318858 332648
rect 322842 332596 322848 332648
rect 322900 332636 322906 332648
rect 375374 332636 375380 332648
rect 322900 332608 375380 332636
rect 322900 332596 322906 332608
rect 375374 332596 375380 332608
rect 375432 332596 375438 332648
rect 378042 332596 378048 332648
rect 378100 332636 378106 332648
rect 412606 332636 412634 332676
rect 430574 332664 430580 332676
rect 430632 332664 430638 332716
rect 378100 332608 412634 332636
rect 378100 332596 378106 332608
rect 429102 332596 429108 332648
rect 429160 332636 429166 332648
rect 429930 332636 429936 332648
rect 429160 332608 429936 332636
rect 429160 332596 429166 332608
rect 429930 332596 429936 332608
rect 429988 332596 429994 332648
rect 434622 332596 434628 332648
rect 434680 332636 434686 332648
rect 487154 332636 487160 332648
rect 434680 332608 487160 332636
rect 434680 332596 434686 332608
rect 487154 332596 487160 332608
rect 487212 332596 487218 332648
rect 489822 332596 489828 332648
rect 489880 332636 489886 332648
rect 542354 332636 542360 332648
rect 489880 332608 542360 332636
rect 489880 332596 489886 332608
rect 542354 332596 542360 332608
rect 542412 332596 542418 332648
rect 37274 329468 37280 329520
rect 37332 329508 37338 329520
rect 38102 329508 38108 329520
rect 37332 329480 38108 329508
rect 37332 329468 37338 329480
rect 38102 329468 38108 329480
rect 38160 329468 38166 329520
rect 149238 329468 149244 329520
rect 149296 329508 149302 329520
rect 149790 329508 149796 329520
rect 149296 329480 149796 329508
rect 149296 329468 149302 329480
rect 149790 329468 149796 329480
rect 149848 329468 149854 329520
rect 233234 329468 233240 329520
rect 233292 329508 233298 329520
rect 234062 329508 234068 329520
rect 233292 329480 234068 329508
rect 233292 329468 233298 329480
rect 234062 329468 234068 329480
rect 234120 329468 234126 329520
rect 267734 329468 267740 329520
rect 267792 329508 267798 329520
rect 267918 329508 267924 329520
rect 267792 329480 267924 329508
rect 267792 329468 267798 329480
rect 267918 329468 267924 329480
rect 267976 329468 267982 329520
rect 295334 329468 295340 329520
rect 295392 329508 295398 329520
rect 295978 329508 295984 329520
rect 295392 329480 295984 329508
rect 295392 329468 295398 329480
rect 295978 329468 295984 329480
rect 296036 329468 296042 329520
rect 379514 329468 379520 329520
rect 379572 329508 379578 329520
rect 379974 329508 379980 329520
rect 379572 329480 379980 329508
rect 379572 329468 379578 329480
rect 379974 329468 379980 329480
rect 380032 329468 380038 329520
rect 407114 329468 407120 329520
rect 407172 329508 407178 329520
rect 407942 329508 407948 329520
rect 407172 329480 407948 329508
rect 407172 329468 407178 329480
rect 407942 329468 407948 329480
rect 408000 329468 408006 329520
rect 491294 329468 491300 329520
rect 491352 329508 491358 329520
rect 492030 329508 492036 329520
rect 491352 329480 492036 329508
rect 491352 329468 491358 329480
rect 492030 329468 492036 329480
rect 492088 329468 492094 329520
rect 463694 325728 463700 325780
rect 463752 325768 463758 325780
rect 464062 325768 464068 325780
rect 463752 325740 464068 325768
rect 463752 325728 463758 325740
rect 464062 325728 464068 325740
rect 464120 325728 464126 325780
rect 574738 324300 574744 324352
rect 574796 324340 574802 324352
rect 580074 324340 580080 324352
rect 574796 324312 580080 324340
rect 574796 324300 574802 324312
rect 580074 324300 580080 324312
rect 580132 324300 580138 324352
rect 99374 314576 99380 314628
rect 99432 314616 99438 314628
rect 99926 314616 99932 314628
rect 99432 314588 99932 314616
rect 99432 314576 99438 314588
rect 99926 314576 99932 314588
rect 99984 314576 99990 314628
rect 183554 314576 183560 314628
rect 183612 314616 183618 314628
rect 184014 314616 184020 314628
rect 183612 314588 184020 314616
rect 183612 314576 183618 314588
rect 184014 314576 184020 314588
rect 184072 314576 184078 314628
rect 211154 314576 211160 314628
rect 211212 314616 211218 314628
rect 211982 314616 211988 314628
rect 211212 314588 211988 314616
rect 211212 314576 211218 314588
rect 211982 314576 211988 314588
rect 212040 314576 212046 314628
rect 71774 313420 71780 313472
rect 71832 313460 71838 313472
rect 72050 313460 72056 313472
rect 71832 313432 72056 313460
rect 71832 313420 71838 313432
rect 72050 313420 72056 313432
rect 72108 313420 72114 313472
rect 15194 311788 15200 311840
rect 15252 311828 15258 311840
rect 36906 311828 36912 311840
rect 15252 311800 36912 311828
rect 15252 311788 15258 311800
rect 36906 311788 36912 311800
rect 36964 311788 36970 311840
rect 38102 311788 38108 311840
rect 38160 311828 38166 311840
rect 64874 311828 64880 311840
rect 38160 311800 64880 311828
rect 38160 311788 38166 311800
rect 64874 311788 64880 311800
rect 64932 311788 64938 311840
rect 65058 311788 65064 311840
rect 65116 311828 65122 311840
rect 92934 311828 92940 311840
rect 65116 311800 92940 311828
rect 65116 311788 65122 311800
rect 92934 311788 92940 311800
rect 92992 311788 92998 311840
rect 93026 311788 93032 311840
rect 93084 311828 93090 311840
rect 120902 311828 120908 311840
rect 93084 311800 120908 311828
rect 93084 311788 93090 311800
rect 120902 311788 120908 311800
rect 120960 311788 120966 311840
rect 121086 311788 121092 311840
rect 121144 311828 121150 311840
rect 148594 311828 148600 311840
rect 121144 311800 148600 311828
rect 121144 311788 121150 311800
rect 148594 311788 148600 311800
rect 148652 311788 148658 311840
rect 149790 311788 149796 311840
rect 149848 311828 149854 311840
rect 176930 311828 176936 311840
rect 149848 311800 176936 311828
rect 149848 311788 149854 311800
rect 176930 311788 176936 311800
rect 176988 311788 176994 311840
rect 177022 311788 177028 311840
rect 177080 311828 177086 311840
rect 204898 311828 204904 311840
rect 177080 311800 204904 311828
rect 177080 311788 177086 311800
rect 204898 311788 204904 311800
rect 204956 311788 204962 311840
rect 205174 311788 205180 311840
rect 205232 311828 205238 311840
rect 232590 311828 232596 311840
rect 205232 311800 232596 311828
rect 205232 311788 205238 311800
rect 232590 311788 232596 311800
rect 232648 311788 232654 311840
rect 234062 311788 234068 311840
rect 234120 311828 234126 311840
rect 260926 311828 260932 311840
rect 234120 311800 260932 311828
rect 234120 311788 234126 311800
rect 260926 311788 260932 311800
rect 260984 311788 260990 311840
rect 261018 311788 261024 311840
rect 261076 311828 261082 311840
rect 288894 311828 288900 311840
rect 261076 311800 288900 311828
rect 261076 311788 261082 311800
rect 288894 311788 288900 311800
rect 288952 311788 288958 311840
rect 289078 311788 289084 311840
rect 289136 311828 289142 311840
rect 316586 311828 316592 311840
rect 289136 311800 316592 311828
rect 289136 311788 289142 311800
rect 316586 311788 316592 311800
rect 316644 311788 316650 311840
rect 317046 311788 317052 311840
rect 317104 311828 317110 311840
rect 344922 311828 344928 311840
rect 317104 311800 344928 311828
rect 317104 311788 317110 311800
rect 344922 311788 344928 311800
rect 344980 311788 344986 311840
rect 345842 311788 345848 311840
rect 345900 311828 345906 311840
rect 372614 311828 372620 311840
rect 345900 311800 372620 311828
rect 345900 311788 345906 311800
rect 372614 311788 372620 311800
rect 372672 311788 372678 311840
rect 373074 311788 373080 311840
rect 373132 311828 373138 311840
rect 400950 311828 400956 311840
rect 373132 311800 400956 311828
rect 373132 311788 373138 311800
rect 400950 311788 400956 311800
rect 401008 311788 401014 311840
rect 401042 311788 401048 311840
rect 401100 311828 401106 311840
rect 428918 311828 428924 311840
rect 401100 311800 428924 311828
rect 401100 311788 401106 311800
rect 428918 311788 428924 311800
rect 428976 311788 428982 311840
rect 429930 311788 429936 311840
rect 429988 311828 429994 311840
rect 456794 311828 456800 311840
rect 429988 311800 456800 311828
rect 429988 311788 429994 311800
rect 456794 311788 456800 311800
rect 456852 311788 456858 311840
rect 457070 311788 457076 311840
rect 457128 311828 457134 311840
rect 484946 311828 484952 311840
rect 457128 311800 484952 311828
rect 457128 311788 457134 311800
rect 484946 311788 484952 311800
rect 485004 311788 485010 311840
rect 485038 311788 485044 311840
rect 485096 311828 485102 311840
rect 512914 311828 512920 311840
rect 485096 311800 512920 311828
rect 485096 311788 485102 311800
rect 512914 311788 512920 311800
rect 512972 311788 512978 311840
rect 513098 311788 513104 311840
rect 513156 311828 513162 311840
rect 540606 311828 540612 311840
rect 513156 311800 540612 311828
rect 513156 311788 513162 311800
rect 540606 311788 540612 311800
rect 540664 311788 540670 311840
rect 541066 311788 541072 311840
rect 541124 311828 541130 311840
rect 568942 311828 568948 311840
rect 541124 311800 568948 311828
rect 541124 311788 541130 311800
rect 568942 311788 568948 311800
rect 569000 311788 569006 311840
rect 26602 311720 26608 311772
rect 26660 311760 26666 311772
rect 38010 311760 38016 311772
rect 26660 311732 38016 311760
rect 26660 311720 26666 311732
rect 38010 311720 38016 311732
rect 38068 311720 38074 311772
rect 44634 311720 44640 311772
rect 44692 311760 44698 311772
rect 65886 311760 65892 311772
rect 44692 311732 65892 311760
rect 44692 311720 44698 311732
rect 65886 311720 65892 311732
rect 65944 311720 65950 311772
rect 82630 311720 82636 311772
rect 82688 311760 82694 311772
rect 99466 311760 99472 311772
rect 82688 311732 99472 311760
rect 82688 311720 82694 311732
rect 99466 311720 99472 311732
rect 99524 311720 99530 311772
rect 128630 311720 128636 311772
rect 128688 311760 128694 311772
rect 149882 311760 149888 311772
rect 128688 311732 149888 311760
rect 128688 311720 128694 311732
rect 149882 311720 149888 311732
rect 149940 311720 149946 311772
rect 166626 311720 166632 311772
rect 166684 311760 166690 311772
rect 183646 311760 183652 311772
rect 166684 311732 183652 311760
rect 166684 311720 166690 311732
rect 183646 311720 183652 311732
rect 183704 311720 183710 311772
rect 194594 311720 194600 311772
rect 194652 311760 194658 311772
rect 211246 311760 211252 311772
rect 194652 311732 211252 311760
rect 194652 311720 194658 311732
rect 211246 311720 211252 311732
rect 211304 311720 211310 311772
rect 222930 311720 222936 311772
rect 222988 311760 222994 311772
rect 233970 311760 233976 311772
rect 222988 311732 233976 311760
rect 222988 311720 222994 311732
rect 233970 311720 233976 311732
rect 234028 311720 234034 311772
rect 240318 311720 240324 311772
rect 240376 311760 240382 311772
rect 261478 311760 261484 311772
rect 240376 311732 261484 311760
rect 240376 311720 240382 311732
rect 261478 311720 261484 311732
rect 261536 311720 261542 311772
rect 278590 311720 278596 311772
rect 278648 311760 278654 311772
rect 295334 311760 295340 311772
rect 278648 311732 295340 311760
rect 278648 311720 278654 311732
rect 295334 311720 295340 311732
rect 295392 311720 295398 311772
rect 306926 311720 306932 311772
rect 306984 311760 306990 311772
rect 318058 311760 318064 311772
rect 306984 311732 318064 311760
rect 306984 311720 306990 311732
rect 318058 311720 318064 311732
rect 318116 311720 318122 311772
rect 324314 311720 324320 311772
rect 324372 311760 324378 311772
rect 345750 311760 345756 311772
rect 324372 311732 345756 311760
rect 324372 311720 324378 311732
rect 345750 311720 345756 311732
rect 345808 311720 345814 311772
rect 362862 311720 362868 311772
rect 362920 311760 362926 311772
rect 379514 311760 379520 311772
rect 362920 311732 379520 311760
rect 362920 311720 362926 311732
rect 379514 311720 379520 311732
rect 379572 311720 379578 311772
rect 390646 311720 390652 311772
rect 390704 311760 390710 311772
rect 407114 311760 407120 311772
rect 390704 311732 407120 311760
rect 390704 311720 390710 311732
rect 407114 311720 407120 311732
rect 407172 311720 407178 311772
rect 418614 311720 418620 311772
rect 418672 311760 418678 311772
rect 429838 311760 429844 311772
rect 418672 311732 429844 311760
rect 418672 311720 418678 311732
rect 429838 311720 429844 311732
rect 429896 311720 429902 311772
rect 436646 311720 436652 311772
rect 436704 311760 436710 311772
rect 457438 311760 457444 311772
rect 436704 311732 457444 311760
rect 436704 311720 436710 311732
rect 457438 311720 457444 311732
rect 457496 311720 457502 311772
rect 474642 311720 474648 311772
rect 474700 311760 474706 311772
rect 491294 311760 491300 311772
rect 474700 311732 491300 311760
rect 474700 311720 474706 311732
rect 491294 311720 491300 311732
rect 491352 311720 491358 311772
rect 502610 311720 502616 311772
rect 502668 311760 502674 311772
rect 514018 311760 514024 311772
rect 502668 311732 514024 311760
rect 502668 311720 502674 311732
rect 514018 311720 514024 311732
rect 514076 311720 514082 311772
rect 520642 311720 520648 311772
rect 520700 311760 520706 311772
rect 541618 311760 541624 311772
rect 520700 311732 541624 311760
rect 520700 311720 520706 311732
rect 541618 311720 541624 311732
rect 541676 311720 541682 311772
rect 54938 311652 54944 311704
rect 54996 311692 55002 311704
rect 72050 311692 72056 311704
rect 54996 311664 72056 311692
rect 54996 311652 55002 311664
rect 72050 311652 72056 311664
rect 72108 311652 72114 311704
rect 138934 311652 138940 311704
rect 138992 311692 138998 311704
rect 149698 311692 149704 311704
rect 138992 311664 149704 311692
rect 138992 311652 138998 311664
rect 149698 311652 149704 311664
rect 149756 311652 149762 311704
rect 250622 311652 250628 311704
rect 250680 311692 250686 311704
rect 267734 311692 267740 311704
rect 250680 311664 267740 311692
rect 250680 311652 250686 311664
rect 267734 311652 267740 311664
rect 267792 311652 267798 311704
rect 334618 311652 334624 311704
rect 334676 311692 334682 311704
rect 345658 311692 345664 311704
rect 334676 311664 345664 311692
rect 334676 311652 334682 311664
rect 345658 311652 345664 311664
rect 345716 311652 345722 311704
rect 446950 311652 446956 311704
rect 447008 311692 447014 311704
rect 463694 311692 463700 311704
rect 447008 311664 463700 311692
rect 447008 311652 447014 311664
rect 463694 311652 463700 311664
rect 463752 311652 463758 311704
rect 530946 311652 530952 311704
rect 531004 311692 531010 311704
rect 547966 311692 547972 311704
rect 531004 311664 547972 311692
rect 531004 311652 531010 311664
rect 547966 311652 547972 311664
rect 548024 311652 548030 311704
rect 558638 311108 558644 311160
rect 558696 311148 558702 311160
rect 568942 311148 568948 311160
rect 558696 311120 568948 311148
rect 558696 311108 558702 311120
rect 568942 311108 568948 311120
rect 569000 311108 569006 311160
rect 548334 309748 548340 309800
rect 548392 309788 548398 309800
rect 569034 309788 569040 309800
rect 548392 309760 569040 309788
rect 548392 309748 548398 309760
rect 569034 309748 569040 309760
rect 569092 309748 569098 309800
rect 100018 309272 100024 309324
rect 100076 309312 100082 309324
rect 120994 309312 121000 309324
rect 100076 309284 121000 309312
rect 100076 309272 100082 309284
rect 120994 309272 121000 309284
rect 121052 309272 121058 309324
rect 268010 309272 268016 309324
rect 268068 309312 268074 309324
rect 289078 309312 289084 309324
rect 268068 309284 289084 309312
rect 268068 309272 268074 309284
rect 289078 309272 289084 309284
rect 289136 309272 289142 309324
rect 380342 309272 380348 309324
rect 380400 309312 380406 309324
rect 401042 309312 401048 309324
rect 380400 309284 401048 309312
rect 380400 309272 380406 309284
rect 401042 309272 401048 309284
rect 401100 309272 401106 309324
rect 464338 309272 464344 309324
rect 464396 309312 464402 309324
rect 485038 309312 485044 309324
rect 464396 309284 485044 309312
rect 464396 309272 464402 309284
rect 485038 309272 485044 309284
rect 485096 309272 485102 309324
rect 36906 309204 36912 309256
rect 36964 309244 36970 309256
rect 54294 309244 54300 309256
rect 36964 309216 54300 309244
rect 36964 309204 36970 309216
rect 54294 309204 54300 309216
rect 54352 309204 54358 309256
rect 65886 309204 65892 309256
rect 65944 309244 65950 309256
rect 81986 309244 81992 309256
rect 65944 309216 81992 309244
rect 65944 309204 65950 309216
rect 81986 309204 81992 309216
rect 82044 309204 82050 309256
rect 92934 309204 92940 309256
rect 92992 309244 92998 309256
rect 110322 309244 110328 309256
rect 92992 309216 110328 309244
rect 92992 309204 92998 309216
rect 110322 309204 110328 309216
rect 110380 309204 110386 309256
rect 176930 309204 176936 309256
rect 176988 309244 176994 309256
rect 194318 309244 194324 309256
rect 176988 309216 194324 309244
rect 176988 309204 176994 309216
rect 194318 309204 194324 309216
rect 194376 309204 194382 309256
rect 261478 309204 261484 309256
rect 261536 309244 261542 309256
rect 278314 309244 278320 309256
rect 261536 309216 278320 309244
rect 261536 309204 261542 309216
rect 278314 309204 278320 309216
rect 278372 309204 278378 309256
rect 317138 309204 317144 309256
rect 317196 309244 317202 309256
rect 334342 309244 334348 309256
rect 317196 309216 334348 309244
rect 317196 309204 317202 309216
rect 334342 309204 334348 309216
rect 334400 309204 334406 309256
rect 372798 309204 372804 309256
rect 372856 309244 372862 309256
rect 390002 309244 390008 309256
rect 372856 309216 390008 309244
rect 372856 309204 372862 309216
rect 390002 309204 390008 309216
rect 390060 309204 390066 309256
rect 457438 309204 457444 309256
rect 457496 309244 457502 309256
rect 473998 309244 474004 309256
rect 457496 309216 474004 309244
rect 457496 309204 457502 309216
rect 473998 309204 474004 309216
rect 474056 309204 474062 309256
rect 15194 309136 15200 309188
rect 15252 309176 15258 309188
rect 26326 309176 26332 309188
rect 15252 309148 26332 309176
rect 15252 309136 15258 309148
rect 26326 309136 26332 309148
rect 26384 309136 26390 309188
rect 38010 309136 38016 309188
rect 38068 309176 38074 309188
rect 64598 309176 64604 309188
rect 38068 309148 64604 309176
rect 38068 309136 38074 309148
rect 64598 309136 64604 309148
rect 64656 309136 64662 309188
rect 72326 309136 72332 309188
rect 72384 309176 72390 309188
rect 93118 309176 93124 309188
rect 72384 309148 93124 309176
rect 72384 309136 72390 309148
rect 93118 309136 93124 309148
rect 93176 309136 93182 309188
rect 121086 309136 121092 309188
rect 121144 309176 121150 309188
rect 138290 309176 138296 309188
rect 121144 309148 138296 309176
rect 121144 309136 121150 309148
rect 138290 309136 138296 309148
rect 138348 309136 138354 309188
rect 156322 309136 156328 309188
rect 156380 309176 156386 309188
rect 177298 309176 177304 309188
rect 156380 309148 177304 309176
rect 156380 309136 156386 309148
rect 177298 309136 177304 309148
rect 177356 309136 177362 309188
rect 184014 309136 184020 309188
rect 184072 309176 184078 309188
rect 204898 309176 204904 309188
rect 184072 309148 204904 309176
rect 184072 309136 184078 309148
rect 204898 309136 204904 309148
rect 204956 309136 204962 309188
rect 209038 309136 209044 309188
rect 209096 309176 209102 309188
rect 222194 309176 222200 309188
rect 209096 309148 222200 309176
rect 209096 309136 209102 309148
rect 222194 309136 222200 309148
rect 222252 309136 222258 309188
rect 232958 309136 232964 309188
rect 233016 309176 233022 309188
rect 250346 309176 250352 309188
rect 233016 309148 250352 309176
rect 233016 309136 233022 309148
rect 250346 309136 250352 309148
rect 250404 309136 250410 309188
rect 288802 309136 288808 309188
rect 288860 309176 288866 309188
rect 306006 309176 306012 309188
rect 288860 309148 306012 309176
rect 288860 309136 288866 309148
rect 306006 309136 306012 309148
rect 306064 309136 306070 309188
rect 317046 309136 317052 309188
rect 317104 309176 317110 309188
rect 344646 309176 344652 309188
rect 317104 309148 344652 309176
rect 317104 309136 317110 309148
rect 344646 309136 344652 309148
rect 344704 309136 344710 309188
rect 352006 309136 352012 309188
rect 352064 309176 352070 309188
rect 373258 309176 373264 309188
rect 352064 309148 373264 309176
rect 352064 309136 352070 309148
rect 373258 309136 373264 309148
rect 373316 309136 373322 309188
rect 401134 309136 401140 309188
rect 401192 309176 401198 309188
rect 418338 309176 418344 309188
rect 401192 309148 418344 309176
rect 401192 309136 401198 309148
rect 418338 309136 418344 309148
rect 418396 309136 418402 309188
rect 429838 309136 429844 309188
rect 429896 309176 429902 309188
rect 456610 309176 456616 309188
rect 429896 309148 456616 309176
rect 429896 309136 429902 309148
rect 456610 309136 456616 309148
rect 456668 309136 456674 309188
rect 484946 309136 484952 309188
rect 485004 309176 485010 309188
rect 502334 309176 502340 309188
rect 485004 309148 502340 309176
rect 485004 309136 485010 309148
rect 502334 309136 502340 309148
rect 502392 309136 502398 309188
rect 512914 309136 512920 309188
rect 512972 309176 512978 309188
rect 530302 309176 530308 309188
rect 512972 309148 530308 309176
rect 512972 309136 512978 309148
rect 530302 309136 530308 309148
rect 530360 309136 530366 309188
rect 120718 306280 120724 306332
rect 120776 306320 120782 306332
rect 121086 306320 121092 306332
rect 120776 306292 121092 306320
rect 120776 306280 120782 306292
rect 121086 306280 121092 306292
rect 121144 306280 121150 306332
rect 568850 306280 568856 306332
rect 568908 306280 568914 306332
rect 36722 306212 36728 306264
rect 36780 306252 36786 306264
rect 36906 306252 36912 306264
rect 36780 306224 36912 306252
rect 36780 306212 36786 306224
rect 36906 306212 36912 306224
rect 36964 306212 36970 306264
rect 120810 306212 120816 306264
rect 120868 306252 120874 306264
rect 120994 306252 121000 306264
rect 120868 306224 121000 306252
rect 120868 306212 120874 306224
rect 120994 306212 121000 306224
rect 121052 306212 121058 306264
rect 288710 306212 288716 306264
rect 288768 306252 288774 306264
rect 288894 306252 288900 306264
rect 288768 306224 288900 306252
rect 288768 306212 288774 306224
rect 288894 306212 288900 306224
rect 288952 306212 288958 306264
rect 568868 306128 568896 306280
rect 568850 306076 568856 306128
rect 568908 306076 568914 306128
rect 36814 305736 36820 305788
rect 36872 305736 36878 305788
rect 484762 305736 484768 305788
rect 484820 305736 484826 305788
rect 512730 305736 512736 305788
rect 512788 305736 512794 305788
rect 36832 305584 36860 305736
rect 316770 305668 316776 305720
rect 316828 305708 316834 305720
rect 317138 305708 317144 305720
rect 316828 305680 317144 305708
rect 316828 305668 316834 305680
rect 317138 305668 317144 305680
rect 317196 305668 317202 305720
rect 400766 305668 400772 305720
rect 400824 305708 400830 305720
rect 401134 305708 401140 305720
rect 400824 305680 401140 305708
rect 400824 305668 400830 305680
rect 401134 305668 401140 305680
rect 401192 305668 401198 305720
rect 36814 305532 36820 305584
rect 36872 305532 36878 305584
rect 484780 305572 484808 305736
rect 484854 305572 484860 305584
rect 484780 305544 484860 305572
rect 484854 305532 484860 305544
rect 484912 305532 484918 305584
rect 512748 305572 512776 305736
rect 512822 305572 512828 305584
rect 512748 305544 512828 305572
rect 512822 305532 512828 305544
rect 512880 305532 512886 305584
rect 512730 304580 512736 304632
rect 512788 304620 512794 304632
rect 512914 304620 512920 304632
rect 512788 304592 512920 304620
rect 512788 304580 512794 304592
rect 512914 304580 512920 304592
rect 512972 304580 512978 304632
rect 568758 304240 568764 304292
rect 568816 304280 568822 304292
rect 568942 304280 568948 304292
rect 568816 304252 568948 304280
rect 568816 304240 568822 304252
rect 568942 304240 568948 304252
rect 569000 304240 569006 304292
rect 204806 303764 204812 303816
rect 204864 303804 204870 303816
rect 204990 303804 204996 303816
rect 204864 303776 204996 303804
rect 204864 303764 204870 303776
rect 204990 303764 204996 303776
rect 205048 303764 205054 303816
rect 204806 303628 204812 303680
rect 204864 303668 204870 303680
rect 209038 303668 209044 303680
rect 204864 303640 209044 303668
rect 204864 303628 204870 303640
rect 209038 303628 209044 303640
rect 209096 303628 209102 303680
rect 484762 302676 484768 302728
rect 484820 302716 484826 302728
rect 484946 302716 484952 302728
rect 484820 302688 484952 302716
rect 484820 302676 484826 302688
rect 484946 302676 484952 302688
rect 485004 302676 485010 302728
rect 92750 301520 92756 301572
rect 92808 301560 92814 301572
rect 92934 301560 92940 301572
rect 92808 301532 92940 301560
rect 92808 301520 92814 301532
rect 92934 301520 92940 301532
rect 92992 301520 92998 301572
rect 232774 301520 232780 301572
rect 232832 301560 232838 301572
rect 232958 301560 232964 301572
rect 232832 301532 232964 301560
rect 232832 301520 232838 301532
rect 232958 301520 232964 301532
rect 233016 301520 233022 301572
rect 316862 301520 316868 301572
rect 316920 301560 316926 301572
rect 317046 301560 317052 301572
rect 316920 301532 317052 301560
rect 316920 301520 316926 301532
rect 317046 301520 317052 301532
rect 317104 301520 317110 301572
rect 372798 301520 372804 301572
rect 372856 301560 372862 301572
rect 372982 301560 372988 301572
rect 372856 301532 372988 301560
rect 372856 301520 372862 301532
rect 372982 301520 372988 301532
rect 373040 301520 373046 301572
rect 176838 297440 176844 297492
rect 176896 297440 176902 297492
rect 400950 297440 400956 297492
rect 401008 297440 401014 297492
rect 176856 297288 176884 297440
rect 400968 297288 400996 297440
rect 176838 297236 176844 297288
rect 176896 297236 176902 297288
rect 400950 297236 400956 297288
rect 401008 297236 401014 297288
rect 3142 292680 3148 292732
rect 3200 292720 3206 292732
rect 6270 292720 6276 292732
rect 3200 292692 6276 292720
rect 3200 292680 3206 292692
rect 6270 292680 6276 292692
rect 6328 292680 6334 292732
rect 176746 292476 176752 292528
rect 176804 292516 176810 292528
rect 176930 292516 176936 292528
rect 176804 292488 176936 292516
rect 176804 292476 176810 292488
rect 176930 292476 176936 292488
rect 176988 292476 176994 292528
rect 400858 292476 400864 292528
rect 400916 292516 400922 292528
rect 401042 292516 401048 292528
rect 400916 292488 401048 292516
rect 400916 292476 400922 292488
rect 401042 292476 401048 292488
rect 401100 292476 401106 292528
rect 64874 291864 64880 291916
rect 64932 291904 64938 291916
rect 65886 291904 65892 291916
rect 64932 291876 65892 291904
rect 64932 291864 64938 291876
rect 65886 291864 65892 291876
rect 65944 291864 65950 291916
rect 289078 289756 289084 289808
rect 289136 289796 289142 289808
rect 295702 289796 295708 289808
rect 289136 289768 295708 289796
rect 289136 289756 289142 289768
rect 295702 289756 295708 289768
rect 295760 289756 295766 289808
rect 93118 289076 93124 289128
rect 93176 289116 93182 289128
rect 99742 289116 99748 289128
rect 93176 289088 99748 289116
rect 93176 289076 93182 289088
rect 99742 289076 99748 289088
rect 99800 289076 99806 289128
rect 120810 289076 120816 289128
rect 120868 289116 120874 289128
rect 127710 289116 127716 289128
rect 120868 289088 127716 289116
rect 120868 289076 120874 289088
rect 127710 289076 127716 289088
rect 127768 289076 127774 289128
rect 177298 289076 177304 289128
rect 177356 289116 177362 289128
rect 183738 289116 183744 289128
rect 177356 289088 183744 289116
rect 177356 289076 177362 289088
rect 183738 289076 183744 289088
rect 183796 289076 183802 289128
rect 373258 289076 373264 289128
rect 373316 289116 373322 289128
rect 379698 289116 379704 289128
rect 373316 289088 379704 289116
rect 373316 289076 373322 289088
rect 379698 289076 379704 289088
rect 379756 289076 379762 289128
rect 400858 289076 400864 289128
rect 400916 289116 400922 289128
rect 407758 289116 407764 289128
rect 400916 289088 407764 289116
rect 400916 289076 400922 289088
rect 407758 289076 407764 289088
rect 407816 289076 407822 289128
rect 204898 288396 204904 288448
rect 204956 288436 204962 288448
rect 211706 288436 211712 288448
rect 204956 288408 211712 288436
rect 204956 288396 204962 288408
rect 211706 288396 211712 288408
rect 211764 288396 211770 288448
rect 485038 288396 485044 288448
rect 485096 288436 485102 288448
rect 491662 288436 491668 288448
rect 485096 288408 491668 288436
rect 485096 288396 485102 288408
rect 491662 288396 491668 288408
rect 491720 288396 491726 288448
rect 547874 286152 547880 286204
rect 547932 286192 547938 286204
rect 548150 286192 548156 286204
rect 547932 286164 548156 286192
rect 547932 286152 547938 286164
rect 548150 286152 548156 286164
rect 548208 286152 548214 286204
rect 15378 284248 15384 284300
rect 15436 284288 15442 284300
rect 43990 284288 43996 284300
rect 15436 284260 43996 284288
rect 15436 284248 15442 284260
rect 43990 284248 43996 284260
rect 44048 284248 44054 284300
rect 138290 284248 138296 284300
rect 138348 284288 138354 284300
rect 176838 284288 176844 284300
rect 138348 284260 176844 284288
rect 138348 284248 138354 284260
rect 176838 284248 176844 284260
rect 176896 284248 176902 284300
rect 194318 284248 194324 284300
rect 194376 284288 194382 284300
rect 232866 284288 232872 284300
rect 194376 284260 232872 284288
rect 194376 284248 194382 284260
rect 232866 284248 232872 284260
rect 232924 284248 232930 284300
rect 238846 284248 238852 284300
rect 238904 284288 238910 284300
rect 238904 284260 248414 284288
rect 238904 284248 238910 284260
rect 26326 284180 26332 284232
rect 26384 284220 26390 284232
rect 38010 284220 38016 284232
rect 26384 284192 38016 284220
rect 26384 284180 26390 284192
rect 38010 284180 38016 284192
rect 38068 284180 38074 284232
rect 42886 284180 42892 284232
rect 42944 284220 42950 284232
rect 71774 284220 71780 284232
rect 42944 284192 71780 284220
rect 42944 284180 42950 284192
rect 71774 284180 71780 284192
rect 71832 284180 71838 284232
rect 110322 284180 110328 284232
rect 110380 284220 110386 284232
rect 148778 284220 148784 284232
rect 110380 284192 148784 284220
rect 110380 284180 110386 284192
rect 148778 284180 148784 284192
rect 148836 284180 148842 284232
rect 166626 284180 166632 284232
rect 166684 284220 166690 284232
rect 204990 284220 204996 284232
rect 166684 284192 204996 284220
rect 166684 284180 166690 284192
rect 204990 284180 204996 284192
rect 205048 284180 205054 284232
rect 211246 284180 211252 284232
rect 211304 284220 211310 284232
rect 240042 284220 240048 284232
rect 211304 284192 240048 284220
rect 211304 284180 211310 284192
rect 240042 284180 240048 284192
rect 240100 284180 240106 284232
rect 248386 284220 248414 284260
rect 295426 284248 295432 284300
rect 295484 284288 295490 284300
rect 324038 284288 324044 284300
rect 295484 284260 324044 284288
rect 295484 284248 295490 284260
rect 324038 284248 324044 284260
rect 324096 284248 324102 284300
rect 334342 284248 334348 284300
rect 334400 284288 334406 284300
rect 372890 284288 372896 284300
rect 334400 284260 372896 284288
rect 334400 284248 334406 284260
rect 372890 284248 372896 284260
rect 372948 284248 372954 284300
rect 390462 284248 390468 284300
rect 390520 284288 390526 284300
rect 428734 284288 428740 284300
rect 390520 284260 428740 284288
rect 390520 284248 390526 284260
rect 428734 284248 428740 284260
rect 428792 284248 428798 284300
rect 434806 284248 434812 284300
rect 434864 284288 434870 284300
rect 434864 284260 441614 284288
rect 434864 284248 434870 284260
rect 268010 284220 268016 284232
rect 248386 284192 268016 284220
rect 268010 284180 268016 284192
rect 268068 284180 268074 284232
rect 278314 284180 278320 284232
rect 278372 284220 278378 284232
rect 316954 284220 316960 284232
rect 278372 284192 316960 284220
rect 278372 284180 278378 284192
rect 316954 284180 316960 284192
rect 317012 284180 317018 284232
rect 323026 284180 323032 284232
rect 323084 284220 323090 284232
rect 352006 284220 352012 284232
rect 323084 284192 352012 284220
rect 323084 284180 323090 284192
rect 352006 284180 352012 284192
rect 352064 284180 352070 284232
rect 362310 284180 362316 284232
rect 362368 284220 362374 284232
rect 400950 284220 400956 284232
rect 362368 284192 400956 284220
rect 362368 284180 362374 284192
rect 400950 284180 400956 284192
rect 401008 284180 401014 284232
rect 407206 284180 407212 284232
rect 407264 284220 407270 284232
rect 436002 284220 436008 284232
rect 407264 284192 436008 284220
rect 407264 284180 407270 284192
rect 436002 284180 436008 284192
rect 436060 284180 436066 284232
rect 441586 284220 441614 284260
rect 491386 284248 491392 284300
rect 491444 284288 491450 284300
rect 519998 284288 520004 284300
rect 491444 284260 520004 284288
rect 491444 284248 491450 284260
rect 519998 284248 520004 284260
rect 520056 284248 520062 284300
rect 530302 284248 530308 284300
rect 530360 284288 530366 284300
rect 568850 284288 568856 284300
rect 530360 284260 568856 284288
rect 530360 284248 530366 284260
rect 568850 284248 568856 284260
rect 568908 284248 568914 284300
rect 463694 284220 463700 284232
rect 441586 284192 463700 284220
rect 463694 284180 463700 284192
rect 463752 284180 463758 284232
rect 474642 284180 474648 284232
rect 474700 284220 474706 284232
rect 512822 284220 512828 284232
rect 474700 284192 512828 284220
rect 474700 284180 474706 284192
rect 512822 284180 512828 284192
rect 512880 284180 512886 284232
rect 518986 284180 518992 284232
rect 519044 284220 519050 284232
rect 547874 284220 547880 284232
rect 519044 284192 547880 284220
rect 519044 284180 519050 284192
rect 547874 284180 547880 284192
rect 547932 284180 547938 284232
rect 82630 284112 82636 284164
rect 82688 284152 82694 284164
rect 120902 284152 120908 284164
rect 82688 284124 120908 284152
rect 82688 284112 82694 284124
rect 120902 284112 120908 284124
rect 120960 284112 120966 284164
rect 127066 284112 127072 284164
rect 127124 284152 127130 284164
rect 156046 284152 156052 284164
rect 127124 284124 156052 284152
rect 127124 284112 127130 284124
rect 156046 284112 156052 284124
rect 156104 284112 156110 284164
rect 250346 284112 250352 284164
rect 250404 284152 250410 284164
rect 288894 284152 288900 284164
rect 250404 284124 288900 284152
rect 250404 284112 250410 284124
rect 288894 284112 288900 284124
rect 288952 284112 288958 284164
rect 306282 284112 306288 284164
rect 306340 284152 306346 284164
rect 316862 284152 316868 284164
rect 306340 284124 316868 284152
rect 306340 284112 306346 284124
rect 316862 284112 316868 284124
rect 316920 284112 316926 284164
rect 418338 284112 418344 284164
rect 418396 284152 418402 284164
rect 429838 284152 429844 284164
rect 418396 284124 429844 284152
rect 418396 284112 418402 284124
rect 429838 284112 429844 284124
rect 429896 284112 429902 284164
rect 446306 284112 446312 284164
rect 446364 284152 446370 284164
rect 484854 284152 484860 284164
rect 446364 284124 484860 284152
rect 446364 284112 446370 284124
rect 484854 284112 484860 284124
rect 484912 284112 484918 284164
rect 502334 284112 502340 284164
rect 502392 284152 502398 284164
rect 540790 284152 540796 284164
rect 502392 284124 540796 284152
rect 502392 284112 502398 284124
rect 540790 284112 540796 284124
rect 540848 284112 540854 284164
rect 548150 284112 548156 284164
rect 548208 284152 548214 284164
rect 557994 284152 558000 284164
rect 548208 284124 558000 284152
rect 548208 284112 548214 284124
rect 557994 284112 558000 284124
rect 558052 284112 558058 284164
rect 54294 284044 54300 284096
rect 54352 284084 54358 284096
rect 92842 284084 92848 284096
rect 54352 284056 92848 284084
rect 54352 284044 54358 284056
rect 92842 284044 92848 284056
rect 92900 284044 92906 284096
rect 15194 283160 15200 283212
rect 15252 283200 15258 283212
rect 16022 283200 16028 283212
rect 15252 283172 16028 283200
rect 15252 283160 15258 283172
rect 16022 283160 16028 283172
rect 16080 283160 16086 283212
rect 26602 282140 26608 282192
rect 26660 282180 26666 282192
rect 36814 282180 36820 282192
rect 26660 282152 36820 282180
rect 26660 282140 26666 282152
rect 36814 282140 36820 282152
rect 36872 282140 36878 282192
rect 38010 281596 38016 281648
rect 38068 281636 38074 281648
rect 44174 281636 44180 281648
rect 38068 281608 44180 281636
rect 38068 281596 38074 281608
rect 44174 281596 44180 281608
rect 44232 281596 44238 281648
rect 71866 281596 71872 281648
rect 71924 281636 71930 281648
rect 110598 281636 110604 281648
rect 71924 281608 110604 281636
rect 71924 281596 71930 281608
rect 110598 281596 110604 281608
rect 110656 281596 110662 281648
rect 211246 281596 211252 281648
rect 211304 281636 211310 281648
rect 250622 281636 250628 281648
rect 211304 281608 250628 281636
rect 211304 281596 211310 281608
rect 250622 281596 250628 281608
rect 250680 281596 250686 281648
rect 295426 281596 295432 281648
rect 295484 281636 295490 281648
rect 334618 281636 334624 281648
rect 295484 281608 334624 281636
rect 295484 281596 295490 281608
rect 334618 281596 334624 281608
rect 334676 281596 334682 281648
rect 407206 281596 407212 281648
rect 407264 281636 407270 281648
rect 446306 281636 446312 281648
rect 407264 281608 446312 281636
rect 407264 281596 407270 281608
rect 446306 281596 446312 281608
rect 446364 281596 446370 281648
rect 491386 281596 491392 281648
rect 491444 281636 491450 281648
rect 530302 281636 530308 281648
rect 491444 281608 530308 281636
rect 491444 281596 491450 281608
rect 530302 281596 530308 281608
rect 530360 281596 530366 281648
rect 15378 281528 15384 281580
rect 15436 281568 15442 281580
rect 54294 281568 54300 281580
rect 15436 281540 54300 281568
rect 15436 281528 15442 281540
rect 54294 281528 54300 281540
rect 54352 281528 54358 281580
rect 99466 281528 99472 281580
rect 99524 281568 99530 281580
rect 138290 281568 138296 281580
rect 99524 281540 138296 281568
rect 99524 281528 99530 281540
rect 138290 281528 138296 281540
rect 138348 281528 138354 281580
rect 149698 281528 149704 281580
rect 149756 281568 149762 281580
rect 166626 281568 166632 281580
rect 149756 281540 166632 281568
rect 149756 281528 149762 281540
rect 166626 281528 166632 281540
rect 166684 281528 166690 281580
rect 183646 281528 183652 281580
rect 183704 281568 183710 281580
rect 222286 281568 222292 281580
rect 183704 281540 222292 281568
rect 183704 281528 183710 281540
rect 222286 281528 222292 281540
rect 222344 281528 222350 281580
rect 267826 281528 267832 281580
rect 267884 281568 267890 281580
rect 306466 281568 306472 281580
rect 267884 281540 306472 281568
rect 267884 281528 267890 281540
rect 306466 281528 306472 281540
rect 306524 281528 306530 281580
rect 318058 281528 318064 281580
rect 318116 281568 318122 281580
rect 324314 281568 324320 281580
rect 318116 281540 324320 281568
rect 318116 281528 318122 281540
rect 324314 281528 324320 281540
rect 324372 281528 324378 281580
rect 345750 281528 345756 281580
rect 345808 281568 345814 281580
rect 362310 281568 362316 281580
rect 345808 281540 362316 281568
rect 345808 281528 345814 281540
rect 362310 281528 362316 281540
rect 362368 281528 362374 281580
rect 379606 281528 379612 281580
rect 379664 281568 379670 281580
rect 418614 281568 418620 281580
rect 379664 281540 418620 281568
rect 379664 281528 379670 281540
rect 418614 281528 418620 281540
rect 418672 281528 418678 281580
rect 429930 281528 429936 281580
rect 429988 281568 429994 281580
rect 436094 281568 436100 281580
rect 429988 281540 436100 281568
rect 429988 281528 429994 281540
rect 436094 281528 436100 281540
rect 436152 281528 436158 281580
rect 463786 281528 463792 281580
rect 463844 281568 463850 281580
rect 502610 281568 502616 281580
rect 463844 281540 502616 281568
rect 463844 281528 463850 281540
rect 502610 281528 502616 281540
rect 502668 281528 502674 281580
rect 541618 281528 541624 281580
rect 541676 281568 541682 281580
rect 558638 281568 558644 281580
rect 541676 281540 558644 281568
rect 541676 281528 541682 281540
rect 558638 281528 558644 281540
rect 558696 281528 558702 281580
rect 233970 280100 233976 280152
rect 234028 280140 234034 280152
rect 240134 280140 240140 280152
rect 234028 280112 240140 280140
rect 234028 280100 234034 280112
rect 240134 280100 240140 280112
rect 240192 280100 240198 280152
rect 205082 279352 205088 279404
rect 205140 279352 205146 279404
rect 205100 279200 205128 279352
rect 205082 279148 205088 279200
rect 205140 279148 205146 279200
rect 42702 278740 42708 278792
rect 42760 278780 42766 278792
rect 95234 278780 95240 278792
rect 42760 278752 95240 278780
rect 42760 278740 42766 278752
rect 95234 278740 95240 278752
rect 95292 278740 95298 278792
rect 97902 278740 97908 278792
rect 97960 278780 97966 278792
rect 150434 278780 150440 278792
rect 97960 278752 150440 278780
rect 97960 278740 97966 278752
rect 150434 278740 150440 278752
rect 150492 278740 150498 278792
rect 154482 278740 154488 278792
rect 154540 278780 154546 278792
rect 207014 278780 207020 278792
rect 154540 278752 207020 278780
rect 154540 278740 154546 278752
rect 207014 278740 207020 278752
rect 207072 278740 207078 278792
rect 209682 278740 209688 278792
rect 209740 278780 209746 278792
rect 262214 278780 262220 278792
rect 209740 278752 262220 278780
rect 209740 278740 209746 278752
rect 262214 278740 262220 278752
rect 262272 278740 262278 278792
rect 266262 278740 266268 278792
rect 266320 278780 266326 278792
rect 318794 278780 318800 278792
rect 266320 278752 318800 278780
rect 266320 278740 266326 278752
rect 318794 278740 318800 278752
rect 318852 278740 318858 278792
rect 322842 278740 322848 278792
rect 322900 278780 322906 278792
rect 375374 278780 375380 278792
rect 322900 278752 375380 278780
rect 322900 278740 322906 278752
rect 375374 278740 375380 278752
rect 375432 278740 375438 278792
rect 378042 278740 378048 278792
rect 378100 278780 378106 278792
rect 430574 278780 430580 278792
rect 378100 278752 430580 278780
rect 378100 278740 378106 278752
rect 430574 278740 430580 278752
rect 430632 278740 430638 278792
rect 434622 278740 434628 278792
rect 434680 278780 434686 278792
rect 487154 278780 487160 278792
rect 434680 278752 487160 278780
rect 434680 278740 434686 278752
rect 487154 278740 487160 278752
rect 487212 278740 487218 278792
rect 489822 278740 489828 278792
rect 489880 278780 489886 278792
rect 542354 278780 542360 278792
rect 489880 278752 542360 278780
rect 489880 278740 489886 278752
rect 542354 278740 542360 278752
rect 542412 278740 542418 278792
rect 149238 278332 149244 278384
rect 149296 278372 149302 278384
rect 149790 278372 149796 278384
rect 149296 278344 149796 278372
rect 149296 278332 149302 278344
rect 149790 278332 149796 278344
rect 149848 278332 149854 278384
rect 71774 272552 71780 272604
rect 71832 272592 71838 272604
rect 71958 272592 71964 272604
rect 71832 272564 71964 272592
rect 71832 272552 71838 272564
rect 71958 272552 71964 272564
rect 72016 272552 72022 272604
rect 99374 272552 99380 272604
rect 99432 272592 99438 272604
rect 99926 272592 99932 272604
rect 99432 272564 99932 272592
rect 99432 272552 99438 272564
rect 99926 272552 99932 272564
rect 99984 272552 99990 272604
rect 183554 272552 183560 272604
rect 183612 272592 183618 272604
rect 184014 272592 184020 272604
rect 183612 272564 184020 272592
rect 183612 272552 183618 272564
rect 184014 272552 184020 272564
rect 184072 272552 184078 272604
rect 211154 272552 211160 272604
rect 211212 272592 211218 272604
rect 211982 272592 211988 272604
rect 211212 272564 211988 272592
rect 211212 272552 211218 272564
rect 211982 272552 211988 272564
rect 212040 272552 212046 272604
rect 267734 272552 267740 272604
rect 267792 272592 267798 272604
rect 267918 272592 267924 272604
rect 267792 272564 267924 272592
rect 267792 272552 267798 272564
rect 267918 272552 267924 272564
rect 267976 272552 267982 272604
rect 295334 272552 295340 272604
rect 295392 272592 295398 272604
rect 295978 272592 295984 272604
rect 295392 272564 295984 272592
rect 295392 272552 295398 272564
rect 295978 272552 295984 272564
rect 296036 272552 296042 272604
rect 379514 272552 379520 272604
rect 379572 272592 379578 272604
rect 379974 272592 379980 272604
rect 379572 272564 379980 272592
rect 379572 272552 379578 272564
rect 379974 272552 379980 272564
rect 380032 272552 380038 272604
rect 407114 272552 407120 272604
rect 407172 272592 407178 272604
rect 407942 272592 407948 272604
rect 407172 272564 407948 272592
rect 407172 272552 407178 272564
rect 407942 272552 407948 272564
rect 408000 272552 408006 272604
rect 463694 272552 463700 272604
rect 463752 272592 463758 272604
rect 464062 272592 464068 272604
rect 463752 272564 464068 272592
rect 463752 272552 463758 272564
rect 464062 272552 464068 272564
rect 464120 272552 464126 272604
rect 491294 272552 491300 272604
rect 491352 272592 491358 272604
rect 492030 272592 492036 272604
rect 491352 272564 492036 272592
rect 491352 272552 491358 272564
rect 492030 272552 492036 272564
rect 492088 272552 492094 272604
rect 15286 256640 15292 256692
rect 15344 256680 15350 256692
rect 36906 256680 36912 256692
rect 15344 256652 36912 256680
rect 15344 256640 15350 256652
rect 36906 256640 36912 256652
rect 36964 256640 36970 256692
rect 37090 256640 37096 256692
rect 37148 256680 37154 256692
rect 64874 256680 64880 256692
rect 37148 256652 64880 256680
rect 37148 256640 37154 256652
rect 64874 256640 64880 256652
rect 64932 256640 64938 256692
rect 65058 256640 65064 256692
rect 65116 256680 65122 256692
rect 92934 256680 92940 256692
rect 65116 256652 92940 256680
rect 65116 256640 65122 256652
rect 92934 256640 92940 256652
rect 92992 256640 92998 256692
rect 93026 256640 93032 256692
rect 93084 256680 93090 256692
rect 120902 256680 120908 256692
rect 93084 256652 120908 256680
rect 93084 256640 93090 256652
rect 120902 256640 120908 256652
rect 120960 256640 120966 256692
rect 121086 256640 121092 256692
rect 121144 256680 121150 256692
rect 148594 256680 148600 256692
rect 121144 256652 148600 256680
rect 121144 256640 121150 256652
rect 148594 256640 148600 256652
rect 148652 256640 148658 256692
rect 149790 256640 149796 256692
rect 149848 256680 149854 256692
rect 176930 256680 176936 256692
rect 149848 256652 176936 256680
rect 149848 256640 149854 256652
rect 176930 256640 176936 256652
rect 176988 256640 176994 256692
rect 177022 256640 177028 256692
rect 177080 256680 177086 256692
rect 204898 256680 204904 256692
rect 177080 256652 204904 256680
rect 177080 256640 177086 256652
rect 204898 256640 204904 256652
rect 204956 256640 204962 256692
rect 205174 256640 205180 256692
rect 205232 256680 205238 256692
rect 232590 256680 232596 256692
rect 205232 256652 232596 256680
rect 205232 256640 205238 256652
rect 232590 256640 232596 256652
rect 232648 256640 232654 256692
rect 233050 256640 233056 256692
rect 233108 256680 233114 256692
rect 260926 256680 260932 256692
rect 233108 256652 260932 256680
rect 233108 256640 233114 256652
rect 260926 256640 260932 256652
rect 260984 256640 260990 256692
rect 261018 256640 261024 256692
rect 261076 256680 261082 256692
rect 288894 256680 288900 256692
rect 261076 256652 288900 256680
rect 261076 256640 261082 256652
rect 288894 256640 288900 256652
rect 288952 256640 288958 256692
rect 289078 256640 289084 256692
rect 289136 256680 289142 256692
rect 316586 256680 316592 256692
rect 289136 256652 316592 256680
rect 289136 256640 289142 256652
rect 316586 256640 316592 256652
rect 316644 256640 316650 256692
rect 317046 256640 317052 256692
rect 317104 256680 317110 256692
rect 344922 256680 344928 256692
rect 317104 256652 344928 256680
rect 317104 256640 317110 256652
rect 344922 256640 344928 256652
rect 344980 256640 344986 256692
rect 345658 256640 345664 256692
rect 345716 256680 345722 256692
rect 372614 256680 372620 256692
rect 345716 256652 372620 256680
rect 345716 256640 345722 256652
rect 372614 256640 372620 256652
rect 372672 256640 372678 256692
rect 373074 256640 373080 256692
rect 373132 256680 373138 256692
rect 400950 256680 400956 256692
rect 373132 256652 400956 256680
rect 373132 256640 373138 256652
rect 400950 256640 400956 256652
rect 401008 256640 401014 256692
rect 401042 256640 401048 256692
rect 401100 256680 401106 256692
rect 428918 256680 428924 256692
rect 401100 256652 428924 256680
rect 401100 256640 401106 256652
rect 428918 256640 428924 256652
rect 428976 256640 428982 256692
rect 429102 256640 429108 256692
rect 429160 256680 429166 256692
rect 456794 256680 456800 256692
rect 429160 256652 456800 256680
rect 429160 256640 429166 256652
rect 456794 256640 456800 256652
rect 456852 256640 456858 256692
rect 457070 256640 457076 256692
rect 457128 256680 457134 256692
rect 484946 256680 484952 256692
rect 457128 256652 484952 256680
rect 457128 256640 457134 256652
rect 484946 256640 484952 256652
rect 485004 256640 485010 256692
rect 485038 256640 485044 256692
rect 485096 256680 485102 256692
rect 512914 256680 512920 256692
rect 485096 256652 512920 256680
rect 485096 256640 485102 256652
rect 512914 256640 512920 256652
rect 512972 256640 512978 256692
rect 513098 256640 513104 256692
rect 513156 256680 513162 256692
rect 540606 256680 540612 256692
rect 513156 256652 540612 256680
rect 513156 256640 513162 256652
rect 540606 256640 540612 256652
rect 540664 256640 540670 256692
rect 541066 256640 541072 256692
rect 541124 256680 541130 256692
rect 568942 256680 568948 256692
rect 541124 256652 568948 256680
rect 541124 256640 541130 256652
rect 568942 256640 568948 256652
rect 569000 256640 569006 256692
rect 26602 256572 26608 256624
rect 26660 256612 26666 256624
rect 38010 256612 38016 256624
rect 26660 256584 38016 256612
rect 26660 256572 26666 256584
rect 38010 256572 38016 256584
rect 38068 256572 38074 256624
rect 54938 256572 54944 256624
rect 54996 256612 55002 256624
rect 71774 256612 71780 256624
rect 54996 256584 71780 256612
rect 54996 256572 55002 256584
rect 71774 256572 71780 256584
rect 71832 256572 71838 256624
rect 82630 256572 82636 256624
rect 82688 256612 82694 256624
rect 99374 256612 99380 256624
rect 82688 256584 99380 256612
rect 82688 256572 82694 256584
rect 99374 256572 99380 256584
rect 99432 256572 99438 256624
rect 128630 256572 128636 256624
rect 128688 256612 128694 256624
rect 149698 256612 149704 256624
rect 128688 256584 149704 256612
rect 128688 256572 128694 256584
rect 149698 256572 149704 256584
rect 149756 256572 149762 256624
rect 166626 256572 166632 256624
rect 166684 256612 166690 256624
rect 183554 256612 183560 256624
rect 166684 256584 183560 256612
rect 166684 256572 166690 256584
rect 183554 256572 183560 256584
rect 183612 256572 183618 256624
rect 194594 256572 194600 256624
rect 194652 256612 194658 256624
rect 211154 256612 211160 256624
rect 194652 256584 211160 256612
rect 194652 256572 194658 256584
rect 211154 256572 211160 256584
rect 211212 256572 211218 256624
rect 222930 256572 222936 256624
rect 222988 256612 222994 256624
rect 233970 256612 233976 256624
rect 222988 256584 233976 256612
rect 222988 256572 222994 256584
rect 233970 256572 233976 256584
rect 234028 256572 234034 256624
rect 250622 256572 250628 256624
rect 250680 256612 250686 256624
rect 267734 256612 267740 256624
rect 250680 256584 267740 256612
rect 250680 256572 250686 256584
rect 267734 256572 267740 256584
rect 267792 256572 267798 256624
rect 278590 256572 278596 256624
rect 278648 256612 278654 256624
rect 295334 256612 295340 256624
rect 278648 256584 295340 256612
rect 278648 256572 278654 256584
rect 295334 256572 295340 256584
rect 295392 256572 295398 256624
rect 306926 256572 306932 256624
rect 306984 256612 306990 256624
rect 318058 256612 318064 256624
rect 306984 256584 318064 256612
rect 306984 256572 306990 256584
rect 318058 256572 318064 256584
rect 318116 256572 318122 256624
rect 324314 256572 324320 256624
rect 324372 256612 324378 256624
rect 345750 256612 345756 256624
rect 324372 256584 345756 256612
rect 324372 256572 324378 256584
rect 345750 256572 345756 256584
rect 345808 256572 345814 256624
rect 362862 256572 362868 256624
rect 362920 256612 362926 256624
rect 379514 256612 379520 256624
rect 362920 256584 379520 256612
rect 362920 256572 362926 256584
rect 379514 256572 379520 256584
rect 379572 256572 379578 256624
rect 390646 256572 390652 256624
rect 390704 256612 390710 256624
rect 407114 256612 407120 256624
rect 390704 256584 407120 256612
rect 390704 256572 390710 256584
rect 407114 256572 407120 256584
rect 407172 256572 407178 256624
rect 418614 256572 418620 256624
rect 418672 256612 418678 256624
rect 429930 256612 429936 256624
rect 418672 256584 429936 256612
rect 418672 256572 418678 256584
rect 429930 256572 429936 256584
rect 429988 256572 429994 256624
rect 446950 256572 446956 256624
rect 447008 256612 447014 256624
rect 463694 256612 463700 256624
rect 447008 256584 463700 256612
rect 447008 256572 447014 256584
rect 463694 256572 463700 256584
rect 463752 256572 463758 256624
rect 474642 256572 474648 256624
rect 474700 256612 474706 256624
rect 491294 256612 491300 256624
rect 474700 256584 491300 256612
rect 474700 256572 474706 256584
rect 491294 256572 491300 256584
rect 491352 256572 491358 256624
rect 520642 256572 520648 256624
rect 520700 256612 520706 256624
rect 541618 256612 541624 256624
rect 520700 256584 541624 256612
rect 520700 256572 520706 256584
rect 541618 256572 541624 256584
rect 541676 256572 541682 256624
rect 138934 256504 138940 256556
rect 138992 256544 138998 256556
rect 155954 256544 155960 256556
rect 138992 256516 155960 256544
rect 138992 256504 138998 256516
rect 155954 256504 155960 256516
rect 156012 256504 156018 256556
rect 334618 256504 334624 256556
rect 334676 256544 334682 256556
rect 351914 256544 351920 256556
rect 334676 256516 351920 256544
rect 334676 256504 334682 256516
rect 351914 256504 351920 256516
rect 351972 256504 351978 256556
rect 530946 256504 530952 256556
rect 531004 256544 531010 256556
rect 547966 256544 547972 256556
rect 531004 256516 547972 256544
rect 531004 256504 531010 256516
rect 547966 256504 547972 256516
rect 548024 256504 548030 256556
rect 558638 256028 558644 256080
rect 558696 256068 558702 256080
rect 568942 256068 568948 256080
rect 558696 256040 568948 256068
rect 558696 256028 558702 256040
rect 568942 256028 568948 256040
rect 569000 256028 569006 256080
rect 548334 255960 548340 256012
rect 548392 256000 548398 256012
rect 569034 256000 569040 256012
rect 548392 255972 569040 256000
rect 548392 255960 548398 255972
rect 569034 255960 569040 255972
rect 569092 255960 569098 256012
rect 100018 255416 100024 255468
rect 100076 255456 100082 255468
rect 121086 255456 121092 255468
rect 100076 255428 121092 255456
rect 100076 255416 100082 255428
rect 121086 255416 121092 255428
rect 121144 255416 121150 255468
rect 268010 255416 268016 255468
rect 268068 255456 268074 255468
rect 289170 255456 289176 255468
rect 268068 255428 289176 255456
rect 268068 255416 268074 255428
rect 289170 255416 289176 255428
rect 289228 255416 289234 255468
rect 380342 255416 380348 255468
rect 380400 255456 380406 255468
rect 401134 255456 401140 255468
rect 380400 255428 401140 255456
rect 380400 255416 380406 255428
rect 401134 255416 401140 255428
rect 401192 255416 401198 255468
rect 464338 255416 464344 255468
rect 464396 255456 464402 255468
rect 485130 255456 485136 255468
rect 464396 255428 485136 255456
rect 464396 255416 464402 255428
rect 485130 255416 485136 255428
rect 485188 255416 485194 255468
rect 37642 255348 37648 255400
rect 37700 255388 37706 255400
rect 54294 255388 54300 255400
rect 37700 255360 54300 255388
rect 37700 255348 37706 255360
rect 54294 255348 54300 255360
rect 54352 255348 54358 255400
rect 65886 255348 65892 255400
rect 65944 255388 65950 255400
rect 81986 255388 81992 255400
rect 65944 255360 81992 255388
rect 65944 255348 65950 255360
rect 81986 255348 81992 255360
rect 82044 255348 82050 255400
rect 92934 255348 92940 255400
rect 92992 255388 92998 255400
rect 110322 255388 110328 255400
rect 92992 255360 110328 255388
rect 92992 255348 92998 255360
rect 110322 255348 110328 255360
rect 110380 255348 110386 255400
rect 177022 255348 177028 255400
rect 177080 255388 177086 255400
rect 194318 255388 194324 255400
rect 177080 255360 194324 255388
rect 177080 255348 177086 255360
rect 194318 255348 194324 255360
rect 194376 255348 194382 255400
rect 261478 255348 261484 255400
rect 261536 255388 261542 255400
rect 278314 255388 278320 255400
rect 261536 255360 278320 255388
rect 261536 255348 261542 255360
rect 278314 255348 278320 255360
rect 278372 255348 278378 255400
rect 317138 255348 317144 255400
rect 317196 255388 317202 255400
rect 334342 255388 334348 255400
rect 317196 255360 334348 255388
rect 317196 255348 317202 255360
rect 334342 255348 334348 255360
rect 334400 255348 334406 255400
rect 372982 255348 372988 255400
rect 373040 255388 373046 255400
rect 390002 255388 390008 255400
rect 373040 255360 390008 255388
rect 373040 255348 373046 255360
rect 390002 255348 390008 255360
rect 390060 255348 390066 255400
rect 457438 255348 457444 255400
rect 457496 255388 457502 255400
rect 473998 255388 474004 255400
rect 457496 255360 474004 255388
rect 457496 255348 457502 255360
rect 473998 255348 474004 255360
rect 474056 255348 474062 255400
rect 15194 255280 15200 255332
rect 15252 255320 15258 255332
rect 26326 255320 26332 255332
rect 15252 255292 26332 255320
rect 15252 255280 15258 255292
rect 26326 255280 26332 255292
rect 26384 255280 26390 255332
rect 38102 255280 38108 255332
rect 38160 255320 38166 255332
rect 64598 255320 64604 255332
rect 38160 255292 64604 255320
rect 38160 255280 38166 255292
rect 64598 255280 64604 255292
rect 64656 255280 64662 255332
rect 72326 255280 72332 255332
rect 72384 255320 72390 255332
rect 93118 255320 93124 255332
rect 72384 255292 93124 255320
rect 72384 255280 72390 255292
rect 93118 255280 93124 255292
rect 93176 255280 93182 255332
rect 120994 255280 121000 255332
rect 121052 255320 121058 255332
rect 138290 255320 138296 255332
rect 121052 255292 138296 255320
rect 121052 255280 121058 255292
rect 138290 255280 138296 255292
rect 138348 255280 138354 255332
rect 156322 255280 156328 255332
rect 156380 255320 156386 255332
rect 177298 255320 177304 255332
rect 156380 255292 177304 255320
rect 156380 255280 156386 255292
rect 177298 255280 177304 255292
rect 177356 255280 177362 255332
rect 184014 255280 184020 255332
rect 184072 255320 184078 255332
rect 204990 255320 204996 255332
rect 184072 255292 204996 255320
rect 184072 255280 184078 255292
rect 204990 255280 204996 255292
rect 205048 255280 205054 255332
rect 208394 255280 208400 255332
rect 208452 255320 208458 255332
rect 222194 255320 222200 255332
rect 208452 255292 222200 255320
rect 208452 255280 208458 255292
rect 222194 255280 222200 255292
rect 222252 255280 222258 255332
rect 232958 255280 232964 255332
rect 233016 255320 233022 255332
rect 250346 255320 250352 255332
rect 233016 255292 250352 255320
rect 233016 255280 233022 255292
rect 250346 255280 250352 255292
rect 250404 255280 250410 255332
rect 289078 255280 289084 255332
rect 289136 255320 289142 255332
rect 306006 255320 306012 255332
rect 289136 255292 306012 255320
rect 289136 255280 289142 255292
rect 306006 255280 306012 255292
rect 306064 255280 306070 255332
rect 317046 255280 317052 255332
rect 317104 255320 317110 255332
rect 344646 255320 344652 255332
rect 317104 255292 344652 255320
rect 317104 255280 317110 255292
rect 344646 255280 344652 255292
rect 344704 255280 344710 255332
rect 352006 255280 352012 255332
rect 352064 255320 352070 255332
rect 373258 255320 373264 255332
rect 352064 255292 373264 255320
rect 352064 255280 352070 255292
rect 373258 255280 373264 255292
rect 373316 255280 373322 255332
rect 401042 255280 401048 255332
rect 401100 255320 401106 255332
rect 418338 255320 418344 255332
rect 401100 255292 418344 255320
rect 401100 255280 401106 255292
rect 418338 255280 418344 255292
rect 418396 255280 418402 255332
rect 429838 255280 429844 255332
rect 429896 255320 429902 255332
rect 456610 255320 456616 255332
rect 429896 255292 456616 255320
rect 429896 255280 429902 255292
rect 456610 255280 456616 255292
rect 456668 255280 456674 255332
rect 485038 255280 485044 255332
rect 485096 255320 485102 255332
rect 502334 255320 502340 255332
rect 485096 255292 502340 255320
rect 485096 255280 485102 255292
rect 502334 255280 502340 255292
rect 502392 255280 502398 255332
rect 513098 255280 513104 255332
rect 513156 255320 513162 255332
rect 530302 255320 530308 255332
rect 513156 255292 530308 255320
rect 513156 255280 513162 255292
rect 530302 255280 530308 255292
rect 530360 255280 530366 255332
rect 36722 252288 36728 252340
rect 36780 252328 36786 252340
rect 37642 252328 37648 252340
rect 36780 252300 37648 252328
rect 36780 252288 36786 252300
rect 37642 252288 37648 252300
rect 37700 252288 37706 252340
rect 120718 252220 120724 252272
rect 120776 252260 120782 252272
rect 120994 252260 121000 252272
rect 120776 252232 121000 252260
rect 120776 252220 120782 252232
rect 120994 252220 121000 252232
rect 121052 252220 121058 252272
rect 204714 252220 204720 252272
rect 204772 252260 204778 252272
rect 204990 252260 204996 252272
rect 204772 252232 204996 252260
rect 204772 252220 204778 252232
rect 204990 252220 204996 252232
rect 205048 252220 205054 252272
rect 400858 252220 400864 252272
rect 400916 252260 400922 252272
rect 401134 252260 401140 252272
rect 400916 252232 401140 252260
rect 400916 252220 400922 252232
rect 401134 252220 401140 252232
rect 401192 252220 401198 252272
rect 120810 252152 120816 252204
rect 120868 252192 120874 252204
rect 121086 252192 121092 252204
rect 120868 252164 121092 252192
rect 120868 252152 120874 252164
rect 121086 252152 121092 252164
rect 121144 252152 121150 252204
rect 512730 252016 512736 252068
rect 512788 252056 512794 252068
rect 513098 252056 513104 252068
rect 512788 252028 513104 252056
rect 512788 252016 512794 252028
rect 513098 252016 513104 252028
rect 513156 252016 513162 252068
rect 316770 251880 316776 251932
rect 316828 251920 316834 251932
rect 317138 251920 317144 251932
rect 316828 251892 317144 251920
rect 316828 251880 316834 251892
rect 317138 251880 317144 251892
rect 317196 251880 317202 251932
rect 232774 251812 232780 251864
rect 232832 251852 232838 251864
rect 232958 251852 232964 251864
rect 232832 251824 232964 251852
rect 232832 251812 232838 251824
rect 232958 251812 232964 251824
rect 233016 251812 233022 251864
rect 316862 251812 316868 251864
rect 316920 251852 316926 251864
rect 317046 251852 317052 251864
rect 316920 251824 317052 251852
rect 316920 251812 316926 251824
rect 317046 251812 317052 251824
rect 317104 251812 317110 251864
rect 92750 251744 92756 251796
rect 92808 251784 92814 251796
rect 92934 251784 92940 251796
rect 92808 251756 92940 251784
rect 92808 251744 92814 251756
rect 92934 251744 92940 251756
rect 92992 251744 92998 251796
rect 176746 251336 176752 251388
rect 176804 251376 176810 251388
rect 177022 251376 177028 251388
rect 176804 251348 177028 251376
rect 176804 251336 176810 251348
rect 177022 251336 177028 251348
rect 177080 251336 177086 251388
rect 484762 251336 484768 251388
rect 484820 251376 484826 251388
rect 485038 251376 485044 251388
rect 484820 251348 485044 251376
rect 484820 251336 484826 251348
rect 485038 251336 485044 251348
rect 485096 251336 485102 251388
rect 288802 251268 288808 251320
rect 288860 251308 288866 251320
rect 289078 251308 289084 251320
rect 288860 251280 289084 251308
rect 288860 251268 288866 251280
rect 289078 251268 289084 251280
rect 289136 251268 289142 251320
rect 204806 250520 204812 250572
rect 204864 250560 204870 250572
rect 208394 250560 208400 250572
rect 204864 250532 208400 250560
rect 204864 250520 204870 250532
rect 208394 250520 208400 250532
rect 208452 250520 208458 250572
rect 372798 250112 372804 250164
rect 372856 250152 372862 250164
rect 372982 250152 372988 250164
rect 372856 250124 372988 250152
rect 372856 250112 372862 250124
rect 372982 250112 372988 250124
rect 373040 250112 373046 250164
rect 400766 249092 400772 249144
rect 400824 249132 400830 249144
rect 401042 249132 401048 249144
rect 400824 249104 401048 249132
rect 400824 249092 400830 249104
rect 401042 249092 401048 249104
rect 401100 249092 401106 249144
rect 568758 249092 568764 249144
rect 568816 249132 568822 249144
rect 568942 249132 568948 249144
rect 568816 249104 568948 249132
rect 568816 249092 568822 249104
rect 568942 249092 568948 249104
rect 569000 249092 569006 249144
rect 3234 240116 3240 240168
rect 3292 240156 3298 240168
rect 14458 240156 14464 240168
rect 3292 240128 14464 240156
rect 3292 240116 3298 240128
rect 14458 240116 14464 240128
rect 14516 240116 14522 240168
rect 64874 235696 64880 235748
rect 64932 235736 64938 235748
rect 65886 235736 65892 235748
rect 64932 235708 65892 235736
rect 64932 235696 64938 235708
rect 65886 235696 65892 235708
rect 65944 235696 65950 235748
rect 204898 235424 204904 235476
rect 204956 235464 204962 235476
rect 211706 235464 211712 235476
rect 204956 235436 211712 235464
rect 204956 235424 204962 235436
rect 211706 235424 211712 235436
rect 211764 235424 211770 235476
rect 485130 235288 485136 235340
rect 485188 235328 485194 235340
rect 491662 235328 491668 235340
rect 485188 235300 491668 235328
rect 485188 235288 485194 235300
rect 491662 235288 491668 235300
rect 491720 235288 491726 235340
rect 93118 235220 93124 235272
rect 93176 235260 93182 235272
rect 99742 235260 99748 235272
rect 93176 235232 99748 235260
rect 93176 235220 93182 235232
rect 99742 235220 99748 235232
rect 99800 235220 99806 235272
rect 120810 235220 120816 235272
rect 120868 235260 120874 235272
rect 127710 235260 127716 235272
rect 120868 235232 127716 235260
rect 120868 235220 120874 235232
rect 127710 235220 127716 235232
rect 127768 235220 127774 235272
rect 177298 235220 177304 235272
rect 177356 235260 177362 235272
rect 183646 235260 183652 235272
rect 177356 235232 183652 235260
rect 177356 235220 177362 235232
rect 183646 235220 183652 235232
rect 183704 235220 183710 235272
rect 373258 235220 373264 235272
rect 373316 235260 373322 235272
rect 379698 235260 379704 235272
rect 373316 235232 379704 235260
rect 373316 235220 373322 235232
rect 379698 235220 379704 235232
rect 379756 235220 379762 235272
rect 400858 235220 400864 235272
rect 400916 235260 400922 235272
rect 407758 235260 407764 235272
rect 400916 235232 407764 235260
rect 400916 235220 400922 235232
rect 407758 235220 407764 235232
rect 407816 235220 407822 235272
rect 289170 235016 289176 235068
rect 289228 235056 289234 235068
rect 295702 235056 295708 235068
rect 289228 235028 295708 235056
rect 289228 235016 289234 235028
rect 295702 235016 295708 235028
rect 295760 235016 295766 235068
rect 42702 233180 42708 233232
rect 42760 233220 42766 233232
rect 95234 233220 95240 233232
rect 42760 233192 95240 233220
rect 42760 233180 42766 233192
rect 95234 233180 95240 233192
rect 95292 233180 95298 233232
rect 97902 233180 97908 233232
rect 97960 233220 97966 233232
rect 150434 233220 150440 233232
rect 97960 233192 150440 233220
rect 97960 233180 97966 233192
rect 150434 233180 150440 233192
rect 150492 233180 150498 233232
rect 154482 233180 154488 233232
rect 154540 233220 154546 233232
rect 207014 233220 207020 233232
rect 154540 233192 207020 233220
rect 154540 233180 154546 233192
rect 207014 233180 207020 233192
rect 207072 233180 207078 233232
rect 209682 233180 209688 233232
rect 209740 233220 209746 233232
rect 262214 233220 262220 233232
rect 209740 233192 262220 233220
rect 209740 233180 209746 233192
rect 262214 233180 262220 233192
rect 262272 233180 262278 233232
rect 266262 233180 266268 233232
rect 266320 233220 266326 233232
rect 318794 233220 318800 233232
rect 266320 233192 318800 233220
rect 266320 233180 266326 233192
rect 318794 233180 318800 233192
rect 318852 233180 318858 233232
rect 322842 233180 322848 233232
rect 322900 233220 322906 233232
rect 375374 233220 375380 233232
rect 322900 233192 375380 233220
rect 322900 233180 322906 233192
rect 375374 233180 375380 233192
rect 375432 233180 375438 233232
rect 378042 233180 378048 233232
rect 378100 233220 378106 233232
rect 430574 233220 430580 233232
rect 378100 233192 430580 233220
rect 378100 233180 378106 233192
rect 430574 233180 430580 233192
rect 430632 233180 430638 233232
rect 434622 233180 434628 233232
rect 434680 233220 434686 233232
rect 487154 233220 487160 233232
rect 434680 233192 487160 233220
rect 434680 233180 434686 233192
rect 487154 233180 487160 233192
rect 487212 233180 487218 233232
rect 489822 233180 489828 233232
rect 489880 233220 489886 233232
rect 542354 233220 542360 233232
rect 489880 233192 542360 233220
rect 489880 233180 489886 233192
rect 542354 233180 542360 233192
rect 542412 233180 542418 233232
rect 547874 232704 547880 232756
rect 547932 232744 547938 232756
rect 548150 232744 548156 232756
rect 547932 232716 548156 232744
rect 547932 232704 547938 232716
rect 548150 232704 548156 232716
rect 548208 232704 548214 232756
rect 38010 231820 38016 231872
rect 38068 231860 38074 231872
rect 580074 231860 580080 231872
rect 38068 231832 580080 231860
rect 38068 231820 38074 231832
rect 580074 231820 580080 231832
rect 580132 231820 580138 231872
rect 15378 230392 15384 230444
rect 15436 230432 15442 230444
rect 43990 230432 43996 230444
rect 15436 230404 43996 230432
rect 15436 230392 15442 230404
rect 43990 230392 43996 230404
rect 44048 230392 44054 230444
rect 138290 230392 138296 230444
rect 138348 230432 138354 230444
rect 176838 230432 176844 230444
rect 138348 230404 176844 230432
rect 138348 230392 138354 230404
rect 176838 230392 176844 230404
rect 176896 230392 176902 230444
rect 194318 230392 194324 230444
rect 194376 230432 194382 230444
rect 232866 230432 232872 230444
rect 194376 230404 232872 230432
rect 194376 230392 194382 230404
rect 232866 230392 232872 230404
rect 232924 230392 232930 230444
rect 238846 230392 238852 230444
rect 238904 230432 238910 230444
rect 238904 230404 248414 230432
rect 238904 230392 238910 230404
rect 26326 230324 26332 230376
rect 26384 230364 26390 230376
rect 38102 230364 38108 230376
rect 26384 230336 38108 230364
rect 26384 230324 26390 230336
rect 38102 230324 38108 230336
rect 38160 230324 38166 230376
rect 42886 230324 42892 230376
rect 42944 230364 42950 230376
rect 71774 230364 71780 230376
rect 42944 230336 71780 230364
rect 42944 230324 42950 230336
rect 71774 230324 71780 230336
rect 71832 230324 71838 230376
rect 110322 230324 110328 230376
rect 110380 230364 110386 230376
rect 148778 230364 148784 230376
rect 110380 230336 148784 230364
rect 110380 230324 110386 230336
rect 148778 230324 148784 230336
rect 148836 230324 148842 230376
rect 166626 230324 166632 230376
rect 166684 230364 166690 230376
rect 204990 230364 204996 230376
rect 166684 230336 204996 230364
rect 166684 230324 166690 230336
rect 204990 230324 204996 230336
rect 205048 230324 205054 230376
rect 211246 230324 211252 230376
rect 211304 230364 211310 230376
rect 240042 230364 240048 230376
rect 211304 230336 240048 230364
rect 211304 230324 211310 230336
rect 240042 230324 240048 230336
rect 240100 230324 240106 230376
rect 248386 230364 248414 230404
rect 295426 230392 295432 230444
rect 295484 230432 295490 230444
rect 324038 230432 324044 230444
rect 295484 230404 324044 230432
rect 295484 230392 295490 230404
rect 324038 230392 324044 230404
rect 324096 230392 324102 230444
rect 334342 230392 334348 230444
rect 334400 230432 334406 230444
rect 372890 230432 372896 230444
rect 334400 230404 372896 230432
rect 334400 230392 334406 230404
rect 372890 230392 372896 230404
rect 372948 230392 372954 230444
rect 390462 230392 390468 230444
rect 390520 230432 390526 230444
rect 428734 230432 428740 230444
rect 390520 230404 428740 230432
rect 390520 230392 390526 230404
rect 428734 230392 428740 230404
rect 428792 230392 428798 230444
rect 434806 230392 434812 230444
rect 434864 230432 434870 230444
rect 434864 230404 441614 230432
rect 434864 230392 434870 230404
rect 268010 230364 268016 230376
rect 248386 230336 268016 230364
rect 268010 230324 268016 230336
rect 268068 230324 268074 230376
rect 278314 230324 278320 230376
rect 278372 230364 278378 230376
rect 316954 230364 316960 230376
rect 278372 230336 316960 230364
rect 278372 230324 278378 230336
rect 316954 230324 316960 230336
rect 317012 230324 317018 230376
rect 323026 230324 323032 230376
rect 323084 230364 323090 230376
rect 352006 230364 352012 230376
rect 323084 230336 352012 230364
rect 323084 230324 323090 230336
rect 352006 230324 352012 230336
rect 352064 230324 352070 230376
rect 362310 230324 362316 230376
rect 362368 230364 362374 230376
rect 400950 230364 400956 230376
rect 362368 230336 400956 230364
rect 362368 230324 362374 230336
rect 400950 230324 400956 230336
rect 401008 230324 401014 230376
rect 407206 230324 407212 230376
rect 407264 230364 407270 230376
rect 436002 230364 436008 230376
rect 407264 230336 436008 230364
rect 407264 230324 407270 230336
rect 436002 230324 436008 230336
rect 436060 230324 436066 230376
rect 441586 230364 441614 230404
rect 491386 230392 491392 230444
rect 491444 230432 491450 230444
rect 519998 230432 520004 230444
rect 491444 230404 520004 230432
rect 491444 230392 491450 230404
rect 519998 230392 520004 230404
rect 520056 230392 520062 230444
rect 530302 230392 530308 230444
rect 530360 230432 530366 230444
rect 568850 230432 568856 230444
rect 530360 230404 568856 230432
rect 530360 230392 530366 230404
rect 568850 230392 568856 230404
rect 568908 230392 568914 230444
rect 463694 230364 463700 230376
rect 441586 230336 463700 230364
rect 463694 230324 463700 230336
rect 463752 230324 463758 230376
rect 474642 230324 474648 230376
rect 474700 230364 474706 230376
rect 512822 230364 512828 230376
rect 474700 230336 512828 230364
rect 474700 230324 474706 230336
rect 512822 230324 512828 230336
rect 512880 230324 512886 230376
rect 548150 230324 548156 230376
rect 548208 230364 548214 230376
rect 557994 230364 558000 230376
rect 548208 230336 558000 230364
rect 548208 230324 548214 230336
rect 557994 230324 558000 230336
rect 558052 230324 558058 230376
rect 82630 230256 82636 230308
rect 82688 230296 82694 230308
rect 120902 230296 120908 230308
rect 82688 230268 120908 230296
rect 82688 230256 82694 230268
rect 120902 230256 120908 230268
rect 120960 230256 120966 230308
rect 127066 230256 127072 230308
rect 127124 230296 127130 230308
rect 156046 230296 156052 230308
rect 127124 230268 156052 230296
rect 127124 230256 127130 230268
rect 156046 230256 156052 230268
rect 156104 230256 156110 230308
rect 250346 230256 250352 230308
rect 250404 230296 250410 230308
rect 288894 230296 288900 230308
rect 250404 230268 288900 230296
rect 250404 230256 250410 230268
rect 288894 230256 288900 230268
rect 288952 230256 288958 230308
rect 306282 230256 306288 230308
rect 306340 230296 306346 230308
rect 316862 230296 316868 230308
rect 306340 230268 316868 230296
rect 306340 230256 306346 230268
rect 316862 230256 316868 230268
rect 316920 230256 316926 230308
rect 418338 230256 418344 230308
rect 418396 230296 418402 230308
rect 429838 230296 429844 230308
rect 418396 230268 429844 230296
rect 418396 230256 418402 230268
rect 429838 230256 429844 230268
rect 429896 230256 429902 230308
rect 446306 230256 446312 230308
rect 446364 230296 446370 230308
rect 484854 230296 484860 230308
rect 446364 230268 484860 230296
rect 446364 230256 446370 230268
rect 484854 230256 484860 230268
rect 484912 230256 484918 230308
rect 502334 230256 502340 230308
rect 502392 230296 502398 230308
rect 540790 230296 540796 230308
rect 502392 230268 540796 230296
rect 502392 230256 502398 230268
rect 540790 230256 540796 230268
rect 540848 230256 540854 230308
rect 54294 230188 54300 230240
rect 54352 230228 54358 230240
rect 92842 230228 92848 230240
rect 54352 230200 92848 230228
rect 54352 230188 54358 230200
rect 92842 230188 92848 230200
rect 92900 230188 92906 230240
rect 518986 230188 518992 230240
rect 519044 230228 519050 230240
rect 547874 230228 547880 230240
rect 519044 230200 547880 230228
rect 519044 230188 519050 230200
rect 547874 230188 547880 230200
rect 547932 230188 547938 230240
rect 26602 228352 26608 228404
rect 26660 228392 26666 228404
rect 36814 228392 36820 228404
rect 26660 228364 36820 228392
rect 26660 228352 26666 228364
rect 36814 228352 36820 228364
rect 36872 228352 36878 228404
rect 15930 227876 15936 227928
rect 15988 227916 15994 227928
rect 54294 227916 54300 227928
rect 15988 227888 54300 227916
rect 15988 227876 15994 227888
rect 54294 227876 54300 227888
rect 54352 227876 54358 227928
rect 149698 227876 149704 227928
rect 149756 227916 149762 227928
rect 166626 227916 166632 227928
rect 149756 227888 166632 227916
rect 149756 227876 149762 227888
rect 166626 227876 166632 227888
rect 166684 227876 166690 227928
rect 407850 227876 407856 227928
rect 407908 227916 407914 227928
rect 446306 227916 446312 227928
rect 407908 227888 446312 227916
rect 407908 227876 407914 227888
rect 446306 227876 446312 227888
rect 446364 227876 446370 227928
rect 491938 227876 491944 227928
rect 491996 227916 492002 227928
rect 491996 227888 499574 227916
rect 491996 227876 492002 227888
rect 65886 227808 65892 227860
rect 65944 227848 65950 227860
rect 82630 227848 82636 227860
rect 65944 227820 82636 227848
rect 65944 227808 65950 227820
rect 82630 227808 82636 227820
rect 82688 227808 82694 227860
rect 99834 227808 99840 227860
rect 99892 227848 99898 227860
rect 138290 227848 138296 227860
rect 99892 227820 138296 227848
rect 99892 227808 99898 227820
rect 138290 227808 138296 227820
rect 138348 227808 138354 227860
rect 149882 227808 149888 227860
rect 149940 227848 149946 227860
rect 156322 227848 156328 227860
rect 149940 227820 156328 227848
rect 149940 227808 149946 227820
rect 156322 227808 156328 227820
rect 156380 227808 156386 227860
rect 211890 227808 211896 227860
rect 211948 227848 211954 227860
rect 250622 227848 250628 227860
rect 211948 227820 250628 227848
rect 211948 227808 211954 227820
rect 250622 227808 250628 227820
rect 250680 227808 250686 227860
rect 261478 227808 261484 227860
rect 261536 227848 261542 227860
rect 278590 227848 278596 227860
rect 261536 227820 278596 227848
rect 261536 227808 261542 227820
rect 278590 227808 278596 227820
rect 278648 227808 278654 227860
rect 295886 227808 295892 227860
rect 295944 227848 295950 227860
rect 334618 227848 334624 227860
rect 295944 227820 334624 227848
rect 295944 227808 295950 227820
rect 334618 227808 334624 227820
rect 334676 227808 334682 227860
rect 379882 227808 379888 227860
rect 379940 227848 379946 227860
rect 418614 227848 418620 227860
rect 379940 227820 418620 227848
rect 379940 227808 379946 227820
rect 418614 227808 418620 227820
rect 418672 227808 418678 227860
rect 429838 227808 429844 227860
rect 429896 227848 429902 227860
rect 436094 227848 436100 227860
rect 429896 227820 436100 227848
rect 429896 227808 429902 227820
rect 436094 227808 436100 227820
rect 436152 227808 436158 227860
rect 458818 227808 458824 227860
rect 458876 227848 458882 227860
rect 474642 227848 474648 227860
rect 458876 227820 474648 227848
rect 458876 227808 458882 227820
rect 474642 227808 474648 227820
rect 474700 227808 474706 227860
rect 486418 227808 486424 227860
rect 486476 227848 486482 227860
rect 492306 227848 492312 227860
rect 486476 227820 492312 227848
rect 486476 227808 486482 227820
rect 492306 227808 492312 227820
rect 492364 227808 492370 227860
rect 499546 227848 499574 227888
rect 530302 227848 530308 227860
rect 499546 227820 530308 227848
rect 530302 227808 530308 227820
rect 530360 227808 530366 227860
rect 38102 227740 38108 227792
rect 38160 227780 38166 227792
rect 44174 227780 44180 227792
rect 38160 227752 44180 227780
rect 38160 227740 38166 227752
rect 44174 227740 44180 227752
rect 44232 227740 44238 227792
rect 71866 227740 71872 227792
rect 71924 227780 71930 227792
rect 110598 227780 110604 227792
rect 71924 227752 110604 227780
rect 71924 227740 71930 227752
rect 110598 227740 110604 227752
rect 110656 227740 110662 227792
rect 183922 227740 183928 227792
rect 183980 227780 183986 227792
rect 222286 227780 222292 227792
rect 183980 227752 222292 227780
rect 183980 227740 183986 227752
rect 222286 227740 222292 227752
rect 222344 227740 222350 227792
rect 233970 227740 233976 227792
rect 234028 227780 234034 227792
rect 240318 227780 240324 227792
rect 234028 227752 240324 227780
rect 234028 227740 234034 227752
rect 240318 227740 240324 227752
rect 240376 227740 240382 227792
rect 267826 227740 267832 227792
rect 267884 227780 267890 227792
rect 306466 227780 306472 227792
rect 267884 227752 306472 227780
rect 267884 227740 267890 227752
rect 306466 227740 306472 227752
rect 306524 227740 306530 227792
rect 318058 227740 318064 227792
rect 318116 227780 318122 227792
rect 324314 227780 324320 227792
rect 318116 227752 324320 227780
rect 318116 227740 318122 227752
rect 324314 227740 324320 227752
rect 324372 227740 324378 227792
rect 345658 227740 345664 227792
rect 345716 227780 345722 227792
rect 362310 227780 362316 227792
rect 345716 227752 362316 227780
rect 345716 227740 345722 227752
rect 362310 227740 362316 227752
rect 362368 227740 362374 227792
rect 378870 227740 378876 227792
rect 378928 227780 378934 227792
rect 390646 227780 390652 227792
rect 378928 227752 390652 227780
rect 378928 227740 378934 227752
rect 390646 227740 390652 227752
rect 390704 227740 390710 227792
rect 402238 227740 402244 227792
rect 402296 227780 402302 227792
rect 408310 227780 408316 227792
rect 402296 227752 408316 227780
rect 402296 227740 402302 227752
rect 408310 227740 408316 227752
rect 408368 227740 408374 227792
rect 460198 227740 460204 227792
rect 460256 227780 460262 227792
rect 464338 227780 464344 227792
rect 460256 227752 464344 227780
rect 460256 227740 460262 227752
rect 464338 227740 464344 227752
rect 464396 227740 464402 227792
rect 502610 227780 502616 227792
rect 464448 227752 502616 227780
rect 463970 227672 463976 227724
rect 464028 227712 464034 227724
rect 464448 227712 464476 227752
rect 502610 227740 502616 227752
rect 502668 227740 502674 227792
rect 514018 227740 514024 227792
rect 514076 227780 514082 227792
rect 520274 227780 520280 227792
rect 514076 227752 520280 227780
rect 514076 227740 514082 227752
rect 520274 227740 520280 227752
rect 520332 227740 520338 227792
rect 541618 227740 541624 227792
rect 541676 227780 541682 227792
rect 558638 227780 558644 227792
rect 541676 227752 558644 227780
rect 541676 227740 541682 227752
rect 558638 227740 558644 227752
rect 558696 227740 558702 227792
rect 464028 227684 464476 227712
rect 464028 227672 464034 227684
rect 15194 227128 15200 227180
rect 15252 227168 15258 227180
rect 16022 227168 16028 227180
rect 15252 227140 16028 227168
rect 15252 227128 15258 227140
rect 16022 227128 16028 227140
rect 16080 227128 16086 227180
rect 205082 225360 205088 225412
rect 205140 225360 205146 225412
rect 205100 225208 205128 225360
rect 345014 225224 345020 225276
rect 345072 225264 345078 225276
rect 347038 225264 347044 225276
rect 345072 225236 347044 225264
rect 345072 225224 345078 225236
rect 347038 225224 347044 225236
rect 347096 225224 347102 225276
rect 205082 225156 205088 225208
rect 205140 225156 205146 225208
rect 434622 225088 434628 225140
rect 434680 225128 434686 225140
rect 487154 225128 487160 225140
rect 434680 225100 487160 225128
rect 434680 225088 434686 225100
rect 487154 225088 487160 225100
rect 487212 225088 487218 225140
rect 322842 225020 322848 225072
rect 322900 225060 322906 225072
rect 375374 225060 375380 225072
rect 322900 225032 375380 225060
rect 322900 225020 322906 225032
rect 375374 225020 375380 225032
rect 375432 225020 375438 225072
rect 405642 225020 405648 225072
rect 405700 225060 405706 225072
rect 458174 225060 458180 225072
rect 405700 225032 458180 225060
rect 405700 225020 405706 225032
rect 458174 225020 458180 225032
rect 458232 225020 458238 225072
rect 293862 224952 293868 225004
rect 293920 224992 293926 225004
rect 346394 224992 346400 225004
rect 293920 224964 346400 224992
rect 293920 224952 293926 224964
rect 346394 224952 346400 224964
rect 346452 224952 346458 225004
rect 348418 224952 348424 225004
rect 348476 224992 348482 225004
rect 352006 224992 352012 225004
rect 348476 224964 352012 224992
rect 348476 224952 348482 224964
rect 352006 224952 352012 224964
rect 352064 224952 352070 225004
rect 429102 224952 429108 225004
rect 429160 224992 429166 225004
rect 429930 224992 429936 225004
rect 429160 224964 429936 224992
rect 429160 224952 429166 224964
rect 429930 224952 429936 224964
rect 429988 224952 429994 225004
rect 37274 222300 37280 222352
rect 37332 222340 37338 222352
rect 38194 222340 38200 222352
rect 37332 222312 38200 222340
rect 37332 222300 37338 222312
rect 38194 222300 38200 222312
rect 38252 222300 38258 222352
rect 99374 222300 99380 222352
rect 99432 222340 99438 222352
rect 99926 222340 99932 222352
rect 99432 222312 99932 222340
rect 99432 222300 99438 222312
rect 99926 222300 99932 222312
rect 99984 222300 99990 222352
rect 183554 222300 183560 222352
rect 183612 222340 183618 222352
rect 184014 222340 184020 222352
rect 183612 222312 184020 222340
rect 183612 222300 183618 222312
rect 184014 222300 184020 222312
rect 184072 222300 184078 222352
rect 211154 222300 211160 222352
rect 211212 222340 211218 222352
rect 211982 222340 211988 222352
rect 211212 222312 211988 222340
rect 211212 222300 211218 222312
rect 211982 222300 211988 222312
rect 212040 222300 212046 222352
rect 267734 222300 267740 222352
rect 267792 222340 267798 222352
rect 267918 222340 267924 222352
rect 267792 222312 267924 222340
rect 267792 222300 267798 222312
rect 267918 222300 267924 222312
rect 267976 222300 267982 222352
rect 295334 222300 295340 222352
rect 295392 222340 295398 222352
rect 295978 222340 295984 222352
rect 295392 222312 295984 222340
rect 295392 222300 295398 222312
rect 295978 222300 295984 222312
rect 296036 222300 296042 222352
rect 379514 222300 379520 222352
rect 379572 222340 379578 222352
rect 379974 222340 379980 222352
rect 379572 222312 379980 222340
rect 379572 222300 379578 222312
rect 379974 222300 379980 222312
rect 380032 222300 380038 222352
rect 71774 221008 71780 221060
rect 71832 221048 71838 221060
rect 71958 221048 71964 221060
rect 71832 221020 71964 221048
rect 71832 221008 71838 221020
rect 71958 221008 71964 221020
rect 72016 221008 72022 221060
rect 233234 220668 233240 220720
rect 233292 220708 233298 220720
rect 234062 220708 234068 220720
rect 233292 220680 234068 220708
rect 233292 220668 233298 220680
rect 234062 220668 234068 220680
rect 234120 220668 234126 220720
rect 149238 220056 149244 220108
rect 149296 220096 149302 220108
rect 149790 220096 149796 220108
rect 149296 220068 149796 220096
rect 149296 220056 149302 220068
rect 149790 220056 149796 220068
rect 149848 220056 149854 220108
rect 15286 202784 15292 202836
rect 15344 202824 15350 202836
rect 36906 202824 36912 202836
rect 15344 202796 36912 202824
rect 15344 202784 15350 202796
rect 36906 202784 36912 202796
rect 36964 202784 36970 202836
rect 38194 202784 38200 202836
rect 38252 202824 38258 202836
rect 64874 202824 64880 202836
rect 38252 202796 64880 202824
rect 38252 202784 38258 202796
rect 64874 202784 64880 202796
rect 64932 202784 64938 202836
rect 65058 202784 65064 202836
rect 65116 202824 65122 202836
rect 92934 202824 92940 202836
rect 65116 202796 92940 202824
rect 65116 202784 65122 202796
rect 92934 202784 92940 202796
rect 92992 202784 92998 202836
rect 93026 202784 93032 202836
rect 93084 202824 93090 202836
rect 120902 202824 120908 202836
rect 93084 202796 120908 202824
rect 93084 202784 93090 202796
rect 120902 202784 120908 202796
rect 120960 202784 120966 202836
rect 121086 202784 121092 202836
rect 121144 202824 121150 202836
rect 148594 202824 148600 202836
rect 121144 202796 148600 202824
rect 121144 202784 121150 202796
rect 148594 202784 148600 202796
rect 148652 202784 148658 202836
rect 149790 202784 149796 202836
rect 149848 202824 149854 202836
rect 176930 202824 176936 202836
rect 149848 202796 176936 202824
rect 149848 202784 149854 202796
rect 176930 202784 176936 202796
rect 176988 202784 176994 202836
rect 177022 202784 177028 202836
rect 177080 202824 177086 202836
rect 204622 202824 204628 202836
rect 177080 202796 204628 202824
rect 177080 202784 177086 202796
rect 204622 202784 204628 202796
rect 204680 202784 204686 202836
rect 205174 202784 205180 202836
rect 205232 202824 205238 202836
rect 232590 202824 232596 202836
rect 205232 202796 232596 202824
rect 205232 202784 205238 202796
rect 232590 202784 232596 202796
rect 232648 202784 232654 202836
rect 234062 202784 234068 202836
rect 234120 202824 234126 202836
rect 260926 202824 260932 202836
rect 234120 202796 260932 202824
rect 234120 202784 234126 202796
rect 260926 202784 260932 202796
rect 260984 202784 260990 202836
rect 261018 202784 261024 202836
rect 261076 202824 261082 202836
rect 288526 202824 288532 202836
rect 261076 202796 288532 202824
rect 261076 202784 261082 202796
rect 288526 202784 288532 202796
rect 288584 202784 288590 202836
rect 289078 202784 289084 202836
rect 289136 202824 289142 202836
rect 316586 202824 316592 202836
rect 289136 202796 316592 202824
rect 289136 202784 289142 202796
rect 316586 202784 316592 202796
rect 316644 202784 316650 202836
rect 317046 202784 317052 202836
rect 317104 202824 317110 202836
rect 344922 202824 344928 202836
rect 317104 202796 344928 202824
rect 317104 202784 317110 202796
rect 344922 202784 344928 202796
rect 344980 202784 344986 202836
rect 347038 202784 347044 202836
rect 347096 202824 347102 202836
rect 372614 202824 372620 202836
rect 347096 202796 372620 202824
rect 347096 202784 347102 202796
rect 372614 202784 372620 202796
rect 372672 202784 372678 202836
rect 373074 202784 373080 202836
rect 373132 202824 373138 202836
rect 400582 202824 400588 202836
rect 373132 202796 400588 202824
rect 373132 202784 373138 202796
rect 400582 202784 400588 202796
rect 400640 202784 400646 202836
rect 401042 202784 401048 202836
rect 401100 202824 401106 202836
rect 428918 202824 428924 202836
rect 401100 202796 428924 202824
rect 401100 202784 401106 202796
rect 428918 202784 428924 202796
rect 428976 202784 428982 202836
rect 429930 202784 429936 202836
rect 429988 202824 429994 202836
rect 456794 202824 456800 202836
rect 429988 202796 456800 202824
rect 429988 202784 429994 202796
rect 456794 202784 456800 202796
rect 456852 202784 456858 202836
rect 457070 202784 457076 202836
rect 457128 202824 457134 202836
rect 484670 202824 484676 202836
rect 457128 202796 484676 202824
rect 457128 202784 457134 202796
rect 484670 202784 484676 202796
rect 484728 202784 484734 202836
rect 485038 202784 485044 202836
rect 485096 202824 485102 202836
rect 512914 202824 512920 202836
rect 485096 202796 512920 202824
rect 485096 202784 485102 202796
rect 512914 202784 512920 202796
rect 512972 202784 512978 202836
rect 513098 202784 513104 202836
rect 513156 202824 513162 202836
rect 540606 202824 540612 202836
rect 513156 202796 540612 202824
rect 513156 202784 513162 202796
rect 540606 202784 540612 202796
rect 540664 202784 540670 202836
rect 541066 202784 541072 202836
rect 541124 202824 541130 202836
rect 568942 202824 568948 202836
rect 541124 202796 568948 202824
rect 541124 202784 541130 202796
rect 568942 202784 568948 202796
rect 569000 202784 569006 202836
rect 26602 202716 26608 202768
rect 26660 202756 26666 202768
rect 38102 202756 38108 202768
rect 26660 202728 38108 202756
rect 26660 202716 26666 202728
rect 38102 202716 38108 202728
rect 38160 202716 38166 202768
rect 44634 202716 44640 202768
rect 44692 202756 44698 202768
rect 65886 202756 65892 202768
rect 44692 202728 65892 202756
rect 44692 202716 44698 202728
rect 65886 202716 65892 202728
rect 65944 202716 65950 202768
rect 82630 202716 82636 202768
rect 82688 202756 82694 202768
rect 99374 202756 99380 202768
rect 82688 202728 99380 202756
rect 82688 202716 82694 202728
rect 99374 202716 99380 202728
rect 99432 202716 99438 202768
rect 128630 202716 128636 202768
rect 128688 202756 128694 202768
rect 149698 202756 149704 202768
rect 128688 202728 149704 202756
rect 128688 202716 128694 202728
rect 149698 202716 149704 202728
rect 149756 202716 149762 202768
rect 166626 202716 166632 202768
rect 166684 202756 166690 202768
rect 183554 202756 183560 202768
rect 166684 202728 183560 202756
rect 166684 202716 166690 202728
rect 183554 202716 183560 202728
rect 183612 202716 183618 202768
rect 194962 202716 194968 202768
rect 195020 202756 195026 202768
rect 211154 202756 211160 202768
rect 195020 202728 211160 202756
rect 195020 202716 195026 202728
rect 211154 202716 211160 202728
rect 211212 202716 211218 202768
rect 222930 202716 222936 202768
rect 222988 202756 222994 202768
rect 233970 202756 233976 202768
rect 222988 202728 233976 202756
rect 222988 202716 222994 202728
rect 233970 202716 233976 202728
rect 234028 202716 234034 202768
rect 240318 202716 240324 202768
rect 240376 202756 240382 202768
rect 261478 202756 261484 202768
rect 240376 202728 261484 202756
rect 240376 202716 240382 202728
rect 261478 202716 261484 202728
rect 261536 202716 261542 202768
rect 278498 202716 278504 202768
rect 278556 202756 278562 202768
rect 295334 202756 295340 202768
rect 278556 202728 295340 202756
rect 278556 202716 278562 202728
rect 295334 202716 295340 202728
rect 295392 202716 295398 202768
rect 306926 202716 306932 202768
rect 306984 202756 306990 202768
rect 318058 202756 318064 202768
rect 306984 202728 318064 202756
rect 306984 202716 306990 202728
rect 318058 202716 318064 202728
rect 318116 202716 318122 202768
rect 324314 202716 324320 202768
rect 324372 202756 324378 202768
rect 345658 202756 345664 202768
rect 324372 202728 345664 202756
rect 324372 202716 324378 202728
rect 345658 202716 345664 202728
rect 345716 202716 345722 202768
rect 352650 202716 352656 202768
rect 352708 202756 352714 202768
rect 378870 202756 378876 202768
rect 352708 202728 378876 202756
rect 352708 202716 352714 202728
rect 378870 202716 378876 202728
rect 378928 202716 378934 202768
rect 390922 202716 390928 202768
rect 390980 202756 390986 202768
rect 402238 202756 402244 202768
rect 390980 202728 402244 202756
rect 390980 202716 390986 202728
rect 402238 202716 402244 202728
rect 402296 202716 402302 202768
rect 418614 202716 418620 202768
rect 418672 202756 418678 202768
rect 429838 202756 429844 202768
rect 418672 202728 429844 202756
rect 418672 202716 418678 202728
rect 429838 202716 429844 202728
rect 429896 202716 429902 202768
rect 436646 202716 436652 202768
rect 436704 202756 436710 202768
rect 458818 202756 458824 202768
rect 436704 202728 458824 202756
rect 436704 202716 436710 202728
rect 458818 202716 458824 202728
rect 458876 202716 458882 202768
rect 474458 202716 474464 202768
rect 474516 202756 474522 202768
rect 486418 202756 486424 202768
rect 474516 202728 486424 202756
rect 474516 202716 474522 202728
rect 486418 202716 486424 202728
rect 486476 202716 486482 202768
rect 502610 202716 502616 202768
rect 502668 202756 502674 202768
rect 514018 202756 514024 202768
rect 502668 202728 514024 202756
rect 502668 202716 502674 202728
rect 514018 202716 514024 202728
rect 514076 202716 514082 202768
rect 520642 202716 520648 202768
rect 520700 202756 520706 202768
rect 541618 202756 541624 202768
rect 520700 202728 541624 202756
rect 520700 202716 520706 202728
rect 541618 202716 541624 202728
rect 541676 202716 541682 202768
rect 54846 202648 54852 202700
rect 54904 202688 54910 202700
rect 71774 202688 71780 202700
rect 54904 202660 71780 202688
rect 54904 202648 54910 202660
rect 71774 202648 71780 202660
rect 71832 202648 71838 202700
rect 138934 202648 138940 202700
rect 138992 202688 138998 202700
rect 149882 202688 149888 202700
rect 138992 202660 149888 202688
rect 138992 202648 138998 202660
rect 149882 202648 149888 202660
rect 149940 202648 149946 202700
rect 250622 202648 250628 202700
rect 250680 202688 250686 202700
rect 267734 202688 267740 202700
rect 250680 202660 267740 202688
rect 250680 202648 250686 202660
rect 267734 202648 267740 202660
rect 267792 202648 267798 202700
rect 334618 202648 334624 202700
rect 334676 202688 334682 202700
rect 348418 202688 348424 202700
rect 334676 202660 348424 202688
rect 334676 202648 334682 202660
rect 348418 202648 348424 202660
rect 348476 202648 348482 202700
rect 362862 202648 362868 202700
rect 362920 202688 362926 202700
rect 379514 202688 379520 202700
rect 362920 202660 379520 202688
rect 362920 202648 362926 202660
rect 379514 202648 379520 202660
rect 379572 202648 379578 202700
rect 446950 202648 446956 202700
rect 447008 202688 447014 202700
rect 460198 202688 460204 202700
rect 447008 202660 460204 202688
rect 447008 202648 447014 202660
rect 460198 202648 460204 202660
rect 460256 202648 460262 202700
rect 530946 202648 530952 202700
rect 531004 202688 531010 202700
rect 547966 202688 547972 202700
rect 531004 202660 547972 202688
rect 531004 202648 531010 202660
rect 547966 202648 547972 202660
rect 548024 202648 548030 202700
rect 558638 202104 558644 202156
rect 558696 202144 558702 202156
rect 568758 202144 568764 202156
rect 558696 202116 568764 202144
rect 558696 202104 558702 202116
rect 568758 202104 568764 202116
rect 568816 202104 568822 202156
rect 548334 200744 548340 200796
rect 548392 200784 548398 200796
rect 569034 200784 569040 200796
rect 548392 200756 569040 200784
rect 548392 200744 548398 200756
rect 569034 200744 569040 200756
rect 569092 200744 569098 200796
rect 156322 200336 156328 200388
rect 156380 200376 156386 200388
rect 177298 200376 177304 200388
rect 156380 200348 177304 200376
rect 156380 200336 156386 200348
rect 177298 200336 177304 200348
rect 177356 200336 177362 200388
rect 92750 200268 92756 200320
rect 92808 200308 92814 200320
rect 110322 200308 110328 200320
rect 92808 200280 110328 200308
rect 92808 200268 92814 200280
rect 110322 200268 110328 200280
rect 110380 200268 110386 200320
rect 120718 200268 120724 200320
rect 120776 200308 120782 200320
rect 138290 200308 138296 200320
rect 120776 200280 138296 200308
rect 120776 200268 120782 200280
rect 138290 200268 138296 200280
rect 138348 200268 138354 200320
rect 149698 200268 149704 200320
rect 149756 200308 149762 200320
rect 165982 200308 165988 200320
rect 149756 200280 165988 200308
rect 149756 200268 149762 200280
rect 165982 200268 165988 200280
rect 166040 200268 166046 200320
rect 184014 200268 184020 200320
rect 184072 200308 184078 200320
rect 204898 200308 204904 200320
rect 184072 200280 204904 200308
rect 184072 200268 184078 200280
rect 204898 200268 204904 200280
rect 204956 200268 204962 200320
rect 464338 200268 464344 200320
rect 464396 200308 464402 200320
rect 485038 200308 485044 200320
rect 464396 200280 485044 200308
rect 464396 200268 464402 200280
rect 485038 200268 485044 200280
rect 485096 200268 485102 200320
rect 36998 200200 37004 200252
rect 37056 200240 37062 200252
rect 54294 200240 54300 200252
rect 37056 200212 54300 200240
rect 37056 200200 37062 200212
rect 54294 200200 54300 200212
rect 54352 200200 54358 200252
rect 65886 200200 65892 200252
rect 65944 200240 65950 200252
rect 81986 200240 81992 200252
rect 65944 200212 81992 200240
rect 65944 200200 65950 200212
rect 81986 200200 81992 200212
rect 82044 200200 82050 200252
rect 100018 200200 100024 200252
rect 100076 200240 100082 200252
rect 120902 200240 120908 200252
rect 100076 200212 120908 200240
rect 100076 200200 100082 200212
rect 120902 200200 120908 200212
rect 120960 200200 120966 200252
rect 176746 200200 176752 200252
rect 176804 200240 176810 200252
rect 194318 200240 194324 200252
rect 176804 200212 194324 200240
rect 176804 200200 176810 200212
rect 194318 200200 194324 200212
rect 194376 200200 194382 200252
rect 261478 200200 261484 200252
rect 261536 200240 261542 200252
rect 278314 200240 278320 200252
rect 261536 200212 278320 200240
rect 261536 200200 261542 200212
rect 278314 200200 278320 200212
rect 278372 200200 278378 200252
rect 288894 200200 288900 200252
rect 288952 200240 288958 200252
rect 306006 200240 306012 200252
rect 288952 200212 306012 200240
rect 288952 200200 288958 200212
rect 306006 200200 306012 200212
rect 306064 200200 306070 200252
rect 316770 200200 316776 200252
rect 316828 200240 316834 200252
rect 334342 200240 334348 200252
rect 316828 200212 334348 200240
rect 316828 200200 316834 200212
rect 334342 200200 334348 200212
rect 334400 200200 334406 200252
rect 372890 200200 372896 200252
rect 372948 200240 372954 200252
rect 390002 200240 390008 200252
rect 372948 200212 390008 200240
rect 372948 200200 372954 200212
rect 390002 200200 390008 200212
rect 390060 200200 390066 200252
rect 400766 200200 400772 200252
rect 400824 200240 400830 200252
rect 418338 200240 418344 200252
rect 400824 200212 418344 200240
rect 400824 200200 400830 200212
rect 418338 200200 418344 200212
rect 418396 200200 418402 200252
rect 457438 200200 457444 200252
rect 457496 200240 457502 200252
rect 473998 200240 474004 200252
rect 457496 200212 474004 200240
rect 457496 200200 457502 200212
rect 473998 200200 474004 200212
rect 474056 200200 474062 200252
rect 15194 200132 15200 200184
rect 15252 200172 15258 200184
rect 26326 200172 26332 200184
rect 15252 200144 26332 200172
rect 15252 200132 15258 200144
rect 26326 200132 26332 200144
rect 26384 200132 26390 200184
rect 38102 200132 38108 200184
rect 38160 200172 38166 200184
rect 64598 200172 64604 200184
rect 38160 200144 64604 200172
rect 38160 200132 38166 200144
rect 64598 200132 64604 200144
rect 64656 200132 64662 200184
rect 72326 200132 72332 200184
rect 72384 200172 72390 200184
rect 93118 200172 93124 200184
rect 72384 200144 93124 200172
rect 72384 200132 72390 200144
rect 93118 200132 93124 200144
rect 93176 200132 93182 200184
rect 94498 200132 94504 200184
rect 94556 200172 94562 200184
rect 120626 200172 120632 200184
rect 94556 200144 120632 200172
rect 94556 200132 94562 200144
rect 120626 200132 120632 200144
rect 120684 200132 120690 200184
rect 120810 200132 120816 200184
rect 120868 200172 120874 200184
rect 148594 200172 148600 200184
rect 120868 200144 148600 200172
rect 120868 200132 120874 200144
rect 148594 200132 148600 200144
rect 148652 200132 148658 200184
rect 149790 200132 149796 200184
rect 149848 200172 149854 200184
rect 176654 200172 176660 200184
rect 149848 200144 176660 200172
rect 149848 200132 149854 200144
rect 176654 200132 176660 200144
rect 176712 200132 176718 200184
rect 204806 200132 204812 200184
rect 204864 200172 204870 200184
rect 222286 200172 222292 200184
rect 204864 200144 222292 200172
rect 204864 200132 204870 200144
rect 222286 200132 222292 200144
rect 222344 200132 222350 200184
rect 232774 200132 232780 200184
rect 232832 200172 232838 200184
rect 250346 200172 250352 200184
rect 232832 200144 250352 200172
rect 232832 200132 232838 200144
rect 250346 200132 250352 200144
rect 250404 200132 250410 200184
rect 268010 200132 268016 200184
rect 268068 200172 268074 200184
rect 289078 200172 289084 200184
rect 268068 200144 289084 200172
rect 268068 200132 268074 200144
rect 289078 200132 289084 200144
rect 289136 200132 289142 200184
rect 290458 200132 290464 200184
rect 290516 200172 290522 200184
rect 316310 200172 316316 200184
rect 290516 200144 316316 200172
rect 290516 200132 290522 200144
rect 316310 200132 316316 200144
rect 316368 200132 316374 200184
rect 318058 200132 318064 200184
rect 318116 200172 318122 200184
rect 344646 200172 344652 200184
rect 318116 200144 344652 200172
rect 318116 200132 318122 200144
rect 344646 200132 344652 200144
rect 344704 200132 344710 200184
rect 352006 200132 352012 200184
rect 352064 200172 352070 200184
rect 373258 200172 373264 200184
rect 352064 200144 373264 200172
rect 352064 200132 352070 200144
rect 373258 200132 373264 200144
rect 373316 200132 373322 200184
rect 380342 200132 380348 200184
rect 380400 200172 380406 200184
rect 400858 200172 400864 200184
rect 380400 200144 400864 200172
rect 380400 200132 380406 200144
rect 400858 200132 400864 200144
rect 400916 200132 400922 200184
rect 429838 200132 429844 200184
rect 429896 200172 429902 200184
rect 456610 200172 456616 200184
rect 429896 200144 456616 200172
rect 429896 200132 429902 200144
rect 456610 200132 456616 200144
rect 456668 200132 456674 200184
rect 484854 200132 484860 200184
rect 484912 200172 484918 200184
rect 502334 200172 502340 200184
rect 484912 200144 502340 200172
rect 484912 200132 484918 200144
rect 502334 200132 502340 200144
rect 502392 200132 502398 200184
rect 512730 200132 512736 200184
rect 512788 200172 512794 200184
rect 530302 200172 530308 200184
rect 512788 200144 530308 200172
rect 512788 200132 512794 200144
rect 530302 200132 530308 200144
rect 530360 200132 530366 200184
rect 547138 200132 547144 200184
rect 547196 200172 547202 200184
rect 557994 200172 558000 200184
rect 547196 200144 558000 200172
rect 547196 200132 547202 200144
rect 557994 200132 558000 200144
rect 558052 200132 558058 200184
rect 92750 198296 92756 198348
rect 92808 198296 92814 198348
rect 232774 198296 232780 198348
rect 232832 198296 232838 198348
rect 400766 198296 400772 198348
rect 400824 198296 400830 198348
rect 400858 198296 400864 198348
rect 400916 198296 400922 198348
rect 512730 198296 512736 198348
rect 512788 198296 512794 198348
rect 568758 198296 568764 198348
rect 568816 198296 568822 198348
rect 92768 198144 92796 198296
rect 204714 198228 204720 198280
rect 204772 198268 204778 198280
rect 204990 198268 204996 198280
rect 204772 198240 204996 198268
rect 204772 198228 204778 198240
rect 204990 198228 204996 198240
rect 205048 198228 205054 198280
rect 232792 198144 232820 198296
rect 400784 198144 400812 198296
rect 400876 198144 400904 198296
rect 512748 198144 512776 198296
rect 568776 198144 568804 198296
rect 92750 198092 92756 198144
rect 92808 198092 92814 198144
rect 232774 198092 232780 198144
rect 232832 198092 232838 198144
rect 400766 198092 400772 198144
rect 400824 198092 400830 198144
rect 400858 198092 400864 198144
rect 400916 198092 400922 198144
rect 512730 198092 512736 198144
rect 512788 198092 512794 198144
rect 568758 198092 568764 198144
rect 568816 198092 568822 198144
rect 36814 195168 36820 195220
rect 36872 195208 36878 195220
rect 36998 195208 37004 195220
rect 36872 195180 37004 195208
rect 36872 195168 36878 195180
rect 36998 195168 37004 195180
rect 37056 195168 37062 195220
rect 569310 191836 569316 191888
rect 569368 191876 569374 191888
rect 580074 191876 580080 191888
rect 569368 191848 580080 191876
rect 569368 191836 569374 191848
rect 580074 191836 580080 191848
rect 580132 191836 580138 191888
rect 2774 187688 2780 187740
rect 2832 187728 2838 187740
rect 5166 187728 5172 187740
rect 2832 187700 5172 187728
rect 2832 187688 2838 187700
rect 5166 187688 5172 187700
rect 5224 187688 5230 187740
rect 64874 185580 64880 185632
rect 64932 185620 64938 185632
rect 65886 185620 65892 185632
rect 64932 185592 65892 185620
rect 64932 185580 64938 185592
rect 65886 185580 65892 185592
rect 65944 185580 65950 185632
rect 289078 182112 289084 182164
rect 289136 182152 289142 182164
rect 295702 182152 295708 182164
rect 289136 182124 295708 182152
rect 289136 182112 289142 182124
rect 295702 182112 295708 182124
rect 295760 182112 295766 182164
rect 93118 181432 93124 181484
rect 93176 181472 93182 181484
rect 99742 181472 99748 181484
rect 93176 181444 99748 181472
rect 93176 181432 93182 181444
rect 99742 181432 99748 181444
rect 99800 181432 99806 181484
rect 120902 181432 120908 181484
rect 120960 181472 120966 181484
rect 127710 181472 127716 181484
rect 120960 181444 127716 181472
rect 120960 181432 120966 181444
rect 127710 181432 127716 181444
rect 127768 181432 127774 181484
rect 177298 181432 177304 181484
rect 177356 181472 177362 181484
rect 183738 181472 183744 181484
rect 177356 181444 183744 181472
rect 177356 181432 177362 181444
rect 183738 181432 183744 181444
rect 183796 181432 183802 181484
rect 373258 181432 373264 181484
rect 373316 181472 373322 181484
rect 379698 181472 379704 181484
rect 373316 181444 379704 181472
rect 373316 181432 373322 181444
rect 379698 181432 379704 181444
rect 379756 181432 379762 181484
rect 400858 181432 400864 181484
rect 400916 181472 400922 181484
rect 407758 181472 407764 181484
rect 400916 181444 407764 181472
rect 400916 181432 400922 181444
rect 407758 181432 407764 181444
rect 407816 181432 407822 181484
rect 204898 180820 204904 180872
rect 204956 180860 204962 180872
rect 211706 180860 211712 180872
rect 204956 180832 211712 180860
rect 204956 180820 204962 180832
rect 211706 180820 211712 180832
rect 211764 180820 211770 180872
rect 485038 180820 485044 180872
rect 485096 180860 485102 180872
rect 491662 180860 491668 180872
rect 485096 180832 491668 180860
rect 485096 180820 485102 180832
rect 491662 180820 491668 180832
rect 491720 180820 491726 180872
rect 42702 179324 42708 179376
rect 42760 179364 42766 179376
rect 95234 179364 95240 179376
rect 42760 179336 95240 179364
rect 42760 179324 42766 179336
rect 95234 179324 95240 179336
rect 95292 179324 95298 179376
rect 97902 179324 97908 179376
rect 97960 179364 97966 179376
rect 150434 179364 150440 179376
rect 97960 179336 150440 179364
rect 97960 179324 97966 179336
rect 150434 179324 150440 179336
rect 150492 179324 150498 179376
rect 154482 179324 154488 179376
rect 154540 179364 154546 179376
rect 207014 179364 207020 179376
rect 154540 179336 207020 179364
rect 154540 179324 154546 179336
rect 207014 179324 207020 179336
rect 207072 179324 207078 179376
rect 209682 179324 209688 179376
rect 209740 179364 209746 179376
rect 262214 179364 262220 179376
rect 209740 179336 262220 179364
rect 209740 179324 209746 179336
rect 262214 179324 262220 179336
rect 262272 179324 262278 179376
rect 266262 179324 266268 179376
rect 266320 179364 266326 179376
rect 318794 179364 318800 179376
rect 266320 179336 318800 179364
rect 266320 179324 266326 179336
rect 318794 179324 318800 179336
rect 318852 179324 318858 179376
rect 322842 179324 322848 179376
rect 322900 179364 322906 179376
rect 375374 179364 375380 179376
rect 322900 179336 375380 179364
rect 322900 179324 322906 179336
rect 375374 179324 375380 179336
rect 375432 179324 375438 179376
rect 378042 179324 378048 179376
rect 378100 179364 378106 179376
rect 430574 179364 430580 179376
rect 378100 179336 430580 179364
rect 378100 179324 378106 179336
rect 430574 179324 430580 179336
rect 430632 179324 430638 179376
rect 434622 179324 434628 179376
rect 434680 179364 434686 179376
rect 487154 179364 487160 179376
rect 434680 179336 487160 179364
rect 434680 179324 434686 179336
rect 487154 179324 487160 179336
rect 487212 179324 487218 179376
rect 489822 179324 489828 179376
rect 489880 179364 489886 179376
rect 542354 179364 542360 179376
rect 489880 179336 542360 179364
rect 489880 179324 489886 179336
rect 542354 179324 542360 179336
rect 542412 179324 542418 179376
rect 288802 178848 288808 178900
rect 288860 178888 288866 178900
rect 288986 178888 288992 178900
rect 288860 178860 288992 178888
rect 288860 178848 288866 178860
rect 288986 178848 288992 178860
rect 289044 178848 289050 178900
rect 372798 178848 372804 178900
rect 372856 178888 372862 178900
rect 372982 178888 372988 178900
rect 372856 178860 372988 178888
rect 372856 178848 372862 178860
rect 372982 178848 372988 178860
rect 373040 178848 373046 178900
rect 484762 178848 484768 178900
rect 484820 178888 484826 178900
rect 484946 178888 484952 178900
rect 484820 178860 484952 178888
rect 484820 178848 484826 178860
rect 484946 178848 484952 178860
rect 485004 178848 485010 178900
rect 547874 178644 547880 178696
rect 547932 178684 547938 178696
rect 548150 178684 548156 178696
rect 547932 178656 548156 178684
rect 547932 178644 547938 178656
rect 548150 178644 548156 178656
rect 548208 178644 548214 178696
rect 15378 176604 15384 176656
rect 15436 176644 15442 176656
rect 43990 176644 43996 176656
rect 15436 176616 43996 176644
rect 15436 176604 15442 176616
rect 43990 176604 43996 176616
rect 44048 176604 44054 176656
rect 110322 176604 110328 176656
rect 110380 176644 110386 176656
rect 120810 176644 120816 176656
rect 110380 176616 120816 176644
rect 110380 176604 110386 176616
rect 120810 176604 120816 176616
rect 120868 176604 120874 176656
rect 166626 176604 166632 176656
rect 166684 176644 166690 176656
rect 204990 176644 204996 176656
rect 166684 176616 204996 176644
rect 166684 176604 166690 176616
rect 204990 176604 204996 176616
rect 205048 176604 205054 176656
rect 211246 176604 211252 176656
rect 211304 176644 211310 176656
rect 240042 176644 240048 176656
rect 211304 176616 240048 176644
rect 211304 176604 211310 176616
rect 240042 176604 240048 176616
rect 240100 176604 240106 176656
rect 295426 176604 295432 176656
rect 295484 176644 295490 176656
rect 324038 176644 324044 176656
rect 295484 176616 324044 176644
rect 295484 176604 295490 176616
rect 324038 176604 324044 176616
rect 324096 176604 324102 176656
rect 334342 176604 334348 176656
rect 334400 176644 334406 176656
rect 372982 176644 372988 176656
rect 334400 176616 372988 176644
rect 334400 176604 334406 176616
rect 372982 176604 372988 176616
rect 373040 176604 373046 176656
rect 390462 176604 390468 176656
rect 390520 176644 390526 176656
rect 428734 176644 428740 176656
rect 390520 176616 428740 176644
rect 390520 176604 390526 176616
rect 428734 176604 428740 176616
rect 428792 176604 428798 176656
rect 434806 176604 434812 176656
rect 434864 176644 434870 176656
rect 434864 176616 441614 176644
rect 434864 176604 434870 176616
rect 26326 176536 26332 176588
rect 26384 176576 26390 176588
rect 38102 176576 38108 176588
rect 26384 176548 38108 176576
rect 26384 176536 26390 176548
rect 38102 176536 38108 176548
rect 38160 176536 38166 176588
rect 42886 176536 42892 176588
rect 42944 176576 42950 176588
rect 71774 176576 71780 176588
rect 42944 176548 71780 176576
rect 42944 176536 42950 176548
rect 71774 176536 71780 176548
rect 71832 176536 71838 176588
rect 82630 176536 82636 176588
rect 82688 176576 82694 176588
rect 94498 176576 94504 176588
rect 82688 176548 94504 176576
rect 82688 176536 82694 176548
rect 94498 176536 94504 176548
rect 94556 176536 94562 176588
rect 138290 176536 138296 176588
rect 138348 176576 138354 176588
rect 149790 176576 149796 176588
rect 138348 176548 149796 176576
rect 138348 176536 138354 176548
rect 149790 176536 149796 176548
rect 149848 176536 149854 176588
rect 194318 176536 194324 176588
rect 194376 176576 194382 176588
rect 232866 176576 232872 176588
rect 194376 176548 232872 176576
rect 194376 176536 194382 176548
rect 232866 176536 232872 176548
rect 232924 176536 232930 176588
rect 238846 176536 238852 176588
rect 238904 176576 238910 176588
rect 268010 176576 268016 176588
rect 238904 176548 268016 176576
rect 238904 176536 238910 176548
rect 268010 176536 268016 176548
rect 268068 176536 268074 176588
rect 278314 176536 278320 176588
rect 278372 176576 278378 176588
rect 290458 176576 290464 176588
rect 278372 176548 290464 176576
rect 278372 176536 278378 176548
rect 290458 176536 290464 176548
rect 290516 176536 290522 176588
rect 306282 176536 306288 176588
rect 306340 176576 306346 176588
rect 318058 176576 318064 176588
rect 306340 176548 318064 176576
rect 306340 176536 306346 176548
rect 318058 176536 318064 176548
rect 318116 176536 318122 176588
rect 323026 176536 323032 176588
rect 323084 176576 323090 176588
rect 352006 176576 352012 176588
rect 323084 176548 352012 176576
rect 323084 176536 323090 176548
rect 352006 176536 352012 176548
rect 352064 176536 352070 176588
rect 362310 176536 362316 176588
rect 362368 176576 362374 176588
rect 400950 176576 400956 176588
rect 362368 176548 400956 176576
rect 362368 176536 362374 176548
rect 400950 176536 400956 176548
rect 401008 176536 401014 176588
rect 407206 176536 407212 176588
rect 407264 176576 407270 176588
rect 436002 176576 436008 176588
rect 407264 176548 436008 176576
rect 407264 176536 407270 176548
rect 436002 176536 436008 176548
rect 436060 176536 436066 176588
rect 441586 176576 441614 176616
rect 491386 176604 491392 176656
rect 491444 176644 491450 176656
rect 519998 176644 520004 176656
rect 491444 176616 520004 176644
rect 491444 176604 491450 176616
rect 519998 176604 520004 176616
rect 520056 176604 520062 176656
rect 530302 176604 530308 176656
rect 530360 176644 530366 176656
rect 568850 176644 568856 176656
rect 530360 176616 568856 176644
rect 530360 176604 530366 176616
rect 568850 176604 568856 176616
rect 568908 176604 568914 176656
rect 463694 176576 463700 176588
rect 441586 176548 463700 176576
rect 463694 176536 463700 176548
rect 463752 176536 463758 176588
rect 474642 176536 474648 176588
rect 474700 176576 474706 176588
rect 512822 176576 512828 176588
rect 474700 176548 512828 176576
rect 474700 176536 474706 176548
rect 512822 176536 512828 176548
rect 512880 176536 512886 176588
rect 518986 176536 518992 176588
rect 519044 176576 519050 176588
rect 547874 176576 547880 176588
rect 519044 176548 547880 176576
rect 519044 176536 519050 176548
rect 547874 176536 547880 176548
rect 547932 176536 547938 176588
rect 54294 176468 54300 176520
rect 54352 176508 54358 176520
rect 92842 176508 92848 176520
rect 54352 176480 92848 176508
rect 54352 176468 54358 176480
rect 92842 176468 92848 176480
rect 92900 176468 92906 176520
rect 127066 176468 127072 176520
rect 127124 176508 127130 176520
rect 156046 176508 156052 176520
rect 127124 176480 156052 176508
rect 127124 176468 127130 176480
rect 156046 176468 156052 176480
rect 156104 176468 156110 176520
rect 250346 176468 250352 176520
rect 250404 176508 250410 176520
rect 288986 176508 288992 176520
rect 250404 176480 288992 176508
rect 250404 176468 250410 176480
rect 288986 176468 288992 176480
rect 289044 176468 289050 176520
rect 418338 176468 418344 176520
rect 418396 176508 418402 176520
rect 429838 176508 429844 176520
rect 418396 176480 429844 176508
rect 418396 176468 418402 176480
rect 429838 176468 429844 176480
rect 429896 176468 429902 176520
rect 446306 176468 446312 176520
rect 446364 176508 446370 176520
rect 484946 176508 484952 176520
rect 446364 176480 484952 176508
rect 446364 176468 446370 176480
rect 484946 176468 484952 176480
rect 485004 176468 485010 176520
rect 502334 176468 502340 176520
rect 502392 176508 502398 176520
rect 502392 176480 528554 176508
rect 502392 176468 502398 176480
rect 528526 176440 528554 176480
rect 540606 176468 540612 176520
rect 540664 176508 540670 176520
rect 547138 176508 547144 176520
rect 540664 176480 547144 176508
rect 540664 176468 540670 176480
rect 547138 176468 547144 176480
rect 547196 176468 547202 176520
rect 548150 176468 548156 176520
rect 548208 176508 548214 176520
rect 557994 176508 558000 176520
rect 548208 176480 558000 176508
rect 548208 176468 548214 176480
rect 557994 176468 558000 176480
rect 558052 176468 558058 176520
rect 540790 176440 540796 176452
rect 528526 176412 540796 176440
rect 540790 176400 540796 176412
rect 540848 176400 540854 176452
rect 15194 175992 15200 176044
rect 15252 176032 15258 176044
rect 16022 176032 16028 176044
rect 15252 176004 16028 176032
rect 15252 175992 15258 176004
rect 16022 175992 16028 176004
rect 16080 175992 16086 176044
rect 26602 174496 26608 174548
rect 26660 174536 26666 174548
rect 36814 174536 36820 174548
rect 26660 174508 36820 174536
rect 26660 174496 26666 174508
rect 36814 174496 36820 174508
rect 36872 174496 36878 174548
rect 15378 174020 15384 174072
rect 15436 174060 15442 174072
rect 54294 174060 54300 174072
rect 15436 174032 54300 174060
rect 15436 174020 15442 174032
rect 54294 174020 54300 174032
rect 54352 174020 54358 174072
rect 66898 174020 66904 174072
rect 66956 174060 66962 174072
rect 82630 174060 82636 174072
rect 66956 174032 82636 174060
rect 66956 174020 66962 174032
rect 82630 174020 82636 174032
rect 82688 174020 82694 174072
rect 149698 174020 149704 174072
rect 149756 174060 149762 174072
rect 166626 174060 166632 174072
rect 149756 174032 166632 174060
rect 149756 174020 149762 174032
rect 166626 174020 166632 174032
rect 166684 174020 166690 174072
rect 200086 174032 209774 174060
rect 71866 173952 71872 174004
rect 71924 173992 71930 174004
rect 110598 173992 110604 174004
rect 71924 173964 110604 173992
rect 71924 173952 71930 173964
rect 110598 173952 110604 173964
rect 110656 173952 110662 174004
rect 122098 173952 122104 174004
rect 122156 173992 122162 174004
rect 128354 173992 128360 174004
rect 122156 173964 128360 173992
rect 122156 173952 122162 173964
rect 128354 173952 128360 173964
rect 128412 173952 128418 174004
rect 177298 173952 177304 174004
rect 177356 173992 177362 174004
rect 194594 173992 194600 174004
rect 177356 173964 194600 173992
rect 177356 173952 177362 173964
rect 194594 173952 194600 173964
rect 194652 173952 194658 174004
rect 36906 173884 36912 173936
rect 36964 173924 36970 173936
rect 43438 173924 43444 173936
rect 36964 173896 43444 173924
rect 36964 173884 36970 173896
rect 43438 173884 43444 173896
rect 43496 173884 43502 173936
rect 99374 173884 99380 173936
rect 99432 173924 99438 173936
rect 138290 173924 138296 173936
rect 99432 173896 138296 173924
rect 99432 173884 99438 173896
rect 138290 173884 138296 173896
rect 138348 173884 138354 173936
rect 178678 173884 178684 173936
rect 178736 173924 178742 173936
rect 184290 173924 184296 173936
rect 178736 173896 184296 173924
rect 178736 173884 178742 173896
rect 184290 173884 184296 173896
rect 184348 173884 184354 173936
rect 200086 173924 200114 174032
rect 209746 173936 209774 174032
rect 211246 174020 211252 174072
rect 211304 174060 211310 174072
rect 211304 174032 219434 174060
rect 211304 174020 211310 174032
rect 211982 173992 211988 174004
rect 209884 173964 211988 173992
rect 184400 173896 200114 173924
rect 183646 173816 183652 173868
rect 183704 173856 183710 173868
rect 184400 173856 184428 173896
rect 206278 173884 206284 173936
rect 206336 173924 206342 173936
rect 206336 173896 209544 173924
rect 209746 173896 209780 173936
rect 206336 173884 206342 173896
rect 183704 173828 184428 173856
rect 209516 173856 209544 173896
rect 209774 173884 209780 173896
rect 209832 173884 209838 173936
rect 209884 173856 209912 173964
rect 211982 173952 211988 173964
rect 212040 173952 212046 174004
rect 219406 173992 219434 174032
rect 374638 174020 374644 174072
rect 374696 174060 374702 174072
rect 380342 174060 380348 174072
rect 374696 174032 380348 174060
rect 374696 174020 374702 174032
rect 380342 174020 380348 174032
rect 380400 174020 380406 174072
rect 407206 174020 407212 174072
rect 407264 174060 407270 174072
rect 407264 174032 412634 174060
rect 407264 174020 407270 174032
rect 250622 173992 250628 174004
rect 219406 173964 250628 173992
rect 250622 173952 250628 173964
rect 250680 173952 250686 174004
rect 262858 173952 262864 174004
rect 262916 173992 262922 174004
rect 262916 173964 267734 173992
rect 262916 173952 262922 173964
rect 209958 173884 209964 173936
rect 210016 173924 210022 173936
rect 222286 173924 222292 173936
rect 210016 173896 222292 173924
rect 210016 173884 210022 173896
rect 222286 173884 222292 173896
rect 222344 173884 222350 173936
rect 234062 173884 234068 173936
rect 234120 173924 234126 173936
rect 240318 173924 240324 173936
rect 234120 173896 240324 173924
rect 234120 173884 234126 173896
rect 240318 173884 240324 173896
rect 240376 173884 240382 173936
rect 264238 173884 264244 173936
rect 264296 173924 264302 173936
rect 267706 173924 267734 173964
rect 267826 173952 267832 174004
rect 267884 173992 267890 174004
rect 306466 173992 306472 174004
rect 267884 173964 306472 173992
rect 267884 173952 267890 173964
rect 306466 173952 306472 173964
rect 306524 173952 306530 174004
rect 318058 173952 318064 174004
rect 318116 173992 318122 174004
rect 324314 173992 324320 174004
rect 318116 173964 324320 173992
rect 318116 173952 318122 173964
rect 324314 173952 324320 173964
rect 324372 173952 324378 174004
rect 345842 173952 345848 174004
rect 345900 173992 345906 174004
rect 362310 173992 362316 174004
rect 345900 173964 362316 173992
rect 345900 173952 345906 173964
rect 362310 173952 362316 173964
rect 362368 173952 362374 174004
rect 373258 173952 373264 174004
rect 373316 173992 373322 174004
rect 390646 173992 390652 174004
rect 373316 173964 390652 173992
rect 373316 173952 373322 173964
rect 390646 173952 390652 173964
rect 390704 173952 390710 174004
rect 402238 173952 402244 174004
rect 402296 173992 402302 174004
rect 408310 173992 408316 174004
rect 402296 173964 408316 173992
rect 402296 173952 402302 173964
rect 408310 173952 408316 173964
rect 408368 173952 408374 174004
rect 412606 173992 412634 174032
rect 491386 174020 491392 174072
rect 491444 174060 491450 174072
rect 492398 174060 492404 174072
rect 491444 174032 492404 174060
rect 491444 174020 491450 174032
rect 492398 174020 492404 174032
rect 492456 174020 492462 174072
rect 530302 174060 530308 174072
rect 509206 174032 530308 174060
rect 446306 173992 446312 174004
rect 412606 173964 446312 173992
rect 446306 173952 446312 173964
rect 446364 173952 446370 174004
rect 463786 173952 463792 174004
rect 463844 173992 463850 174004
rect 502610 173992 502616 174004
rect 463844 173964 502616 173992
rect 463844 173952 463850 173964
rect 502610 173952 502616 173964
rect 502668 173952 502674 174004
rect 278590 173924 278596 173936
rect 264296 173896 267596 173924
rect 267706 173896 278596 173924
rect 264296 173884 264302 173896
rect 209516 173828 209912 173856
rect 267568 173856 267596 173896
rect 278590 173884 278596 173896
rect 278648 173884 278654 173936
rect 295334 173884 295340 173936
rect 295392 173924 295398 173936
rect 334618 173924 334624 173936
rect 295392 173896 334624 173924
rect 295392 173884 295398 173896
rect 334618 173884 334624 173896
rect 334676 173884 334682 173936
rect 345750 173884 345756 173936
rect 345808 173924 345814 173936
rect 352006 173924 352012 173936
rect 345808 173896 352012 173924
rect 345808 173884 345814 173896
rect 352006 173884 352012 173896
rect 352064 173884 352070 173936
rect 379606 173884 379612 173936
rect 379664 173924 379670 173936
rect 418614 173924 418620 173936
rect 379664 173896 418620 173924
rect 379664 173884 379670 173896
rect 418614 173884 418620 173896
rect 418672 173884 418678 173936
rect 429930 173884 429936 173936
rect 429988 173924 429994 173936
rect 436094 173924 436100 173936
rect 429988 173896 436100 173924
rect 429988 173884 429994 173896
rect 436094 173884 436100 173896
rect 436152 173884 436158 173936
rect 457438 173884 457444 173936
rect 457496 173924 457502 173936
rect 474642 173924 474648 173936
rect 457496 173896 474648 173924
rect 457496 173884 457502 173896
rect 474642 173884 474648 173896
rect 474700 173884 474706 173936
rect 486418 173884 486424 173936
rect 486476 173924 486482 173936
rect 492306 173924 492312 173936
rect 486476 173896 492312 173924
rect 486476 173884 486482 173896
rect 492306 173884 492312 173896
rect 492364 173884 492370 173936
rect 492398 173884 492404 173936
rect 492456 173924 492462 173936
rect 509206 173924 509234 174032
rect 530302 174020 530308 174032
rect 530360 174020 530366 174072
rect 541618 174020 541624 174072
rect 541676 174060 541682 174072
rect 558638 174060 558644 174072
rect 541676 174032 558644 174060
rect 541676 174020 541682 174032
rect 558638 174020 558644 174032
rect 558696 174020 558702 174072
rect 492456 173896 509234 173924
rect 492456 173884 492462 173896
rect 514018 173884 514024 173936
rect 514076 173924 514082 173936
rect 520274 173924 520280 173936
rect 514076 173896 518894 173924
rect 514076 173884 514082 173896
rect 267918 173856 267924 173868
rect 267568 173828 267924 173856
rect 183704 173816 183710 173828
rect 267918 173816 267924 173828
rect 267976 173816 267982 173868
rect 518866 173856 518894 173896
rect 519096 173896 520280 173924
rect 519096 173856 519124 173896
rect 520274 173884 520280 173896
rect 520332 173884 520338 173936
rect 518866 173828 519124 173856
rect 148962 172048 148968 172100
rect 149020 172088 149026 172100
rect 153838 172088 153844 172100
rect 149020 172060 153844 172088
rect 149020 172048 149026 172060
rect 153838 172048 153844 172060
rect 153896 172048 153902 172100
rect 238662 171436 238668 171488
rect 238720 171476 238726 171488
rect 291194 171476 291200 171488
rect 238720 171448 291200 171476
rect 238720 171436 238726 171448
rect 291194 171436 291200 171448
rect 291252 171436 291258 171488
rect 462222 171436 462228 171488
rect 462280 171476 462286 171488
rect 514754 171476 514760 171488
rect 462280 171448 514760 171476
rect 462280 171436 462286 171448
rect 514754 171436 514760 171448
rect 514812 171436 514818 171488
rect 205082 171368 205088 171420
rect 205140 171368 205146 171420
rect 209682 171368 209688 171420
rect 209740 171408 209746 171420
rect 262214 171408 262220 171420
rect 209740 171380 262220 171408
rect 209740 171368 209746 171380
rect 262214 171368 262220 171380
rect 262272 171368 262278 171420
rect 434622 171368 434628 171420
rect 434680 171408 434686 171420
rect 487154 171408 487160 171420
rect 434680 171380 487160 171408
rect 434680 171368 434686 171380
rect 487154 171368 487160 171380
rect 487212 171368 487218 171420
rect 205100 171216 205128 171368
rect 541158 171232 541164 171284
rect 541216 171272 541222 171284
rect 544378 171272 544384 171284
rect 541216 171244 544384 171272
rect 541216 171232 541222 171244
rect 544378 171232 544384 171244
rect 544436 171232 544442 171284
rect 40678 171164 40684 171216
rect 40736 171204 40742 171216
rect 44174 171204 44180 171216
rect 40736 171176 44180 171204
rect 40736 171164 40742 171176
rect 44174 171164 44180 171176
rect 44232 171164 44238 171216
rect 71130 171164 71136 171216
rect 71188 171204 71194 171216
rect 71958 171204 71964 171216
rect 71188 171176 71964 171204
rect 71188 171164 71194 171176
rect 71958 171164 71964 171176
rect 72016 171164 72022 171216
rect 205082 171164 205088 171216
rect 205140 171164 205146 171216
rect 429102 171164 429108 171216
rect 429160 171204 429166 171216
rect 429838 171204 429844 171216
rect 429160 171176 429844 171204
rect 429160 171164 429166 171176
rect 429838 171164 429844 171176
rect 429896 171164 429902 171216
rect 13538 171096 13544 171148
rect 13596 171136 13602 171148
rect 66254 171136 66260 171148
rect 13596 171108 66260 171136
rect 13596 171096 13602 171108
rect 66254 171096 66260 171108
rect 66312 171096 66318 171148
rect 70302 171096 70308 171148
rect 70360 171136 70366 171148
rect 122834 171136 122840 171148
rect 70360 171108 122840 171136
rect 70360 171096 70366 171108
rect 122834 171096 122840 171108
rect 122892 171096 122898 171148
rect 233234 166268 233240 166320
rect 233292 166308 233298 166320
rect 233970 166308 233976 166320
rect 233292 166280 233976 166308
rect 233292 166268 233298 166280
rect 233970 166268 233976 166280
rect 234028 166268 234034 166320
rect 463694 166268 463700 166320
rect 463752 166308 463758 166320
rect 464062 166308 464068 166320
rect 463752 166280 464068 166308
rect 463752 166268 463758 166280
rect 464062 166268 464068 166280
rect 464120 166268 464126 166320
rect 93118 153824 93124 153876
rect 93176 153864 93182 153876
rect 99466 153864 99472 153876
rect 93176 153836 99472 153864
rect 93176 153824 93182 153836
rect 99466 153824 99472 153836
rect 99524 153824 99530 153876
rect 289170 153688 289176 153740
rect 289228 153728 289234 153740
rect 295426 153728 295432 153740
rect 289228 153700 295432 153728
rect 289228 153688 289234 153700
rect 295426 153688 295432 153700
rect 295484 153688 295490 153740
rect 569402 151784 569408 151836
rect 569460 151824 569466 151836
rect 580074 151824 580080 151836
rect 569460 151796 580080 151824
rect 569460 151784 569466 151796
rect 580074 151784 580080 151796
rect 580132 151784 580138 151836
rect 2774 149336 2780 149388
rect 2832 149376 2838 149388
rect 5258 149376 5264 149388
rect 2832 149348 5264 149376
rect 2832 149336 2838 149348
rect 5258 149336 5264 149348
rect 5316 149336 5322 149388
rect 15286 148996 15292 149048
rect 15344 149036 15350 149048
rect 36906 149036 36912 149048
rect 15344 149008 36912 149036
rect 15344 148996 15350 149008
rect 36906 148996 36912 149008
rect 36964 148996 36970 149048
rect 65058 148996 65064 149048
rect 65116 149036 65122 149048
rect 92934 149036 92940 149048
rect 65116 149008 92940 149036
rect 65116 148996 65122 149008
rect 92934 148996 92940 149008
rect 92992 148996 92998 149048
rect 93026 148996 93032 149048
rect 93084 149036 93090 149048
rect 120902 149036 120908 149048
rect 93084 149008 120908 149036
rect 93084 148996 93090 149008
rect 120902 148996 120908 149008
rect 120960 148996 120966 149048
rect 121086 148996 121092 149048
rect 121144 149036 121150 149048
rect 148594 149036 148600 149048
rect 121144 149008 148600 149036
rect 121144 148996 121150 149008
rect 148594 148996 148600 149008
rect 148652 148996 148658 149048
rect 153838 148996 153844 149048
rect 153896 149036 153902 149048
rect 176930 149036 176936 149048
rect 153896 149008 176936 149036
rect 153896 148996 153902 149008
rect 176930 148996 176936 149008
rect 176988 148996 176994 149048
rect 177022 148996 177028 149048
rect 177080 149036 177086 149048
rect 204898 149036 204904 149048
rect 177080 149008 204904 149036
rect 177080 148996 177086 149008
rect 204898 148996 204904 149008
rect 204956 148996 204962 149048
rect 205174 148996 205180 149048
rect 205232 149036 205238 149048
rect 232590 149036 232596 149048
rect 205232 149008 232596 149036
rect 205232 148996 205238 149008
rect 232590 148996 232596 149008
rect 232648 148996 232654 149048
rect 233970 148996 233976 149048
rect 234028 149036 234034 149048
rect 260926 149036 260932 149048
rect 234028 149008 260932 149036
rect 234028 148996 234034 149008
rect 260926 148996 260932 149008
rect 260984 148996 260990 149048
rect 261018 148996 261024 149048
rect 261076 149036 261082 149048
rect 288894 149036 288900 149048
rect 261076 149008 288900 149036
rect 261076 148996 261082 149008
rect 288894 148996 288900 149008
rect 288952 148996 288958 149048
rect 289078 148996 289084 149048
rect 289136 149036 289142 149048
rect 316586 149036 316592 149048
rect 289136 149008 316592 149036
rect 289136 148996 289142 149008
rect 316586 148996 316592 149008
rect 316644 148996 316650 149048
rect 317046 148996 317052 149048
rect 317104 149036 317110 149048
rect 344922 149036 344928 149048
rect 317104 149008 344928 149036
rect 317104 148996 317110 149008
rect 344922 148996 344928 149008
rect 344980 148996 344986 149048
rect 345658 148996 345664 149048
rect 345716 149036 345722 149048
rect 372614 149036 372620 149048
rect 345716 149008 372620 149036
rect 345716 148996 345722 149008
rect 372614 148996 372620 149008
rect 372672 148996 372678 149048
rect 373074 148996 373080 149048
rect 373132 149036 373138 149048
rect 400950 149036 400956 149048
rect 373132 149008 400956 149036
rect 373132 148996 373138 149008
rect 400950 148996 400956 149008
rect 401008 148996 401014 149048
rect 401042 148996 401048 149048
rect 401100 149036 401106 149048
rect 428918 149036 428924 149048
rect 401100 149008 428924 149036
rect 401100 148996 401106 149008
rect 428918 148996 428924 149008
rect 428976 148996 428982 149048
rect 429838 148996 429844 149048
rect 429896 149036 429902 149048
rect 456794 149036 456800 149048
rect 429896 149008 456800 149036
rect 429896 148996 429902 149008
rect 456794 148996 456800 149008
rect 456852 148996 456858 149048
rect 457070 148996 457076 149048
rect 457128 149036 457134 149048
rect 484946 149036 484952 149048
rect 457128 149008 484952 149036
rect 457128 148996 457134 149008
rect 484946 148996 484952 149008
rect 485004 148996 485010 149048
rect 485038 148996 485044 149048
rect 485096 149036 485102 149048
rect 512914 149036 512920 149048
rect 485096 149008 512920 149036
rect 485096 148996 485102 149008
rect 512914 148996 512920 149008
rect 512972 148996 512978 149048
rect 513098 148996 513104 149048
rect 513156 149036 513162 149048
rect 540606 149036 540612 149048
rect 513156 149008 540612 149036
rect 513156 148996 513162 149008
rect 540606 148996 540612 149008
rect 540664 148996 540670 149048
rect 544378 148996 544384 149048
rect 544436 149036 544442 149048
rect 568942 149036 568948 149048
rect 544436 149008 568948 149036
rect 544436 148996 544442 149008
rect 568942 148996 568948 149008
rect 569000 148996 569006 149048
rect 26602 148928 26608 148980
rect 26660 148968 26666 148980
rect 40678 148968 40684 148980
rect 26660 148940 40684 148968
rect 26660 148928 26666 148940
rect 40678 148928 40684 148940
rect 40736 148928 40742 148980
rect 43438 148928 43444 148980
rect 43496 148968 43502 148980
rect 64874 148968 64880 148980
rect 43496 148940 64880 148968
rect 43496 148928 43502 148940
rect 64874 148928 64880 148940
rect 64932 148928 64938 148980
rect 82630 148928 82636 148980
rect 82688 148968 82694 148980
rect 93118 148968 93124 148980
rect 82688 148940 93124 148968
rect 82688 148928 82694 148940
rect 93118 148928 93124 148940
rect 93176 148928 93182 148980
rect 110598 148928 110604 148980
rect 110656 148968 110662 148980
rect 122098 148968 122104 148980
rect 110656 148940 122104 148968
rect 110656 148928 110662 148940
rect 122098 148928 122104 148940
rect 122156 148928 122162 148980
rect 128630 148928 128636 148980
rect 128688 148968 128694 148980
rect 149698 148968 149704 148980
rect 128688 148940 149704 148968
rect 128688 148928 128694 148940
rect 149698 148928 149704 148940
rect 149756 148928 149762 148980
rect 156322 148928 156328 148980
rect 156380 148968 156386 148980
rect 177298 148968 177304 148980
rect 156380 148940 177304 148968
rect 156380 148928 156386 148940
rect 177298 148928 177304 148940
rect 177356 148928 177362 148980
rect 194594 148928 194600 148980
rect 194652 148968 194658 148980
rect 206278 148968 206284 148980
rect 194652 148940 206284 148968
rect 194652 148928 194658 148940
rect 206278 148928 206284 148940
rect 206336 148928 206342 148980
rect 222930 148928 222936 148980
rect 222988 148968 222994 148980
rect 234062 148968 234068 148980
rect 222988 148940 234068 148968
rect 222988 148928 222994 148940
rect 234062 148928 234068 148940
rect 234120 148928 234126 148980
rect 240318 148928 240324 148980
rect 240376 148968 240382 148980
rect 262858 148968 262864 148980
rect 240376 148940 262864 148968
rect 240376 148928 240382 148940
rect 262858 148928 262864 148940
rect 262916 148928 262922 148980
rect 278590 148928 278596 148980
rect 278648 148968 278654 148980
rect 289170 148968 289176 148980
rect 278648 148940 289176 148968
rect 278648 148928 278654 148940
rect 289170 148928 289176 148940
rect 289228 148928 289234 148980
rect 306926 148928 306932 148980
rect 306984 148968 306990 148980
rect 318058 148968 318064 148980
rect 306984 148940 318064 148968
rect 306984 148928 306990 148940
rect 318058 148928 318064 148940
rect 318116 148928 318122 148980
rect 324314 148928 324320 148980
rect 324372 148968 324378 148980
rect 345842 148968 345848 148980
rect 324372 148940 345848 148968
rect 324372 148928 324378 148940
rect 345842 148928 345848 148940
rect 345900 148928 345906 148980
rect 352650 148928 352656 148980
rect 352708 148968 352714 148980
rect 373258 148968 373264 148980
rect 352708 148940 373264 148968
rect 352708 148928 352714 148940
rect 373258 148928 373264 148940
rect 373316 148928 373322 148980
rect 390646 148928 390652 148980
rect 390704 148968 390710 148980
rect 402238 148968 402244 148980
rect 390704 148940 402244 148968
rect 390704 148928 390710 148940
rect 402238 148928 402244 148940
rect 402296 148928 402302 148980
rect 418614 148928 418620 148980
rect 418672 148968 418678 148980
rect 429930 148968 429936 148980
rect 418672 148940 429936 148968
rect 418672 148928 418678 148940
rect 429930 148928 429936 148940
rect 429988 148928 429994 148980
rect 436646 148928 436652 148980
rect 436704 148968 436710 148980
rect 457438 148968 457444 148980
rect 436704 148940 457444 148968
rect 436704 148928 436710 148940
rect 457438 148928 457444 148940
rect 457496 148928 457502 148980
rect 474642 148928 474648 148980
rect 474700 148968 474706 148980
rect 486418 148968 486424 148980
rect 474700 148940 486424 148968
rect 474700 148928 474706 148940
rect 486418 148928 486424 148940
rect 486476 148928 486482 148980
rect 502610 148928 502616 148980
rect 502668 148968 502674 148980
rect 514018 148968 514024 148980
rect 502668 148940 514024 148968
rect 502668 148928 502674 148940
rect 514018 148928 514024 148940
rect 514076 148928 514082 148980
rect 520642 148928 520648 148980
rect 520700 148968 520706 148980
rect 541618 148968 541624 148980
rect 520700 148940 541624 148968
rect 520700 148928 520706 148940
rect 541618 148928 541624 148940
rect 541676 148928 541682 148980
rect 54846 148860 54852 148912
rect 54904 148900 54910 148912
rect 71130 148900 71136 148912
rect 54904 148872 71136 148900
rect 54904 148860 54910 148872
rect 71130 148860 71136 148872
rect 71188 148860 71194 148912
rect 138934 148860 138940 148912
rect 138992 148900 138998 148912
rect 155218 148900 155224 148912
rect 138992 148872 155224 148900
rect 138992 148860 138998 148872
rect 155218 148860 155224 148872
rect 155276 148860 155282 148912
rect 166626 148860 166632 148912
rect 166684 148900 166690 148912
rect 178678 148900 178684 148912
rect 166684 148872 178684 148900
rect 166684 148860 166690 148872
rect 178678 148860 178684 148872
rect 178736 148860 178742 148912
rect 250622 148860 250628 148912
rect 250680 148900 250686 148912
rect 264238 148900 264244 148912
rect 250680 148872 264244 148900
rect 250680 148860 250686 148872
rect 264238 148860 264244 148872
rect 264296 148860 264302 148912
rect 334618 148860 334624 148912
rect 334676 148900 334682 148912
rect 345750 148900 345756 148912
rect 334676 148872 345756 148900
rect 334676 148860 334682 148872
rect 345750 148860 345756 148872
rect 345808 148860 345814 148912
rect 362862 148860 362868 148912
rect 362920 148900 362926 148912
rect 374638 148900 374644 148912
rect 362920 148872 374644 148900
rect 362920 148860 362926 148872
rect 374638 148860 374644 148872
rect 374696 148860 374702 148912
rect 446950 148860 446956 148912
rect 447008 148900 447014 148912
rect 463694 148900 463700 148912
rect 447008 148872 463700 148900
rect 447008 148860 447014 148872
rect 463694 148860 463700 148872
rect 463752 148860 463758 148912
rect 530946 148860 530952 148912
rect 531004 148900 531010 148912
rect 547138 148900 547144 148912
rect 531004 148872 547144 148900
rect 531004 148860 531010 148872
rect 547138 148860 547144 148872
rect 547196 148860 547202 148912
rect 44634 148792 44640 148844
rect 44692 148832 44698 148844
rect 66898 148832 66904 148844
rect 44692 148804 66904 148832
rect 44692 148792 44698 148804
rect 66898 148792 66904 148804
rect 66956 148792 66962 148844
rect 558638 148316 558644 148368
rect 558696 148356 558702 148368
rect 568942 148356 568948 148368
rect 558696 148328 568948 148356
rect 558696 148316 558702 148328
rect 568942 148316 568948 148328
rect 569000 148316 569006 148368
rect 548334 146888 548340 146940
rect 548392 146928 548398 146940
rect 569034 146928 569040 146940
rect 548392 146900 569040 146928
rect 548392 146888 548398 146900
rect 569034 146888 569040 146900
rect 569092 146888 569098 146940
rect 156322 146480 156328 146532
rect 156380 146520 156386 146532
rect 180058 146520 180064 146532
rect 156380 146492 180064 146520
rect 156380 146480 156386 146492
rect 180058 146480 180064 146492
rect 180116 146480 180122 146532
rect 184014 146480 184020 146532
rect 184072 146520 184078 146532
rect 204898 146520 204904 146532
rect 184072 146492 204904 146520
rect 184072 146480 184078 146492
rect 204898 146480 204904 146492
rect 204956 146480 204962 146532
rect 268010 146480 268016 146532
rect 268068 146520 268074 146532
rect 289078 146520 289084 146532
rect 268068 146492 289084 146520
rect 268068 146480 268074 146492
rect 289078 146480 289084 146492
rect 289136 146480 289142 146532
rect 176838 146412 176844 146464
rect 176896 146452 176902 146464
rect 194318 146452 194324 146464
rect 176896 146424 194324 146452
rect 176896 146412 176902 146424
rect 194318 146412 194324 146424
rect 194376 146412 194382 146464
rect 262858 146412 262864 146464
rect 262916 146452 262922 146464
rect 278314 146452 278320 146464
rect 262916 146424 278320 146452
rect 262916 146412 262922 146424
rect 278314 146412 278320 146424
rect 278372 146412 278378 146464
rect 380342 146412 380348 146464
rect 380400 146452 380406 146464
rect 401042 146452 401048 146464
rect 380400 146424 401048 146452
rect 380400 146412 380406 146424
rect 401042 146412 401048 146424
rect 401100 146412 401106 146464
rect 38194 146344 38200 146396
rect 38252 146384 38258 146396
rect 54294 146384 54300 146396
rect 38252 146356 54300 146384
rect 38252 146344 38258 146356
rect 54294 146344 54300 146356
rect 54352 146344 54358 146396
rect 65886 146344 65892 146396
rect 65944 146384 65950 146396
rect 81986 146384 81992 146396
rect 65944 146356 81992 146384
rect 65944 146344 65950 146356
rect 81986 146344 81992 146356
rect 82044 146344 82050 146396
rect 92934 146344 92940 146396
rect 92992 146384 92998 146396
rect 110322 146384 110328 146396
rect 92992 146356 110328 146384
rect 92992 146344 92998 146356
rect 110322 146344 110328 146356
rect 110380 146344 110386 146396
rect 120994 146344 121000 146396
rect 121052 146384 121058 146396
rect 138290 146384 138296 146396
rect 121052 146356 138296 146384
rect 121052 146344 121058 146356
rect 138290 146344 138296 146356
rect 138348 146344 138354 146396
rect 155218 146344 155224 146396
rect 155276 146384 155282 146396
rect 165982 146384 165988 146396
rect 155276 146356 165988 146384
rect 155276 146344 155282 146356
rect 165982 146344 165988 146356
rect 166040 146344 166046 146396
rect 204806 146344 204812 146396
rect 204864 146384 204870 146396
rect 222194 146384 222200 146396
rect 204864 146356 222200 146384
rect 204864 146344 204870 146356
rect 222194 146344 222200 146356
rect 222252 146344 222258 146396
rect 232774 146344 232780 146396
rect 232832 146384 232838 146396
rect 250346 146384 250352 146396
rect 232832 146356 250352 146384
rect 232832 146344 232838 146356
rect 250346 146344 250352 146356
rect 250404 146344 250410 146396
rect 288802 146344 288808 146396
rect 288860 146384 288866 146396
rect 306006 146384 306012 146396
rect 288860 146356 306012 146384
rect 288860 146344 288866 146356
rect 306006 146344 306012 146356
rect 306064 146344 306070 146396
rect 316770 146344 316776 146396
rect 316828 146384 316834 146396
rect 334342 146384 334348 146396
rect 316828 146356 334348 146384
rect 316828 146344 316834 146356
rect 334342 146344 334348 146356
rect 334400 146344 334406 146396
rect 372890 146344 372896 146396
rect 372948 146384 372954 146396
rect 390002 146384 390008 146396
rect 372948 146356 390008 146384
rect 372948 146344 372954 146356
rect 390002 146344 390008 146356
rect 390060 146344 390066 146396
rect 457438 146344 457444 146396
rect 457496 146384 457502 146396
rect 473998 146384 474004 146396
rect 457496 146356 474004 146384
rect 457496 146344 457502 146356
rect 473998 146344 474004 146356
rect 474056 146344 474062 146396
rect 484854 146344 484860 146396
rect 484912 146384 484918 146396
rect 502334 146384 502340 146396
rect 484912 146356 502340 146384
rect 484912 146344 484918 146356
rect 502334 146344 502340 146356
rect 502392 146344 502398 146396
rect 512730 146344 512736 146396
rect 512788 146384 512794 146396
rect 530302 146384 530308 146396
rect 512788 146356 530308 146384
rect 512788 146344 512794 146356
rect 530302 146344 530308 146356
rect 530360 146344 530366 146396
rect 15286 146276 15292 146328
rect 15344 146316 15350 146328
rect 26326 146316 26332 146328
rect 15344 146288 26332 146316
rect 15344 146276 15350 146288
rect 26326 146276 26332 146288
rect 26384 146276 26390 146328
rect 38102 146276 38108 146328
rect 38160 146316 38166 146328
rect 64598 146316 64604 146328
rect 38160 146288 64604 146316
rect 38160 146276 38166 146288
rect 64598 146276 64604 146288
rect 64656 146276 64662 146328
rect 72326 146276 72332 146328
rect 72384 146316 72390 146328
rect 93118 146316 93124 146328
rect 72384 146288 93124 146316
rect 72384 146276 72390 146288
rect 93118 146276 93124 146288
rect 93176 146276 93182 146328
rect 100018 146276 100024 146328
rect 100076 146316 100082 146328
rect 121086 146316 121092 146328
rect 100076 146288 121092 146316
rect 100076 146276 100082 146288
rect 121086 146276 121092 146288
rect 121144 146276 121150 146328
rect 122098 146276 122104 146328
rect 122156 146316 122162 146328
rect 148594 146316 148600 146328
rect 122156 146288 148600 146316
rect 122156 146276 122162 146288
rect 148594 146276 148600 146288
rect 148652 146276 148658 146328
rect 178678 146276 178684 146328
rect 178736 146316 178742 146328
rect 204622 146316 204628 146328
rect 178736 146288 204628 146316
rect 178736 146276 178742 146288
rect 204622 146276 204628 146288
rect 204680 146276 204686 146328
rect 206278 146276 206284 146328
rect 206336 146316 206342 146328
rect 232314 146316 232320 146328
rect 206336 146288 232320 146316
rect 206336 146276 206342 146288
rect 232314 146276 232320 146288
rect 232372 146276 232378 146328
rect 233970 146276 233976 146328
rect 234028 146316 234034 146328
rect 260650 146316 260656 146328
rect 234028 146288 260656 146316
rect 234028 146276 234034 146288
rect 260650 146276 260656 146288
rect 260708 146276 260714 146328
rect 261478 146276 261484 146328
rect 261536 146316 261542 146328
rect 288618 146316 288624 146328
rect 261536 146288 288624 146316
rect 261536 146276 261542 146288
rect 288618 146276 288624 146288
rect 288676 146276 288682 146328
rect 290458 146276 290464 146328
rect 290516 146316 290522 146328
rect 316310 146316 316316 146328
rect 290516 146288 316316 146316
rect 290516 146276 290522 146288
rect 316310 146276 316316 146288
rect 316368 146276 316374 146328
rect 316862 146276 316868 146328
rect 316920 146316 316926 146328
rect 344646 146316 344652 146328
rect 316920 146288 344652 146316
rect 316920 146276 316926 146288
rect 344646 146276 344652 146288
rect 344704 146276 344710 146328
rect 352006 146276 352012 146328
rect 352064 146316 352070 146328
rect 373258 146316 373264 146328
rect 352064 146288 373264 146316
rect 352064 146276 352070 146288
rect 373258 146276 373264 146288
rect 373316 146276 373322 146328
rect 401134 146276 401140 146328
rect 401192 146316 401198 146328
rect 418338 146316 418344 146328
rect 401192 146288 418344 146316
rect 401192 146276 401198 146288
rect 418338 146276 418344 146288
rect 418396 146276 418402 146328
rect 429838 146276 429844 146328
rect 429896 146316 429902 146328
rect 456610 146316 456616 146328
rect 429896 146288 456616 146316
rect 429896 146276 429902 146288
rect 456610 146276 456616 146288
rect 456668 146276 456674 146328
rect 464338 146276 464344 146328
rect 464396 146316 464402 146328
rect 485038 146316 485044 146328
rect 464396 146288 485044 146316
rect 464396 146276 464402 146288
rect 485038 146276 485044 146288
rect 485096 146276 485102 146328
rect 486418 146276 486424 146328
rect 486476 146316 486482 146328
rect 512638 146316 512644 146328
rect 486476 146288 512644 146316
rect 486476 146276 486482 146288
rect 512638 146276 512644 146288
rect 512696 146276 512702 146328
rect 514018 146276 514024 146328
rect 514076 146316 514082 146328
rect 540606 146316 540612 146328
rect 514076 146288 540612 146316
rect 514076 146276 514082 146288
rect 540606 146276 540612 146288
rect 540664 146276 540670 146328
rect 547138 146276 547144 146328
rect 547196 146316 547202 146328
rect 557994 146316 558000 146328
rect 547196 146288 558000 146316
rect 547196 146276 547202 146288
rect 557994 146276 558000 146288
rect 558052 146276 558058 146328
rect 120718 144236 120724 144288
rect 120776 144276 120782 144288
rect 120994 144276 121000 144288
rect 120776 144248 121000 144276
rect 120776 144236 120782 144248
rect 120994 144236 121000 144248
rect 121052 144236 121058 144288
rect 92750 144168 92756 144220
rect 92808 144208 92814 144220
rect 92934 144208 92940 144220
rect 92808 144180 92940 144208
rect 92808 144168 92814 144180
rect 92934 144168 92940 144180
rect 92992 144168 92998 144220
rect 400766 144168 400772 144220
rect 400824 144208 400830 144220
rect 401134 144208 401140 144220
rect 400824 144180 401140 144208
rect 400824 144168 400830 144180
rect 401134 144168 401140 144180
rect 401192 144168 401198 144220
rect 120810 144100 120816 144152
rect 120868 144140 120874 144152
rect 121086 144140 121092 144152
rect 120868 144112 121092 144140
rect 120868 144100 120874 144112
rect 121086 144100 121092 144112
rect 121144 144100 121150 144152
rect 400858 144100 400864 144152
rect 400916 144140 400922 144152
rect 401042 144140 401048 144152
rect 400916 144112 401048 144140
rect 400916 144100 400922 144112
rect 401042 144100 401048 144112
rect 401100 144100 401106 144152
rect 154482 143624 154488 143676
rect 154540 143664 154546 143676
rect 207014 143664 207020 143676
rect 154540 143636 207020 143664
rect 154540 143624 154546 143636
rect 207014 143624 207020 143636
rect 207072 143624 207078 143676
rect 182082 143556 182088 143608
rect 182140 143596 182146 143608
rect 234706 143596 234712 143608
rect 182140 143568 234712 143596
rect 182140 143556 182146 143568
rect 234706 143556 234712 143568
rect 234764 143556 234770 143608
rect 568758 142808 568764 142860
rect 568816 142848 568822 142860
rect 568942 142848 568948 142860
rect 568816 142820 568948 142848
rect 568816 142808 568822 142820
rect 568942 142808 568948 142820
rect 569000 142808 569006 142860
rect 3326 136688 3332 136740
rect 3384 136728 3390 136740
rect 7558 136728 7564 136740
rect 3384 136700 7564 136728
rect 3384 136688 3390 136700
rect 7558 136688 7564 136700
rect 7616 136688 7622 136740
rect 64874 128596 64880 128648
rect 64932 128636 64938 128648
rect 65886 128636 65892 128648
rect 64932 128608 65892 128636
rect 64932 128596 64938 128608
rect 65886 128596 65892 128608
rect 65944 128596 65950 128648
rect 204898 128256 204904 128308
rect 204956 128296 204962 128308
rect 211706 128296 211712 128308
rect 204956 128268 211712 128296
rect 204956 128256 204962 128268
rect 211706 128256 211712 128268
rect 211764 128256 211770 128308
rect 485038 128256 485044 128308
rect 485096 128296 485102 128308
rect 491662 128296 491668 128308
rect 485096 128268 491668 128296
rect 485096 128256 485102 128268
rect 491662 128256 491668 128268
rect 491720 128256 491726 128308
rect 289078 127984 289084 128036
rect 289136 128024 289142 128036
rect 295702 128024 295708 128036
rect 289136 127996 295708 128024
rect 289136 127984 289142 127996
rect 295702 127984 295708 127996
rect 295760 127984 295766 128036
rect 93118 127576 93124 127628
rect 93176 127616 93182 127628
rect 99742 127616 99748 127628
rect 93176 127588 99748 127616
rect 93176 127576 93182 127588
rect 99742 127576 99748 127588
rect 99800 127576 99806 127628
rect 120810 127576 120816 127628
rect 120868 127616 120874 127628
rect 127710 127616 127716 127628
rect 120868 127588 127716 127616
rect 120868 127576 120874 127588
rect 127710 127576 127716 127588
rect 127768 127576 127774 127628
rect 373258 127576 373264 127628
rect 373316 127616 373322 127628
rect 379698 127616 379704 127628
rect 373316 127588 379704 127616
rect 373316 127576 373322 127588
rect 379698 127576 379704 127588
rect 379756 127576 379762 127628
rect 400858 127576 400864 127628
rect 400916 127616 400922 127628
rect 407758 127616 407764 127628
rect 400916 127588 407764 127616
rect 400916 127576 400922 127588
rect 407758 127576 407764 127588
rect 407816 127576 407822 127628
rect 42702 125536 42708 125588
rect 42760 125576 42766 125588
rect 95234 125576 95240 125588
rect 42760 125548 95240 125576
rect 42760 125536 42766 125548
rect 95234 125536 95240 125548
rect 95292 125536 95298 125588
rect 97902 125536 97908 125588
rect 97960 125576 97966 125588
rect 150434 125576 150440 125588
rect 97960 125548 150440 125576
rect 97960 125536 97966 125548
rect 150434 125536 150440 125548
rect 150492 125536 150498 125588
rect 238662 125536 238668 125588
rect 238720 125576 238726 125588
rect 291194 125576 291200 125588
rect 238720 125548 291200 125576
rect 238720 125536 238726 125548
rect 291194 125536 291200 125548
rect 291252 125536 291258 125588
rect 293862 125536 293868 125588
rect 293920 125576 293926 125588
rect 346394 125576 346400 125588
rect 293920 125548 346400 125576
rect 293920 125536 293926 125548
rect 346394 125536 346400 125548
rect 346452 125536 346458 125588
rect 350442 125536 350448 125588
rect 350500 125576 350506 125588
rect 402974 125576 402980 125588
rect 350500 125548 402980 125576
rect 350500 125536 350506 125548
rect 402974 125536 402980 125548
rect 403032 125536 403038 125588
rect 405642 125536 405648 125588
rect 405700 125576 405706 125588
rect 458174 125576 458180 125588
rect 405700 125548 458180 125576
rect 405700 125536 405706 125548
rect 458174 125536 458180 125548
rect 458232 125536 458238 125588
rect 462222 125536 462228 125588
rect 462280 125576 462286 125588
rect 514754 125576 514760 125588
rect 462280 125548 514760 125576
rect 462280 125536 462286 125548
rect 514754 125536 514760 125548
rect 514812 125536 514818 125588
rect 518802 125536 518808 125588
rect 518860 125576 518866 125588
rect 571334 125576 571340 125588
rect 518860 125548 571340 125576
rect 518860 125536 518866 125548
rect 571334 125536 571340 125548
rect 571392 125536 571398 125588
rect 176746 124856 176752 124908
rect 176804 124856 176810 124908
rect 372798 124856 372804 124908
rect 372856 124856 372862 124908
rect 484762 124856 484768 124908
rect 484820 124856 484826 124908
rect 176764 124704 176792 124856
rect 372816 124704 372844 124856
rect 484780 124704 484808 124856
rect 15286 124652 15292 124704
rect 15344 124692 15350 124704
rect 16114 124692 16120 124704
rect 15344 124664 16120 124692
rect 15344 124652 15350 124664
rect 16114 124652 16120 124664
rect 16172 124652 16178 124704
rect 36538 124652 36544 124704
rect 36596 124692 36602 124704
rect 38194 124692 38200 124704
rect 36596 124664 38200 124692
rect 36596 124652 36602 124664
rect 38194 124652 38200 124664
rect 38252 124652 38258 124704
rect 176746 124652 176752 124704
rect 176804 124652 176810 124704
rect 372798 124652 372804 124704
rect 372856 124652 372862 124704
rect 484762 124652 484768 124704
rect 484820 124652 484826 124704
rect 547874 124652 547880 124704
rect 547932 124692 547938 124704
rect 548150 124692 548156 124704
rect 547932 124664 548156 124692
rect 547932 124652 547938 124664
rect 548150 124652 548156 124664
rect 548208 124652 548214 124704
rect 110322 122748 110328 122800
rect 110380 122788 110386 122800
rect 122098 122788 122104 122800
rect 110380 122760 122104 122788
rect 110380 122748 110386 122760
rect 122098 122748 122104 122760
rect 122156 122748 122162 122800
rect 138290 122748 138296 122800
rect 138348 122788 138354 122800
rect 176746 122788 176752 122800
rect 138348 122760 176752 122788
rect 138348 122748 138354 122760
rect 176746 122748 176752 122760
rect 176804 122748 176810 122800
rect 180058 122748 180064 122800
rect 180116 122788 180122 122800
rect 184014 122788 184020 122800
rect 180116 122760 184020 122788
rect 180116 122748 180122 122760
rect 184014 122748 184020 122760
rect 184072 122748 184078 122800
rect 194318 122748 194324 122800
rect 194376 122788 194382 122800
rect 206278 122788 206284 122800
rect 194376 122760 206284 122788
rect 194376 122748 194382 122760
rect 206278 122748 206284 122760
rect 206336 122748 206342 122800
rect 211246 122748 211252 122800
rect 211304 122788 211310 122800
rect 240042 122788 240048 122800
rect 211304 122760 240048 122788
rect 211304 122748 211310 122760
rect 240042 122748 240048 122760
rect 240100 122748 240106 122800
rect 260650 122748 260656 122800
rect 260708 122788 260714 122800
rect 262858 122788 262864 122800
rect 260708 122760 262864 122788
rect 260708 122748 260714 122760
rect 262858 122748 262864 122760
rect 262916 122748 262922 122800
rect 278314 122748 278320 122800
rect 278372 122788 278378 122800
rect 290458 122788 290464 122800
rect 278372 122760 290464 122788
rect 278372 122748 278378 122760
rect 290458 122748 290464 122760
rect 290516 122748 290522 122800
rect 295426 122748 295432 122800
rect 295484 122788 295490 122800
rect 324038 122788 324044 122800
rect 295484 122760 324044 122788
rect 295484 122748 295490 122760
rect 324038 122748 324044 122760
rect 324096 122748 324102 122800
rect 334342 122748 334348 122800
rect 334400 122788 334406 122800
rect 372798 122788 372804 122800
rect 334400 122760 372804 122788
rect 334400 122748 334406 122760
rect 372798 122748 372804 122760
rect 372856 122748 372862 122800
rect 390462 122748 390468 122800
rect 390520 122788 390526 122800
rect 428734 122788 428740 122800
rect 390520 122760 428740 122788
rect 390520 122748 390526 122760
rect 428734 122748 428740 122760
rect 428792 122748 428798 122800
rect 434806 122748 434812 122800
rect 434864 122788 434870 122800
rect 434864 122760 441614 122788
rect 434864 122748 434870 122760
rect 26326 122680 26332 122732
rect 26384 122720 26390 122732
rect 38102 122720 38108 122732
rect 26384 122692 38108 122720
rect 26384 122680 26390 122692
rect 38102 122680 38108 122692
rect 38160 122680 38166 122732
rect 42886 122680 42892 122732
rect 42944 122720 42950 122732
rect 71774 122720 71780 122732
rect 42944 122692 71780 122720
rect 42944 122680 42950 122692
rect 71774 122680 71780 122692
rect 71832 122680 71838 122732
rect 82630 122680 82636 122732
rect 82688 122720 82694 122732
rect 120902 122720 120908 122732
rect 82688 122692 120908 122720
rect 82688 122680 82694 122692
rect 120902 122680 120908 122692
rect 120960 122680 120966 122732
rect 127066 122680 127072 122732
rect 127124 122720 127130 122732
rect 155954 122720 155960 122732
rect 127124 122692 155960 122720
rect 127124 122680 127130 122692
rect 155954 122680 155960 122692
rect 156012 122680 156018 122732
rect 166626 122680 166632 122732
rect 166684 122720 166690 122732
rect 178678 122720 178684 122732
rect 166684 122692 178684 122720
rect 166684 122680 166690 122692
rect 178678 122680 178684 122692
rect 178736 122680 178742 122732
rect 222654 122680 222660 122732
rect 222712 122720 222718 122732
rect 233970 122720 233976 122732
rect 222712 122692 233976 122720
rect 222712 122680 222718 122692
rect 233970 122680 233976 122692
rect 234028 122680 234034 122732
rect 250346 122680 250352 122732
rect 250404 122720 250410 122732
rect 261478 122720 261484 122732
rect 250404 122692 261484 122720
rect 250404 122680 250410 122692
rect 261478 122680 261484 122692
rect 261536 122680 261542 122732
rect 306282 122680 306288 122732
rect 306340 122720 306346 122732
rect 316862 122720 316868 122732
rect 306340 122692 316868 122720
rect 306340 122680 306346 122692
rect 316862 122680 316868 122692
rect 316920 122680 316926 122732
rect 323026 122680 323032 122732
rect 323084 122720 323090 122732
rect 352006 122720 352012 122732
rect 323084 122692 352012 122720
rect 323084 122680 323090 122692
rect 352006 122680 352012 122692
rect 352064 122680 352070 122732
rect 362310 122680 362316 122732
rect 362368 122720 362374 122732
rect 400950 122720 400956 122732
rect 362368 122692 400956 122720
rect 362368 122680 362374 122692
rect 400950 122680 400956 122692
rect 401008 122680 401014 122732
rect 407206 122680 407212 122732
rect 407264 122720 407270 122732
rect 436002 122720 436008 122732
rect 407264 122692 436008 122720
rect 407264 122680 407270 122692
rect 436002 122680 436008 122692
rect 436060 122680 436066 122732
rect 441586 122720 441614 122760
rect 491386 122748 491392 122800
rect 491444 122788 491450 122800
rect 519998 122788 520004 122800
rect 491444 122760 520004 122788
rect 491444 122748 491450 122760
rect 519998 122748 520004 122760
rect 520056 122748 520062 122800
rect 530302 122748 530308 122800
rect 530360 122788 530366 122800
rect 568850 122788 568856 122800
rect 530360 122760 568856 122788
rect 530360 122748 530366 122760
rect 568850 122748 568856 122760
rect 568908 122748 568914 122800
rect 463786 122720 463792 122732
rect 441586 122692 463792 122720
rect 463786 122680 463792 122692
rect 463844 122680 463850 122732
rect 474642 122680 474648 122732
rect 474700 122720 474706 122732
rect 486418 122720 486424 122732
rect 474700 122692 486424 122720
rect 474700 122680 474706 122692
rect 486418 122680 486424 122692
rect 486476 122680 486482 122732
rect 502334 122680 502340 122732
rect 502392 122720 502398 122732
rect 514018 122720 514024 122732
rect 502392 122692 514024 122720
rect 502392 122680 502398 122692
rect 514018 122680 514024 122692
rect 514076 122680 514082 122732
rect 540606 122680 540612 122732
rect 540664 122720 540670 122732
rect 547138 122720 547144 122732
rect 540664 122692 547144 122720
rect 540664 122680 540670 122692
rect 547138 122680 547144 122692
rect 547196 122680 547202 122732
rect 548150 122680 548156 122732
rect 548208 122720 548214 122732
rect 557994 122720 558000 122732
rect 548208 122692 558000 122720
rect 548208 122680 548214 122692
rect 557994 122680 558000 122692
rect 558052 122680 558058 122732
rect 15378 122612 15384 122664
rect 15436 122652 15442 122664
rect 43990 122652 43996 122664
rect 15436 122624 43996 122652
rect 15436 122612 15442 122624
rect 43990 122612 43996 122624
rect 44048 122612 44054 122664
rect 54294 122612 54300 122664
rect 54352 122652 54358 122664
rect 92842 122652 92848 122664
rect 54352 122624 92848 122652
rect 54352 122612 54358 122624
rect 92842 122612 92848 122624
rect 92900 122612 92906 122664
rect 148594 122612 148600 122664
rect 148652 122652 148658 122664
rect 155218 122652 155224 122664
rect 148652 122624 155224 122652
rect 148652 122612 148658 122624
rect 155218 122612 155224 122624
rect 155276 122612 155282 122664
rect 238846 122612 238852 122664
rect 238904 122652 238910 122664
rect 268010 122652 268016 122664
rect 238904 122624 268016 122652
rect 238904 122612 238910 122624
rect 268010 122612 268016 122624
rect 268068 122612 268074 122664
rect 418338 122612 418344 122664
rect 418396 122652 418402 122664
rect 429838 122652 429844 122664
rect 418396 122624 429844 122652
rect 418396 122612 418402 122624
rect 429838 122612 429844 122624
rect 429896 122612 429902 122664
rect 446306 122612 446312 122664
rect 446364 122652 446370 122664
rect 484762 122652 484768 122664
rect 446364 122624 484768 122652
rect 446364 122612 446370 122624
rect 484762 122612 484768 122624
rect 484820 122612 484826 122664
rect 518986 122544 518992 122596
rect 519044 122584 519050 122596
rect 547874 122584 547880 122596
rect 519044 122556 547880 122584
rect 519044 122544 519050 122556
rect 547874 122544 547880 122556
rect 547932 122544 547938 122596
rect 26602 120708 26608 120760
rect 26660 120748 26666 120760
rect 36722 120748 36728 120760
rect 26660 120720 36728 120748
rect 26660 120708 26666 120720
rect 36722 120708 36728 120720
rect 36780 120708 36786 120760
rect 15562 120232 15568 120284
rect 15620 120272 15626 120284
rect 54294 120272 54300 120284
rect 15620 120244 54300 120272
rect 15620 120232 15626 120244
rect 54294 120232 54300 120244
rect 54352 120232 54358 120284
rect 149698 120232 149704 120284
rect 149756 120272 149762 120284
rect 166626 120272 166632 120284
rect 149756 120244 166632 120272
rect 149756 120232 149762 120244
rect 166626 120232 166632 120244
rect 166684 120232 166690 120284
rect 211154 120232 211160 120284
rect 211212 120272 211218 120284
rect 250622 120272 250628 120284
rect 211212 120244 250628 120272
rect 211212 120232 211218 120244
rect 250622 120232 250628 120244
rect 250680 120232 250686 120284
rect 295426 120232 295432 120284
rect 295484 120272 295490 120284
rect 295484 120244 296714 120272
rect 295484 120232 295490 120244
rect 71774 120164 71780 120216
rect 71832 120204 71838 120216
rect 110598 120204 110604 120216
rect 71832 120176 110604 120204
rect 71832 120164 71838 120176
rect 110598 120164 110604 120176
rect 110656 120164 110662 120216
rect 122098 120164 122104 120216
rect 122156 120204 122162 120216
rect 128354 120204 128360 120216
rect 122156 120176 128360 120204
rect 122156 120164 122162 120176
rect 128354 120164 128360 120176
rect 128412 120164 128418 120216
rect 149790 120164 149796 120216
rect 149848 120204 149854 120216
rect 156322 120204 156328 120216
rect 149848 120176 156328 120204
rect 149848 120164 149854 120176
rect 156322 120164 156328 120176
rect 156380 120164 156386 120216
rect 183554 120164 183560 120216
rect 183612 120204 183618 120216
rect 222286 120204 222292 120216
rect 183612 120176 222292 120204
rect 183612 120164 183618 120176
rect 222286 120164 222292 120176
rect 222344 120164 222350 120216
rect 262858 120164 262864 120216
rect 262916 120204 262922 120216
rect 278222 120204 278228 120216
rect 262916 120176 278228 120204
rect 262916 120164 262922 120176
rect 278222 120164 278228 120176
rect 278280 120164 278286 120216
rect 290458 120164 290464 120216
rect 290516 120204 290522 120216
rect 295978 120204 295984 120216
rect 290516 120176 295984 120204
rect 290516 120164 290522 120176
rect 295978 120164 295984 120176
rect 296036 120164 296042 120216
rect 296686 120204 296714 120244
rect 407206 120232 407212 120284
rect 407264 120272 407270 120284
rect 407264 120244 412634 120272
rect 407264 120232 407270 120244
rect 334618 120204 334624 120216
rect 296686 120176 334624 120204
rect 334618 120164 334624 120176
rect 334676 120164 334682 120216
rect 378870 120164 378876 120216
rect 378928 120204 378934 120216
rect 390738 120204 390744 120216
rect 378928 120176 390744 120204
rect 378928 120164 378934 120176
rect 390738 120164 390744 120176
rect 390796 120164 390802 120216
rect 402238 120164 402244 120216
rect 402296 120204 402302 120216
rect 408310 120204 408316 120216
rect 402296 120176 408316 120204
rect 402296 120164 402302 120176
rect 408310 120164 408316 120176
rect 408368 120164 408374 120216
rect 412606 120204 412634 120244
rect 429838 120232 429844 120284
rect 429896 120272 429902 120284
rect 436094 120272 436100 120284
rect 429896 120244 436100 120272
rect 429896 120232 429902 120244
rect 436094 120232 436100 120244
rect 436152 120232 436158 120284
rect 491386 120232 491392 120284
rect 491444 120272 491450 120284
rect 491444 120244 499574 120272
rect 491444 120232 491450 120244
rect 446306 120204 446312 120216
rect 412606 120176 446312 120204
rect 446306 120164 446312 120176
rect 446364 120164 446370 120216
rect 457438 120164 457444 120216
rect 457496 120204 457502 120216
rect 474366 120204 474372 120216
rect 457496 120176 474372 120204
rect 457496 120164 457502 120176
rect 474366 120164 474372 120176
rect 474424 120164 474430 120216
rect 486418 120164 486424 120216
rect 486476 120204 486482 120216
rect 492306 120204 492312 120216
rect 486476 120176 492312 120204
rect 486476 120164 486482 120176
rect 492306 120164 492312 120176
rect 492364 120164 492370 120216
rect 499546 120204 499574 120244
rect 541618 120232 541624 120284
rect 541676 120272 541682 120284
rect 558638 120272 558644 120284
rect 541676 120244 558644 120272
rect 541676 120232 541682 120244
rect 558638 120232 558644 120244
rect 558696 120232 558702 120284
rect 530302 120204 530308 120216
rect 499546 120176 530308 120204
rect 530302 120164 530308 120176
rect 530360 120164 530366 120216
rect 36906 120096 36912 120148
rect 36964 120136 36970 120148
rect 43438 120136 43444 120148
rect 36964 120108 43444 120136
rect 36964 120096 36970 120108
rect 43438 120096 43444 120108
rect 43496 120096 43502 120148
rect 65886 120096 65892 120148
rect 65944 120136 65950 120148
rect 82630 120136 82636 120148
rect 65944 120108 82636 120136
rect 65944 120096 65950 120108
rect 82630 120096 82636 120108
rect 82688 120096 82694 120148
rect 99374 120096 99380 120148
rect 99432 120136 99438 120148
rect 138290 120136 138296 120148
rect 99432 120108 138296 120136
rect 99432 120096 99438 120108
rect 138290 120096 138296 120108
rect 138348 120096 138354 120148
rect 233970 120096 233976 120148
rect 234028 120136 234034 120148
rect 240318 120136 240324 120148
rect 234028 120108 240324 120136
rect 234028 120096 234034 120108
rect 240318 120096 240324 120108
rect 240376 120096 240382 120148
rect 267826 120096 267832 120148
rect 267884 120136 267890 120148
rect 306466 120136 306472 120148
rect 267884 120108 306472 120136
rect 267884 120096 267890 120108
rect 306466 120096 306472 120108
rect 306524 120096 306530 120148
rect 345658 120096 345664 120148
rect 345716 120136 345722 120148
rect 362310 120136 362316 120148
rect 345716 120108 362316 120136
rect 345716 120096 345722 120108
rect 362310 120096 362316 120108
rect 362368 120096 362374 120148
rect 379514 120096 379520 120148
rect 379572 120136 379578 120148
rect 418614 120136 418620 120148
rect 379572 120108 418620 120136
rect 379572 120096 379578 120108
rect 418614 120096 418620 120108
rect 418672 120096 418678 120148
rect 458818 120096 458824 120148
rect 458876 120136 458882 120148
rect 464062 120136 464068 120148
rect 458876 120108 464068 120136
rect 458876 120096 458882 120108
rect 464062 120096 464068 120108
rect 464120 120096 464126 120148
rect 502610 120136 502616 120148
rect 464172 120108 502616 120136
rect 463786 120028 463792 120080
rect 463844 120068 463850 120080
rect 464172 120068 464200 120108
rect 502610 120096 502616 120108
rect 502668 120096 502674 120148
rect 514018 120096 514024 120148
rect 514076 120136 514082 120148
rect 520274 120136 520280 120148
rect 514076 120108 520280 120136
rect 514076 120096 514082 120108
rect 520274 120096 520280 120108
rect 520332 120096 520338 120148
rect 463844 120040 464200 120068
rect 463844 120028 463850 120040
rect 205082 117376 205088 117428
rect 205140 117376 205146 117428
rect 293862 117376 293868 117428
rect 293920 117416 293926 117428
rect 346394 117416 346400 117428
rect 293920 117388 346400 117416
rect 293920 117376 293926 117388
rect 346394 117376 346400 117388
rect 346452 117376 346458 117428
rect 40678 117240 40684 117292
rect 40736 117280 40742 117292
rect 44082 117280 44088 117292
rect 40736 117252 44088 117280
rect 40736 117240 40742 117252
rect 44082 117240 44088 117252
rect 44140 117240 44146 117292
rect 205100 117224 205128 117376
rect 238662 117308 238668 117360
rect 238720 117348 238726 117360
rect 291194 117348 291200 117360
rect 238720 117320 291200 117348
rect 238720 117308 238726 117320
rect 291194 117308 291200 117320
rect 291252 117308 291258 117360
rect 322842 117308 322848 117360
rect 322900 117348 322906 117360
rect 375374 117348 375380 117360
rect 322900 117320 375380 117348
rect 322900 117308 322906 117320
rect 375374 117308 375380 117320
rect 375432 117308 375438 117360
rect 434622 117308 434628 117360
rect 434680 117348 434686 117360
rect 487154 117348 487160 117360
rect 434680 117320 487160 117348
rect 434680 117308 434686 117320
rect 487154 117308 487160 117320
rect 487212 117308 487218 117360
rect 264238 117240 264244 117292
rect 264296 117280 264302 117292
rect 267918 117280 267924 117292
rect 264296 117252 267924 117280
rect 264296 117240 264302 117252
rect 267918 117240 267924 117252
rect 267976 117240 267982 117292
rect 345014 117240 345020 117292
rect 345072 117280 345078 117292
rect 347038 117280 347044 117292
rect 345072 117252 347044 117280
rect 345072 117240 345078 117252
rect 347038 117240 347044 117252
rect 347096 117240 347102 117292
rect 348418 117240 348424 117292
rect 348476 117280 348482 117292
rect 352006 117280 352012 117292
rect 348476 117252 352012 117280
rect 348476 117240 348482 117252
rect 352006 117240 352012 117252
rect 352064 117240 352070 117292
rect 429102 117240 429108 117292
rect 429160 117280 429166 117292
rect 429930 117280 429936 117292
rect 429160 117252 429936 117280
rect 429160 117240 429166 117252
rect 429930 117240 429936 117252
rect 429988 117240 429994 117292
rect 541158 117240 541164 117292
rect 541216 117280 541222 117292
rect 544378 117280 544384 117292
rect 541216 117252 544384 117280
rect 541216 117240 541222 117252
rect 544378 117240 544384 117252
rect 544436 117240 544442 117292
rect 205082 117172 205088 117224
rect 205140 117172 205146 117224
rect 149238 115200 149244 115252
rect 149296 115240 149302 115252
rect 149882 115240 149888 115252
rect 149296 115212 149888 115240
rect 149296 115200 149302 115212
rect 149882 115200 149888 115212
rect 149940 115200 149946 115252
rect 233234 114520 233240 114572
rect 233292 114560 233298 114572
rect 234062 114560 234068 114572
rect 233292 114532 234068 114560
rect 233292 114520 233298 114532
rect 234062 114520 234068 114532
rect 234120 114520 234126 114572
rect 569494 111800 569500 111852
rect 569552 111840 569558 111852
rect 580074 111840 580080 111852
rect 569552 111812 580080 111840
rect 569552 111800 569558 111812
rect 580074 111800 580080 111812
rect 580132 111800 580138 111852
rect 99374 100240 99380 100292
rect 99432 100280 99438 100292
rect 99926 100280 99932 100292
rect 99432 100252 99932 100280
rect 99432 100240 99438 100252
rect 99926 100240 99932 100252
rect 99984 100240 99990 100292
rect 183554 100240 183560 100292
rect 183612 100280 183618 100292
rect 184014 100280 184020 100292
rect 183612 100252 184020 100280
rect 183612 100240 183618 100252
rect 184014 100240 184020 100252
rect 184072 100240 184078 100292
rect 211154 100240 211160 100292
rect 211212 100280 211218 100292
rect 211982 100280 211988 100292
rect 211212 100252 211988 100280
rect 211212 100240 211218 100252
rect 211982 100240 211988 100252
rect 212040 100240 212046 100292
rect 379514 100240 379520 100292
rect 379572 100280 379578 100292
rect 379974 100280 379980 100292
rect 379572 100252 379980 100280
rect 379572 100240 379578 100252
rect 379974 100240 379980 100252
rect 380032 100240 380038 100292
rect 71774 97520 71780 97572
rect 71832 97560 71838 97572
rect 72418 97560 72424 97572
rect 71832 97532 72424 97560
rect 71832 97520 71838 97532
rect 72418 97520 72424 97532
rect 72476 97520 72482 97572
rect 15194 95140 15200 95192
rect 15252 95180 15258 95192
rect 36906 95180 36912 95192
rect 15252 95152 36912 95180
rect 15252 95140 15258 95152
rect 36906 95140 36912 95152
rect 36964 95140 36970 95192
rect 65058 95140 65064 95192
rect 65116 95180 65122 95192
rect 92934 95180 92940 95192
rect 65116 95152 92940 95180
rect 65116 95140 65122 95152
rect 92934 95140 92940 95152
rect 92992 95140 92998 95192
rect 93026 95140 93032 95192
rect 93084 95180 93090 95192
rect 120902 95180 120908 95192
rect 93084 95152 120908 95180
rect 93084 95140 93090 95152
rect 120902 95140 120908 95152
rect 120960 95140 120966 95192
rect 121086 95140 121092 95192
rect 121144 95180 121150 95192
rect 148594 95180 148600 95192
rect 121144 95152 148600 95180
rect 121144 95140 121150 95152
rect 148594 95140 148600 95152
rect 148652 95140 148658 95192
rect 149882 95140 149888 95192
rect 149940 95180 149946 95192
rect 176930 95180 176936 95192
rect 149940 95152 176936 95180
rect 149940 95140 149946 95152
rect 176930 95140 176936 95152
rect 176988 95140 176994 95192
rect 177022 95140 177028 95192
rect 177080 95180 177086 95192
rect 204898 95180 204904 95192
rect 177080 95152 204904 95180
rect 177080 95140 177086 95152
rect 204898 95140 204904 95152
rect 204956 95140 204962 95192
rect 205174 95140 205180 95192
rect 205232 95180 205238 95192
rect 232590 95180 232596 95192
rect 205232 95152 232596 95180
rect 205232 95140 205238 95152
rect 232590 95140 232596 95152
rect 232648 95140 232654 95192
rect 234062 95140 234068 95192
rect 234120 95180 234126 95192
rect 260926 95180 260932 95192
rect 234120 95152 260932 95180
rect 234120 95140 234126 95152
rect 260926 95140 260932 95152
rect 260984 95140 260990 95192
rect 261018 95140 261024 95192
rect 261076 95180 261082 95192
rect 288894 95180 288900 95192
rect 261076 95152 288900 95180
rect 261076 95140 261082 95152
rect 288894 95140 288900 95152
rect 288952 95140 288958 95192
rect 289078 95140 289084 95192
rect 289136 95180 289142 95192
rect 316586 95180 316592 95192
rect 289136 95152 316592 95180
rect 289136 95140 289142 95152
rect 316586 95140 316592 95152
rect 316644 95140 316650 95192
rect 318058 95140 318064 95192
rect 318116 95180 318122 95192
rect 344922 95180 344928 95192
rect 318116 95152 344928 95180
rect 318116 95140 318122 95152
rect 344922 95140 344928 95152
rect 344980 95140 344986 95192
rect 347038 95140 347044 95192
rect 347096 95180 347102 95192
rect 372614 95180 372620 95192
rect 347096 95152 372620 95180
rect 347096 95140 347102 95152
rect 372614 95140 372620 95152
rect 372672 95140 372678 95192
rect 373074 95140 373080 95192
rect 373132 95180 373138 95192
rect 400950 95180 400956 95192
rect 373132 95152 400956 95180
rect 373132 95140 373138 95152
rect 400950 95140 400956 95152
rect 401008 95140 401014 95192
rect 401042 95140 401048 95192
rect 401100 95180 401106 95192
rect 428918 95180 428924 95192
rect 401100 95152 428924 95180
rect 401100 95140 401106 95152
rect 428918 95140 428924 95152
rect 428976 95140 428982 95192
rect 429930 95140 429936 95192
rect 429988 95180 429994 95192
rect 456794 95180 456800 95192
rect 429988 95152 456800 95180
rect 429988 95140 429994 95152
rect 456794 95140 456800 95152
rect 456852 95140 456858 95192
rect 457070 95140 457076 95192
rect 457128 95180 457134 95192
rect 484946 95180 484952 95192
rect 457128 95152 484952 95180
rect 457128 95140 457134 95152
rect 484946 95140 484952 95152
rect 485004 95140 485010 95192
rect 485038 95140 485044 95192
rect 485096 95180 485102 95192
rect 512914 95180 512920 95192
rect 485096 95152 512920 95180
rect 485096 95140 485102 95152
rect 512914 95140 512920 95152
rect 512972 95140 512978 95192
rect 513098 95140 513104 95192
rect 513156 95180 513162 95192
rect 540606 95180 540612 95192
rect 513156 95152 540612 95180
rect 513156 95140 513162 95152
rect 540606 95140 540612 95152
rect 540664 95140 540670 95192
rect 544378 95140 544384 95192
rect 544436 95180 544442 95192
rect 568942 95180 568948 95192
rect 544436 95152 568948 95180
rect 544436 95140 544442 95152
rect 568942 95140 568948 95152
rect 569000 95140 569006 95192
rect 26602 95072 26608 95124
rect 26660 95112 26666 95124
rect 40678 95112 40684 95124
rect 26660 95084 40684 95112
rect 26660 95072 26666 95084
rect 40678 95072 40684 95084
rect 40736 95072 40742 95124
rect 43438 95072 43444 95124
rect 43496 95112 43502 95124
rect 64874 95112 64880 95124
rect 43496 95084 64880 95112
rect 43496 95072 43502 95084
rect 64874 95072 64880 95084
rect 64932 95072 64938 95124
rect 82630 95072 82636 95124
rect 82688 95112 82694 95124
rect 99466 95112 99472 95124
rect 82688 95084 99472 95112
rect 82688 95072 82694 95084
rect 99466 95072 99472 95084
rect 99524 95072 99530 95124
rect 110598 95072 110604 95124
rect 110656 95112 110662 95124
rect 122098 95112 122104 95124
rect 110656 95084 122104 95112
rect 110656 95072 110662 95084
rect 122098 95072 122104 95084
rect 122156 95072 122162 95124
rect 128630 95072 128636 95124
rect 128688 95112 128694 95124
rect 149698 95112 149704 95124
rect 128688 95084 149704 95112
rect 128688 95072 128694 95084
rect 149698 95072 149704 95084
rect 149756 95072 149762 95124
rect 166626 95072 166632 95124
rect 166684 95112 166690 95124
rect 183646 95112 183652 95124
rect 166684 95084 183652 95112
rect 166684 95072 166690 95084
rect 183646 95072 183652 95084
rect 183704 95072 183710 95124
rect 194594 95072 194600 95124
rect 194652 95112 194658 95124
rect 211246 95112 211252 95124
rect 194652 95084 211252 95112
rect 194652 95072 194658 95084
rect 211246 95072 211252 95084
rect 211304 95072 211310 95124
rect 222930 95072 222936 95124
rect 222988 95112 222994 95124
rect 233970 95112 233976 95124
rect 222988 95084 233976 95112
rect 222988 95072 222994 95084
rect 233970 95072 233976 95084
rect 234028 95072 234034 95124
rect 240318 95072 240324 95124
rect 240376 95112 240382 95124
rect 262858 95112 262864 95124
rect 240376 95084 262864 95112
rect 240376 95072 240382 95084
rect 262858 95072 262864 95084
rect 262916 95072 262922 95124
rect 278590 95072 278596 95124
rect 278648 95112 278654 95124
rect 290458 95112 290464 95124
rect 278648 95084 290464 95112
rect 278648 95072 278654 95084
rect 290458 95072 290464 95084
rect 290516 95072 290522 95124
rect 324314 95072 324320 95124
rect 324372 95112 324378 95124
rect 345658 95112 345664 95124
rect 324372 95084 345664 95112
rect 324372 95072 324378 95084
rect 345658 95072 345664 95084
rect 345716 95072 345722 95124
rect 352650 95072 352656 95124
rect 352708 95112 352714 95124
rect 378870 95112 378876 95124
rect 352708 95084 378876 95112
rect 352708 95072 352714 95084
rect 378870 95072 378876 95084
rect 378928 95072 378934 95124
rect 390646 95072 390652 95124
rect 390704 95112 390710 95124
rect 402238 95112 402244 95124
rect 390704 95084 402244 95112
rect 390704 95072 390710 95084
rect 402238 95072 402244 95084
rect 402296 95072 402302 95124
rect 418614 95072 418620 95124
rect 418672 95112 418678 95124
rect 429838 95112 429844 95124
rect 418672 95084 429844 95112
rect 418672 95072 418678 95084
rect 429838 95072 429844 95084
rect 429896 95072 429902 95124
rect 436646 95072 436652 95124
rect 436704 95112 436710 95124
rect 457438 95112 457444 95124
rect 436704 95084 457444 95112
rect 436704 95072 436710 95084
rect 457438 95072 457444 95084
rect 457496 95072 457502 95124
rect 474642 95072 474648 95124
rect 474700 95112 474706 95124
rect 486418 95112 486424 95124
rect 474700 95084 486424 95112
rect 474700 95072 474706 95084
rect 486418 95072 486424 95084
rect 486476 95072 486482 95124
rect 502610 95072 502616 95124
rect 502668 95112 502674 95124
rect 514018 95112 514024 95124
rect 502668 95084 514024 95112
rect 502668 95072 502674 95084
rect 514018 95072 514024 95084
rect 514076 95072 514082 95124
rect 520642 95072 520648 95124
rect 520700 95112 520706 95124
rect 541618 95112 541624 95124
rect 520700 95084 541624 95112
rect 520700 95072 520706 95084
rect 541618 95072 541624 95084
rect 541676 95072 541682 95124
rect 54938 95004 54944 95056
rect 54996 95044 55002 95056
rect 72142 95044 72148 95056
rect 54996 95016 72148 95044
rect 54996 95004 55002 95016
rect 72142 95004 72148 95016
rect 72200 95004 72206 95056
rect 138934 95004 138940 95056
rect 138992 95044 138998 95056
rect 149790 95044 149796 95056
rect 138992 95016 149796 95044
rect 138992 95004 138998 95016
rect 149790 95004 149796 95016
rect 149848 95004 149854 95056
rect 250622 95004 250628 95056
rect 250680 95044 250686 95056
rect 264238 95044 264244 95056
rect 250680 95016 264244 95044
rect 250680 95004 250686 95016
rect 264238 95004 264244 95016
rect 264296 95004 264302 95056
rect 334618 95004 334624 95056
rect 334676 95044 334682 95056
rect 348418 95044 348424 95056
rect 334676 95016 348424 95044
rect 334676 95004 334682 95016
rect 348418 95004 348424 95016
rect 348476 95004 348482 95056
rect 362862 95004 362868 95056
rect 362920 95044 362926 95056
rect 379606 95044 379612 95056
rect 362920 95016 379612 95044
rect 362920 95004 362926 95016
rect 379606 95004 379612 95016
rect 379664 95004 379670 95056
rect 446950 95004 446956 95056
rect 447008 95044 447014 95056
rect 458818 95044 458824 95056
rect 447008 95016 458824 95044
rect 447008 95004 447014 95016
rect 458818 95004 458824 95016
rect 458876 95004 458882 95056
rect 530946 95004 530952 95056
rect 531004 95044 531010 95056
rect 547138 95044 547144 95056
rect 531004 95016 547144 95044
rect 531004 95004 531010 95016
rect 547138 95004 547144 95016
rect 547196 95004 547202 95056
rect 44634 94936 44640 94988
rect 44692 94976 44698 94988
rect 65886 94976 65892 94988
rect 44692 94948 65892 94976
rect 44692 94936 44698 94948
rect 65886 94936 65892 94948
rect 65944 94936 65950 94988
rect 558638 94460 558644 94512
rect 558696 94500 558702 94512
rect 568758 94500 568764 94512
rect 558696 94472 568764 94500
rect 558696 94460 558702 94472
rect 568758 94460 568764 94472
rect 568816 94460 568822 94512
rect 548334 93100 548340 93152
rect 548392 93140 548398 93152
rect 569034 93140 569040 93152
rect 548392 93112 569040 93140
rect 548392 93100 548398 93112
rect 569034 93100 569040 93112
rect 569092 93100 569098 93152
rect 100018 92692 100024 92744
rect 100076 92732 100082 92744
rect 120810 92732 120816 92744
rect 100076 92704 120816 92732
rect 100076 92692 100082 92704
rect 120810 92692 120816 92704
rect 120868 92692 120874 92744
rect 184014 92692 184020 92744
rect 184072 92732 184078 92744
rect 204898 92732 204904 92744
rect 184072 92704 204904 92732
rect 184072 92692 184078 92704
rect 204898 92692 204904 92704
rect 204956 92692 204962 92744
rect 268010 92692 268016 92744
rect 268068 92732 268074 92744
rect 289078 92732 289084 92744
rect 268068 92704 289084 92732
rect 268068 92692 268074 92704
rect 289078 92692 289084 92704
rect 289136 92692 289142 92744
rect 65886 92624 65892 92676
rect 65944 92664 65950 92676
rect 81986 92664 81992 92676
rect 65944 92636 81992 92664
rect 65944 92624 65950 92636
rect 81986 92624 81992 92636
rect 82044 92624 82050 92676
rect 92750 92624 92756 92676
rect 92808 92664 92814 92676
rect 110322 92664 110328 92676
rect 92808 92636 110328 92664
rect 92808 92624 92814 92636
rect 110322 92624 110328 92636
rect 110380 92624 110386 92676
rect 149790 92624 149796 92676
rect 149848 92664 149854 92676
rect 165982 92664 165988 92676
rect 149848 92636 165988 92664
rect 149848 92624 149854 92636
rect 165982 92624 165988 92636
rect 166040 92624 166046 92676
rect 176746 92624 176752 92676
rect 176804 92664 176810 92676
rect 194318 92664 194324 92676
rect 176804 92636 194324 92664
rect 176804 92624 176810 92636
rect 194318 92624 194324 92636
rect 194376 92624 194382 92676
rect 261570 92624 261576 92676
rect 261628 92664 261634 92676
rect 278314 92664 278320 92676
rect 261628 92636 278320 92664
rect 261628 92624 261634 92636
rect 278314 92624 278320 92636
rect 278372 92624 278378 92676
rect 345750 92624 345756 92676
rect 345808 92664 345814 92676
rect 362310 92664 362316 92676
rect 345808 92636 362316 92664
rect 345808 92624 345814 92636
rect 362310 92624 362316 92636
rect 362368 92624 362374 92676
rect 372798 92624 372804 92676
rect 372856 92664 372862 92676
rect 390002 92664 390008 92676
rect 372856 92636 390008 92664
rect 372856 92624 372862 92636
rect 390002 92624 390008 92636
rect 390060 92624 390066 92676
rect 458818 92624 458824 92676
rect 458876 92664 458882 92676
rect 473998 92664 474004 92676
rect 458876 92636 474004 92664
rect 458876 92624 458882 92636
rect 473998 92624 474004 92636
rect 474056 92624 474062 92676
rect 36906 92556 36912 92608
rect 36964 92596 36970 92608
rect 54294 92596 54300 92608
rect 36964 92568 54300 92596
rect 36964 92556 36970 92568
rect 54294 92556 54300 92568
rect 54352 92556 54358 92608
rect 72326 92556 72332 92608
rect 72384 92596 72390 92608
rect 93118 92596 93124 92608
rect 72384 92568 93124 92596
rect 72384 92556 72390 92568
rect 93118 92556 93124 92568
rect 93176 92556 93182 92608
rect 120718 92556 120724 92608
rect 120776 92596 120782 92608
rect 138290 92596 138296 92608
rect 120776 92568 138296 92596
rect 120776 92556 120782 92568
rect 138290 92556 138296 92568
rect 138348 92556 138354 92608
rect 156322 92556 156328 92608
rect 156380 92596 156386 92608
rect 180058 92596 180064 92608
rect 156380 92568 180064 92596
rect 156380 92556 156386 92568
rect 180058 92556 180064 92568
rect 180116 92556 180122 92608
rect 204806 92556 204812 92608
rect 204864 92596 204870 92608
rect 222194 92596 222200 92608
rect 204864 92568 222200 92596
rect 204864 92556 204870 92568
rect 222194 92556 222200 92568
rect 222252 92556 222258 92608
rect 232774 92556 232780 92608
rect 232832 92596 232838 92608
rect 250346 92596 250352 92608
rect 232832 92568 250352 92596
rect 232832 92556 232838 92568
rect 250346 92556 250352 92568
rect 250404 92556 250410 92608
rect 288802 92556 288808 92608
rect 288860 92596 288866 92608
rect 306006 92596 306012 92608
rect 288860 92568 306012 92596
rect 288860 92556 288866 92568
rect 306006 92556 306012 92568
rect 306064 92556 306070 92608
rect 316770 92556 316776 92608
rect 316828 92596 316834 92608
rect 334342 92596 334348 92608
rect 316828 92568 334348 92596
rect 316828 92556 316834 92568
rect 334342 92556 334348 92568
rect 334400 92556 334406 92608
rect 352006 92556 352012 92608
rect 352064 92596 352070 92608
rect 376018 92596 376024 92608
rect 352064 92568 376024 92596
rect 352064 92556 352070 92568
rect 376018 92556 376024 92568
rect 376076 92556 376082 92608
rect 380342 92556 380348 92608
rect 380400 92596 380406 92608
rect 400858 92596 400864 92608
rect 380400 92568 400864 92596
rect 380400 92556 380406 92568
rect 400858 92556 400864 92568
rect 400916 92556 400922 92608
rect 435358 92556 435364 92608
rect 435416 92596 435422 92608
rect 446306 92596 446312 92608
rect 435416 92568 446312 92596
rect 435416 92556 435422 92568
rect 446306 92556 446312 92568
rect 446364 92556 446370 92608
rect 464338 92556 464344 92608
rect 464396 92596 464402 92608
rect 485038 92596 485044 92608
rect 464396 92568 485044 92596
rect 464396 92556 464402 92568
rect 485038 92556 485044 92568
rect 485096 92556 485102 92608
rect 512914 92556 512920 92608
rect 512972 92596 512978 92608
rect 530302 92596 530308 92608
rect 512972 92568 530308 92596
rect 512972 92556 512978 92568
rect 530302 92556 530308 92568
rect 530360 92556 530366 92608
rect 541710 92556 541716 92608
rect 541768 92596 541774 92608
rect 557994 92596 558000 92608
rect 541768 92568 558000 92596
rect 541768 92556 541774 92568
rect 557994 92556 558000 92568
rect 558052 92556 558058 92608
rect 15194 92488 15200 92540
rect 15252 92528 15258 92540
rect 26326 92528 26332 92540
rect 15252 92500 26332 92528
rect 15252 92488 15258 92500
rect 26326 92488 26332 92500
rect 26384 92488 26390 92540
rect 38102 92488 38108 92540
rect 38160 92528 38166 92540
rect 64598 92528 64604 92540
rect 38160 92500 64604 92528
rect 38160 92488 38166 92500
rect 64598 92488 64604 92500
rect 64656 92488 64662 92540
rect 66898 92488 66904 92540
rect 66956 92528 66962 92540
rect 92474 92528 92480 92540
rect 66956 92500 92480 92528
rect 66956 92488 66962 92500
rect 92474 92488 92480 92500
rect 92532 92488 92538 92540
rect 94498 92488 94504 92540
rect 94556 92528 94562 92540
rect 120626 92528 120632 92540
rect 94556 92500 120632 92528
rect 94556 92488 94562 92500
rect 120626 92488 120632 92500
rect 120684 92488 120690 92540
rect 122098 92488 122104 92540
rect 122156 92528 122162 92540
rect 148594 92528 148600 92540
rect 122156 92500 148600 92528
rect 122156 92488 122162 92500
rect 148594 92488 148600 92500
rect 148652 92488 148658 92540
rect 149698 92488 149704 92540
rect 149756 92528 149762 92540
rect 176654 92528 176660 92540
rect 149756 92500 176660 92528
rect 149756 92488 149762 92500
rect 176654 92488 176660 92500
rect 176712 92488 176718 92540
rect 178678 92488 178684 92540
rect 178736 92528 178742 92540
rect 204622 92528 204628 92540
rect 178736 92500 204628 92528
rect 178736 92488 178742 92500
rect 204622 92488 204628 92500
rect 204680 92488 204686 92540
rect 206278 92488 206284 92540
rect 206336 92528 206342 92540
rect 232314 92528 232320 92540
rect 206336 92500 232320 92528
rect 206336 92488 206342 92500
rect 232314 92488 232320 92500
rect 232372 92488 232378 92540
rect 233970 92488 233976 92540
rect 234028 92528 234034 92540
rect 260650 92528 260656 92540
rect 234028 92500 260656 92528
rect 234028 92488 234034 92500
rect 260650 92488 260656 92500
rect 260708 92488 260714 92540
rect 261478 92488 261484 92540
rect 261536 92528 261542 92540
rect 288618 92528 288624 92540
rect 261536 92500 288624 92528
rect 261536 92488 261542 92500
rect 288618 92488 288624 92500
rect 288676 92488 288682 92540
rect 290458 92488 290464 92540
rect 290516 92528 290522 92540
rect 316310 92528 316316 92540
rect 290516 92500 316316 92528
rect 290516 92488 290522 92500
rect 316310 92488 316316 92500
rect 316368 92488 316374 92540
rect 316862 92488 316868 92540
rect 316920 92528 316926 92540
rect 344646 92528 344652 92540
rect 316920 92500 344652 92528
rect 316920 92488 316926 92500
rect 344646 92488 344652 92500
rect 344704 92488 344710 92540
rect 345658 92488 345664 92540
rect 345716 92528 345722 92540
rect 372614 92528 372620 92540
rect 345716 92500 372620 92528
rect 345716 92488 345722 92500
rect 372614 92488 372620 92500
rect 372672 92488 372678 92540
rect 374638 92488 374644 92540
rect 374696 92528 374702 92540
rect 400306 92528 400312 92540
rect 374696 92500 400312 92528
rect 374696 92488 374702 92500
rect 400306 92488 400312 92500
rect 400364 92488 400370 92540
rect 400766 92488 400772 92540
rect 400824 92528 400830 92540
rect 418338 92528 418344 92540
rect 400824 92500 418344 92528
rect 400824 92488 400830 92500
rect 418338 92488 418344 92500
rect 418396 92488 418402 92540
rect 429838 92488 429844 92540
rect 429896 92528 429902 92540
rect 456610 92528 456616 92540
rect 429896 92500 456616 92528
rect 429896 92488 429902 92500
rect 456610 92488 456616 92500
rect 456668 92488 456674 92540
rect 457438 92488 457444 92540
rect 457496 92528 457502 92540
rect 484394 92528 484400 92540
rect 457496 92500 484400 92528
rect 457496 92488 457502 92500
rect 484394 92488 484400 92500
rect 484452 92488 484458 92540
rect 484762 92488 484768 92540
rect 484820 92528 484826 92540
rect 502334 92528 502340 92540
rect 484820 92500 502340 92528
rect 484820 92488 484826 92500
rect 502334 92488 502340 92500
rect 502392 92488 502398 92540
rect 514018 92488 514024 92540
rect 514076 92528 514082 92540
rect 540606 92528 540612 92540
rect 514076 92500 540612 92528
rect 514076 92488 514082 92500
rect 540606 92488 540612 92500
rect 540664 92488 540670 92540
rect 541618 92488 541624 92540
rect 541676 92528 541682 92540
rect 568574 92528 568580 92540
rect 541676 92500 568580 92528
rect 541676 92488 541682 92500
rect 568574 92488 568580 92500
rect 568632 92488 568638 92540
rect 209682 89700 209688 89752
rect 209740 89740 209746 89752
rect 262214 89740 262220 89752
rect 209740 89712 262220 89740
rect 209740 89700 209746 89712
rect 262214 89700 262220 89712
rect 262272 89700 262278 89752
rect 405642 89700 405648 89752
rect 405700 89740 405706 89752
rect 458174 89740 458180 89752
rect 405700 89712 458180 89740
rect 405700 89700 405706 89712
rect 458174 89700 458180 89712
rect 458232 89700 458238 89752
rect 489822 89700 489828 89752
rect 489880 89740 489886 89752
rect 542354 89740 542360 89752
rect 489880 89712 542360 89740
rect 489880 89700 489886 89712
rect 542354 89700 542360 89712
rect 542412 89700 542418 89752
rect 434714 87184 434720 87236
rect 434772 87224 434778 87236
rect 435726 87224 435732 87236
rect 434772 87196 435732 87224
rect 434772 87184 434778 87196
rect 435726 87184 435732 87196
rect 435784 87184 435790 87236
rect 36814 85008 36820 85060
rect 36872 85048 36878 85060
rect 36998 85048 37004 85060
rect 36872 85020 37004 85048
rect 36872 85008 36878 85020
rect 36998 85008 37004 85020
rect 37056 85008 37062 85060
rect 512822 85008 512828 85060
rect 512880 85048 512886 85060
rect 513006 85048 513012 85060
rect 512880 85020 513012 85048
rect 512880 85008 512886 85020
rect 513006 85008 513012 85020
rect 513064 85008 513070 85060
rect 3326 84600 3332 84652
rect 3384 84640 3390 84652
rect 9030 84640 9036 84652
rect 3384 84612 9036 84640
rect 3384 84600 3390 84612
rect 9030 84600 9036 84612
rect 9088 84600 9094 84652
rect 36814 77256 36820 77308
rect 36872 77296 36878 77308
rect 36998 77296 37004 77308
rect 36872 77268 37004 77296
rect 36872 77256 36878 77268
rect 36998 77256 37004 77268
rect 37056 77256 37062 77308
rect 512822 77256 512828 77308
rect 512880 77296 512886 77308
rect 513006 77296 513012 77308
rect 512880 77268 513012 77296
rect 512880 77256 512886 77268
rect 513006 77256 513012 77268
rect 513064 77256 513070 77308
rect 93118 73788 93124 73840
rect 93176 73828 93182 73840
rect 99742 73828 99748 73840
rect 93176 73800 99748 73828
rect 93176 73788 93182 73800
rect 99742 73788 99748 73800
rect 99800 73788 99806 73840
rect 120810 73788 120816 73840
rect 120868 73828 120874 73840
rect 127710 73828 127716 73840
rect 120868 73800 127716 73828
rect 120868 73788 120874 73800
rect 127710 73788 127716 73800
rect 127768 73788 127774 73840
rect 400858 73788 400864 73840
rect 400916 73828 400922 73840
rect 407758 73828 407764 73840
rect 400916 73800 407764 73828
rect 400916 73788 400922 73800
rect 407758 73788 407764 73800
rect 407816 73788 407822 73840
rect 485038 73652 485044 73704
rect 485096 73692 485102 73704
rect 491662 73692 491668 73704
rect 485096 73664 491668 73692
rect 485096 73652 485102 73664
rect 491662 73652 491668 73664
rect 491720 73652 491726 73704
rect 204898 73448 204904 73500
rect 204956 73488 204962 73500
rect 211706 73488 211712 73500
rect 204956 73460 211712 73488
rect 204956 73448 204962 73460
rect 211706 73448 211712 73460
rect 211764 73448 211770 73500
rect 289078 73176 289084 73228
rect 289136 73216 289142 73228
rect 295702 73216 295708 73228
rect 289136 73188 295708 73216
rect 289136 73176 289142 73188
rect 295702 73176 295708 73188
rect 295760 73176 295766 73228
rect 64874 72564 64880 72616
rect 64932 72604 64938 72616
rect 65886 72604 65892 72616
rect 64932 72576 65892 72604
rect 64932 72564 64938 72576
rect 65886 72564 65892 72576
rect 65944 72564 65950 72616
rect 261018 72292 261024 72344
rect 261076 72332 261082 72344
rect 261570 72332 261576 72344
rect 261076 72304 261576 72332
rect 261076 72292 261082 72304
rect 261570 72292 261576 72304
rect 261628 72292 261634 72344
rect 148962 71680 148968 71732
rect 149020 71720 149026 71732
rect 149790 71720 149796 71732
rect 149020 71692 149796 71720
rect 149020 71680 149026 71692
rect 149790 71680 149796 71692
rect 149848 71680 149854 71732
rect 344922 71680 344928 71732
rect 344980 71720 344986 71732
rect 345750 71720 345756 71732
rect 344980 71692 345756 71720
rect 344980 71680 344986 71692
rect 345750 71680 345756 71692
rect 345808 71680 345814 71732
rect 540882 71680 540888 71732
rect 540940 71720 540946 71732
rect 541710 71720 541716 71732
rect 540940 71692 541716 71720
rect 540940 71680 540946 71692
rect 541710 71680 541716 71692
rect 541768 71680 541774 71732
rect 547874 70660 547880 70712
rect 547932 70700 547938 70712
rect 548150 70700 548156 70712
rect 547932 70672 548156 70700
rect 547932 70660 547938 70672
rect 548150 70660 548156 70672
rect 548208 70660 548214 70712
rect 15194 69640 15200 69692
rect 15252 69680 15258 69692
rect 16022 69680 16028 69692
rect 15252 69652 16028 69680
rect 15252 69640 15258 69652
rect 16022 69640 16028 69652
rect 16080 69640 16086 69692
rect 15378 68960 15384 69012
rect 15436 69000 15442 69012
rect 43990 69000 43996 69012
rect 15436 68972 43996 69000
rect 15436 68960 15442 68972
rect 43990 68960 43996 68972
rect 44048 68960 44054 69012
rect 82630 68960 82636 69012
rect 82688 69000 82694 69012
rect 94498 69000 94504 69012
rect 82688 68972 94504 69000
rect 82688 68960 82694 68972
rect 94498 68960 94504 68972
rect 94556 68960 94562 69012
rect 110322 68960 110328 69012
rect 110380 69000 110386 69012
rect 122098 69000 122104 69012
rect 110380 68972 122104 69000
rect 110380 68960 110386 68972
rect 122098 68960 122104 68972
rect 122156 68960 122162 69012
rect 166626 68960 166632 69012
rect 166684 69000 166690 69012
rect 178678 69000 178684 69012
rect 166684 68972 178684 69000
rect 166684 68960 166690 68972
rect 178678 68960 178684 68972
rect 178736 68960 178742 69012
rect 180058 68960 180064 69012
rect 180116 69000 180122 69012
rect 184014 69000 184020 69012
rect 180116 68972 184020 69000
rect 180116 68960 180122 68972
rect 184014 68960 184020 68972
rect 184072 68960 184078 69012
rect 194318 68960 194324 69012
rect 194376 69000 194382 69012
rect 206278 69000 206284 69012
rect 194376 68972 206284 69000
rect 194376 68960 194382 68972
rect 206278 68960 206284 68972
rect 206336 68960 206342 69012
rect 211246 68960 211252 69012
rect 211304 69000 211310 69012
rect 240042 69000 240048 69012
rect 211304 68972 240048 69000
rect 211304 68960 211310 68972
rect 240042 68960 240048 68972
rect 240100 68960 240106 69012
rect 278314 68960 278320 69012
rect 278372 69000 278378 69012
rect 290458 69000 290464 69012
rect 278372 68972 290464 69000
rect 278372 68960 278378 68972
rect 290458 68960 290464 68972
rect 290516 68960 290522 69012
rect 295426 68960 295432 69012
rect 295484 69000 295490 69012
rect 324038 69000 324044 69012
rect 295484 68972 324044 69000
rect 295484 68960 295490 68972
rect 324038 68960 324044 68972
rect 324096 68960 324102 69012
rect 362310 68960 362316 69012
rect 362368 69000 362374 69012
rect 374638 69000 374644 69012
rect 362368 68972 374644 69000
rect 362368 68960 362374 68972
rect 374638 68960 374644 68972
rect 374696 68960 374702 69012
rect 376018 68960 376024 69012
rect 376076 69000 376082 69012
rect 379698 69000 379704 69012
rect 376076 68972 379704 69000
rect 376076 68960 376082 68972
rect 379698 68960 379704 68972
rect 379756 68960 379762 69012
rect 428642 68960 428648 69012
rect 428700 69000 428706 69012
rect 435358 69000 435364 69012
rect 428700 68972 435364 69000
rect 428700 68960 428706 68972
rect 435358 68960 435364 68972
rect 435416 68960 435422 69012
rect 456610 68960 456616 69012
rect 456668 69000 456674 69012
rect 458818 69000 458824 69012
rect 456668 68972 458824 69000
rect 456668 68960 456674 68972
rect 458818 68960 458824 68972
rect 458876 68960 458882 69012
rect 474642 68960 474648 69012
rect 474700 69000 474706 69012
rect 512822 69000 512828 69012
rect 474700 68972 512828 69000
rect 474700 68960 474706 68972
rect 512822 68960 512828 68972
rect 512880 68960 512886 69012
rect 548150 68960 548156 69012
rect 548208 69000 548214 69012
rect 557994 69000 558000 69012
rect 548208 68972 558000 69000
rect 548208 68960 548214 68972
rect 557994 68960 558000 68972
rect 558052 68960 558058 69012
rect 26326 68892 26332 68944
rect 26384 68932 26390 68944
rect 38102 68932 38108 68944
rect 26384 68904 38108 68932
rect 26384 68892 26390 68904
rect 38102 68892 38108 68904
rect 38160 68892 38166 68944
rect 54294 68892 54300 68944
rect 54352 68932 54358 68944
rect 66898 68932 66904 68944
rect 54352 68904 66904 68932
rect 54352 68892 54358 68904
rect 66898 68892 66904 68904
rect 66956 68892 66962 68944
rect 138290 68892 138296 68944
rect 138348 68932 138354 68944
rect 149698 68932 149704 68944
rect 138348 68904 149704 68932
rect 138348 68892 138354 68904
rect 149698 68892 149704 68904
rect 149756 68892 149762 68944
rect 222654 68892 222660 68944
rect 222712 68932 222718 68944
rect 233970 68932 233976 68944
rect 222712 68904 233976 68932
rect 222712 68892 222718 68904
rect 233970 68892 233976 68904
rect 234028 68892 234034 68944
rect 250346 68892 250352 68944
rect 250404 68932 250410 68944
rect 261478 68932 261484 68944
rect 250404 68904 261484 68932
rect 250404 68892 250410 68904
rect 261478 68892 261484 68904
rect 261536 68892 261542 68944
rect 306282 68892 306288 68944
rect 306340 68932 306346 68944
rect 316862 68932 316868 68944
rect 306340 68904 316868 68932
rect 306340 68892 306346 68904
rect 316862 68892 316868 68904
rect 316920 68892 316926 68944
rect 334342 68892 334348 68944
rect 334400 68932 334406 68944
rect 345658 68932 345664 68944
rect 334400 68904 345664 68932
rect 334400 68892 334406 68904
rect 345658 68892 345664 68904
rect 345716 68892 345722 68944
rect 407206 68892 407212 68944
rect 407264 68932 407270 68944
rect 436002 68932 436008 68944
rect 407264 68904 436008 68932
rect 407264 68892 407270 68904
rect 436002 68892 436008 68904
rect 436060 68892 436066 68944
rect 446306 68892 446312 68944
rect 446364 68932 446370 68944
rect 457438 68932 457444 68944
rect 446364 68904 457444 68932
rect 446364 68892 446370 68904
rect 457438 68892 457444 68904
rect 457496 68892 457502 68944
rect 491386 68892 491392 68944
rect 491444 68932 491450 68944
rect 519998 68932 520004 68944
rect 491444 68904 520004 68932
rect 491444 68892 491450 68904
rect 519998 68892 520004 68904
rect 520056 68892 520062 68944
rect 530302 68892 530308 68944
rect 530360 68932 530366 68944
rect 541618 68932 541624 68944
rect 530360 68904 541624 68932
rect 530360 68892 530366 68904
rect 541618 68892 541624 68904
rect 541676 68892 541682 68944
rect 42886 68824 42892 68876
rect 42944 68864 42950 68876
rect 71774 68864 71780 68876
rect 42944 68836 71780 68864
rect 42944 68824 42950 68836
rect 71774 68824 71780 68836
rect 71832 68824 71838 68876
rect 127066 68824 127072 68876
rect 127124 68864 127130 68876
rect 156046 68864 156052 68876
rect 127124 68836 156052 68864
rect 127124 68824 127130 68836
rect 156046 68824 156052 68836
rect 156104 68824 156110 68876
rect 238846 68824 238852 68876
rect 238904 68864 238910 68876
rect 268010 68864 268016 68876
rect 238904 68836 268016 68864
rect 238904 68824 238910 68836
rect 268010 68824 268016 68836
rect 268068 68824 268074 68876
rect 323026 68824 323032 68876
rect 323084 68864 323090 68876
rect 352006 68864 352012 68876
rect 323084 68836 352012 68864
rect 323084 68824 323090 68836
rect 352006 68824 352012 68836
rect 352064 68824 352070 68876
rect 418338 68824 418344 68876
rect 418396 68864 418402 68876
rect 429838 68864 429844 68876
rect 418396 68836 429844 68864
rect 418396 68824 418402 68836
rect 429838 68824 429844 68836
rect 429896 68824 429902 68876
rect 434714 68824 434720 68876
rect 434772 68864 434778 68876
rect 463694 68864 463700 68876
rect 434772 68836 463700 68864
rect 434772 68824 434778 68836
rect 463694 68824 463700 68836
rect 463752 68824 463758 68876
rect 502334 68824 502340 68876
rect 502392 68864 502398 68876
rect 514018 68864 514024 68876
rect 502392 68836 514024 68864
rect 502392 68824 502398 68836
rect 514018 68824 514024 68836
rect 514076 68824 514082 68876
rect 518894 68824 518900 68876
rect 518952 68864 518958 68876
rect 547874 68864 547880 68876
rect 518952 68836 547880 68864
rect 518952 68824 518958 68836
rect 547874 68824 547880 68836
rect 547932 68824 547938 68876
rect 390462 68756 390468 68808
rect 390520 68796 390526 68808
rect 428734 68796 428740 68808
rect 390520 68768 428740 68796
rect 390520 68756 390526 68768
rect 428734 68756 428740 68768
rect 428792 68756 428798 68808
rect 26602 66852 26608 66904
rect 26660 66892 26666 66904
rect 36814 66892 36820 66904
rect 26660 66864 36820 66892
rect 26660 66852 26666 66864
rect 36814 66852 36820 66864
rect 36872 66852 36878 66904
rect 15378 66376 15384 66428
rect 15436 66416 15442 66428
rect 54294 66416 54300 66428
rect 15436 66388 54300 66416
rect 15436 66376 15442 66388
rect 54294 66376 54300 66388
rect 54352 66376 54358 66428
rect 211246 66376 211252 66428
rect 211304 66416 211310 66428
rect 250622 66416 250628 66428
rect 211304 66388 250628 66416
rect 211304 66376 211310 66388
rect 250622 66376 250628 66388
rect 250680 66376 250686 66428
rect 345658 66376 345664 66428
rect 345716 66416 345722 66428
rect 362310 66416 362316 66428
rect 345716 66388 362316 66416
rect 345716 66376 345722 66388
rect 362310 66376 362316 66388
rect 362368 66376 362374 66428
rect 374638 66376 374644 66428
rect 374696 66416 374702 66428
rect 380342 66416 380348 66428
rect 374696 66388 380348 66416
rect 374696 66376 374702 66388
rect 380342 66376 380348 66388
rect 380400 66376 380406 66428
rect 491386 66376 491392 66428
rect 491444 66416 491450 66428
rect 491444 66388 499574 66416
rect 491444 66376 491450 66388
rect 65886 66308 65892 66360
rect 65944 66348 65950 66360
rect 82630 66348 82636 66360
rect 65944 66320 82636 66348
rect 65944 66308 65950 66320
rect 82630 66308 82636 66320
rect 82688 66308 82694 66360
rect 99466 66308 99472 66360
rect 99524 66348 99530 66360
rect 138290 66348 138296 66360
rect 99524 66320 138296 66348
rect 99524 66308 99530 66320
rect 138290 66308 138296 66320
rect 138348 66308 138354 66360
rect 149698 66308 149704 66360
rect 149756 66348 149762 66360
rect 156322 66348 156328 66360
rect 149756 66320 156328 66348
rect 149756 66308 149762 66320
rect 156322 66308 156328 66320
rect 156380 66308 156386 66360
rect 183646 66308 183652 66360
rect 183704 66348 183710 66360
rect 222378 66348 222384 66360
rect 183704 66320 222384 66348
rect 183704 66308 183710 66320
rect 222378 66308 222384 66320
rect 222436 66308 222442 66360
rect 267826 66308 267832 66360
rect 267884 66348 267890 66360
rect 306374 66348 306380 66360
rect 267884 66320 306380 66348
rect 267884 66308 267890 66320
rect 306374 66308 306380 66320
rect 306432 66308 306438 66360
rect 318058 66308 318064 66360
rect 318116 66348 318122 66360
rect 324314 66348 324320 66360
rect 318116 66320 324320 66348
rect 318116 66308 318122 66320
rect 324314 66308 324320 66320
rect 324372 66308 324378 66360
rect 373258 66308 373264 66360
rect 373316 66348 373322 66360
rect 390646 66348 390652 66360
rect 373316 66320 390652 66348
rect 373316 66308 373322 66320
rect 390646 66308 390652 66320
rect 390704 66308 390710 66360
rect 407114 66308 407120 66360
rect 407172 66348 407178 66360
rect 446306 66348 446312 66360
rect 407172 66320 446312 66348
rect 407172 66308 407178 66320
rect 446306 66308 446312 66320
rect 446364 66308 446370 66360
rect 457438 66308 457444 66360
rect 457496 66348 457502 66360
rect 474642 66348 474648 66360
rect 457496 66320 474648 66348
rect 457496 66308 457502 66320
rect 474642 66308 474648 66320
rect 474700 66308 474706 66360
rect 486418 66308 486424 66360
rect 486476 66348 486482 66360
rect 492306 66348 492312 66360
rect 486476 66320 492312 66348
rect 486476 66308 486482 66320
rect 492306 66308 492312 66320
rect 492364 66308 492370 66360
rect 499546 66348 499574 66388
rect 530302 66348 530308 66360
rect 499546 66320 530308 66348
rect 530302 66308 530308 66320
rect 530360 66308 530366 66360
rect 36906 66240 36912 66292
rect 36964 66280 36970 66292
rect 43438 66280 43444 66292
rect 36964 66252 43444 66280
rect 36964 66240 36970 66252
rect 43438 66240 43444 66252
rect 43496 66240 43502 66292
rect 71866 66240 71872 66292
rect 71924 66280 71930 66292
rect 110598 66280 110604 66292
rect 71924 66252 110604 66280
rect 71924 66240 71930 66252
rect 110598 66240 110604 66252
rect 110656 66240 110662 66292
rect 122098 66240 122104 66292
rect 122156 66280 122162 66292
rect 128354 66280 128360 66292
rect 122156 66252 128360 66280
rect 122156 66240 122162 66252
rect 128354 66240 128360 66252
rect 128412 66240 128418 66292
rect 149882 66240 149888 66292
rect 149940 66280 149946 66292
rect 166626 66280 166632 66292
rect 149940 66252 166632 66280
rect 149940 66240 149946 66252
rect 166626 66240 166632 66252
rect 166684 66240 166690 66292
rect 182818 66240 182824 66292
rect 182876 66280 182882 66292
rect 194594 66280 194600 66292
rect 182876 66252 194600 66280
rect 182876 66240 182882 66252
rect 194594 66240 194600 66252
rect 194652 66240 194658 66292
rect 206278 66240 206284 66292
rect 206336 66280 206342 66292
rect 211982 66280 211988 66292
rect 206336 66252 211988 66280
rect 206336 66240 206342 66252
rect 211982 66240 211988 66252
rect 212040 66240 212046 66292
rect 234062 66240 234068 66292
rect 234120 66280 234126 66292
rect 240318 66280 240324 66292
rect 234120 66252 240324 66280
rect 234120 66240 234126 66252
rect 240318 66240 240324 66252
rect 240376 66240 240382 66292
rect 261478 66240 261484 66292
rect 261536 66280 261542 66292
rect 278590 66280 278596 66292
rect 261536 66252 278596 66280
rect 261536 66240 261542 66252
rect 278590 66240 278596 66252
rect 278648 66240 278654 66292
rect 295426 66240 295432 66292
rect 295484 66280 295490 66292
rect 334618 66280 334624 66292
rect 295484 66252 334624 66280
rect 295484 66240 295490 66252
rect 334618 66240 334624 66252
rect 334676 66240 334682 66292
rect 379606 66240 379612 66292
rect 379664 66280 379670 66292
rect 418614 66280 418620 66292
rect 379664 66252 418620 66280
rect 379664 66240 379670 66252
rect 418614 66240 418620 66252
rect 418672 66240 418678 66292
rect 458818 66240 458824 66292
rect 458876 66280 458882 66292
rect 464338 66280 464344 66292
rect 458876 66252 464344 66280
rect 458876 66240 458882 66252
rect 464338 66240 464344 66252
rect 464396 66240 464402 66292
rect 502610 66280 502616 66292
rect 464448 66252 502616 66280
rect 463786 66172 463792 66224
rect 463844 66212 463850 66224
rect 464448 66212 464476 66252
rect 502610 66240 502616 66252
rect 502668 66240 502674 66292
rect 514018 66240 514024 66292
rect 514076 66280 514082 66292
rect 520274 66280 520280 66292
rect 514076 66252 520280 66280
rect 514076 66240 514082 66252
rect 520274 66240 520280 66252
rect 520332 66240 520338 66292
rect 541618 66240 541624 66292
rect 541676 66280 541682 66292
rect 558638 66280 558644 66292
rect 541676 66252 558644 66280
rect 541676 66240 541682 66252
rect 558638 66240 558644 66252
rect 558696 66240 558702 66292
rect 463844 66184 464476 66212
rect 463844 66172 463850 66184
rect 348418 63520 348424 63572
rect 348476 63560 348482 63572
rect 352006 63560 352012 63572
rect 348476 63532 352012 63560
rect 348476 63520 348482 63532
rect 352006 63520 352012 63532
rect 352064 63520 352070 63572
rect 205082 63384 205088 63436
rect 205140 63384 205146 63436
rect 40678 63248 40684 63300
rect 40736 63288 40742 63300
rect 43990 63288 43996 63300
rect 40736 63260 43996 63288
rect 40736 63248 40742 63260
rect 43990 63248 43996 63260
rect 44048 63248 44054 63300
rect 205100 63232 205128 63384
rect 345014 63248 345020 63300
rect 345072 63288 345078 63300
rect 347038 63288 347044 63300
rect 345072 63260 347044 63288
rect 345072 63248 345078 63260
rect 347038 63248 347044 63260
rect 347096 63248 347102 63300
rect 429102 63248 429108 63300
rect 429160 63288 429166 63300
rect 429838 63288 429844 63300
rect 429160 63260 429844 63288
rect 429160 63248 429166 63260
rect 429838 63248 429844 63260
rect 429896 63248 429902 63300
rect 205082 63180 205088 63232
rect 205140 63180 205146 63232
rect 93118 61344 93124 61396
rect 93176 61384 93182 61396
rect 99926 61384 99932 61396
rect 93176 61356 99932 61384
rect 93176 61344 93182 61356
rect 99926 61344 99932 61356
rect 99984 61344 99990 61396
rect 177298 61344 177304 61396
rect 177356 61384 177362 61396
rect 184014 61384 184020 61396
rect 177356 61356 184020 61384
rect 177356 61344 177362 61356
rect 184014 61344 184020 61356
rect 184072 61344 184078 61396
rect 65978 60732 65984 60784
rect 66036 60772 66042 60784
rect 71958 60772 71964 60784
rect 66036 60744 71964 60772
rect 66036 60732 66042 60744
rect 71958 60732 71964 60744
rect 72016 60732 72022 60784
rect 261570 60732 261576 60784
rect 261628 60772 261634 60784
rect 267918 60772 267924 60784
rect 261628 60744 267924 60772
rect 261628 60732 261634 60744
rect 267918 60732 267924 60744
rect 267976 60732 267982 60784
rect 289170 60732 289176 60784
rect 289228 60772 289234 60784
rect 295978 60772 295984 60784
rect 289228 60744 295984 60772
rect 289228 60732 289234 60744
rect 295978 60732 295984 60744
rect 296036 60732 296042 60784
rect 541710 60732 541716 60784
rect 541768 60772 541774 60784
rect 548058 60772 548064 60784
rect 541768 60744 548064 60772
rect 541768 60732 541774 60744
rect 548058 60732 548064 60744
rect 548116 60732 548122 60784
rect 149238 59236 149244 59288
rect 149296 59276 149302 59288
rect 149790 59276 149796 59288
rect 149296 59248 149796 59276
rect 149296 59236 149302 59248
rect 149790 59236 149796 59248
rect 149848 59236 149854 59288
rect 233234 59236 233240 59288
rect 233292 59276 233298 59288
rect 233970 59276 233976 59288
rect 233292 59248 233976 59276
rect 233292 59236 233298 59248
rect 233970 59236 233976 59248
rect 234028 59236 234034 59288
rect 407114 50328 407120 50380
rect 407172 50368 407178 50380
rect 407942 50368 407948 50380
rect 407172 50340 407948 50368
rect 407172 50328 407178 50340
rect 407942 50328 407948 50340
rect 408000 50328 408006 50380
rect 2958 44140 2964 44192
rect 3016 44180 3022 44192
rect 11882 44180 11888 44192
rect 3016 44152 11888 44180
rect 3016 44140 3022 44152
rect 11882 44140 11888 44152
rect 11940 44140 11946 44192
rect 489822 44072 489828 44124
rect 489880 44112 489886 44124
rect 542354 44112 542360 44124
rect 489880 44084 542360 44112
rect 489880 44072 489886 44084
rect 542354 44072 542360 44084
rect 542412 44072 542418 44124
rect 15286 41352 15292 41404
rect 15344 41392 15350 41404
rect 36906 41392 36912 41404
rect 15344 41364 36912 41392
rect 15344 41352 15350 41364
rect 36906 41352 36912 41364
rect 36964 41352 36970 41404
rect 65058 41352 65064 41404
rect 65116 41392 65122 41404
rect 92934 41392 92940 41404
rect 65116 41364 92940 41392
rect 65116 41352 65122 41364
rect 92934 41352 92940 41364
rect 92992 41352 92998 41404
rect 93026 41352 93032 41404
rect 93084 41392 93090 41404
rect 120902 41392 120908 41404
rect 93084 41364 120908 41392
rect 93084 41352 93090 41364
rect 120902 41352 120908 41364
rect 120960 41352 120966 41404
rect 121086 41352 121092 41404
rect 121144 41392 121150 41404
rect 148594 41392 148600 41404
rect 121144 41364 148600 41392
rect 121144 41352 121150 41364
rect 148594 41352 148600 41364
rect 148652 41352 148658 41404
rect 149790 41352 149796 41404
rect 149848 41392 149854 41404
rect 176930 41392 176936 41404
rect 149848 41364 176936 41392
rect 149848 41352 149854 41364
rect 176930 41352 176936 41364
rect 176988 41352 176994 41404
rect 177022 41352 177028 41404
rect 177080 41392 177086 41404
rect 204898 41392 204904 41404
rect 177080 41364 204904 41392
rect 177080 41352 177086 41364
rect 204898 41352 204904 41364
rect 204956 41352 204962 41404
rect 205174 41352 205180 41404
rect 205232 41392 205238 41404
rect 232590 41392 232596 41404
rect 205232 41364 232596 41392
rect 205232 41352 205238 41364
rect 232590 41352 232596 41364
rect 232648 41352 232654 41404
rect 233970 41352 233976 41404
rect 234028 41392 234034 41404
rect 260926 41392 260932 41404
rect 234028 41364 260932 41392
rect 234028 41352 234034 41364
rect 260926 41352 260932 41364
rect 260984 41352 260990 41404
rect 261018 41352 261024 41404
rect 261076 41392 261082 41404
rect 288894 41392 288900 41404
rect 261076 41364 288900 41392
rect 261076 41352 261082 41364
rect 288894 41352 288900 41364
rect 288952 41352 288958 41404
rect 289078 41352 289084 41404
rect 289136 41392 289142 41404
rect 316586 41392 316592 41404
rect 289136 41364 316592 41392
rect 289136 41352 289142 41364
rect 316586 41352 316592 41364
rect 316644 41352 316650 41404
rect 317046 41352 317052 41404
rect 317104 41392 317110 41404
rect 344922 41392 344928 41404
rect 317104 41364 344928 41392
rect 317104 41352 317110 41364
rect 344922 41352 344928 41364
rect 344980 41352 344986 41404
rect 347038 41352 347044 41404
rect 347096 41392 347102 41404
rect 372614 41392 372620 41404
rect 347096 41364 372620 41392
rect 347096 41352 347102 41364
rect 372614 41352 372620 41364
rect 372672 41352 372678 41404
rect 373074 41352 373080 41404
rect 373132 41392 373138 41404
rect 400950 41392 400956 41404
rect 373132 41364 400956 41392
rect 373132 41352 373138 41364
rect 400950 41352 400956 41364
rect 401008 41352 401014 41404
rect 401042 41352 401048 41404
rect 401100 41392 401106 41404
rect 428918 41392 428924 41404
rect 401100 41364 428924 41392
rect 401100 41352 401106 41364
rect 428918 41352 428924 41364
rect 428976 41352 428982 41404
rect 429838 41352 429844 41404
rect 429896 41392 429902 41404
rect 456794 41392 456800 41404
rect 429896 41364 456800 41392
rect 429896 41352 429902 41364
rect 456794 41352 456800 41364
rect 456852 41352 456858 41404
rect 457070 41352 457076 41404
rect 457128 41392 457134 41404
rect 484946 41392 484952 41404
rect 457128 41364 484952 41392
rect 457128 41352 457134 41364
rect 484946 41352 484952 41364
rect 485004 41352 485010 41404
rect 485038 41352 485044 41404
rect 485096 41392 485102 41404
rect 512914 41392 512920 41404
rect 485096 41364 512920 41392
rect 485096 41352 485102 41364
rect 512914 41352 512920 41364
rect 512972 41352 512978 41404
rect 513098 41352 513104 41404
rect 513156 41392 513162 41404
rect 540606 41392 540612 41404
rect 513156 41364 540612 41392
rect 513156 41352 513162 41364
rect 540606 41352 540612 41364
rect 540664 41352 540670 41404
rect 541066 41352 541072 41404
rect 541124 41392 541130 41404
rect 568942 41392 568948 41404
rect 541124 41364 568948 41392
rect 541124 41352 541130 41364
rect 568942 41352 568948 41364
rect 569000 41352 569006 41404
rect 26602 41284 26608 41336
rect 26660 41324 26666 41336
rect 40678 41324 40684 41336
rect 26660 41296 40684 41324
rect 26660 41284 26666 41296
rect 40678 41284 40684 41296
rect 40736 41284 40742 41336
rect 43438 41284 43444 41336
rect 43496 41324 43502 41336
rect 64874 41324 64880 41336
rect 43496 41296 64880 41324
rect 43496 41284 43502 41296
rect 64874 41284 64880 41296
rect 64932 41284 64938 41336
rect 82630 41284 82636 41336
rect 82688 41324 82694 41336
rect 93118 41324 93124 41336
rect 82688 41296 93124 41324
rect 82688 41284 82694 41296
rect 93118 41284 93124 41296
rect 93176 41284 93182 41336
rect 110598 41284 110604 41336
rect 110656 41324 110662 41336
rect 122098 41324 122104 41336
rect 110656 41296 122104 41324
rect 110656 41284 110662 41296
rect 122098 41284 122104 41296
rect 122156 41284 122162 41336
rect 128630 41284 128636 41336
rect 128688 41324 128694 41336
rect 149882 41324 149888 41336
rect 128688 41296 149888 41324
rect 128688 41284 128694 41296
rect 149882 41284 149888 41296
rect 149940 41284 149946 41336
rect 156322 41284 156328 41336
rect 156380 41324 156386 41336
rect 182818 41324 182824 41336
rect 156380 41296 182824 41324
rect 156380 41284 156386 41296
rect 182818 41284 182824 41296
rect 182876 41284 182882 41336
rect 194594 41284 194600 41336
rect 194652 41324 194658 41336
rect 206278 41324 206284 41336
rect 194652 41296 206284 41324
rect 194652 41284 194658 41296
rect 206278 41284 206284 41296
rect 206336 41284 206342 41336
rect 222930 41284 222936 41336
rect 222988 41324 222994 41336
rect 234062 41324 234068 41336
rect 222988 41296 234068 41324
rect 222988 41284 222994 41296
rect 234062 41284 234068 41296
rect 234120 41284 234126 41336
rect 240318 41284 240324 41336
rect 240376 41324 240382 41336
rect 261478 41324 261484 41336
rect 240376 41296 261484 41324
rect 240376 41284 240382 41296
rect 261478 41284 261484 41296
rect 261536 41284 261542 41336
rect 278590 41284 278596 41336
rect 278648 41324 278654 41336
rect 289170 41324 289176 41336
rect 278648 41296 289176 41324
rect 278648 41284 278654 41296
rect 289170 41284 289176 41296
rect 289228 41284 289234 41336
rect 306926 41284 306932 41336
rect 306984 41324 306990 41336
rect 318058 41324 318064 41336
rect 306984 41296 318064 41324
rect 306984 41284 306990 41296
rect 318058 41284 318064 41296
rect 318116 41284 318122 41336
rect 324314 41284 324320 41336
rect 324372 41324 324378 41336
rect 345658 41324 345664 41336
rect 324372 41296 345664 41324
rect 324372 41284 324378 41296
rect 345658 41284 345664 41296
rect 345716 41284 345722 41336
rect 352650 41284 352656 41336
rect 352708 41324 352714 41336
rect 373258 41324 373264 41336
rect 352708 41296 373264 41324
rect 352708 41284 352714 41296
rect 373258 41284 373264 41296
rect 373316 41284 373322 41336
rect 390646 41284 390652 41336
rect 390704 41324 390710 41336
rect 407206 41324 407212 41336
rect 390704 41296 407212 41324
rect 390704 41284 390710 41296
rect 407206 41284 407212 41296
rect 407264 41284 407270 41336
rect 418614 41284 418620 41336
rect 418672 41324 418678 41336
rect 436094 41324 436100 41336
rect 418672 41296 436100 41324
rect 418672 41284 418678 41296
rect 436094 41284 436100 41296
rect 436152 41284 436158 41336
rect 436646 41284 436652 41336
rect 436704 41324 436710 41336
rect 457438 41324 457444 41336
rect 436704 41296 457444 41324
rect 436704 41284 436710 41296
rect 457438 41284 457444 41296
rect 457496 41284 457502 41336
rect 474642 41284 474648 41336
rect 474700 41324 474706 41336
rect 486418 41324 486424 41336
rect 474700 41296 486424 41324
rect 474700 41284 474706 41296
rect 486418 41284 486424 41296
rect 486476 41284 486482 41336
rect 502610 41284 502616 41336
rect 502668 41324 502674 41336
rect 514018 41324 514024 41336
rect 502668 41296 514024 41324
rect 502668 41284 502674 41296
rect 514018 41284 514024 41296
rect 514076 41284 514082 41336
rect 520642 41284 520648 41336
rect 520700 41324 520706 41336
rect 541618 41324 541624 41336
rect 520700 41296 541624 41324
rect 520700 41284 520706 41296
rect 541618 41284 541624 41296
rect 541676 41284 541682 41336
rect 54938 41216 54944 41268
rect 54996 41256 55002 41268
rect 65978 41256 65984 41268
rect 54996 41228 65984 41256
rect 54996 41216 55002 41228
rect 65978 41216 65984 41228
rect 66036 41216 66042 41268
rect 138934 41216 138940 41268
rect 138992 41256 138998 41268
rect 149698 41256 149704 41268
rect 138992 41228 149704 41256
rect 138992 41216 138998 41228
rect 149698 41216 149704 41228
rect 149756 41216 149762 41268
rect 166626 41216 166632 41268
rect 166684 41256 166690 41268
rect 177298 41256 177304 41268
rect 166684 41228 177304 41256
rect 166684 41216 166690 41228
rect 177298 41216 177304 41228
rect 177356 41216 177362 41268
rect 250622 41216 250628 41268
rect 250680 41256 250686 41268
rect 261570 41256 261576 41268
rect 250680 41228 261576 41256
rect 250680 41216 250686 41228
rect 261570 41216 261576 41228
rect 261628 41216 261634 41268
rect 334618 41216 334624 41268
rect 334676 41256 334682 41268
rect 348418 41256 348424 41268
rect 334676 41228 348424 41256
rect 334676 41216 334682 41228
rect 348418 41216 348424 41228
rect 348476 41216 348482 41268
rect 362862 41216 362868 41268
rect 362920 41256 362926 41268
rect 374638 41256 374644 41268
rect 362920 41228 374644 41256
rect 362920 41216 362926 41228
rect 374638 41216 374644 41228
rect 374696 41216 374702 41268
rect 446950 41216 446956 41268
rect 447008 41256 447014 41268
rect 458818 41256 458824 41268
rect 447008 41228 458824 41256
rect 447008 41216 447014 41228
rect 458818 41216 458824 41228
rect 458876 41216 458882 41268
rect 530946 41216 530952 41268
rect 531004 41256 531010 41268
rect 541710 41256 541716 41268
rect 531004 41228 541716 41256
rect 531004 41216 531010 41228
rect 541710 41216 541716 41228
rect 541768 41216 541774 41268
rect 44634 41148 44640 41200
rect 44692 41188 44698 41200
rect 65886 41188 65892 41200
rect 44692 41160 65892 41188
rect 44692 41148 44698 41160
rect 65886 41148 65892 41160
rect 65944 41148 65950 41200
rect 558638 40672 558644 40724
rect 558696 40712 558702 40724
rect 568850 40712 568856 40724
rect 558696 40684 568856 40712
rect 558696 40672 558702 40684
rect 568850 40672 568856 40684
rect 568908 40672 568914 40724
rect 46934 39380 46940 39432
rect 46992 39420 46998 39432
rect 205082 39420 205088 39432
rect 46992 39392 205088 39420
rect 46992 39380 46998 39392
rect 205082 39380 205088 39392
rect 205140 39380 205146 39432
rect 548334 39380 548340 39432
rect 548392 39420 548398 39432
rect 569034 39420 569040 39432
rect 548392 39392 569040 39420
rect 548392 39380 548398 39392
rect 569034 39380 569040 39392
rect 569092 39380 569098 39432
rect 4982 39312 4988 39364
rect 5040 39352 5046 39364
rect 41782 39352 41788 39364
rect 5040 39324 41788 39352
rect 5040 39312 5046 39324
rect 41782 39312 41788 39324
rect 41840 39312 41846 39364
rect 61102 39312 61108 39364
rect 61160 39352 61166 39364
rect 569310 39352 569316 39364
rect 61160 39324 569316 39352
rect 61160 39312 61166 39324
rect 569310 39312 569316 39324
rect 569368 39312 569374 39364
rect 156322 38836 156328 38888
rect 156380 38876 156386 38888
rect 180058 38876 180064 38888
rect 156380 38848 180064 38876
rect 156380 38836 156386 38848
rect 180058 38836 180064 38848
rect 180116 38836 180122 38888
rect 352006 38836 352012 38888
rect 352064 38876 352070 38888
rect 373258 38876 373264 38888
rect 352064 38848 373264 38876
rect 352064 38836 352070 38848
rect 373258 38836 373264 38848
rect 373316 38836 373322 38888
rect 100018 38768 100024 38820
rect 100076 38808 100082 38820
rect 120994 38808 121000 38820
rect 100076 38780 121000 38808
rect 100076 38768 100082 38780
rect 120994 38768 121000 38780
rect 121052 38768 121058 38820
rect 176838 38768 176844 38820
rect 176896 38808 176902 38820
rect 194318 38808 194324 38820
rect 176896 38780 194324 38808
rect 176896 38768 176902 38780
rect 194318 38768 194324 38780
rect 194376 38768 194382 38820
rect 268010 38768 268016 38820
rect 268068 38808 268074 38820
rect 289078 38808 289084 38820
rect 268068 38780 289084 38808
rect 268068 38768 268074 38780
rect 289078 38768 289084 38780
rect 289136 38768 289142 38820
rect 345658 38768 345664 38820
rect 345716 38808 345722 38820
rect 362310 38808 362316 38820
rect 345716 38780 362316 38808
rect 345716 38768 345722 38780
rect 362310 38768 362316 38780
rect 362368 38768 362374 38820
rect 56594 38700 56600 38752
rect 56652 38740 56658 38752
rect 92474 38740 92480 38752
rect 56652 38712 92480 38740
rect 56652 38700 56658 38712
rect 92474 38700 92480 38712
rect 92532 38700 92538 38752
rect 92750 38700 92756 38752
rect 92808 38740 92814 38752
rect 110322 38740 110328 38752
rect 92808 38712 110328 38740
rect 92808 38700 92814 38712
rect 110322 38700 110328 38712
rect 110380 38700 110386 38752
rect 155218 38700 155224 38752
rect 155276 38740 155282 38752
rect 165982 38740 165988 38752
rect 155276 38712 165988 38740
rect 155276 38700 155282 38712
rect 165982 38700 165988 38712
rect 166040 38700 166046 38752
rect 184014 38700 184020 38752
rect 184072 38740 184078 38752
rect 204898 38740 204904 38752
rect 184072 38712 204904 38740
rect 184072 38700 184078 38712
rect 204898 38700 204904 38712
rect 204956 38700 204962 38752
rect 261478 38700 261484 38752
rect 261536 38740 261542 38752
rect 278314 38740 278320 38752
rect 261536 38712 278320 38740
rect 261536 38700 261542 38712
rect 278314 38700 278320 38712
rect 278372 38700 278378 38752
rect 317138 38700 317144 38752
rect 317196 38740 317202 38752
rect 334342 38740 334348 38752
rect 317196 38712 334348 38740
rect 317196 38700 317202 38712
rect 334342 38700 334348 38712
rect 334400 38700 334406 38752
rect 372798 38700 372804 38752
rect 372856 38740 372862 38752
rect 390002 38740 390008 38752
rect 372856 38712 390008 38740
rect 372856 38700 372862 38712
rect 390002 38700 390008 38712
rect 390060 38700 390066 38752
rect 401042 38700 401048 38752
rect 401100 38740 401106 38752
rect 418338 38740 418344 38752
rect 401100 38712 418344 38740
rect 401100 38700 401106 38712
rect 418338 38700 418344 38712
rect 418396 38700 418402 38752
rect 457438 38700 457444 38752
rect 457496 38740 457502 38752
rect 473998 38740 474004 38752
rect 457496 38712 474004 38740
rect 457496 38700 457502 38712
rect 473998 38700 474004 38712
rect 474056 38700 474062 38752
rect 484854 38700 484860 38752
rect 484912 38740 484918 38752
rect 502334 38740 502340 38752
rect 484912 38712 502340 38740
rect 484912 38700 484918 38712
rect 502334 38700 502340 38712
rect 502392 38700 502398 38752
rect 512730 38700 512736 38752
rect 512788 38740 512794 38752
rect 530302 38740 530308 38752
rect 512788 38712 530308 38740
rect 512788 38700 512794 38712
rect 530302 38700 530308 38712
rect 530360 38700 530366 38752
rect 13722 38632 13728 38684
rect 13780 38672 13786 38684
rect 81986 38672 81992 38684
rect 13780 38644 81992 38672
rect 13780 38632 13786 38644
rect 81986 38632 81992 38644
rect 82044 38632 82050 38684
rect 121086 38632 121092 38684
rect 121144 38672 121150 38684
rect 138290 38672 138296 38684
rect 121144 38644 138296 38672
rect 121144 38632 121150 38644
rect 138290 38632 138296 38644
rect 138348 38632 138354 38684
rect 178678 38632 178684 38684
rect 178736 38672 178742 38684
rect 204622 38672 204628 38684
rect 178736 38644 204628 38672
rect 178736 38632 178742 38644
rect 204622 38632 204628 38644
rect 204680 38632 204686 38684
rect 204806 38632 204812 38684
rect 204864 38672 204870 38684
rect 222194 38672 222200 38684
rect 204864 38644 222200 38672
rect 204864 38632 204870 38644
rect 222194 38632 222200 38644
rect 222252 38632 222258 38684
rect 233970 38632 233976 38684
rect 234028 38672 234034 38684
rect 260650 38672 260656 38684
rect 234028 38644 260656 38672
rect 234028 38632 234034 38644
rect 260650 38632 260656 38644
rect 260708 38632 260714 38684
rect 288894 38632 288900 38684
rect 288952 38672 288958 38684
rect 306006 38672 306012 38684
rect 288952 38644 306012 38672
rect 288952 38632 288958 38644
rect 306006 38632 306012 38644
rect 306064 38632 306070 38684
rect 317046 38632 317052 38684
rect 317104 38672 317110 38684
rect 344646 38672 344652 38684
rect 317104 38644 344652 38672
rect 317104 38632 317110 38644
rect 344646 38632 344652 38644
rect 344704 38632 344710 38684
rect 345750 38632 345756 38684
rect 345808 38672 345814 38684
rect 372614 38672 372620 38684
rect 345808 38644 372620 38672
rect 345808 38632 345814 38644
rect 372614 38632 372620 38644
rect 372672 38632 372678 38684
rect 380342 38632 380348 38684
rect 380400 38672 380406 38684
rect 401134 38672 401140 38684
rect 380400 38644 401140 38672
rect 380400 38632 380406 38644
rect 401134 38632 401140 38644
rect 401192 38632 401198 38684
rect 402238 38632 402244 38684
rect 402296 38672 402302 38684
rect 428642 38672 428648 38684
rect 402296 38644 428648 38672
rect 402296 38632 402302 38644
rect 428642 38632 428648 38644
rect 428700 38632 428706 38684
rect 428734 38632 428740 38684
rect 428792 38672 428798 38684
rect 446306 38672 446312 38684
rect 428792 38644 446312 38672
rect 428792 38632 428798 38644
rect 446306 38632 446312 38644
rect 446364 38632 446370 38684
rect 464338 38632 464344 38684
rect 464396 38672 464402 38684
rect 485038 38672 485044 38684
rect 464396 38644 485044 38672
rect 464396 38632 464402 38644
rect 485038 38632 485044 38644
rect 485096 38632 485102 38684
rect 486418 38632 486424 38684
rect 486476 38672 486482 38684
rect 512638 38672 512644 38684
rect 486476 38644 512644 38672
rect 486476 38632 486482 38644
rect 512638 38632 512644 38644
rect 512696 38632 512702 38684
rect 512822 38632 512828 38684
rect 512880 38672 512886 38684
rect 540606 38672 540612 38684
rect 512880 38644 540612 38672
rect 512880 38632 512886 38644
rect 540606 38632 540612 38644
rect 540664 38632 540670 38684
rect 26970 38564 26976 38616
rect 27028 38604 27034 38616
rect 37918 38604 37924 38616
rect 27028 38576 37924 38604
rect 27028 38564 27034 38576
rect 37918 38564 37924 38576
rect 37976 38564 37982 38616
rect 14458 38496 14464 38548
rect 14516 38536 14522 38548
rect 38562 38536 38568 38548
rect 14516 38508 38568 38536
rect 14516 38496 14522 38508
rect 38562 38496 38568 38508
rect 38620 38496 38626 38548
rect 3970 38428 3976 38480
rect 4028 38468 4034 38480
rect 33410 38468 33416 38480
rect 4028 38440 33416 38468
rect 4028 38428 4034 38440
rect 33410 38428 33416 38440
rect 33468 38428 33474 38480
rect 57882 38428 57888 38480
rect 57940 38468 57946 38480
rect 65794 38468 65800 38480
rect 57940 38440 65800 38468
rect 57940 38428 57946 38440
rect 65794 38428 65800 38440
rect 65852 38428 65858 38480
rect 11698 38360 11704 38412
rect 11756 38400 11762 38412
rect 22462 38400 22468 38412
rect 11756 38372 22468 38400
rect 11756 38360 11762 38372
rect 22462 38360 22468 38372
rect 22520 38360 22526 38412
rect 23750 38360 23756 38412
rect 23808 38400 23814 38412
rect 152458 38400 152464 38412
rect 23808 38372 152464 38400
rect 23808 38360 23814 38372
rect 152458 38360 152464 38372
rect 152516 38360 152522 38412
rect 19242 38292 19248 38344
rect 19300 38332 19306 38344
rect 234614 38332 234620 38344
rect 19300 38304 234620 38332
rect 19300 38292 19306 38304
rect 234614 38292 234620 38304
rect 234672 38292 234678 38344
rect 3418 38224 3424 38276
rect 3476 38264 3482 38276
rect 54662 38264 54668 38276
rect 3476 38236 54668 38264
rect 3476 38224 3482 38236
rect 54662 38224 54668 38236
rect 54720 38224 54726 38276
rect 64598 38224 64604 38276
rect 64656 38264 64662 38276
rect 569494 38264 569500 38276
rect 64656 38236 569500 38264
rect 64656 38224 64662 38236
rect 569494 38224 569500 38236
rect 569552 38224 569558 38276
rect 10318 38156 10324 38208
rect 10376 38196 10382 38208
rect 30190 38196 30196 38208
rect 10376 38168 30196 38196
rect 10376 38156 10382 38168
rect 30190 38156 30196 38168
rect 30248 38156 30254 38208
rect 32122 38156 32128 38208
rect 32180 38196 32186 38208
rect 545758 38196 545764 38208
rect 32180 38168 545764 38196
rect 32180 38156 32186 38168
rect 545758 38156 545764 38168
rect 545816 38156 545822 38208
rect 5166 38088 5172 38140
rect 5224 38128 5230 38140
rect 45002 38128 45008 38140
rect 5224 38100 45008 38128
rect 5224 38088 5230 38100
rect 45002 38088 45008 38100
rect 45060 38088 45066 38140
rect 51442 38088 51448 38140
rect 51500 38128 51506 38140
rect 569402 38128 569408 38140
rect 51500 38100 569408 38128
rect 51500 38088 51506 38100
rect 569402 38088 569408 38100
rect 569460 38088 569466 38140
rect 4798 38020 4804 38072
rect 4856 38060 4862 38072
rect 20530 38060 20536 38072
rect 4856 38032 20536 38060
rect 4856 38020 4862 38032
rect 20530 38020 20536 38032
rect 20588 38020 20594 38072
rect 25682 38020 25688 38072
rect 25740 38060 25746 38072
rect 580626 38060 580632 38072
rect 25740 38032 580632 38060
rect 25740 38020 25746 38032
rect 580626 38020 580632 38032
rect 580684 38020 580690 38072
rect 17310 37952 17316 38004
rect 17368 37992 17374 38004
rect 580442 37992 580448 38004
rect 17368 37964 580448 37992
rect 17368 37952 17374 37964
rect 580442 37952 580448 37964
rect 580500 37952 580506 38004
rect 16022 37884 16028 37936
rect 16080 37924 16086 37936
rect 580902 37924 580908 37936
rect 16080 37896 580908 37924
rect 16080 37884 16086 37896
rect 580902 37884 580908 37896
rect 580960 37884 580966 37936
rect 35342 37340 35348 37392
rect 35400 37380 35406 37392
rect 38010 37380 38016 37392
rect 35400 37352 38016 37380
rect 35400 37340 35406 37352
rect 38010 37340 38016 37352
rect 38068 37340 38074 37392
rect 40034 37340 40040 37392
rect 40092 37380 40098 37392
rect 48222 37380 48228 37392
rect 40092 37352 48228 37380
rect 40092 37340 40098 37352
rect 48222 37340 48228 37352
rect 48280 37340 48286 37392
rect 59814 37340 59820 37392
rect 59872 37380 59878 37392
rect 65702 37380 65708 37392
rect 59872 37352 65708 37380
rect 59872 37340 59878 37352
rect 65702 37340 65708 37352
rect 65760 37340 65766 37392
rect 36630 37272 36636 37324
rect 36688 37312 36694 37324
rect 95234 37312 95240 37324
rect 36688 37284 95240 37312
rect 36688 37272 36694 37284
rect 95234 37272 95240 37284
rect 95292 37272 95298 37324
rect 64506 36796 64512 36848
rect 64564 36836 64570 36848
rect 95878 36836 95884 36848
rect 64564 36808 95884 36836
rect 64564 36796 64570 36808
rect 95878 36796 95884 36808
rect 95936 36796 95942 36848
rect 64230 36728 64236 36780
rect 64288 36768 64294 36780
rect 569218 36768 569224 36780
rect 64288 36740 569224 36768
rect 64288 36728 64294 36740
rect 569218 36728 569224 36740
rect 569276 36728 569282 36780
rect 64414 36660 64420 36712
rect 64472 36700 64478 36712
rect 580350 36700 580356 36712
rect 64472 36672 580356 36700
rect 64472 36660 64478 36672
rect 580350 36660 580356 36672
rect 580408 36660 580414 36712
rect 64322 36592 64328 36644
rect 64380 36632 64386 36644
rect 580534 36632 580540 36644
rect 64380 36604 580540 36632
rect 64380 36592 64386 36604
rect 580534 36592 580540 36604
rect 580592 36592 580598 36644
rect 13538 36524 13544 36576
rect 13596 36564 13602 36576
rect 580810 36564 580816 36576
rect 13596 36536 580816 36564
rect 13596 36524 13602 36536
rect 580810 36524 580816 36536
rect 580868 36524 580874 36576
rect 120718 36252 120724 36304
rect 120776 36292 120782 36304
rect 121086 36292 121092 36304
rect 120776 36264 121092 36292
rect 120776 36252 120782 36264
rect 121086 36252 121092 36264
rect 121144 36252 121150 36304
rect 316862 36184 316868 36236
rect 316920 36224 316926 36236
rect 317046 36224 317052 36236
rect 316920 36196 317052 36224
rect 316920 36184 316926 36196
rect 317046 36184 317052 36196
rect 317104 36184 317110 36236
rect 400766 36184 400772 36236
rect 400824 36224 400830 36236
rect 401042 36224 401048 36236
rect 400824 36196 401048 36224
rect 400824 36184 400830 36196
rect 401042 36184 401048 36196
rect 401100 36184 401106 36236
rect 120810 36116 120816 36168
rect 120868 36156 120874 36168
rect 120994 36156 121000 36168
rect 120868 36128 121000 36156
rect 120868 36116 120874 36128
rect 120994 36116 121000 36128
rect 121052 36116 121058 36168
rect 316770 36116 316776 36168
rect 316828 36156 316834 36168
rect 317138 36156 317144 36168
rect 316828 36128 317144 36156
rect 316828 36116 316834 36128
rect 317138 36116 317144 36128
rect 317196 36116 317202 36168
rect 400858 36116 400864 36168
rect 400916 36156 400922 36168
rect 401134 36156 401140 36168
rect 400916 36128 401140 36156
rect 400916 36116 400922 36128
rect 401134 36116 401140 36128
rect 401192 36116 401198 36168
rect 39850 36048 39856 36100
rect 39908 36088 39914 36100
rect 61378 36088 61384 36100
rect 39908 36060 61384 36088
rect 39908 36048 39914 36060
rect 61378 36048 61384 36060
rect 61436 36048 61442 36100
rect 3418 35980 3424 36032
rect 3476 36020 3482 36032
rect 43438 36020 43444 36032
rect 3476 35992 43444 36020
rect 3476 35980 3482 35992
rect 43438 35980 43444 35992
rect 43496 35980 43502 36032
rect 50522 35980 50528 36032
rect 50580 36020 50586 36032
rect 61470 36020 61476 36032
rect 50580 35992 61476 36020
rect 50580 35980 50586 35992
rect 61470 35980 61476 35992
rect 61528 35980 61534 36032
rect 28718 35912 28724 35964
rect 28776 35952 28782 35964
rect 580902 35952 580908 35964
rect 28776 35924 580908 35952
rect 28776 35912 28782 35924
rect 580902 35912 580908 35924
rect 580960 35912 580966 35964
rect 3786 35164 3792 35216
rect 3844 35204 3850 35216
rect 61286 35204 61292 35216
rect 3844 35176 61292 35204
rect 3844 35164 3850 35176
rect 61286 35164 61292 35176
rect 61344 35164 61350 35216
rect 3326 31696 3332 31748
rect 3384 31736 3390 31748
rect 12434 31736 12440 31748
rect 3384 31708 12440 31736
rect 3384 31696 3390 31708
rect 12434 31696 12440 31708
rect 12492 31696 12498 31748
rect 64322 31016 64328 31068
rect 64380 31056 64386 31068
rect 64598 31056 64604 31068
rect 64380 31028 64604 31056
rect 64380 31016 64386 31028
rect 64598 31016 64604 31028
rect 64656 31016 64662 31068
rect 63494 27072 63500 27124
rect 63552 27112 63558 27124
rect 65610 27112 65616 27124
rect 63552 27084 65616 27112
rect 63552 27072 63558 27084
rect 65610 27072 65616 27084
rect 65668 27072 65674 27124
rect 5074 23400 5080 23452
rect 5132 23440 5138 23452
rect 12434 23440 12440 23452
rect 5132 23412 12440 23440
rect 5132 23400 5138 23412
rect 12434 23400 12440 23412
rect 12492 23400 12498 23452
rect 6178 22040 6184 22092
rect 6236 22080 6242 22092
rect 12434 22080 12440 22092
rect 6236 22052 12440 22080
rect 6236 22040 6242 22052
rect 12434 22040 12440 22052
rect 12492 22040 12498 22092
rect 176746 21360 176752 21412
rect 176804 21400 176810 21412
rect 176930 21400 176936 21412
rect 176804 21372 176936 21400
rect 176804 21360 176810 21372
rect 176930 21360 176936 21372
rect 176988 21360 176994 21412
rect 484762 21360 484768 21412
rect 484820 21400 484826 21412
rect 484946 21400 484952 21412
rect 484820 21372 484952 21400
rect 484820 21360 484826 21372
rect 484946 21360 484952 21372
rect 485004 21360 485010 21412
rect 7558 20612 7564 20664
rect 7616 20652 7622 20664
rect 12434 20652 12440 20664
rect 7616 20624 12440 20652
rect 7616 20612 7622 20624
rect 12434 20612 12440 20624
rect 12492 20612 12498 20664
rect 63494 19252 63500 19304
rect 63552 19292 63558 19304
rect 69658 19292 69664 19304
rect 63552 19264 69664 19292
rect 63552 19252 63558 19264
rect 69658 19252 69664 19264
rect 69716 19252 69722 19304
rect 289078 18640 289084 18692
rect 289136 18680 289142 18692
rect 295702 18680 295708 18692
rect 289136 18652 295708 18680
rect 289136 18640 289142 18652
rect 295702 18640 295708 18652
rect 295760 18640 295766 18692
rect 120810 18572 120816 18624
rect 120868 18612 120874 18624
rect 127710 18612 127716 18624
rect 120868 18584 127716 18612
rect 120868 18572 120874 18584
rect 127710 18572 127716 18584
rect 127768 18572 127774 18624
rect 373258 18572 373264 18624
rect 373316 18612 373322 18624
rect 379698 18612 379704 18624
rect 373316 18584 379704 18612
rect 373316 18572 373322 18584
rect 379698 18572 379704 18584
rect 379756 18572 379762 18624
rect 400858 18572 400864 18624
rect 400916 18612 400922 18624
rect 407758 18612 407764 18624
rect 400916 18584 407764 18612
rect 400916 18572 400922 18584
rect 407758 18572 407764 18584
rect 407816 18572 407822 18624
rect 204898 17960 204904 18012
rect 204956 18000 204962 18012
rect 211706 18000 211712 18012
rect 204956 17972 211712 18000
rect 204956 17960 204962 17972
rect 211706 17960 211712 17972
rect 211764 17960 211770 18012
rect 485038 17960 485044 18012
rect 485096 18000 485102 18012
rect 491662 18000 491668 18012
rect 485096 17972 491668 18000
rect 485096 17960 485102 17972
rect 491662 17960 491668 17972
rect 491720 17960 491726 18012
rect 6270 17892 6276 17944
rect 6328 17932 6334 17944
rect 12434 17932 12440 17944
rect 6328 17904 12440 17932
rect 6328 17892 6334 17904
rect 12434 17892 12440 17904
rect 12492 17892 12498 17944
rect 288526 16668 288532 16720
rect 288584 16708 288590 16720
rect 288894 16708 288900 16720
rect 288584 16680 288900 16708
rect 288584 16668 288590 16680
rect 288894 16668 288900 16680
rect 288952 16668 288958 16720
rect 568482 16668 568488 16720
rect 568540 16708 568546 16720
rect 569034 16708 569040 16720
rect 568540 16680 569040 16708
rect 568540 16668 568546 16680
rect 569034 16668 569040 16680
rect 569092 16668 569098 16720
rect 3786 16532 3792 16584
rect 3844 16572 3850 16584
rect 63586 16572 63592 16584
rect 3844 16544 63592 16572
rect 3844 16532 3850 16544
rect 63586 16532 63592 16544
rect 63644 16532 63650 16584
rect 4890 15104 4896 15156
rect 4948 15144 4954 15156
rect 35342 15144 35348 15156
rect 4948 15116 35348 15144
rect 4948 15104 4954 15116
rect 35342 15104 35348 15116
rect 35400 15104 35406 15156
rect 41782 15104 41788 15156
rect 41840 15144 41846 15156
rect 429194 15144 429200 15156
rect 41840 15116 429200 15144
rect 41840 15104 41846 15116
rect 429194 15104 429200 15116
rect 429252 15104 429258 15156
rect 5258 15036 5264 15088
rect 5316 15076 5322 15088
rect 22462 15076 22468 15088
rect 5316 15048 22468 15076
rect 5316 15036 5322 15048
rect 22462 15036 22468 15048
rect 22520 15036 22526 15088
rect 52730 15036 52736 15088
rect 52788 15076 52794 15088
rect 233878 15076 233884 15088
rect 52788 15048 233884 15076
rect 52788 15036 52794 15048
rect 233878 15036 233884 15048
rect 233936 15036 233942 15088
rect 23750 14968 23756 15020
rect 23808 15008 23814 15020
rect 65518 15008 65524 15020
rect 23808 14980 65524 15008
rect 23808 14968 23814 14980
rect 65518 14968 65524 14980
rect 65576 14968 65582 15020
rect 48222 14900 48228 14952
rect 48280 14940 48286 14952
rect 71038 14940 71044 14952
rect 48280 14912 71044 14940
rect 48280 14900 48286 14912
rect 71038 14900 71044 14912
rect 71096 14900 71102 14952
rect 9030 13744 9036 13796
rect 9088 13784 9094 13796
rect 16022 13784 16028 13796
rect 9088 13756 16028 13784
rect 9088 13744 9094 13756
rect 16022 13744 16028 13756
rect 16080 13744 16086 13796
rect 148594 13744 148600 13796
rect 148652 13784 148658 13796
rect 155218 13784 155224 13796
rect 148652 13756 155224 13784
rect 148652 13744 148658 13756
rect 155218 13744 155224 13756
rect 155276 13744 155282 13796
rect 166626 13744 166632 13796
rect 166684 13784 166690 13796
rect 178678 13784 178684 13796
rect 166684 13756 178684 13784
rect 166684 13744 166690 13756
rect 178678 13744 178684 13756
rect 178736 13744 178742 13796
rect 180058 13744 180064 13796
rect 180116 13784 180122 13796
rect 184014 13784 184020 13796
rect 180116 13756 184020 13784
rect 180116 13744 180122 13756
rect 184014 13744 184020 13756
rect 184072 13744 184078 13796
rect 222654 13744 222660 13796
rect 222712 13784 222718 13796
rect 233970 13784 233976 13796
rect 222712 13756 233976 13784
rect 222712 13744 222718 13756
rect 233970 13744 233976 13756
rect 234028 13744 234034 13796
rect 306282 13744 306288 13796
rect 306340 13784 306346 13796
rect 316862 13784 316868 13796
rect 306340 13756 316868 13784
rect 306340 13744 306346 13756
rect 316862 13744 316868 13756
rect 316920 13744 316926 13796
rect 390462 13744 390468 13796
rect 390520 13784 390526 13796
rect 402238 13784 402244 13796
rect 390520 13756 402244 13784
rect 390520 13744 390526 13756
rect 402238 13744 402244 13756
rect 402296 13744 402302 13796
rect 474642 13744 474648 13796
rect 474700 13784 474706 13796
rect 486418 13784 486424 13796
rect 474700 13756 486424 13784
rect 474700 13744 474706 13756
rect 486418 13744 486424 13756
rect 486476 13744 486482 13796
rect 502334 13744 502340 13796
rect 502392 13784 502398 13796
rect 512822 13784 512828 13796
rect 502392 13756 512828 13784
rect 502392 13744 502398 13756
rect 512822 13744 512828 13756
rect 512880 13744 512886 13796
rect 547874 13744 547880 13796
rect 547932 13784 547938 13796
rect 557994 13784 558000 13796
rect 547932 13756 558000 13784
rect 547932 13744 547938 13756
rect 557994 13744 558000 13756
rect 558052 13744 558058 13796
rect 17310 13676 17316 13728
rect 17368 13716 17374 13728
rect 574738 13716 574744 13728
rect 17368 13688 574744 13716
rect 17368 13676 17374 13688
rect 574738 13676 574744 13688
rect 574796 13676 574802 13728
rect 3510 13608 3516 13660
rect 3568 13648 3574 13660
rect 28902 13648 28908 13660
rect 3568 13620 28908 13648
rect 3568 13608 3574 13620
rect 28902 13608 28908 13620
rect 28960 13608 28966 13660
rect 32122 13608 32128 13660
rect 32180 13648 32186 13660
rect 580074 13648 580080 13660
rect 32180 13620 580080 13648
rect 32180 13608 32186 13620
rect 580074 13608 580080 13620
rect 580132 13608 580138 13660
rect 4062 13540 4068 13592
rect 4120 13580 4126 13592
rect 25682 13580 25688 13592
rect 4120 13552 25688 13580
rect 4120 13540 4126 13552
rect 25682 13540 25688 13552
rect 25740 13540 25746 13592
rect 36630 13540 36636 13592
rect 36688 13580 36694 13592
rect 580718 13580 580724 13592
rect 36688 13552 580724 13580
rect 36688 13540 36694 13552
rect 580718 13540 580724 13552
rect 580776 13540 580782 13592
rect 43070 13472 43076 13524
rect 43128 13512 43134 13524
rect 580166 13512 580172 13524
rect 43128 13484 580172 13512
rect 43128 13472 43134 13484
rect 580166 13472 580172 13484
rect 580224 13472 580230 13524
rect 3694 13404 3700 13456
rect 3752 13444 3758 13456
rect 57882 13444 57888 13456
rect 3752 13416 57888 13444
rect 3752 13404 3758 13416
rect 57882 13404 57888 13416
rect 57940 13404 57946 13456
rect 59814 13404 59820 13456
rect 59872 13444 59878 13456
rect 580258 13444 580264 13456
rect 59872 13416 580264 13444
rect 59872 13404 59878 13416
rect 580258 13404 580264 13416
rect 580316 13404 580322 13456
rect 19242 13336 19248 13388
rect 19300 13376 19306 13388
rect 518158 13376 518164 13388
rect 19300 13348 518164 13376
rect 19300 13336 19306 13348
rect 518158 13336 518164 13348
rect 518216 13336 518222 13388
rect 519998 13376 520004 13388
rect 518866 13348 520004 13376
rect 26970 13268 26976 13320
rect 27028 13308 27034 13320
rect 378778 13308 378784 13320
rect 27028 13280 378784 13308
rect 27028 13268 27034 13280
rect 378778 13268 378784 13280
rect 378836 13268 378842 13320
rect 407206 13268 407212 13320
rect 407264 13308 407270 13320
rect 436002 13308 436008 13320
rect 407264 13280 436008 13308
rect 407264 13268 407270 13280
rect 436002 13268 436008 13280
rect 436060 13268 436066 13320
rect 446306 13268 446312 13320
rect 446364 13308 446370 13320
rect 484946 13308 484952 13320
rect 446364 13280 484952 13308
rect 446364 13268 446370 13280
rect 484946 13268 484952 13280
rect 485004 13268 485010 13320
rect 491386 13268 491392 13320
rect 491444 13308 491450 13320
rect 518866 13308 518894 13348
rect 519998 13336 520004 13348
rect 520056 13336 520062 13388
rect 530302 13336 530308 13388
rect 530360 13376 530366 13388
rect 568942 13376 568948 13388
rect 530360 13348 568948 13376
rect 530360 13336 530366 13348
rect 568942 13336 568948 13348
rect 569000 13336 569006 13388
rect 491444 13280 518894 13308
rect 491444 13268 491450 13280
rect 518986 13268 518992 13320
rect 519044 13308 519050 13320
rect 547966 13308 547972 13320
rect 519044 13280 547972 13308
rect 519044 13268 519050 13280
rect 547966 13268 547972 13280
rect 548024 13268 548030 13320
rect 6914 13200 6920 13252
rect 6972 13240 6978 13252
rect 55950 13240 55956 13252
rect 6972 13212 55956 13240
rect 6972 13200 6978 13212
rect 55950 13200 55956 13212
rect 56008 13200 56014 13252
rect 82630 13200 82636 13252
rect 82688 13240 82694 13252
rect 120902 13240 120908 13252
rect 82688 13212 120908 13240
rect 82688 13200 82694 13212
rect 120902 13200 120908 13212
rect 120960 13200 120966 13252
rect 138290 13200 138296 13252
rect 138348 13240 138354 13252
rect 176930 13240 176936 13252
rect 138348 13212 176936 13240
rect 138348 13200 138354 13212
rect 176930 13200 176936 13212
rect 176988 13200 176994 13252
rect 194318 13200 194324 13252
rect 194376 13240 194382 13252
rect 232774 13240 232780 13252
rect 194376 13212 232780 13240
rect 194376 13200 194382 13212
rect 232774 13200 232780 13212
rect 232832 13200 232838 13252
rect 238846 13200 238852 13252
rect 238904 13240 238910 13252
rect 238904 13212 248414 13240
rect 238904 13200 238910 13212
rect 11790 13132 11796 13184
rect 11848 13172 11854 13184
rect 54662 13172 54668 13184
rect 11848 13144 54668 13172
rect 11848 13132 11854 13144
rect 54662 13132 54668 13144
rect 54720 13132 54726 13184
rect 71866 13132 71872 13184
rect 71924 13172 71930 13184
rect 100018 13172 100024 13184
rect 71924 13144 100024 13172
rect 71924 13132 71930 13144
rect 100018 13132 100024 13144
rect 100076 13132 100082 13184
rect 110322 13132 110328 13184
rect 110380 13172 110386 13184
rect 148778 13172 148784 13184
rect 110380 13144 148784 13172
rect 110380 13132 110386 13144
rect 148778 13132 148784 13144
rect 148836 13132 148842 13184
rect 211246 13132 211252 13184
rect 211304 13172 211310 13184
rect 240042 13172 240048 13184
rect 211304 13144 240048 13172
rect 211304 13132 211310 13144
rect 240042 13132 240048 13144
rect 240100 13132 240106 13184
rect 248386 13172 248414 13212
rect 250346 13200 250352 13252
rect 250404 13240 250410 13252
rect 288802 13240 288808 13252
rect 250404 13212 288808 13240
rect 250404 13200 250410 13212
rect 288802 13200 288808 13212
rect 288860 13200 288866 13252
rect 295426 13200 295432 13252
rect 295484 13240 295490 13252
rect 295484 13212 320036 13240
rect 295484 13200 295490 13212
rect 268010 13172 268016 13184
rect 248386 13144 268016 13172
rect 268010 13132 268016 13144
rect 268068 13132 268074 13184
rect 278314 13132 278320 13184
rect 278372 13172 278378 13184
rect 316954 13172 316960 13184
rect 278372 13144 316960 13172
rect 278372 13132 278378 13144
rect 316954 13132 316960 13144
rect 317012 13132 317018 13184
rect 320008 13172 320036 13212
rect 323026 13200 323032 13252
rect 323084 13240 323090 13252
rect 352006 13240 352012 13252
rect 323084 13212 352012 13240
rect 323084 13200 323090 13212
rect 352006 13200 352012 13212
rect 352064 13200 352070 13252
rect 362310 13200 362316 13252
rect 362368 13240 362374 13252
rect 400950 13240 400956 13252
rect 362368 13212 400956 13240
rect 362368 13200 362374 13212
rect 400950 13200 400956 13212
rect 401008 13200 401014 13252
rect 434806 13200 434812 13252
rect 434864 13240 434870 13252
rect 463694 13240 463700 13252
rect 434864 13212 463700 13240
rect 434864 13200 434870 13212
rect 463694 13200 463700 13212
rect 463752 13200 463758 13252
rect 324038 13172 324044 13184
rect 320008 13144 324044 13172
rect 324038 13132 324044 13144
rect 324096 13132 324102 13184
rect 334342 13132 334348 13184
rect 334400 13172 334406 13184
rect 345750 13172 345756 13184
rect 334400 13144 345756 13172
rect 334400 13132 334406 13144
rect 345750 13132 345756 13144
rect 345808 13132 345814 13184
rect 1394 13064 1400 13116
rect 1452 13104 1458 13116
rect 33410 13104 33416 13116
rect 1452 13076 33416 13104
rect 1452 13064 1458 13076
rect 33410 13064 33416 13076
rect 33468 13064 33474 13116
rect 38562 13064 38568 13116
rect 38620 13104 38626 13116
rect 72050 13104 72056 13116
rect 38620 13076 72056 13104
rect 38620 13064 38626 13076
rect 72050 13064 72056 13076
rect 72108 13064 72114 13116
rect 127066 13064 127072 13116
rect 127124 13104 127130 13116
rect 156046 13104 156052 13116
rect 127124 13076 156052 13104
rect 127124 13064 127130 13076
rect 156046 13064 156052 13076
rect 156104 13064 156110 13116
rect 8938 12996 8944 13048
rect 8996 13036 9002 13048
rect 30190 13036 30196 13048
rect 8996 13008 30196 13036
rect 8996 12996 9002 13008
rect 30190 12996 30196 13008
rect 30248 12996 30254 13048
rect 39850 12996 39856 13048
rect 39908 13036 39914 13048
rect 68278 13036 68284 13048
rect 39908 13008 68284 13036
rect 39908 12996 39914 13008
rect 68278 12996 68284 13008
rect 68336 12996 68342 13048
rect 20530 12928 20536 12980
rect 20588 12968 20594 12980
rect 578878 12968 578884 12980
rect 20588 12940 578884 12968
rect 20588 12928 20594 12940
rect 578878 12928 578884 12940
rect 578936 12928 578942 12980
rect 3602 12860 3608 12912
rect 3660 12900 3666 12912
rect 46290 12900 46296 12912
rect 3660 12872 46296 12900
rect 3660 12860 3666 12872
rect 46290 12860 46296 12872
rect 46348 12860 46354 12912
rect 3878 12792 3884 12844
rect 3936 12832 3942 12844
rect 51442 12832 51448 12844
rect 3936 12804 51448 12832
rect 3936 12792 3942 12804
rect 51442 12792 51448 12804
rect 51500 12792 51506 12844
rect 64230 3680 64236 3732
rect 64288 3720 64294 3732
rect 125870 3720 125876 3732
rect 64288 3692 125876 3720
rect 64288 3680 64294 3692
rect 125870 3680 125876 3692
rect 125928 3680 125934 3732
rect 64138 3612 64144 3664
rect 64196 3652 64202 3664
rect 126974 3652 126980 3664
rect 64196 3624 126980 3652
rect 64196 3612 64202 3624
rect 126974 3612 126980 3624
rect 127032 3612 127038 3664
rect 61470 3544 61476 3596
rect 61528 3584 61534 3596
rect 132954 3584 132960 3596
rect 61528 3556 132960 3584
rect 61528 3544 61534 3556
rect 132954 3544 132960 3556
rect 133012 3544 133018 3596
rect 13722 3476 13728 3528
rect 13780 3516 13786 3528
rect 129366 3516 129372 3528
rect 13780 3488 129372 3516
rect 13780 3476 13786 3488
rect 129366 3476 129372 3488
rect 129424 3476 129430 3528
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 48314 3448 48320 3460
rect 624 3420 48320 3448
rect 624 3408 630 3420
rect 48314 3408 48320 3420
rect 48372 3408 48378 3460
rect 61378 3408 61384 3460
rect 61436 3448 61442 3460
rect 136450 3448 136456 3460
rect 61436 3420 136456 3448
rect 61436 3408 61442 3420
rect 136450 3408 136456 3420
rect 136508 3408 136514 3460
<< via1 >>
rect 37924 700748 37976 700800
rect 105452 700748 105504 700800
rect 65616 700680 65668 700732
rect 267648 700680 267700 700732
rect 65708 700612 65760 700664
rect 332508 700612 332560 700664
rect 95884 700544 95936 700596
rect 364984 700544 365036 700596
rect 13452 700476 13504 700528
rect 300124 700476 300176 700528
rect 378784 700476 378836 700528
rect 397460 700476 397512 700528
rect 71044 700408 71096 700460
rect 170312 700408 170364 700460
rect 205088 700408 205140 700460
rect 494796 700408 494848 700460
rect 65524 700340 65576 700392
rect 137836 700340 137888 700392
rect 152464 700340 152516 700392
rect 462320 700340 462372 700392
rect 518164 700340 518216 700392
rect 527180 700340 527232 700392
rect 65800 700272 65852 700324
rect 202788 700272 202840 700324
rect 233884 700272 233936 700324
rect 559656 700272 559708 700324
rect 68284 699660 68336 699712
rect 72976 699660 73028 699712
rect 100024 687352 100076 687404
rect 121092 687352 121144 687404
rect 268016 687352 268068 687404
rect 289084 687352 289136 687404
rect 380348 687352 380400 687404
rect 401140 687352 401192 687404
rect 464344 687352 464396 687404
rect 485044 687352 485096 687404
rect 36912 687284 36964 687336
rect 54300 687284 54352 687336
rect 65892 687284 65944 687336
rect 81992 687284 82044 687336
rect 92940 687284 92992 687336
rect 110328 687284 110380 687336
rect 176936 687284 176988 687336
rect 194324 687284 194376 687336
rect 261484 687284 261536 687336
rect 278320 687284 278372 687336
rect 317144 687284 317196 687336
rect 334348 687284 334400 687336
rect 372988 687284 373040 687336
rect 390008 687284 390060 687336
rect 457444 687284 457496 687336
rect 474004 687284 474056 687336
rect 15292 687216 15344 687268
rect 26332 687216 26384 687268
rect 39304 687216 39356 687268
rect 64604 687216 64656 687268
rect 72332 687216 72384 687268
rect 93124 687216 93176 687268
rect 121000 687216 121052 687268
rect 138296 687216 138348 687268
rect 156328 687216 156380 687268
rect 177304 687216 177356 687268
rect 184020 687216 184072 687268
rect 204720 687216 204772 687268
rect 209044 687216 209096 687268
rect 222200 687216 222252 687268
rect 232964 687216 233016 687268
rect 250352 687216 250404 687268
rect 288992 687216 289044 687268
rect 306012 687216 306064 687268
rect 317052 687216 317104 687268
rect 344652 687216 344704 687268
rect 352012 687216 352064 687268
rect 373264 687216 373316 687268
rect 401048 687216 401100 687268
rect 418344 687216 418396 687268
rect 429844 687216 429896 687268
rect 456616 687216 456668 687268
rect 484952 687216 485004 687268
rect 502340 687216 502392 687268
rect 512920 687216 512972 687268
rect 530308 687216 530360 687268
rect 92756 684224 92808 684276
rect 92940 684224 92992 684276
rect 120724 684224 120776 684276
rect 121000 684224 121052 684276
rect 204720 684224 204772 684276
rect 204996 684224 205048 684276
rect 232780 684224 232832 684276
rect 232964 684224 233016 684276
rect 316868 684224 316920 684276
rect 317052 684224 317104 684276
rect 372804 684224 372856 684276
rect 372988 684224 373040 684276
rect 400772 684224 400824 684276
rect 401048 684224 401100 684276
rect 120816 684156 120868 684208
rect 121092 684156 121144 684208
rect 316776 684156 316828 684208
rect 317144 684156 317196 684208
rect 400864 684156 400916 684208
rect 401140 684156 401192 684208
rect 176752 683272 176804 683324
rect 288808 683136 288860 683188
rect 484860 683136 484912 683188
rect 512828 683136 512880 683188
rect 176844 683068 176896 683120
rect 288900 682932 288952 682984
rect 484860 682932 484912 682984
rect 512828 682932 512880 682984
rect 512736 682592 512788 682644
rect 512920 682592 512972 682644
rect 204812 681708 204864 681760
rect 209044 681708 209096 681760
rect 288808 681028 288860 681080
rect 288992 681028 289044 681080
rect 176752 679464 176804 679516
rect 176936 679464 176988 679516
rect 484768 677900 484820 677952
rect 484952 677900 485004 677952
rect 64880 669060 64932 669112
rect 65892 669060 65944 669112
rect 36820 668584 36872 668636
rect 37004 668584 37056 668636
rect 204904 667836 204956 667888
rect 211712 667836 211764 667888
rect 485044 667836 485096 667888
rect 491668 667836 491720 667888
rect 289084 667360 289136 667412
rect 295708 667360 295760 667412
rect 93124 667156 93176 667208
rect 99748 667156 99800 667208
rect 120816 667156 120868 667208
rect 127716 667156 127768 667208
rect 177304 667156 177356 667208
rect 183652 667156 183704 667208
rect 373264 667156 373316 667208
rect 379704 667156 379756 667208
rect 400864 667156 400916 667208
rect 407764 667156 407816 667208
rect 42708 665116 42760 665168
rect 95240 665116 95292 665168
rect 97908 665116 97960 665168
rect 150440 665116 150492 665168
rect 154488 665116 154540 665168
rect 207020 665116 207072 665168
rect 209688 665116 209740 665168
rect 262220 665116 262272 665168
rect 266268 665116 266320 665168
rect 318800 665116 318852 665168
rect 322848 665116 322900 665168
rect 375380 665116 375432 665168
rect 378048 665116 378100 665168
rect 430580 665116 430632 665168
rect 434628 665116 434680 665168
rect 487160 665116 487212 665168
rect 489828 665116 489880 665168
rect 542360 665116 542412 665168
rect 15292 664708 15344 664760
rect 16120 664708 16172 664760
rect 36544 664708 36596 664760
rect 36912 664708 36964 664760
rect 15384 662328 15436 662380
rect 43628 662328 43680 662380
rect 138664 662328 138716 662380
rect 176844 662328 176896 662380
rect 194324 662328 194376 662380
rect 232872 662328 232924 662380
rect 238852 662328 238904 662380
rect 26332 662260 26384 662312
rect 39304 662260 39356 662312
rect 42892 662260 42944 662312
rect 71780 662260 71832 662312
rect 82636 662260 82688 662312
rect 120908 662260 120960 662312
rect 127072 662260 127124 662312
rect 155960 662260 156012 662312
rect 166632 662260 166684 662312
rect 204996 662260 205048 662312
rect 211252 662260 211304 662312
rect 239772 662260 239824 662312
rect 295432 662328 295484 662380
rect 323676 662328 323728 662380
rect 334624 662328 334676 662380
rect 372896 662328 372948 662380
rect 390468 662328 390520 662380
rect 428740 662328 428792 662380
rect 434812 662328 434864 662380
rect 268016 662260 268068 662312
rect 278320 662260 278372 662312
rect 316960 662260 317012 662312
rect 323032 662260 323084 662312
rect 352012 662260 352064 662312
rect 362316 662260 362368 662312
rect 400956 662260 401008 662312
rect 407212 662260 407264 662312
rect 436008 662260 436060 662312
rect 491392 662328 491444 662380
rect 520004 662328 520056 662380
rect 530308 662328 530360 662380
rect 568764 662328 568816 662380
rect 463792 662260 463844 662312
rect 474648 662260 474700 662312
rect 512828 662260 512880 662312
rect 518992 662260 519044 662312
rect 547880 662260 547932 662312
rect 54576 662192 54628 662244
rect 92848 662192 92900 662244
rect 110328 662192 110380 662244
rect 148784 662192 148836 662244
rect 250720 662192 250772 662244
rect 288900 662192 288952 662244
rect 306288 662192 306340 662244
rect 316868 662192 316920 662244
rect 418344 662192 418396 662244
rect 429844 662192 429896 662244
rect 446312 662192 446364 662244
rect 484860 662192 484912 662244
rect 502340 662192 502392 662244
rect 540796 662192 540848 662244
rect 13636 661648 13688 661700
rect 558000 661648 558052 661700
rect 26608 660288 26660 660340
rect 36820 660288 36872 660340
rect 38016 659744 38068 659796
rect 44180 659744 44232 659796
rect 71872 659744 71924 659796
rect 110604 659744 110656 659796
rect 211252 659744 211304 659796
rect 250628 659744 250680 659796
rect 295432 659744 295484 659796
rect 334624 659744 334676 659796
rect 407212 659744 407264 659796
rect 446312 659744 446364 659796
rect 491392 659744 491444 659796
rect 530308 659744 530360 659796
rect 15568 659676 15620 659728
rect 54300 659676 54352 659728
rect 99472 659676 99524 659728
rect 138296 659676 138348 659728
rect 149796 659676 149848 659728
rect 166632 659676 166684 659728
rect 183652 659676 183704 659728
rect 222292 659676 222344 659728
rect 233976 659676 234028 659728
rect 240324 659676 240376 659728
rect 267832 659676 267884 659728
rect 306472 659676 306524 659728
rect 318064 659676 318116 659728
rect 324320 659676 324372 659728
rect 345756 659676 345808 659728
rect 362316 659676 362368 659728
rect 379612 659676 379664 659728
rect 418620 659676 418672 659728
rect 429844 659676 429896 659728
rect 436100 659676 436152 659728
rect 463792 659676 463844 659728
rect 502616 659676 502668 659728
rect 541624 659676 541676 659728
rect 558644 659676 558696 659728
rect 205088 657296 205140 657348
rect 205088 657092 205140 657144
rect 3516 656888 3568 656940
rect 11704 656888 11756 656940
rect 42708 656888 42760 656940
rect 95240 656888 95292 656940
rect 97908 656888 97960 656940
rect 150440 656888 150492 656940
rect 154488 656888 154540 656940
rect 207020 656888 207072 656940
rect 209688 656888 209740 656940
rect 262220 656888 262272 656940
rect 266268 656888 266320 656940
rect 318800 656888 318852 656940
rect 322848 656888 322900 656940
rect 375380 656888 375432 656940
rect 378048 656888 378100 656940
rect 430580 656888 430632 656940
rect 434628 656888 434680 656940
rect 487160 656888 487212 656940
rect 489828 656888 489880 656940
rect 542360 656888 542412 656940
rect 71780 655664 71832 655716
rect 71964 655664 72016 655716
rect 99380 655664 99432 655716
rect 99932 655664 99984 655716
rect 183560 655664 183612 655716
rect 184020 655664 184072 655716
rect 211160 655664 211212 655716
rect 211988 655664 212040 655716
rect 267740 655664 267792 655716
rect 267924 655664 267976 655716
rect 295340 655664 295392 655716
rect 295984 655664 296036 655716
rect 379520 655664 379572 655716
rect 379980 655664 380032 655716
rect 407120 655664 407172 655716
rect 407948 655664 408000 655716
rect 463700 655664 463752 655716
rect 464068 655664 464120 655716
rect 491300 655664 491352 655716
rect 492036 655664 492088 655716
rect 15200 634720 15252 634772
rect 36912 634720 36964 634772
rect 37096 634720 37148 634772
rect 64880 634720 64932 634772
rect 65064 634720 65116 634772
rect 92940 634720 92992 634772
rect 93032 634720 93084 634772
rect 120908 634720 120960 634772
rect 121092 634720 121144 634772
rect 148600 634720 148652 634772
rect 149704 634720 149756 634772
rect 176936 634720 176988 634772
rect 177028 634720 177080 634772
rect 204904 634720 204956 634772
rect 205180 634720 205232 634772
rect 232596 634720 232648 634772
rect 233056 634720 233108 634772
rect 260932 634720 260984 634772
rect 261024 634720 261076 634772
rect 288900 634720 288952 634772
rect 289084 634720 289136 634772
rect 316592 634720 316644 634772
rect 317052 634720 317104 634772
rect 344928 634720 344980 634772
rect 345664 634720 345716 634772
rect 372620 634720 372672 634772
rect 373080 634720 373132 634772
rect 400956 634720 401008 634772
rect 401048 634720 401100 634772
rect 428924 634720 428976 634772
rect 429108 634720 429160 634772
rect 456800 634720 456852 634772
rect 457076 634720 457128 634772
rect 484952 634720 485004 634772
rect 485044 634720 485096 634772
rect 512920 634720 512972 634772
rect 513104 634720 513156 634772
rect 540612 634720 540664 634772
rect 541072 634720 541124 634772
rect 568948 634720 569000 634772
rect 26608 634652 26660 634704
rect 38016 634652 38068 634704
rect 54944 634652 54996 634704
rect 71780 634652 71832 634704
rect 82636 634652 82688 634704
rect 99380 634652 99432 634704
rect 128636 634652 128688 634704
rect 149796 634652 149848 634704
rect 166632 634652 166684 634704
rect 183560 634652 183612 634704
rect 194600 634652 194652 634704
rect 211160 634652 211212 634704
rect 222936 634652 222988 634704
rect 233976 634652 234028 634704
rect 250628 634652 250680 634704
rect 267740 634652 267792 634704
rect 278596 634652 278648 634704
rect 295340 634652 295392 634704
rect 306932 634652 306984 634704
rect 318064 634652 318116 634704
rect 324320 634652 324372 634704
rect 345756 634652 345808 634704
rect 362868 634652 362920 634704
rect 379520 634652 379572 634704
rect 390652 634652 390704 634704
rect 407120 634652 407172 634704
rect 418620 634652 418672 634704
rect 429844 634652 429896 634704
rect 446956 634652 447008 634704
rect 463700 634652 463752 634704
rect 474648 634652 474700 634704
rect 491300 634652 491352 634704
rect 520648 634652 520700 634704
rect 541624 634652 541676 634704
rect 138940 634584 138992 634636
rect 155960 634584 156012 634636
rect 334624 634584 334676 634636
rect 351920 634584 351972 634636
rect 530952 634584 531004 634636
rect 547972 634584 548024 634636
rect 558644 634040 558696 634092
rect 568948 634040 569000 634092
rect 548340 632680 548392 632732
rect 569040 632680 569092 632732
rect 100024 632204 100076 632256
rect 121092 632204 121144 632256
rect 184020 632204 184072 632256
rect 204904 632204 204956 632256
rect 268016 632204 268068 632256
rect 289084 632204 289136 632256
rect 380348 632204 380400 632256
rect 401140 632204 401192 632256
rect 464344 632204 464396 632256
rect 485044 632204 485096 632256
rect 37096 632136 37148 632188
rect 54300 632136 54352 632188
rect 65892 632136 65944 632188
rect 81992 632136 82044 632188
rect 92848 632136 92900 632188
rect 110328 632136 110380 632188
rect 176844 632136 176896 632188
rect 194324 632136 194376 632188
rect 261484 632136 261536 632188
rect 278320 632136 278372 632188
rect 317144 632136 317196 632188
rect 334348 632136 334400 632188
rect 372988 632136 373040 632188
rect 390008 632136 390060 632188
rect 457444 632136 457496 632188
rect 474004 632136 474056 632188
rect 2780 632068 2832 632120
rect 4804 632068 4856 632120
rect 15292 632068 15344 632120
rect 26332 632068 26384 632120
rect 39304 632068 39356 632120
rect 64604 632068 64656 632120
rect 72332 632068 72384 632120
rect 93124 632068 93176 632120
rect 121000 632068 121052 632120
rect 138296 632068 138348 632120
rect 156328 632068 156380 632120
rect 177304 632068 177356 632120
rect 204812 632068 204864 632120
rect 222200 632068 222252 632120
rect 232964 632068 233016 632120
rect 250352 632068 250404 632120
rect 288900 632068 288952 632120
rect 306012 632068 306064 632120
rect 317052 632068 317104 632120
rect 344652 632068 344704 632120
rect 352012 632068 352064 632120
rect 373264 632068 373316 632120
rect 401048 632068 401100 632120
rect 418344 632068 418396 632120
rect 429844 632068 429896 632120
rect 456616 632068 456668 632120
rect 484860 632068 484912 632120
rect 502340 632068 502392 632120
rect 514852 632068 514904 632120
rect 530308 632068 530360 632120
rect 36728 630232 36780 630284
rect 37096 630232 37148 630284
rect 120724 630232 120776 630284
rect 121000 630232 121052 630284
rect 204720 630232 204772 630284
rect 204996 630232 205048 630284
rect 120816 630164 120868 630216
rect 121092 630164 121144 630216
rect 400864 630164 400916 630216
rect 401140 630164 401192 630216
rect 316776 628668 316828 628720
rect 317144 628668 317196 628720
rect 232780 628600 232832 628652
rect 232964 628600 233016 628652
rect 316868 628600 316920 628652
rect 317052 628600 317104 628652
rect 372804 628600 372856 628652
rect 372988 628600 373040 628652
rect 400772 628600 400824 628652
rect 401048 628600 401100 628652
rect 512736 628600 512788 628652
rect 514852 628600 514904 628652
rect 568764 625812 568816 625864
rect 568948 625812 569000 625864
rect 92756 613980 92808 614032
rect 92940 613980 92992 614032
rect 93124 613368 93176 613420
rect 99748 613368 99800 613420
rect 120816 613368 120868 613420
rect 127716 613368 127768 613420
rect 177304 613368 177356 613420
rect 183652 613368 183704 613420
rect 373264 613368 373316 613420
rect 379704 613368 379756 613420
rect 400864 613368 400916 613420
rect 407764 613368 407816 613420
rect 64880 613096 64932 613148
rect 65892 613096 65944 613148
rect 204904 613096 204956 613148
rect 211712 613096 211764 613148
rect 485044 613096 485096 613148
rect 491668 613096 491720 613148
rect 289084 612756 289136 612808
rect 295708 612756 295760 612808
rect 42708 611260 42760 611312
rect 95240 611260 95292 611312
rect 97908 611260 97960 611312
rect 150440 611260 150492 611312
rect 154488 611260 154540 611312
rect 207020 611260 207072 611312
rect 209688 611260 209740 611312
rect 262220 611260 262272 611312
rect 266268 611260 266320 611312
rect 318800 611260 318852 611312
rect 322848 611260 322900 611312
rect 375380 611260 375432 611312
rect 378048 611260 378100 611312
rect 430580 611260 430632 611312
rect 434628 611260 434680 611312
rect 487160 611260 487212 611312
rect 489828 611260 489880 611312
rect 542360 611260 542412 611312
rect 176752 610784 176804 610836
rect 176936 610784 176988 610836
rect 288808 610784 288860 610836
rect 288992 610784 289044 610836
rect 484768 610784 484820 610836
rect 484952 610784 485004 610836
rect 547880 610648 547932 610700
rect 548156 610648 548208 610700
rect 15292 610104 15344 610156
rect 15936 609900 15988 609952
rect 15384 608540 15436 608592
rect 43996 608540 44048 608592
rect 138296 608540 138348 608592
rect 176936 608540 176988 608592
rect 194324 608540 194376 608592
rect 232872 608540 232924 608592
rect 238852 608540 238904 608592
rect 26332 608472 26384 608524
rect 39304 608472 39356 608524
rect 42892 608472 42944 608524
rect 71780 608472 71832 608524
rect 110328 608472 110380 608524
rect 148784 608472 148836 608524
rect 166632 608472 166684 608524
rect 204996 608472 205048 608524
rect 211252 608472 211304 608524
rect 240048 608472 240100 608524
rect 295432 608540 295484 608592
rect 324044 608540 324096 608592
rect 334348 608540 334400 608592
rect 372896 608540 372948 608592
rect 390468 608540 390520 608592
rect 428740 608540 428792 608592
rect 434812 608540 434864 608592
rect 268016 608472 268068 608524
rect 278320 608472 278372 608524
rect 316960 608472 317012 608524
rect 323032 608472 323084 608524
rect 352012 608472 352064 608524
rect 362316 608472 362368 608524
rect 400956 608472 401008 608524
rect 407212 608472 407264 608524
rect 436008 608472 436060 608524
rect 491392 608540 491444 608592
rect 520004 608540 520056 608592
rect 530308 608540 530360 608592
rect 568856 608540 568908 608592
rect 463700 608472 463752 608524
rect 474648 608472 474700 608524
rect 512828 608472 512880 608524
rect 548156 608472 548208 608524
rect 558000 608472 558052 608524
rect 82636 608404 82688 608456
rect 120908 608404 120960 608456
rect 127072 608404 127124 608456
rect 156052 608404 156104 608456
rect 250352 608404 250404 608456
rect 288992 608404 289044 608456
rect 306288 608404 306340 608456
rect 316868 608404 316920 608456
rect 418344 608404 418396 608456
rect 429844 608404 429896 608456
rect 446312 608404 446364 608456
rect 484952 608404 485004 608456
rect 502340 608404 502392 608456
rect 540796 608404 540848 608456
rect 54300 608336 54352 608388
rect 92940 608336 92992 608388
rect 518992 608336 519044 608388
rect 547880 608336 547932 608388
rect 26608 606432 26660 606484
rect 36820 606432 36872 606484
rect 15384 605956 15436 606008
rect 54300 605956 54352 606008
rect 2780 605888 2832 605940
rect 4896 605888 4948 605940
rect 71872 605888 71924 605940
rect 110604 605888 110656 605940
rect 149888 605888 149940 605940
rect 156328 605888 156380 605940
rect 211252 605888 211304 605940
rect 250628 605888 250680 605940
rect 267832 605888 267884 605940
rect 306380 605888 306432 605940
rect 318064 605888 318116 605940
rect 324320 605888 324372 605940
rect 345756 605888 345808 605940
rect 362316 605888 362368 605940
rect 407212 605888 407264 605940
rect 446312 605888 446364 605940
rect 463792 605888 463844 605940
rect 502616 605888 502668 605940
rect 514024 605888 514076 605940
rect 520280 605888 520332 605940
rect 38108 605820 38160 605872
rect 44180 605820 44232 605872
rect 65892 605820 65944 605872
rect 82636 605820 82688 605872
rect 99380 605820 99432 605872
rect 138296 605820 138348 605872
rect 149796 605820 149848 605872
rect 166632 605820 166684 605872
rect 183560 605820 183612 605872
rect 222384 605820 222436 605872
rect 234068 605820 234120 605872
rect 240324 605820 240376 605872
rect 261484 605820 261536 605872
rect 278596 605820 278648 605872
rect 295340 605820 295392 605872
rect 334624 605820 334676 605872
rect 345664 605820 345716 605872
rect 352012 605820 352064 605872
rect 379520 605820 379572 605872
rect 418620 605820 418672 605872
rect 429936 605820 429988 605872
rect 436100 605820 436152 605872
rect 457444 605820 457496 605872
rect 474648 605820 474700 605872
rect 491300 605820 491352 605872
rect 530308 605820 530360 605872
rect 541624 605820 541676 605872
rect 558644 605820 558696 605872
rect 205088 603304 205140 603356
rect 345020 603236 345072 603288
rect 345848 603236 345900 603288
rect 205088 603100 205140 603152
rect 429108 603100 429160 603152
rect 429844 603100 429896 603152
rect 37280 599700 37332 599752
rect 38016 599700 38068 599752
rect 71780 599700 71832 599752
rect 71964 599700 72016 599752
rect 211160 599700 211212 599752
rect 211988 599700 212040 599752
rect 233240 599700 233292 599752
rect 233976 599700 234028 599752
rect 267740 599700 267792 599752
rect 267924 599700 267976 599752
rect 407120 599700 407172 599752
rect 407948 599700 408000 599752
rect 463700 599700 463752 599752
rect 464068 599700 464120 599752
rect 93124 585760 93176 585812
rect 99472 585760 99524 585812
rect 177120 585760 177172 585812
rect 183652 585760 183704 585812
rect 373172 585760 373224 585812
rect 379612 585760 379664 585812
rect 289728 585148 289780 585200
rect 295432 585148 295484 585200
rect 485136 585148 485188 585200
rect 491392 585148 491444 585200
rect 15200 580932 15252 580984
rect 36912 580932 36964 580984
rect 38016 580932 38068 580984
rect 64880 580932 64932 580984
rect 65064 580932 65116 580984
rect 92940 580932 92992 580984
rect 93032 580932 93084 580984
rect 120908 580932 120960 580984
rect 121092 580932 121144 580984
rect 148600 580932 148652 580984
rect 149704 580932 149756 580984
rect 176936 580932 176988 580984
rect 177028 580932 177080 580984
rect 204904 580932 204956 580984
rect 205180 580932 205232 580984
rect 232596 580932 232648 580984
rect 233976 580932 234028 580984
rect 260932 580932 260984 580984
rect 261024 580932 261076 580984
rect 288900 580932 288952 580984
rect 289084 580932 289136 580984
rect 316592 580932 316644 580984
rect 317052 580932 317104 580984
rect 344928 580932 344980 580984
rect 345848 580932 345900 580984
rect 372620 580932 372672 580984
rect 373080 580932 373132 580984
rect 400956 580932 401008 580984
rect 401048 580932 401100 580984
rect 428924 580932 428976 580984
rect 429844 580932 429896 580984
rect 456800 580932 456852 580984
rect 457076 580932 457128 580984
rect 484952 580932 485004 580984
rect 485044 580932 485096 580984
rect 512920 580932 512972 580984
rect 513104 580932 513156 580984
rect 540612 580932 540664 580984
rect 541072 580932 541124 580984
rect 568948 580932 569000 580984
rect 26608 580864 26660 580916
rect 38108 580864 38160 580916
rect 44640 580864 44692 580916
rect 65892 580864 65944 580916
rect 82636 580864 82688 580916
rect 93124 580864 93176 580916
rect 128636 580864 128688 580916
rect 149796 580864 149848 580916
rect 166632 580864 166684 580916
rect 177120 580864 177172 580916
rect 194600 580864 194652 580916
rect 211160 580864 211212 580916
rect 222936 580864 222988 580916
rect 234068 580864 234120 580916
rect 240324 580864 240376 580916
rect 261484 580864 261536 580916
rect 278596 580864 278648 580916
rect 289728 580864 289780 580916
rect 306932 580864 306984 580916
rect 318064 580864 318116 580916
rect 324320 580864 324372 580916
rect 345756 580864 345808 580916
rect 362868 580864 362920 580916
rect 373172 580864 373224 580916
rect 390652 580864 390704 580916
rect 407120 580864 407172 580916
rect 418620 580864 418672 580916
rect 429936 580864 429988 580916
rect 436652 580864 436704 580916
rect 457444 580864 457496 580916
rect 474648 580864 474700 580916
rect 485136 580864 485188 580916
rect 502616 580864 502668 580916
rect 514024 580864 514076 580916
rect 520648 580864 520700 580916
rect 541624 580864 541676 580916
rect 54852 580796 54904 580848
rect 71780 580796 71832 580848
rect 138940 580796 138992 580848
rect 149888 580796 149940 580848
rect 250628 580796 250680 580848
rect 267740 580796 267792 580848
rect 334624 580796 334676 580848
rect 345664 580796 345716 580848
rect 446956 580796 447008 580848
rect 463700 580796 463752 580848
rect 530952 580796 531004 580848
rect 547972 580796 548024 580848
rect 558644 580252 558696 580304
rect 568764 580252 568816 580304
rect 548340 578892 548392 578944
rect 569040 578892 569092 578944
rect 100024 578348 100076 578400
rect 121000 578348 121052 578400
rect 184020 578348 184072 578400
rect 204904 578348 204956 578400
rect 36912 578280 36964 578332
rect 53932 578280 53984 578332
rect 65892 578280 65944 578332
rect 81992 578280 82044 578332
rect 92848 578280 92900 578332
rect 110328 578280 110380 578332
rect 176752 578280 176804 578332
rect 194324 578280 194376 578332
rect 261484 578280 261536 578332
rect 278320 578280 278372 578332
rect 288900 578280 288952 578332
rect 306012 578280 306064 578332
rect 316776 578280 316828 578332
rect 333980 578280 334032 578332
rect 372896 578280 372948 578332
rect 390008 578280 390060 578332
rect 400772 578280 400824 578332
rect 418344 578280 418396 578332
rect 457444 578280 457496 578332
rect 474004 578280 474056 578332
rect 484860 578280 484912 578332
rect 502340 578280 502392 578332
rect 15292 578212 15344 578264
rect 26332 578212 26384 578264
rect 39304 578212 39356 578264
rect 64236 578212 64288 578264
rect 72332 578212 72384 578264
rect 93124 578212 93176 578264
rect 121092 578212 121144 578264
rect 138020 578212 138072 578264
rect 156328 578212 156380 578264
rect 177304 578212 177356 578264
rect 204812 578212 204864 578264
rect 222200 578212 222252 578264
rect 232780 578212 232832 578264
rect 250076 578212 250128 578264
rect 268016 578212 268068 578264
rect 289084 578212 289136 578264
rect 316868 578212 316920 578264
rect 344284 578212 344336 578264
rect 352012 578212 352064 578264
rect 373264 578212 373316 578264
rect 380348 578212 380400 578264
rect 400864 578212 400916 578264
rect 429844 578212 429896 578264
rect 456616 578212 456668 578264
rect 464344 578212 464396 578264
rect 485044 578212 485096 578264
rect 512736 578212 512788 578264
rect 530308 578212 530360 578264
rect 176752 576376 176804 576428
rect 232780 576376 232832 576428
rect 316776 576376 316828 576428
rect 316868 576376 316920 576428
rect 400772 576376 400824 576428
rect 400864 576376 400916 576428
rect 512736 576376 512788 576428
rect 568764 576376 568816 576428
rect 120724 576240 120776 576292
rect 121092 576240 121144 576292
rect 204720 576240 204772 576292
rect 204996 576240 205048 576292
rect 176752 576172 176804 576224
rect 232780 576172 232832 576224
rect 316776 576172 316828 576224
rect 316868 576172 316920 576224
rect 400772 576172 400824 576224
rect 400864 576172 400916 576224
rect 512736 576172 512788 576224
rect 568764 576172 568816 576224
rect 36820 571208 36872 571260
rect 37004 571208 37056 571260
rect 120908 567944 120960 567996
rect 120908 567740 120960 567792
rect 120816 565088 120868 565140
rect 121000 565088 121052 565140
rect 64880 562300 64932 562352
rect 65892 562300 65944 562352
rect 289084 560192 289136 560244
rect 295708 560192 295760 560244
rect 93124 559512 93176 559564
rect 99748 559512 99800 559564
rect 120816 559512 120868 559564
rect 127716 559512 127768 559564
rect 177304 559512 177356 559564
rect 183744 559512 183796 559564
rect 373264 559512 373316 559564
rect 379704 559512 379756 559564
rect 400864 559512 400916 559564
rect 407764 559512 407816 559564
rect 204904 558900 204956 558952
rect 211712 558900 211764 558952
rect 485044 558900 485096 558952
rect 491668 558900 491720 558952
rect 42708 557472 42760 557524
rect 95240 557472 95292 557524
rect 97908 557472 97960 557524
rect 150440 557472 150492 557524
rect 154488 557472 154540 557524
rect 207020 557472 207072 557524
rect 209688 557472 209740 557524
rect 262220 557472 262272 557524
rect 266268 557472 266320 557524
rect 318800 557472 318852 557524
rect 322848 557472 322900 557524
rect 375380 557472 375432 557524
rect 378048 557472 378100 557524
rect 430580 557472 430632 557524
rect 434628 557472 434680 557524
rect 487160 557472 487212 557524
rect 489828 557472 489880 557524
rect 542360 557472 542412 557524
rect 288808 556792 288860 556844
rect 288992 556792 289044 556844
rect 372804 556792 372856 556844
rect 372988 556792 373040 556844
rect 484768 556792 484820 556844
rect 484952 556792 485004 556844
rect 87420 556588 87472 556640
rect 92756 556588 92808 556640
rect 547880 556112 547932 556164
rect 548156 556112 548208 556164
rect 15384 554684 15436 554736
rect 43996 554684 44048 554736
rect 138296 554684 138348 554736
rect 176844 554684 176896 554736
rect 194324 554684 194376 554736
rect 232872 554684 232924 554736
rect 238852 554684 238904 554736
rect 26332 554616 26384 554668
rect 39304 554616 39356 554668
rect 42892 554616 42944 554668
rect 71780 554616 71832 554668
rect 110328 554616 110380 554668
rect 148784 554616 148836 554668
rect 166632 554616 166684 554668
rect 204996 554616 205048 554668
rect 211252 554616 211304 554668
rect 240048 554616 240100 554668
rect 295432 554684 295484 554736
rect 324044 554684 324096 554736
rect 334348 554684 334400 554736
rect 372988 554684 373040 554736
rect 390468 554684 390520 554736
rect 428740 554684 428792 554736
rect 434812 554684 434864 554736
rect 268016 554616 268068 554668
rect 278320 554616 278372 554668
rect 316960 554616 317012 554668
rect 323032 554616 323084 554668
rect 352012 554616 352064 554668
rect 362316 554616 362368 554668
rect 400956 554616 401008 554668
rect 407212 554616 407264 554668
rect 436008 554616 436060 554668
rect 491392 554684 491444 554736
rect 520004 554684 520056 554736
rect 530308 554684 530360 554736
rect 568856 554684 568908 554736
rect 463700 554616 463752 554668
rect 474648 554616 474700 554668
rect 512828 554616 512880 554668
rect 548156 554616 548208 554668
rect 558000 554616 558052 554668
rect 82636 554548 82688 554600
rect 120908 554548 120960 554600
rect 127072 554548 127124 554600
rect 156052 554548 156104 554600
rect 250352 554548 250404 554600
rect 288992 554548 289044 554600
rect 306288 554548 306340 554600
rect 316868 554548 316920 554600
rect 418344 554548 418396 554600
rect 429844 554548 429896 554600
rect 446312 554548 446364 554600
rect 484952 554548 485004 554600
rect 502340 554548 502392 554600
rect 540796 554548 540848 554600
rect 54300 554480 54352 554532
rect 87420 554480 87472 554532
rect 518992 554480 519044 554532
rect 547880 554480 547932 554532
rect 3608 553392 3660 553444
rect 10324 553392 10376 553444
rect 15292 553324 15344 553376
rect 16028 553324 16080 553376
rect 26608 552644 26660 552696
rect 36820 552644 36872 552696
rect 15568 552168 15620 552220
rect 54300 552168 54352 552220
rect 429844 552168 429896 552220
rect 436100 552168 436152 552220
rect 71780 552100 71832 552152
rect 110604 552100 110656 552152
rect 149888 552100 149940 552152
rect 156328 552100 156380 552152
rect 211160 552100 211212 552152
rect 250628 552100 250680 552152
rect 261484 552100 261536 552152
rect 278596 552100 278648 552152
rect 295340 552100 295392 552152
rect 334624 552100 334676 552152
rect 345756 552100 345808 552152
rect 362316 552100 362368 552152
rect 407120 552100 407172 552152
rect 446312 552100 446364 552152
rect 457444 552100 457496 552152
rect 474648 552100 474700 552152
rect 491300 552100 491352 552152
rect 530308 552100 530360 552152
rect 38016 552032 38068 552084
rect 44180 552032 44232 552084
rect 65892 552032 65944 552084
rect 82636 552032 82688 552084
rect 99380 552032 99432 552084
rect 138296 552032 138348 552084
rect 149796 552032 149848 552084
rect 166632 552032 166684 552084
rect 183560 552032 183612 552084
rect 222292 552032 222344 552084
rect 267740 552032 267792 552084
rect 306472 552032 306524 552084
rect 318064 552032 318116 552084
rect 324320 552032 324372 552084
rect 345848 552032 345900 552084
rect 352012 552032 352064 552084
rect 379520 552032 379572 552084
rect 418620 552032 418672 552084
rect 463700 552032 463752 552084
rect 502616 552032 502668 552084
rect 541624 552032 541676 552084
rect 558644 552032 558696 552084
rect 233976 550536 234028 550588
rect 240140 550536 240192 550588
rect 514024 550536 514076 550588
rect 520280 550536 520332 550588
rect 205088 549312 205140 549364
rect 429108 549244 429160 549296
rect 429936 549244 429988 549296
rect 205088 549108 205140 549160
rect 37280 548496 37332 548548
rect 38108 548496 38160 548548
rect 233240 548496 233292 548548
rect 234068 548496 234120 548548
rect 71780 533604 71832 533656
rect 72056 533604 72108 533656
rect 99380 533604 99432 533656
rect 99932 533604 99984 533656
rect 183560 533604 183612 533656
rect 184020 533604 184072 533656
rect 211160 533604 211212 533656
rect 211988 533604 212040 533656
rect 267740 533604 267792 533656
rect 268016 533604 268068 533656
rect 295340 533604 295392 533656
rect 295984 533604 296036 533656
rect 379520 533604 379572 533656
rect 379980 533604 380032 533656
rect 407120 533604 407172 533656
rect 407948 533604 408000 533656
rect 463700 533604 463752 533656
rect 464068 533604 464120 533656
rect 491300 531904 491352 531956
rect 492036 531904 492088 531956
rect 2964 527144 3016 527196
rect 6184 527144 6236 527196
rect 15200 527076 15252 527128
rect 36912 527076 36964 527128
rect 38108 527076 38160 527128
rect 64880 527076 64932 527128
rect 65064 527076 65116 527128
rect 92940 527076 92992 527128
rect 93032 527076 93084 527128
rect 120908 527076 120960 527128
rect 121092 527076 121144 527128
rect 148600 527076 148652 527128
rect 149704 527076 149756 527128
rect 176936 527076 176988 527128
rect 177028 527076 177080 527128
rect 204904 527076 204956 527128
rect 205180 527076 205232 527128
rect 232596 527076 232648 527128
rect 234068 527076 234120 527128
rect 260932 527076 260984 527128
rect 261024 527076 261076 527128
rect 288900 527076 288952 527128
rect 289084 527076 289136 527128
rect 316592 527076 316644 527128
rect 317052 527076 317104 527128
rect 344928 527076 344980 527128
rect 345664 527076 345716 527128
rect 372620 527076 372672 527128
rect 373080 527076 373132 527128
rect 400956 527076 401008 527128
rect 401048 527076 401100 527128
rect 428924 527076 428976 527128
rect 429936 527076 429988 527128
rect 456800 527076 456852 527128
rect 457076 527076 457128 527128
rect 484952 527076 485004 527128
rect 485044 527076 485096 527128
rect 512920 527076 512972 527128
rect 513104 527076 513156 527128
rect 540612 527076 540664 527128
rect 541072 527076 541124 527128
rect 568948 527076 569000 527128
rect 26608 527008 26660 527060
rect 38016 527008 38068 527060
rect 44640 527008 44692 527060
rect 65892 527008 65944 527060
rect 82636 527008 82688 527060
rect 99472 527008 99524 527060
rect 128636 527008 128688 527060
rect 149796 527008 149848 527060
rect 166632 527008 166684 527060
rect 183652 527008 183704 527060
rect 194600 527008 194652 527060
rect 211252 527008 211304 527060
rect 222936 527008 222988 527060
rect 233976 527008 234028 527060
rect 240324 527008 240376 527060
rect 261484 527008 261536 527060
rect 278596 527008 278648 527060
rect 295432 527008 295484 527060
rect 306932 527008 306984 527060
rect 318064 527008 318116 527060
rect 324320 527008 324372 527060
rect 345756 527008 345808 527060
rect 362868 527008 362920 527060
rect 379612 527008 379664 527060
rect 390652 527008 390704 527060
rect 407212 527008 407264 527060
rect 418620 527008 418672 527060
rect 429844 527008 429896 527060
rect 436652 527008 436704 527060
rect 457444 527008 457496 527060
rect 474648 527008 474700 527060
rect 491392 527008 491444 527060
rect 502616 527008 502668 527060
rect 514024 527008 514076 527060
rect 520648 527008 520700 527060
rect 541624 527008 541676 527060
rect 54944 526940 54996 526992
rect 71872 526940 71924 526992
rect 138940 526940 138992 526992
rect 149888 526940 149940 526992
rect 250628 526940 250680 526992
rect 267832 526940 267884 526992
rect 334624 526940 334676 526992
rect 345848 526940 345900 526992
rect 446956 526940 447008 526992
rect 463792 526940 463844 526992
rect 530952 526940 531004 526992
rect 547972 526940 548024 526992
rect 558644 526396 558696 526448
rect 568948 526396 569000 526448
rect 548340 525036 548392 525088
rect 569040 525036 569092 525088
rect 184020 524560 184072 524612
rect 204904 524560 204956 524612
rect 464344 524560 464396 524612
rect 485044 524560 485096 524612
rect 37096 524492 37148 524544
rect 54300 524492 54352 524544
rect 65892 524492 65944 524544
rect 81992 524492 82044 524544
rect 92848 524492 92900 524544
rect 110328 524492 110380 524544
rect 121000 524492 121052 524544
rect 138296 524492 138348 524544
rect 177028 524492 177080 524544
rect 194324 524492 194376 524544
rect 261484 524492 261536 524544
rect 278320 524492 278372 524544
rect 288992 524492 289044 524544
rect 306012 524492 306064 524544
rect 317144 524492 317196 524544
rect 334348 524492 334400 524544
rect 372988 524492 373040 524544
rect 390008 524492 390060 524544
rect 401048 524492 401100 524544
rect 418344 524492 418396 524544
rect 457444 524492 457496 524544
rect 474004 524492 474056 524544
rect 15292 524424 15344 524476
rect 26332 524424 26384 524476
rect 38016 524424 38068 524476
rect 64604 524424 64656 524476
rect 72332 524424 72384 524476
rect 93124 524424 93176 524476
rect 100024 524424 100076 524476
rect 121092 524424 121144 524476
rect 156328 524424 156380 524476
rect 177304 524424 177356 524476
rect 204812 524424 204864 524476
rect 222200 524424 222252 524476
rect 232964 524424 233016 524476
rect 250352 524424 250404 524476
rect 268016 524424 268068 524476
rect 289084 524424 289136 524476
rect 317052 524424 317104 524476
rect 344652 524424 344704 524476
rect 352012 524424 352064 524476
rect 373264 524424 373316 524476
rect 380348 524424 380400 524476
rect 401140 524424 401192 524476
rect 429844 524424 429896 524476
rect 456616 524424 456668 524476
rect 484860 524424 484912 524476
rect 502340 524424 502392 524476
rect 514484 524424 514536 524476
rect 530308 524424 530360 524476
rect 36728 522248 36780 522300
rect 37096 522248 37148 522300
rect 120724 522248 120776 522300
rect 121000 522248 121052 522300
rect 204720 522248 204772 522300
rect 204996 522248 205048 522300
rect 512736 522248 512788 522300
rect 514484 522248 514536 522300
rect 568856 522248 568908 522300
rect 120816 522180 120868 522232
rect 121092 522180 121144 522232
rect 400864 522180 400916 522232
rect 401140 522180 401192 522232
rect 568856 522044 568908 522096
rect 176844 521976 176896 522028
rect 177028 521976 177080 522028
rect 316776 521704 316828 521756
rect 317144 521704 317196 521756
rect 372804 521704 372856 521756
rect 372988 521704 373040 521756
rect 400772 521704 400824 521756
rect 401048 521704 401100 521756
rect 232780 521636 232832 521688
rect 232964 521636 233016 521688
rect 316868 521636 316920 521688
rect 317052 521636 317104 521688
rect 288900 519664 288952 519716
rect 288900 519460 288952 519512
rect 154488 518848 154540 518900
rect 155868 518848 155920 518900
rect 462228 518848 462280 518900
rect 463884 518848 463936 518900
rect 92756 507152 92808 507204
rect 92940 507152 92992 507204
rect 204904 505928 204956 505980
rect 211712 505928 211764 505980
rect 93124 505724 93176 505776
rect 99748 505724 99800 505776
rect 120816 505724 120868 505776
rect 127716 505724 127768 505776
rect 177304 505724 177356 505776
rect 183652 505724 183704 505776
rect 373264 505724 373316 505776
rect 379704 505724 379756 505776
rect 400864 505724 400916 505776
rect 407764 505724 407816 505776
rect 289084 505588 289136 505640
rect 295708 505588 295760 505640
rect 485044 505520 485096 505572
rect 491668 505520 491720 505572
rect 64880 503208 64932 503260
rect 65892 503208 65944 503260
rect 484768 502800 484820 502852
rect 484952 502800 485004 502852
rect 547880 502664 547932 502716
rect 548156 502664 548208 502716
rect 15384 500896 15436 500948
rect 43996 500896 44048 500948
rect 138296 500896 138348 500948
rect 176844 500896 176896 500948
rect 194324 500896 194376 500948
rect 232872 500896 232924 500948
rect 238852 500896 238904 500948
rect 26332 500828 26384 500880
rect 38016 500828 38068 500880
rect 42892 500828 42944 500880
rect 71780 500828 71832 500880
rect 110328 500828 110380 500880
rect 148784 500828 148836 500880
rect 166632 500828 166684 500880
rect 204996 500828 205048 500880
rect 211252 500828 211304 500880
rect 240048 500828 240100 500880
rect 295432 500896 295484 500948
rect 324044 500896 324096 500948
rect 334348 500896 334400 500948
rect 372896 500896 372948 500948
rect 390468 500896 390520 500948
rect 428740 500896 428792 500948
rect 434812 500896 434864 500948
rect 268016 500828 268068 500880
rect 278320 500828 278372 500880
rect 316960 500828 317012 500880
rect 323032 500828 323084 500880
rect 352012 500828 352064 500880
rect 362316 500828 362368 500880
rect 400956 500828 401008 500880
rect 407212 500828 407264 500880
rect 436008 500828 436060 500880
rect 491392 500896 491444 500948
rect 520004 500896 520056 500948
rect 530308 500896 530360 500948
rect 568856 500896 568908 500948
rect 463700 500828 463752 500880
rect 474648 500828 474700 500880
rect 512828 500828 512880 500880
rect 548156 500828 548208 500880
rect 558000 500828 558052 500880
rect 82636 500760 82688 500812
rect 120908 500760 120960 500812
rect 127072 500760 127124 500812
rect 156052 500760 156104 500812
rect 250352 500760 250404 500812
rect 288900 500760 288952 500812
rect 306288 500760 306340 500812
rect 316868 500760 316920 500812
rect 418344 500760 418396 500812
rect 429844 500760 429896 500812
rect 446312 500760 446364 500812
rect 484952 500760 485004 500812
rect 502340 500760 502392 500812
rect 540796 500760 540848 500812
rect 54300 500692 54352 500744
rect 92940 500692 92992 500744
rect 518992 500692 519044 500744
rect 547880 500692 547932 500744
rect 26608 498788 26660 498840
rect 36820 498788 36872 498840
rect 15936 498312 15988 498364
rect 54300 498312 54352 498364
rect 65892 498244 65944 498296
rect 82636 498244 82688 498296
rect 99380 498244 99432 498296
rect 138296 498244 138348 498296
rect 149704 498244 149756 498296
rect 156328 498244 156380 498296
rect 211160 498244 211212 498296
rect 250628 498244 250680 498296
rect 267740 498244 267792 498296
rect 306472 498244 306524 498296
rect 318064 498244 318116 498296
rect 324320 498244 324372 498296
rect 345848 498244 345900 498296
rect 362316 498244 362368 498296
rect 407120 498244 407172 498296
rect 446312 498244 446364 498296
rect 457444 498244 457496 498296
rect 474648 498244 474700 498296
rect 491300 498244 491352 498296
rect 530308 498244 530360 498296
rect 38108 498176 38160 498228
rect 44180 498176 44232 498228
rect 71780 498176 71832 498228
rect 110604 498176 110656 498228
rect 149888 498176 149940 498228
rect 166632 498176 166684 498228
rect 183560 498176 183612 498228
rect 222292 498176 222344 498228
rect 234068 498176 234120 498228
rect 240324 498176 240376 498228
rect 261484 498176 261536 498228
rect 278596 498176 278648 498228
rect 295340 498176 295392 498228
rect 334624 498176 334676 498228
rect 345756 498176 345808 498228
rect 352012 498176 352064 498228
rect 379520 498176 379572 498228
rect 418620 498176 418672 498228
rect 429936 498176 429988 498228
rect 436100 498176 436152 498228
rect 463700 498176 463752 498228
rect 502616 498176 502668 498228
rect 514024 498176 514076 498228
rect 520280 498176 520332 498228
rect 541624 498176 541676 498228
rect 558644 498176 558696 498228
rect 15292 497360 15344 497412
rect 16028 497360 16080 497412
rect 205088 495320 205140 495372
rect 429108 495184 429160 495236
rect 429844 495184 429896 495236
rect 205088 495116 205140 495168
rect 37280 492532 37332 492584
rect 38016 492532 38068 492584
rect 149244 492532 149296 492584
rect 149796 492532 149848 492584
rect 233240 492532 233292 492584
rect 233976 492532 234028 492584
rect 463700 485052 463752 485104
rect 463976 485052 464028 485104
rect 99380 477640 99432 477692
rect 99932 477640 99984 477692
rect 183560 477640 183612 477692
rect 184020 477640 184072 477692
rect 211160 477640 211212 477692
rect 211988 477640 212040 477692
rect 267740 477640 267792 477692
rect 268016 477640 268068 477692
rect 295340 477640 295392 477692
rect 295984 477640 296036 477692
rect 379520 477640 379572 477692
rect 379980 477640 380032 477692
rect 407120 477640 407172 477692
rect 407948 477640 408000 477692
rect 491300 477640 491352 477692
rect 492036 477640 492088 477692
rect 71780 475668 71832 475720
rect 72056 475668 72108 475720
rect 15200 473288 15252 473340
rect 36912 473288 36964 473340
rect 38016 473288 38068 473340
rect 64880 473288 64932 473340
rect 65064 473288 65116 473340
rect 92940 473288 92992 473340
rect 93032 473288 93084 473340
rect 120908 473288 120960 473340
rect 121092 473288 121144 473340
rect 148600 473288 148652 473340
rect 149796 473288 149848 473340
rect 176936 473288 176988 473340
rect 177028 473288 177080 473340
rect 204904 473288 204956 473340
rect 205180 473288 205232 473340
rect 232596 473288 232648 473340
rect 233976 473288 234028 473340
rect 260932 473288 260984 473340
rect 261024 473288 261076 473340
rect 288900 473288 288952 473340
rect 289084 473288 289136 473340
rect 316592 473288 316644 473340
rect 317052 473288 317104 473340
rect 344928 473288 344980 473340
rect 345664 473288 345716 473340
rect 372620 473288 372672 473340
rect 373080 473288 373132 473340
rect 400956 473288 401008 473340
rect 401048 473288 401100 473340
rect 428924 473288 428976 473340
rect 429844 473288 429896 473340
rect 456800 473288 456852 473340
rect 457076 473288 457128 473340
rect 484952 473288 485004 473340
rect 485044 473288 485096 473340
rect 512920 473288 512972 473340
rect 513104 473288 513156 473340
rect 540612 473288 540664 473340
rect 541072 473288 541124 473340
rect 568948 473288 569000 473340
rect 26608 473220 26660 473272
rect 38108 473220 38160 473272
rect 44640 473220 44692 473272
rect 65892 473220 65944 473272
rect 82636 473220 82688 473272
rect 99472 473220 99524 473272
rect 128636 473220 128688 473272
rect 149888 473220 149940 473272
rect 166632 473220 166684 473272
rect 183652 473220 183704 473272
rect 194600 473220 194652 473272
rect 211252 473220 211304 473272
rect 222936 473220 222988 473272
rect 234068 473220 234120 473272
rect 240324 473220 240376 473272
rect 261484 473220 261536 473272
rect 278596 473220 278648 473272
rect 295432 473220 295484 473272
rect 306932 473220 306984 473272
rect 318064 473220 318116 473272
rect 324320 473220 324372 473272
rect 345848 473220 345900 473272
rect 362868 473220 362920 473272
rect 379612 473220 379664 473272
rect 390652 473220 390704 473272
rect 407212 473220 407264 473272
rect 418620 473220 418672 473272
rect 429936 473220 429988 473272
rect 436652 473220 436704 473272
rect 457444 473220 457496 473272
rect 474648 473220 474700 473272
rect 491392 473220 491444 473272
rect 502616 473220 502668 473272
rect 514024 473220 514076 473272
rect 520648 473220 520700 473272
rect 541624 473220 541676 473272
rect 54944 473152 54996 473204
rect 71872 473152 71924 473204
rect 138940 473152 138992 473204
rect 149704 473152 149756 473204
rect 250628 473152 250680 473204
rect 267924 473152 267976 473204
rect 334624 473152 334676 473204
rect 345756 473152 345808 473204
rect 446956 473152 447008 473204
rect 463792 473152 463844 473204
rect 530952 473152 531004 473204
rect 547972 473152 548024 473204
rect 558644 472608 558696 472660
rect 568764 472608 568816 472660
rect 548340 471248 548392 471300
rect 569040 471248 569092 471300
rect 100024 470772 100076 470824
rect 120816 470772 120868 470824
rect 184020 470772 184072 470824
rect 204904 470772 204956 470824
rect 268016 470772 268068 470824
rect 289084 470772 289136 470824
rect 380348 470772 380400 470824
rect 400864 470772 400916 470824
rect 464344 470772 464396 470824
rect 485044 470772 485096 470824
rect 92848 470704 92900 470756
rect 110328 470704 110380 470756
rect 176844 470704 176896 470756
rect 194324 470704 194376 470756
rect 261576 470704 261628 470756
rect 278320 470704 278372 470756
rect 372896 470704 372948 470756
rect 390008 470704 390060 470756
rect 457536 470704 457588 470756
rect 474004 470704 474056 470756
rect 72332 470636 72384 470688
rect 93124 470636 93176 470688
rect 120724 470636 120776 470688
rect 138296 470636 138348 470688
rect 156328 470636 156380 470688
rect 177304 470636 177356 470688
rect 204812 470636 204864 470688
rect 222292 470636 222344 470688
rect 232780 470636 232832 470688
rect 250352 470636 250404 470688
rect 288900 470636 288952 470688
rect 306012 470636 306064 470688
rect 316776 470636 316828 470688
rect 334348 470636 334400 470688
rect 352012 470636 352064 470688
rect 373264 470636 373316 470688
rect 400772 470636 400824 470688
rect 418344 470636 418396 470688
rect 484860 470636 484912 470688
rect 502340 470636 502392 470688
rect 512736 470636 512788 470688
rect 530308 470636 530360 470688
rect 15292 470568 15344 470620
rect 26332 470568 26384 470620
rect 36728 470568 36780 470620
rect 54300 470568 54352 470620
rect 69664 470568 69716 470620
rect 579988 470568 580040 470620
rect 36728 468392 36780 468444
rect 120724 468392 120776 468444
rect 120816 468392 120868 468444
rect 232780 468392 232832 468444
rect 316776 468392 316828 468444
rect 400772 468392 400824 468444
rect 400864 468392 400916 468444
rect 512736 468392 512788 468444
rect 568764 468392 568816 468444
rect 204720 468256 204772 468308
rect 204996 468256 205048 468308
rect 36728 468188 36780 468240
rect 120724 468188 120776 468240
rect 120816 468188 120868 468240
rect 232780 468188 232832 468240
rect 316776 468188 316828 468240
rect 400772 468188 400824 468240
rect 400864 468188 400916 468240
rect 512736 468188 512788 468240
rect 568764 468188 568816 468240
rect 289084 452548 289136 452600
rect 295708 452548 295760 452600
rect 92756 451936 92808 451988
rect 92940 451936 92992 451988
rect 93124 451868 93176 451920
rect 99748 451868 99800 451920
rect 120816 451868 120868 451920
rect 127716 451868 127768 451920
rect 177304 451868 177356 451920
rect 183744 451868 183796 451920
rect 373264 451868 373316 451920
rect 379704 451868 379756 451920
rect 400864 451868 400916 451920
rect 407764 451868 407816 451920
rect 204904 451256 204956 451308
rect 211712 451256 211764 451308
rect 485044 451256 485096 451308
rect 491668 451256 491720 451308
rect 2780 448808 2832 448860
rect 4988 448808 5040 448860
rect 176752 448808 176804 448860
rect 176936 448808 176988 448860
rect 288808 448808 288860 448860
rect 288992 448808 289044 448860
rect 372804 448808 372856 448860
rect 372988 448808 373040 448860
rect 484768 448808 484820 448860
rect 484952 448808 485004 448860
rect 547880 448400 547932 448452
rect 548156 448400 548208 448452
rect 15292 448128 15344 448180
rect 16120 448128 16172 448180
rect 15476 445680 15528 445732
rect 43996 445680 44048 445732
rect 54300 445680 54352 445732
rect 92940 445680 92992 445732
rect 110328 445680 110380 445732
rect 148784 445680 148836 445732
rect 194324 445680 194376 445732
rect 232872 445680 232924 445732
rect 238852 445680 238904 445732
rect 26332 445612 26384 445664
rect 64788 445612 64840 445664
rect 82636 445612 82688 445664
rect 120908 445612 120960 445664
rect 138296 445612 138348 445664
rect 176936 445612 176988 445664
rect 211252 445612 211304 445664
rect 240048 445612 240100 445664
rect 295432 445680 295484 445732
rect 324044 445680 324096 445732
rect 334348 445680 334400 445732
rect 372988 445680 373040 445732
rect 390468 445680 390520 445732
rect 428740 445680 428792 445732
rect 434812 445680 434864 445732
rect 268016 445612 268068 445664
rect 306288 445612 306340 445664
rect 344744 445612 344796 445664
rect 362316 445612 362368 445664
rect 400956 445612 401008 445664
rect 407212 445612 407264 445664
rect 436008 445612 436060 445664
rect 491392 445680 491444 445732
rect 520004 445680 520056 445732
rect 530308 445680 530360 445732
rect 568856 445680 568908 445732
rect 463700 445612 463752 445664
rect 474648 445612 474700 445664
rect 512828 445612 512880 445664
rect 518992 445612 519044 445664
rect 547880 445612 547932 445664
rect 42892 445544 42944 445596
rect 71780 445544 71832 445596
rect 127072 445544 127124 445596
rect 156052 445544 156104 445596
rect 166632 445544 166684 445596
rect 204996 445544 205048 445596
rect 278320 445544 278372 445596
rect 316868 445544 316920 445596
rect 323032 445544 323084 445596
rect 352012 445544 352064 445596
rect 446312 445544 446364 445596
rect 484952 445544 485004 445596
rect 502340 445544 502392 445596
rect 540796 445544 540848 445596
rect 548156 445544 548208 445596
rect 558000 445544 558052 445596
rect 250352 445476 250404 445528
rect 288992 445476 289044 445528
rect 26608 445000 26660 445052
rect 36820 445000 36872 445052
rect 15384 444456 15436 444508
rect 54300 444456 54352 444508
rect 65892 444456 65944 444508
rect 82636 444456 82688 444508
rect 99472 444456 99524 444508
rect 138296 444456 138348 444508
rect 149888 444456 149940 444508
rect 156328 444456 156380 444508
rect 211160 444456 211212 444508
rect 250628 444456 250680 444508
rect 261484 444456 261536 444508
rect 278596 444456 278648 444508
rect 295432 444456 295484 444508
rect 334624 444456 334676 444508
rect 345848 444456 345900 444508
rect 362316 444456 362368 444508
rect 407120 444456 407172 444508
rect 446312 444456 446364 444508
rect 457444 444456 457496 444508
rect 474648 444456 474700 444508
rect 491392 444456 491444 444508
rect 530308 444456 530360 444508
rect 71872 444388 71924 444440
rect 110604 444388 110656 444440
rect 149796 444388 149848 444440
rect 166632 444388 166684 444440
rect 183652 444388 183704 444440
rect 222292 444388 222344 444440
rect 267832 444388 267884 444440
rect 306472 444388 306524 444440
rect 318064 444388 318116 444440
rect 324320 444388 324372 444440
rect 345664 444388 345716 444440
rect 352012 444388 352064 444440
rect 379612 444388 379664 444440
rect 418620 444388 418672 444440
rect 463792 444388 463844 444440
rect 502616 444388 502668 444440
rect 514024 444388 514076 444440
rect 520280 444388 520332 444440
rect 541624 444388 541676 444440
rect 558644 444388 558696 444440
rect 429108 441600 429160 441652
rect 429844 441600 429896 441652
rect 205088 441328 205140 441380
rect 345020 441192 345072 441244
rect 345756 441192 345808 441244
rect 205088 441124 205140 441176
rect 93124 439492 93176 439544
rect 99932 439492 99984 439544
rect 177304 439492 177356 439544
rect 184020 439492 184072 439544
rect 373264 439492 373316 439544
rect 379980 439492 380032 439544
rect 457536 439492 457588 439544
rect 464068 439492 464120 439544
rect 37096 438880 37148 438932
rect 44180 438880 44232 438932
rect 65984 438880 66036 438932
rect 71964 438880 72016 438932
rect 261576 438880 261628 438932
rect 267924 438880 267976 438932
rect 289176 438880 289228 438932
rect 295984 438880 296036 438932
rect 485136 438880 485188 438932
rect 492036 438880 492088 438932
rect 37280 436568 37332 436620
rect 38016 436568 38068 436620
rect 233240 436568 233292 436620
rect 233976 436568 234028 436620
rect 211160 427116 211212 427168
rect 211988 427116 212040 427168
rect 407120 427116 407172 427168
rect 407948 427116 408000 427168
rect 15200 419432 15252 419484
rect 36912 419432 36964 419484
rect 38016 419432 38068 419484
rect 64880 419432 64932 419484
rect 65064 419432 65116 419484
rect 92940 419432 92992 419484
rect 93032 419432 93084 419484
rect 120908 419432 120960 419484
rect 121092 419432 121144 419484
rect 148600 419432 148652 419484
rect 149704 419432 149756 419484
rect 176936 419432 176988 419484
rect 177028 419432 177080 419484
rect 204904 419432 204956 419484
rect 205180 419432 205232 419484
rect 232596 419432 232648 419484
rect 233976 419432 234028 419484
rect 260932 419432 260984 419484
rect 261024 419432 261076 419484
rect 288900 419432 288952 419484
rect 289084 419432 289136 419484
rect 316592 419432 316644 419484
rect 317052 419432 317104 419484
rect 344928 419432 344980 419484
rect 345756 419432 345808 419484
rect 372620 419432 372672 419484
rect 373080 419432 373132 419484
rect 400956 419432 401008 419484
rect 401048 419432 401100 419484
rect 428924 419432 428976 419484
rect 429844 419432 429896 419484
rect 456800 419432 456852 419484
rect 457076 419432 457128 419484
rect 484952 419432 485004 419484
rect 485044 419432 485096 419484
rect 512920 419432 512972 419484
rect 513104 419432 513156 419484
rect 540612 419432 540664 419484
rect 541072 419432 541124 419484
rect 568948 419432 569000 419484
rect 26608 419364 26660 419416
rect 37096 419364 37148 419416
rect 44640 419364 44692 419416
rect 65892 419364 65944 419416
rect 82636 419364 82688 419416
rect 93124 419364 93176 419416
rect 128636 419364 128688 419416
rect 149796 419364 149848 419416
rect 166632 419364 166684 419416
rect 177304 419364 177356 419416
rect 194600 419364 194652 419416
rect 211252 419364 211304 419416
rect 222936 419364 222988 419416
rect 240140 419364 240192 419416
rect 240324 419364 240376 419416
rect 261484 419364 261536 419416
rect 278596 419364 278648 419416
rect 289176 419364 289228 419416
rect 306932 419364 306984 419416
rect 318064 419364 318116 419416
rect 324320 419364 324372 419416
rect 345848 419364 345900 419416
rect 362868 419364 362920 419416
rect 373264 419364 373316 419416
rect 390652 419364 390704 419416
rect 407212 419364 407264 419416
rect 418620 419364 418672 419416
rect 436100 419364 436152 419416
rect 436652 419364 436704 419416
rect 457444 419364 457496 419416
rect 474648 419364 474700 419416
rect 485136 419364 485188 419416
rect 502616 419364 502668 419416
rect 514024 419364 514076 419416
rect 520648 419364 520700 419416
rect 541624 419364 541676 419416
rect 54944 419296 54996 419348
rect 65984 419296 66036 419348
rect 138940 419296 138992 419348
rect 149888 419296 149940 419348
rect 250628 419296 250680 419348
rect 261576 419296 261628 419348
rect 334624 419296 334676 419348
rect 345664 419296 345716 419348
rect 446956 419296 447008 419348
rect 457536 419296 457588 419348
rect 530952 419296 531004 419348
rect 547972 419296 548024 419348
rect 558644 418752 558696 418804
rect 568948 418752 569000 418804
rect 548340 417392 548392 417444
rect 569040 417392 569092 417444
rect 100024 416916 100076 416968
rect 121092 416916 121144 416968
rect 268016 416916 268068 416968
rect 289084 416916 289136 416968
rect 380348 416916 380400 416968
rect 401140 416916 401192 416968
rect 464344 416916 464396 416968
rect 485044 416916 485096 416968
rect 92848 416848 92900 416900
rect 110328 416848 110380 416900
rect 176844 416848 176896 416900
rect 194324 416848 194376 416900
rect 204812 416848 204864 416900
rect 222200 416848 222252 416900
rect 261484 416848 261536 416900
rect 278320 416848 278372 416900
rect 372896 416848 372948 416900
rect 390008 416848 390060 416900
rect 457444 416848 457496 416900
rect 474004 416848 474056 416900
rect 15292 416780 15344 416832
rect 26332 416780 26384 416832
rect 36912 416780 36964 416832
rect 54300 416780 54352 416832
rect 72332 416780 72384 416832
rect 93124 416780 93176 416832
rect 121000 416780 121052 416832
rect 138296 416780 138348 416832
rect 156328 416780 156380 416832
rect 177304 416780 177356 416832
rect 184020 416780 184072 416832
rect 204904 416780 204956 416832
rect 232964 416780 233016 416832
rect 250352 416780 250404 416832
rect 288900 416780 288952 416832
rect 306012 416780 306064 416832
rect 316960 416780 317012 416832
rect 334348 416780 334400 416832
rect 352012 416780 352064 416832
rect 373264 416780 373316 416832
rect 401048 416780 401100 416832
rect 418344 416780 418396 416832
rect 484860 416780 484912 416832
rect 502340 416780 502392 416832
rect 512920 416780 512972 416832
rect 530308 416780 530360 416832
rect 120724 414264 120776 414316
rect 121000 414264 121052 414316
rect 232780 414264 232832 414316
rect 232964 414264 233016 414316
rect 400772 414264 400824 414316
rect 401048 414264 401100 414316
rect 36728 414196 36780 414248
rect 36912 414196 36964 414248
rect 120816 414196 120868 414248
rect 121092 414196 121144 414248
rect 204720 414196 204772 414248
rect 204996 414196 205048 414248
rect 400864 414196 400916 414248
rect 401140 414196 401192 414248
rect 512736 412836 512788 412888
rect 512920 412836 512972 412888
rect 36820 412768 36872 412820
rect 316868 412768 316920 412820
rect 512828 412768 512880 412820
rect 36820 412564 36872 412616
rect 316868 412564 316920 412616
rect 512828 412564 512880 412616
rect 568764 410864 568816 410916
rect 568948 410864 569000 410916
rect 3148 410184 3200 410236
rect 8944 410184 8996 410236
rect 316776 408688 316828 408740
rect 316960 408688 317012 408740
rect 3332 397468 3384 397520
rect 11796 397468 11848 397520
rect 204904 397400 204956 397452
rect 211712 397400 211764 397452
rect 485044 397400 485096 397452
rect 491668 397400 491720 397452
rect 93124 396720 93176 396772
rect 99748 396720 99800 396772
rect 120816 396720 120868 396772
rect 127716 396720 127768 396772
rect 177304 396720 177356 396772
rect 183652 396720 183704 396772
rect 373264 396720 373316 396772
rect 379704 396720 379756 396772
rect 400864 396720 400916 396772
rect 407764 396720 407816 396772
rect 289084 396448 289136 396500
rect 295708 396448 295760 396500
rect 92756 394816 92808 394868
rect 176752 394816 176804 394868
rect 288808 394816 288860 394868
rect 372804 394816 372856 394868
rect 484768 394816 484820 394868
rect 15292 394680 15344 394732
rect 16120 394680 16172 394732
rect 547880 394680 547932 394732
rect 548156 394680 548208 394732
rect 92756 394612 92808 394664
rect 176752 394612 176804 394664
rect 288808 394612 288860 394664
rect 372804 394612 372856 394664
rect 484768 394612 484820 394664
rect 15384 391892 15436 391944
rect 43996 391892 44048 391944
rect 54300 391892 54352 391944
rect 92756 391892 92808 391944
rect 138296 391892 138348 391944
rect 176752 391892 176804 391944
rect 194324 391892 194376 391944
rect 232872 391892 232924 391944
rect 238852 391892 238904 391944
rect 26332 391824 26384 391876
rect 64788 391824 64840 391876
rect 82636 391824 82688 391876
rect 120908 391824 120960 391876
rect 127072 391824 127124 391876
rect 155960 391824 156012 391876
rect 166632 391824 166684 391876
rect 204996 391824 205048 391876
rect 211252 391824 211304 391876
rect 240048 391824 240100 391876
rect 295432 391892 295484 391944
rect 324044 391892 324096 391944
rect 334348 391892 334400 391944
rect 372804 391892 372856 391944
rect 390468 391892 390520 391944
rect 428740 391892 428792 391944
rect 434812 391892 434864 391944
rect 268016 391824 268068 391876
rect 306288 391824 306340 391876
rect 344744 391824 344796 391876
rect 362316 391824 362368 391876
rect 400956 391824 401008 391876
rect 407212 391824 407264 391876
rect 436008 391824 436060 391876
rect 491392 391892 491444 391944
rect 520004 391892 520056 391944
rect 530308 391892 530360 391944
rect 568856 391892 568908 391944
rect 463792 391824 463844 391876
rect 474648 391824 474700 391876
rect 512828 391824 512880 391876
rect 548156 391824 548208 391876
rect 558000 391824 558052 391876
rect 42892 391756 42944 391808
rect 71780 391756 71832 391808
rect 110328 391756 110380 391808
rect 148784 391756 148836 391808
rect 278320 391756 278372 391808
rect 316868 391756 316920 391808
rect 323032 391756 323084 391808
rect 352012 391756 352064 391808
rect 446312 391756 446364 391808
rect 484768 391756 484820 391808
rect 502340 391756 502392 391808
rect 540796 391756 540848 391808
rect 250352 391688 250404 391740
rect 288808 391688 288860 391740
rect 518992 391688 519044 391740
rect 547880 391688 547932 391740
rect 26608 389784 26660 389836
rect 36820 389784 36872 389836
rect 15384 389308 15436 389360
rect 54300 389308 54352 389360
rect 65892 389240 65944 389292
rect 82636 389240 82688 389292
rect 99472 389240 99524 389292
rect 138296 389240 138348 389292
rect 149704 389240 149756 389292
rect 156328 389240 156380 389292
rect 211252 389240 211304 389292
rect 250628 389240 250680 389292
rect 261484 389240 261536 389292
rect 278596 389240 278648 389292
rect 295432 389240 295484 389292
rect 334624 389240 334676 389292
rect 345756 389240 345808 389292
rect 362316 389240 362368 389292
rect 407212 389240 407264 389292
rect 446312 389240 446364 389292
rect 457444 389240 457496 389292
rect 474648 389240 474700 389292
rect 491392 389240 491444 389292
rect 530308 389240 530360 389292
rect 38016 389172 38068 389224
rect 44180 389172 44232 389224
rect 71780 389172 71832 389224
rect 110604 389172 110656 389224
rect 149796 389172 149848 389224
rect 166632 389172 166684 389224
rect 183560 389172 183612 389224
rect 222292 389172 222344 389224
rect 233976 389172 234028 389224
rect 240324 389172 240376 389224
rect 267832 389172 267884 389224
rect 306472 389172 306524 389224
rect 318064 389172 318116 389224
rect 324320 389172 324372 389224
rect 345664 389172 345716 389224
rect 352012 389172 352064 389224
rect 379612 389172 379664 389224
rect 418620 389172 418672 389224
rect 429844 389172 429896 389224
rect 436100 389172 436152 389224
rect 463700 389172 463752 389224
rect 502616 389172 502668 389224
rect 514024 389172 514076 389224
rect 520280 389172 520332 389224
rect 541624 389172 541676 389224
rect 558644 389172 558696 389224
rect 205088 387336 205140 387388
rect 345020 387200 345072 387252
rect 345848 387200 345900 387252
rect 205088 387132 205140 387184
rect 429108 386384 429160 386436
rect 429936 386384 429988 386436
rect 37280 385432 37332 385484
rect 38108 385432 38160 385484
rect 99380 385432 99432 385484
rect 99932 385432 99984 385484
rect 149244 385432 149296 385484
rect 149888 385432 149940 385484
rect 211160 385432 211212 385484
rect 211988 385432 212040 385484
rect 233240 385432 233292 385484
rect 234068 385432 234120 385484
rect 295340 385432 295392 385484
rect 295984 385432 296036 385484
rect 379520 385432 379572 385484
rect 379980 385432 380032 385484
rect 407120 385432 407172 385484
rect 407948 385432 408000 385484
rect 491300 385432 491352 385484
rect 492036 385432 492088 385484
rect 267740 384752 267792 384804
rect 267924 384752 267976 384804
rect 463700 378768 463752 378820
rect 463976 378768 464028 378820
rect 569224 378156 569276 378208
rect 579804 378156 579856 378208
rect 183560 370540 183612 370592
rect 184020 370540 184072 370592
rect 42708 368432 42760 368484
rect 95240 368432 95292 368484
rect 97908 368432 97960 368484
rect 150440 368432 150492 368484
rect 154488 368432 154540 368484
rect 207020 368432 207072 368484
rect 209688 368432 209740 368484
rect 262220 368432 262272 368484
rect 266268 368432 266320 368484
rect 318800 368432 318852 368484
rect 322848 368432 322900 368484
rect 375380 368432 375432 368484
rect 378048 368432 378100 368484
rect 430580 368432 430632 368484
rect 434628 368432 434680 368484
rect 487160 368432 487212 368484
rect 489828 368432 489880 368484
rect 542360 368432 542412 368484
rect 71780 367684 71832 367736
rect 72056 367684 72108 367736
rect 15200 365644 15252 365696
rect 36912 365644 36964 365696
rect 38108 365644 38160 365696
rect 64880 365644 64932 365696
rect 65064 365644 65116 365696
rect 92940 365644 92992 365696
rect 93032 365644 93084 365696
rect 120908 365644 120960 365696
rect 121092 365644 121144 365696
rect 148600 365644 148652 365696
rect 149888 365644 149940 365696
rect 176936 365644 176988 365696
rect 177028 365644 177080 365696
rect 204904 365644 204956 365696
rect 205180 365644 205232 365696
rect 232596 365644 232648 365696
rect 234068 365644 234120 365696
rect 260932 365644 260984 365696
rect 261024 365644 261076 365696
rect 288900 365644 288952 365696
rect 289084 365644 289136 365696
rect 316592 365644 316644 365696
rect 317052 365644 317104 365696
rect 344928 365644 344980 365696
rect 345848 365644 345900 365696
rect 372620 365644 372672 365696
rect 373080 365644 373132 365696
rect 400956 365644 401008 365696
rect 401048 365644 401100 365696
rect 428924 365644 428976 365696
rect 429936 365644 429988 365696
rect 456800 365644 456852 365696
rect 457076 365644 457128 365696
rect 484952 365644 485004 365696
rect 485044 365644 485096 365696
rect 512920 365644 512972 365696
rect 513104 365644 513156 365696
rect 540612 365644 540664 365696
rect 541072 365644 541124 365696
rect 568948 365644 569000 365696
rect 26608 365576 26660 365628
rect 38016 365576 38068 365628
rect 44640 365576 44692 365628
rect 65892 365576 65944 365628
rect 82636 365576 82688 365628
rect 99380 365576 99432 365628
rect 128636 365576 128688 365628
rect 149796 365576 149848 365628
rect 166632 365576 166684 365628
rect 183652 365576 183704 365628
rect 194600 365576 194652 365628
rect 211160 365576 211212 365628
rect 222936 365576 222988 365628
rect 233976 365576 234028 365628
rect 240324 365576 240376 365628
rect 261484 365576 261536 365628
rect 278596 365576 278648 365628
rect 295340 365576 295392 365628
rect 306932 365576 306984 365628
rect 318064 365576 318116 365628
rect 324320 365576 324372 365628
rect 345756 365576 345808 365628
rect 362868 365576 362920 365628
rect 379520 365576 379572 365628
rect 390652 365576 390704 365628
rect 407120 365576 407172 365628
rect 418620 365576 418672 365628
rect 429844 365576 429896 365628
rect 436652 365576 436704 365628
rect 457444 365576 457496 365628
rect 474648 365576 474700 365628
rect 491300 365576 491352 365628
rect 502616 365576 502668 365628
rect 514024 365576 514076 365628
rect 520648 365576 520700 365628
rect 541624 365576 541676 365628
rect 54944 365508 54996 365560
rect 71872 365508 71924 365560
rect 138940 365508 138992 365560
rect 149704 365508 149756 365560
rect 250628 365508 250680 365560
rect 267740 365508 267792 365560
rect 334624 365508 334676 365560
rect 345664 365508 345716 365560
rect 446956 365508 447008 365560
rect 463792 365508 463844 365560
rect 530952 365508 531004 365560
rect 547972 365508 548024 365560
rect 558644 364964 558696 365016
rect 568764 364964 568816 365016
rect 548340 363604 548392 363656
rect 569040 363604 569092 363656
rect 100024 363060 100076 363112
rect 121092 363060 121144 363112
rect 184020 363060 184072 363112
rect 204904 363060 204956 363112
rect 464344 363060 464396 363112
rect 485044 363060 485096 363112
rect 36912 362992 36964 363044
rect 54300 362992 54352 363044
rect 65892 362992 65944 363044
rect 81992 362992 82044 363044
rect 92848 362992 92900 363044
rect 110328 362992 110380 363044
rect 176844 362992 176896 363044
rect 194324 362992 194376 363044
rect 261484 362992 261536 363044
rect 278320 362992 278372 363044
rect 288900 362992 288952 363044
rect 306012 362992 306064 363044
rect 317144 362992 317196 363044
rect 334348 362992 334400 363044
rect 372896 362992 372948 363044
rect 390008 362992 390060 363044
rect 401048 362992 401100 363044
rect 418344 362992 418396 363044
rect 457444 362992 457496 363044
rect 474004 362992 474056 363044
rect 15292 362924 15344 362976
rect 26332 362924 26384 362976
rect 38016 362924 38068 362976
rect 64604 362924 64656 362976
rect 72332 362924 72384 362976
rect 93124 362924 93176 362976
rect 121000 362924 121052 362976
rect 138296 362924 138348 362976
rect 156328 362924 156380 362976
rect 177304 362924 177356 362976
rect 204812 362924 204864 362976
rect 222200 362924 222252 362976
rect 232964 362924 233016 362976
rect 250352 362924 250404 362976
rect 268016 362924 268068 362976
rect 289084 362924 289136 362976
rect 317052 362924 317104 362976
rect 344652 362924 344704 362976
rect 352012 362924 352064 362976
rect 373264 362924 373316 362976
rect 380348 362924 380400 362976
rect 401140 362924 401192 362976
rect 429844 362924 429896 362976
rect 456616 362924 456668 362976
rect 484952 362924 485004 362976
rect 502340 362924 502392 362976
rect 512920 362924 512972 362976
rect 530308 362924 530360 362976
rect 568764 360408 568816 360460
rect 120724 360204 120776 360256
rect 121000 360204 121052 360256
rect 204720 360204 204772 360256
rect 204996 360204 205048 360256
rect 400864 360204 400916 360256
rect 401140 360204 401192 360256
rect 568764 360204 568816 360256
rect 120816 360136 120868 360188
rect 121092 360136 121144 360188
rect 316776 358844 316828 358896
rect 317144 358844 317196 358896
rect 400772 358844 400824 358896
rect 401048 358844 401100 358896
rect 232780 358776 232832 358828
rect 232964 358776 233016 358828
rect 316868 358776 316920 358828
rect 317052 358776 317104 358828
rect 36820 355376 36872 355428
rect 37004 355376 37056 355428
rect 484860 355376 484912 355428
rect 512828 355376 512880 355428
rect 513012 355376 513064 355428
rect 484860 355172 484912 355224
rect 484768 352248 484820 352300
rect 484952 352248 485004 352300
rect 36820 347760 36872 347812
rect 37004 347760 37056 347812
rect 512828 347760 512880 347812
rect 513012 347760 513064 347812
rect 92756 345652 92808 345704
rect 92940 345652 92992 345704
rect 372804 345652 372856 345704
rect 372988 345652 373040 345704
rect 2780 345176 2832 345228
rect 5080 345176 5132 345228
rect 64880 342864 64932 342916
rect 65892 342864 65944 342916
rect 93124 342864 93176 342916
rect 99748 342864 99800 342916
rect 120816 342864 120868 342916
rect 127716 342864 127768 342916
rect 177304 342864 177356 342916
rect 183652 342864 183704 342916
rect 373264 342864 373316 342916
rect 379704 342864 379756 342916
rect 400864 342864 400916 342916
rect 407764 342864 407816 342916
rect 204904 342592 204956 342644
rect 211712 342592 211764 342644
rect 485044 342592 485096 342644
rect 491668 342592 491720 342644
rect 289084 342524 289136 342576
rect 295708 342524 295760 342576
rect 288808 340892 288860 340944
rect 288992 340892 289044 340944
rect 176752 340824 176804 340876
rect 176936 340824 176988 340876
rect 547880 340688 547932 340740
rect 548156 340688 548208 340740
rect 15292 340144 15344 340196
rect 15936 339940 15988 339992
rect 15384 338036 15436 338088
rect 43996 338036 44048 338088
rect 138296 338036 138348 338088
rect 176936 338036 176988 338088
rect 194324 338036 194376 338088
rect 232872 338036 232924 338088
rect 238852 338036 238904 338088
rect 26332 337968 26384 338020
rect 38016 337968 38068 338020
rect 42892 337968 42944 338020
rect 71780 337968 71832 338020
rect 110328 337968 110380 338020
rect 148784 337968 148836 338020
rect 166632 337968 166684 338020
rect 204996 337968 205048 338020
rect 211252 337968 211304 338020
rect 240048 337968 240100 338020
rect 295432 338036 295484 338088
rect 324044 338036 324096 338088
rect 334348 338036 334400 338088
rect 372988 338036 373040 338088
rect 390468 338036 390520 338088
rect 428740 338036 428792 338088
rect 434812 338036 434864 338088
rect 268016 337968 268068 338020
rect 278320 337968 278372 338020
rect 316960 337968 317012 338020
rect 323032 337968 323084 338020
rect 352012 337968 352064 338020
rect 362316 337968 362368 338020
rect 400956 337968 401008 338020
rect 407212 337968 407264 338020
rect 436008 337968 436060 338020
rect 491392 338036 491444 338088
rect 520004 338036 520056 338088
rect 530308 338036 530360 338088
rect 568856 338036 568908 338088
rect 463700 337968 463752 338020
rect 474648 337968 474700 338020
rect 512828 337968 512880 338020
rect 548156 337968 548208 338020
rect 558000 337968 558052 338020
rect 82636 337900 82688 337952
rect 120908 337900 120960 337952
rect 127072 337900 127124 337952
rect 156052 337900 156104 337952
rect 250352 337900 250404 337952
rect 288992 337900 289044 337952
rect 306288 337900 306340 337952
rect 316868 337900 316920 337952
rect 418344 337900 418396 337952
rect 429844 337900 429896 337952
rect 446312 337900 446364 337952
rect 484860 337900 484912 337952
rect 502340 337900 502392 337952
rect 540796 337900 540848 337952
rect 54300 337832 54352 337884
rect 92940 337832 92992 337884
rect 518992 337832 519044 337884
rect 547880 337832 547932 337884
rect 26608 335996 26660 336048
rect 36820 335996 36872 336048
rect 15384 335452 15436 335504
rect 54300 335452 54352 335504
rect 429844 335452 429896 335504
rect 436100 335452 436152 335504
rect 71780 335384 71832 335436
rect 110604 335384 110656 335436
rect 149704 335384 149756 335436
rect 156328 335384 156380 335436
rect 211160 335384 211212 335436
rect 250628 335384 250680 335436
rect 267832 335384 267884 335436
rect 306380 335384 306432 335436
rect 318064 335384 318116 335436
rect 324320 335384 324372 335436
rect 345756 335384 345808 335436
rect 362316 335384 362368 335436
rect 407212 335384 407264 335436
rect 446312 335384 446364 335436
rect 457444 335384 457496 335436
rect 474648 335384 474700 335436
rect 491392 335384 491444 335436
rect 530308 335384 530360 335436
rect 38016 335316 38068 335368
rect 44180 335316 44232 335368
rect 65892 335316 65944 335368
rect 82636 335316 82688 335368
rect 99380 335316 99432 335368
rect 138296 335316 138348 335368
rect 149888 335316 149940 335368
rect 166632 335316 166684 335368
rect 183560 335316 183612 335368
rect 222384 335316 222436 335368
rect 233976 335316 234028 335368
rect 240324 335316 240376 335368
rect 261484 335316 261536 335368
rect 278596 335316 278648 335368
rect 295432 335316 295484 335368
rect 334624 335316 334676 335368
rect 345664 335316 345716 335368
rect 352012 335316 352064 335368
rect 379612 335316 379664 335368
rect 418620 335316 418672 335368
rect 463792 335316 463844 335368
rect 502616 335316 502668 335368
rect 514024 335316 514076 335368
rect 520280 335316 520332 335368
rect 541624 335316 541676 335368
rect 558644 335316 558696 335368
rect 205088 333344 205140 333396
rect 345020 333208 345072 333260
rect 345848 333208 345900 333260
rect 205088 333140 205140 333192
rect 42708 332596 42760 332648
rect 95240 332596 95292 332648
rect 97908 332596 97960 332648
rect 150440 332596 150492 332648
rect 154488 332596 154540 332648
rect 207020 332596 207072 332648
rect 209688 332596 209740 332648
rect 262220 332596 262272 332648
rect 266268 332596 266320 332648
rect 318800 332596 318852 332648
rect 322848 332596 322900 332648
rect 375380 332596 375432 332648
rect 378048 332596 378100 332648
rect 430580 332664 430632 332716
rect 429108 332596 429160 332648
rect 429936 332596 429988 332648
rect 434628 332596 434680 332648
rect 487160 332596 487212 332648
rect 489828 332596 489880 332648
rect 542360 332596 542412 332648
rect 37280 329468 37332 329520
rect 38108 329468 38160 329520
rect 149244 329468 149296 329520
rect 149796 329468 149848 329520
rect 233240 329468 233292 329520
rect 234068 329468 234120 329520
rect 267740 329468 267792 329520
rect 267924 329468 267976 329520
rect 295340 329468 295392 329520
rect 295984 329468 296036 329520
rect 379520 329468 379572 329520
rect 379980 329468 380032 329520
rect 407120 329468 407172 329520
rect 407948 329468 408000 329520
rect 491300 329468 491352 329520
rect 492036 329468 492088 329520
rect 463700 325728 463752 325780
rect 464068 325728 464120 325780
rect 574744 324300 574796 324352
rect 580080 324300 580132 324352
rect 99380 314576 99432 314628
rect 99932 314576 99984 314628
rect 183560 314576 183612 314628
rect 184020 314576 184072 314628
rect 211160 314576 211212 314628
rect 211988 314576 212040 314628
rect 71780 313420 71832 313472
rect 72056 313420 72108 313472
rect 15200 311788 15252 311840
rect 36912 311788 36964 311840
rect 38108 311788 38160 311840
rect 64880 311788 64932 311840
rect 65064 311788 65116 311840
rect 92940 311788 92992 311840
rect 93032 311788 93084 311840
rect 120908 311788 120960 311840
rect 121092 311788 121144 311840
rect 148600 311788 148652 311840
rect 149796 311788 149848 311840
rect 176936 311788 176988 311840
rect 177028 311788 177080 311840
rect 204904 311788 204956 311840
rect 205180 311788 205232 311840
rect 232596 311788 232648 311840
rect 234068 311788 234120 311840
rect 260932 311788 260984 311840
rect 261024 311788 261076 311840
rect 288900 311788 288952 311840
rect 289084 311788 289136 311840
rect 316592 311788 316644 311840
rect 317052 311788 317104 311840
rect 344928 311788 344980 311840
rect 345848 311788 345900 311840
rect 372620 311788 372672 311840
rect 373080 311788 373132 311840
rect 400956 311788 401008 311840
rect 401048 311788 401100 311840
rect 428924 311788 428976 311840
rect 429936 311788 429988 311840
rect 456800 311788 456852 311840
rect 457076 311788 457128 311840
rect 484952 311788 485004 311840
rect 485044 311788 485096 311840
rect 512920 311788 512972 311840
rect 513104 311788 513156 311840
rect 540612 311788 540664 311840
rect 541072 311788 541124 311840
rect 568948 311788 569000 311840
rect 26608 311720 26660 311772
rect 38016 311720 38068 311772
rect 44640 311720 44692 311772
rect 65892 311720 65944 311772
rect 82636 311720 82688 311772
rect 99472 311720 99524 311772
rect 128636 311720 128688 311772
rect 149888 311720 149940 311772
rect 166632 311720 166684 311772
rect 183652 311720 183704 311772
rect 194600 311720 194652 311772
rect 211252 311720 211304 311772
rect 222936 311720 222988 311772
rect 233976 311720 234028 311772
rect 240324 311720 240376 311772
rect 261484 311720 261536 311772
rect 278596 311720 278648 311772
rect 295340 311720 295392 311772
rect 306932 311720 306984 311772
rect 318064 311720 318116 311772
rect 324320 311720 324372 311772
rect 345756 311720 345808 311772
rect 362868 311720 362920 311772
rect 379520 311720 379572 311772
rect 390652 311720 390704 311772
rect 407120 311720 407172 311772
rect 418620 311720 418672 311772
rect 429844 311720 429896 311772
rect 436652 311720 436704 311772
rect 457444 311720 457496 311772
rect 474648 311720 474700 311772
rect 491300 311720 491352 311772
rect 502616 311720 502668 311772
rect 514024 311720 514076 311772
rect 520648 311720 520700 311772
rect 541624 311720 541676 311772
rect 54944 311652 54996 311704
rect 72056 311652 72108 311704
rect 138940 311652 138992 311704
rect 149704 311652 149756 311704
rect 250628 311652 250680 311704
rect 267740 311652 267792 311704
rect 334624 311652 334676 311704
rect 345664 311652 345716 311704
rect 446956 311652 447008 311704
rect 463700 311652 463752 311704
rect 530952 311652 531004 311704
rect 547972 311652 548024 311704
rect 558644 311108 558696 311160
rect 568948 311108 569000 311160
rect 548340 309748 548392 309800
rect 569040 309748 569092 309800
rect 100024 309272 100076 309324
rect 121000 309272 121052 309324
rect 268016 309272 268068 309324
rect 289084 309272 289136 309324
rect 380348 309272 380400 309324
rect 401048 309272 401100 309324
rect 464344 309272 464396 309324
rect 485044 309272 485096 309324
rect 36912 309204 36964 309256
rect 54300 309204 54352 309256
rect 65892 309204 65944 309256
rect 81992 309204 82044 309256
rect 92940 309204 92992 309256
rect 110328 309204 110380 309256
rect 176936 309204 176988 309256
rect 194324 309204 194376 309256
rect 261484 309204 261536 309256
rect 278320 309204 278372 309256
rect 317144 309204 317196 309256
rect 334348 309204 334400 309256
rect 372804 309204 372856 309256
rect 390008 309204 390060 309256
rect 457444 309204 457496 309256
rect 474004 309204 474056 309256
rect 15200 309136 15252 309188
rect 26332 309136 26384 309188
rect 38016 309136 38068 309188
rect 64604 309136 64656 309188
rect 72332 309136 72384 309188
rect 93124 309136 93176 309188
rect 121092 309136 121144 309188
rect 138296 309136 138348 309188
rect 156328 309136 156380 309188
rect 177304 309136 177356 309188
rect 184020 309136 184072 309188
rect 204904 309136 204956 309188
rect 209044 309136 209096 309188
rect 222200 309136 222252 309188
rect 232964 309136 233016 309188
rect 250352 309136 250404 309188
rect 288808 309136 288860 309188
rect 306012 309136 306064 309188
rect 317052 309136 317104 309188
rect 344652 309136 344704 309188
rect 352012 309136 352064 309188
rect 373264 309136 373316 309188
rect 401140 309136 401192 309188
rect 418344 309136 418396 309188
rect 429844 309136 429896 309188
rect 456616 309136 456668 309188
rect 484952 309136 485004 309188
rect 502340 309136 502392 309188
rect 512920 309136 512972 309188
rect 530308 309136 530360 309188
rect 120724 306280 120776 306332
rect 121092 306280 121144 306332
rect 568856 306280 568908 306332
rect 36728 306212 36780 306264
rect 36912 306212 36964 306264
rect 120816 306212 120868 306264
rect 121000 306212 121052 306264
rect 288716 306212 288768 306264
rect 288900 306212 288952 306264
rect 568856 306076 568908 306128
rect 36820 305736 36872 305788
rect 484768 305736 484820 305788
rect 512736 305736 512788 305788
rect 316776 305668 316828 305720
rect 317144 305668 317196 305720
rect 400772 305668 400824 305720
rect 401140 305668 401192 305720
rect 36820 305532 36872 305584
rect 484860 305532 484912 305584
rect 512828 305532 512880 305584
rect 512736 304580 512788 304632
rect 512920 304580 512972 304632
rect 568764 304240 568816 304292
rect 568948 304240 569000 304292
rect 204812 303764 204864 303816
rect 204996 303764 205048 303816
rect 204812 303628 204864 303680
rect 209044 303628 209096 303680
rect 484768 302676 484820 302728
rect 484952 302676 485004 302728
rect 92756 301520 92808 301572
rect 92940 301520 92992 301572
rect 232780 301520 232832 301572
rect 232964 301520 233016 301572
rect 316868 301520 316920 301572
rect 317052 301520 317104 301572
rect 372804 301520 372856 301572
rect 372988 301520 373040 301572
rect 176844 297440 176896 297492
rect 400956 297440 401008 297492
rect 176844 297236 176896 297288
rect 400956 297236 401008 297288
rect 3148 292680 3200 292732
rect 6276 292680 6328 292732
rect 176752 292476 176804 292528
rect 176936 292476 176988 292528
rect 400864 292476 400916 292528
rect 401048 292476 401100 292528
rect 64880 291864 64932 291916
rect 65892 291864 65944 291916
rect 289084 289756 289136 289808
rect 295708 289756 295760 289808
rect 93124 289076 93176 289128
rect 99748 289076 99800 289128
rect 120816 289076 120868 289128
rect 127716 289076 127768 289128
rect 177304 289076 177356 289128
rect 183744 289076 183796 289128
rect 373264 289076 373316 289128
rect 379704 289076 379756 289128
rect 400864 289076 400916 289128
rect 407764 289076 407816 289128
rect 204904 288396 204956 288448
rect 211712 288396 211764 288448
rect 485044 288396 485096 288448
rect 491668 288396 491720 288448
rect 547880 286152 547932 286204
rect 548156 286152 548208 286204
rect 15384 284248 15436 284300
rect 43996 284248 44048 284300
rect 138296 284248 138348 284300
rect 176844 284248 176896 284300
rect 194324 284248 194376 284300
rect 232872 284248 232924 284300
rect 238852 284248 238904 284300
rect 26332 284180 26384 284232
rect 38016 284180 38068 284232
rect 42892 284180 42944 284232
rect 71780 284180 71832 284232
rect 110328 284180 110380 284232
rect 148784 284180 148836 284232
rect 166632 284180 166684 284232
rect 204996 284180 205048 284232
rect 211252 284180 211304 284232
rect 240048 284180 240100 284232
rect 295432 284248 295484 284300
rect 324044 284248 324096 284300
rect 334348 284248 334400 284300
rect 372896 284248 372948 284300
rect 390468 284248 390520 284300
rect 428740 284248 428792 284300
rect 434812 284248 434864 284300
rect 268016 284180 268068 284232
rect 278320 284180 278372 284232
rect 316960 284180 317012 284232
rect 323032 284180 323084 284232
rect 352012 284180 352064 284232
rect 362316 284180 362368 284232
rect 400956 284180 401008 284232
rect 407212 284180 407264 284232
rect 436008 284180 436060 284232
rect 491392 284248 491444 284300
rect 520004 284248 520056 284300
rect 530308 284248 530360 284300
rect 568856 284248 568908 284300
rect 463700 284180 463752 284232
rect 474648 284180 474700 284232
rect 512828 284180 512880 284232
rect 518992 284180 519044 284232
rect 547880 284180 547932 284232
rect 82636 284112 82688 284164
rect 120908 284112 120960 284164
rect 127072 284112 127124 284164
rect 156052 284112 156104 284164
rect 250352 284112 250404 284164
rect 288900 284112 288952 284164
rect 306288 284112 306340 284164
rect 316868 284112 316920 284164
rect 418344 284112 418396 284164
rect 429844 284112 429896 284164
rect 446312 284112 446364 284164
rect 484860 284112 484912 284164
rect 502340 284112 502392 284164
rect 540796 284112 540848 284164
rect 548156 284112 548208 284164
rect 558000 284112 558052 284164
rect 54300 284044 54352 284096
rect 92848 284044 92900 284096
rect 15200 283160 15252 283212
rect 16028 283160 16080 283212
rect 26608 282140 26660 282192
rect 36820 282140 36872 282192
rect 38016 281596 38068 281648
rect 44180 281596 44232 281648
rect 71872 281596 71924 281648
rect 110604 281596 110656 281648
rect 211252 281596 211304 281648
rect 250628 281596 250680 281648
rect 295432 281596 295484 281648
rect 334624 281596 334676 281648
rect 407212 281596 407264 281648
rect 446312 281596 446364 281648
rect 491392 281596 491444 281648
rect 530308 281596 530360 281648
rect 15384 281528 15436 281580
rect 54300 281528 54352 281580
rect 99472 281528 99524 281580
rect 138296 281528 138348 281580
rect 149704 281528 149756 281580
rect 166632 281528 166684 281580
rect 183652 281528 183704 281580
rect 222292 281528 222344 281580
rect 267832 281528 267884 281580
rect 306472 281528 306524 281580
rect 318064 281528 318116 281580
rect 324320 281528 324372 281580
rect 345756 281528 345808 281580
rect 362316 281528 362368 281580
rect 379612 281528 379664 281580
rect 418620 281528 418672 281580
rect 429936 281528 429988 281580
rect 436100 281528 436152 281580
rect 463792 281528 463844 281580
rect 502616 281528 502668 281580
rect 541624 281528 541676 281580
rect 558644 281528 558696 281580
rect 233976 280100 234028 280152
rect 240140 280100 240192 280152
rect 205088 279352 205140 279404
rect 205088 279148 205140 279200
rect 42708 278740 42760 278792
rect 95240 278740 95292 278792
rect 97908 278740 97960 278792
rect 150440 278740 150492 278792
rect 154488 278740 154540 278792
rect 207020 278740 207072 278792
rect 209688 278740 209740 278792
rect 262220 278740 262272 278792
rect 266268 278740 266320 278792
rect 318800 278740 318852 278792
rect 322848 278740 322900 278792
rect 375380 278740 375432 278792
rect 378048 278740 378100 278792
rect 430580 278740 430632 278792
rect 434628 278740 434680 278792
rect 487160 278740 487212 278792
rect 489828 278740 489880 278792
rect 542360 278740 542412 278792
rect 149244 278332 149296 278384
rect 149796 278332 149848 278384
rect 71780 272552 71832 272604
rect 71964 272552 72016 272604
rect 99380 272552 99432 272604
rect 99932 272552 99984 272604
rect 183560 272552 183612 272604
rect 184020 272552 184072 272604
rect 211160 272552 211212 272604
rect 211988 272552 212040 272604
rect 267740 272552 267792 272604
rect 267924 272552 267976 272604
rect 295340 272552 295392 272604
rect 295984 272552 296036 272604
rect 379520 272552 379572 272604
rect 379980 272552 380032 272604
rect 407120 272552 407172 272604
rect 407948 272552 408000 272604
rect 463700 272552 463752 272604
rect 464068 272552 464120 272604
rect 491300 272552 491352 272604
rect 492036 272552 492088 272604
rect 15292 256640 15344 256692
rect 36912 256640 36964 256692
rect 37096 256640 37148 256692
rect 64880 256640 64932 256692
rect 65064 256640 65116 256692
rect 92940 256640 92992 256692
rect 93032 256640 93084 256692
rect 120908 256640 120960 256692
rect 121092 256640 121144 256692
rect 148600 256640 148652 256692
rect 149796 256640 149848 256692
rect 176936 256640 176988 256692
rect 177028 256640 177080 256692
rect 204904 256640 204956 256692
rect 205180 256640 205232 256692
rect 232596 256640 232648 256692
rect 233056 256640 233108 256692
rect 260932 256640 260984 256692
rect 261024 256640 261076 256692
rect 288900 256640 288952 256692
rect 289084 256640 289136 256692
rect 316592 256640 316644 256692
rect 317052 256640 317104 256692
rect 344928 256640 344980 256692
rect 345664 256640 345716 256692
rect 372620 256640 372672 256692
rect 373080 256640 373132 256692
rect 400956 256640 401008 256692
rect 401048 256640 401100 256692
rect 428924 256640 428976 256692
rect 429108 256640 429160 256692
rect 456800 256640 456852 256692
rect 457076 256640 457128 256692
rect 484952 256640 485004 256692
rect 485044 256640 485096 256692
rect 512920 256640 512972 256692
rect 513104 256640 513156 256692
rect 540612 256640 540664 256692
rect 541072 256640 541124 256692
rect 568948 256640 569000 256692
rect 26608 256572 26660 256624
rect 38016 256572 38068 256624
rect 54944 256572 54996 256624
rect 71780 256572 71832 256624
rect 82636 256572 82688 256624
rect 99380 256572 99432 256624
rect 128636 256572 128688 256624
rect 149704 256572 149756 256624
rect 166632 256572 166684 256624
rect 183560 256572 183612 256624
rect 194600 256572 194652 256624
rect 211160 256572 211212 256624
rect 222936 256572 222988 256624
rect 233976 256572 234028 256624
rect 250628 256572 250680 256624
rect 267740 256572 267792 256624
rect 278596 256572 278648 256624
rect 295340 256572 295392 256624
rect 306932 256572 306984 256624
rect 318064 256572 318116 256624
rect 324320 256572 324372 256624
rect 345756 256572 345808 256624
rect 362868 256572 362920 256624
rect 379520 256572 379572 256624
rect 390652 256572 390704 256624
rect 407120 256572 407172 256624
rect 418620 256572 418672 256624
rect 429936 256572 429988 256624
rect 446956 256572 447008 256624
rect 463700 256572 463752 256624
rect 474648 256572 474700 256624
rect 491300 256572 491352 256624
rect 520648 256572 520700 256624
rect 541624 256572 541676 256624
rect 138940 256504 138992 256556
rect 155960 256504 156012 256556
rect 334624 256504 334676 256556
rect 351920 256504 351972 256556
rect 530952 256504 531004 256556
rect 547972 256504 548024 256556
rect 558644 256028 558696 256080
rect 568948 256028 569000 256080
rect 548340 255960 548392 256012
rect 569040 255960 569092 256012
rect 100024 255416 100076 255468
rect 121092 255416 121144 255468
rect 268016 255416 268068 255468
rect 289176 255416 289228 255468
rect 380348 255416 380400 255468
rect 401140 255416 401192 255468
rect 464344 255416 464396 255468
rect 485136 255416 485188 255468
rect 37648 255348 37700 255400
rect 54300 255348 54352 255400
rect 65892 255348 65944 255400
rect 81992 255348 82044 255400
rect 92940 255348 92992 255400
rect 110328 255348 110380 255400
rect 177028 255348 177080 255400
rect 194324 255348 194376 255400
rect 261484 255348 261536 255400
rect 278320 255348 278372 255400
rect 317144 255348 317196 255400
rect 334348 255348 334400 255400
rect 372988 255348 373040 255400
rect 390008 255348 390060 255400
rect 457444 255348 457496 255400
rect 474004 255348 474056 255400
rect 15200 255280 15252 255332
rect 26332 255280 26384 255332
rect 38108 255280 38160 255332
rect 64604 255280 64656 255332
rect 72332 255280 72384 255332
rect 93124 255280 93176 255332
rect 121000 255280 121052 255332
rect 138296 255280 138348 255332
rect 156328 255280 156380 255332
rect 177304 255280 177356 255332
rect 184020 255280 184072 255332
rect 204996 255280 205048 255332
rect 208400 255280 208452 255332
rect 222200 255280 222252 255332
rect 232964 255280 233016 255332
rect 250352 255280 250404 255332
rect 289084 255280 289136 255332
rect 306012 255280 306064 255332
rect 317052 255280 317104 255332
rect 344652 255280 344704 255332
rect 352012 255280 352064 255332
rect 373264 255280 373316 255332
rect 401048 255280 401100 255332
rect 418344 255280 418396 255332
rect 429844 255280 429896 255332
rect 456616 255280 456668 255332
rect 485044 255280 485096 255332
rect 502340 255280 502392 255332
rect 513104 255280 513156 255332
rect 530308 255280 530360 255332
rect 36728 252288 36780 252340
rect 37648 252288 37700 252340
rect 120724 252220 120776 252272
rect 121000 252220 121052 252272
rect 204720 252220 204772 252272
rect 204996 252220 205048 252272
rect 400864 252220 400916 252272
rect 401140 252220 401192 252272
rect 120816 252152 120868 252204
rect 121092 252152 121144 252204
rect 512736 252016 512788 252068
rect 513104 252016 513156 252068
rect 316776 251880 316828 251932
rect 317144 251880 317196 251932
rect 232780 251812 232832 251864
rect 232964 251812 233016 251864
rect 316868 251812 316920 251864
rect 317052 251812 317104 251864
rect 92756 251744 92808 251796
rect 92940 251744 92992 251796
rect 176752 251336 176804 251388
rect 177028 251336 177080 251388
rect 484768 251336 484820 251388
rect 485044 251336 485096 251388
rect 288808 251268 288860 251320
rect 289084 251268 289136 251320
rect 204812 250520 204864 250572
rect 208400 250520 208452 250572
rect 372804 250112 372856 250164
rect 372988 250112 373040 250164
rect 400772 249092 400824 249144
rect 401048 249092 401100 249144
rect 568764 249092 568816 249144
rect 568948 249092 569000 249144
rect 3240 240116 3292 240168
rect 14464 240116 14516 240168
rect 64880 235696 64932 235748
rect 65892 235696 65944 235748
rect 204904 235424 204956 235476
rect 211712 235424 211764 235476
rect 485136 235288 485188 235340
rect 491668 235288 491720 235340
rect 93124 235220 93176 235272
rect 99748 235220 99800 235272
rect 120816 235220 120868 235272
rect 127716 235220 127768 235272
rect 177304 235220 177356 235272
rect 183652 235220 183704 235272
rect 373264 235220 373316 235272
rect 379704 235220 379756 235272
rect 400864 235220 400916 235272
rect 407764 235220 407816 235272
rect 289176 235016 289228 235068
rect 295708 235016 295760 235068
rect 42708 233180 42760 233232
rect 95240 233180 95292 233232
rect 97908 233180 97960 233232
rect 150440 233180 150492 233232
rect 154488 233180 154540 233232
rect 207020 233180 207072 233232
rect 209688 233180 209740 233232
rect 262220 233180 262272 233232
rect 266268 233180 266320 233232
rect 318800 233180 318852 233232
rect 322848 233180 322900 233232
rect 375380 233180 375432 233232
rect 378048 233180 378100 233232
rect 430580 233180 430632 233232
rect 434628 233180 434680 233232
rect 487160 233180 487212 233232
rect 489828 233180 489880 233232
rect 542360 233180 542412 233232
rect 547880 232704 547932 232756
rect 548156 232704 548208 232756
rect 38016 231820 38068 231872
rect 580080 231820 580132 231872
rect 15384 230392 15436 230444
rect 43996 230392 44048 230444
rect 138296 230392 138348 230444
rect 176844 230392 176896 230444
rect 194324 230392 194376 230444
rect 232872 230392 232924 230444
rect 238852 230392 238904 230444
rect 26332 230324 26384 230376
rect 38108 230324 38160 230376
rect 42892 230324 42944 230376
rect 71780 230324 71832 230376
rect 110328 230324 110380 230376
rect 148784 230324 148836 230376
rect 166632 230324 166684 230376
rect 204996 230324 205048 230376
rect 211252 230324 211304 230376
rect 240048 230324 240100 230376
rect 295432 230392 295484 230444
rect 324044 230392 324096 230444
rect 334348 230392 334400 230444
rect 372896 230392 372948 230444
rect 390468 230392 390520 230444
rect 428740 230392 428792 230444
rect 434812 230392 434864 230444
rect 268016 230324 268068 230376
rect 278320 230324 278372 230376
rect 316960 230324 317012 230376
rect 323032 230324 323084 230376
rect 352012 230324 352064 230376
rect 362316 230324 362368 230376
rect 400956 230324 401008 230376
rect 407212 230324 407264 230376
rect 436008 230324 436060 230376
rect 491392 230392 491444 230444
rect 520004 230392 520056 230444
rect 530308 230392 530360 230444
rect 568856 230392 568908 230444
rect 463700 230324 463752 230376
rect 474648 230324 474700 230376
rect 512828 230324 512880 230376
rect 548156 230324 548208 230376
rect 558000 230324 558052 230376
rect 82636 230256 82688 230308
rect 120908 230256 120960 230308
rect 127072 230256 127124 230308
rect 156052 230256 156104 230308
rect 250352 230256 250404 230308
rect 288900 230256 288952 230308
rect 306288 230256 306340 230308
rect 316868 230256 316920 230308
rect 418344 230256 418396 230308
rect 429844 230256 429896 230308
rect 446312 230256 446364 230308
rect 484860 230256 484912 230308
rect 502340 230256 502392 230308
rect 540796 230256 540848 230308
rect 54300 230188 54352 230240
rect 92848 230188 92900 230240
rect 518992 230188 519044 230240
rect 547880 230188 547932 230240
rect 26608 228352 26660 228404
rect 36820 228352 36872 228404
rect 15936 227876 15988 227928
rect 54300 227876 54352 227928
rect 149704 227876 149756 227928
rect 166632 227876 166684 227928
rect 407856 227876 407908 227928
rect 446312 227876 446364 227928
rect 491944 227876 491996 227928
rect 65892 227808 65944 227860
rect 82636 227808 82688 227860
rect 99840 227808 99892 227860
rect 138296 227808 138348 227860
rect 149888 227808 149940 227860
rect 156328 227808 156380 227860
rect 211896 227808 211948 227860
rect 250628 227808 250680 227860
rect 261484 227808 261536 227860
rect 278596 227808 278648 227860
rect 295892 227808 295944 227860
rect 334624 227808 334676 227860
rect 379888 227808 379940 227860
rect 418620 227808 418672 227860
rect 429844 227808 429896 227860
rect 436100 227808 436152 227860
rect 458824 227808 458876 227860
rect 474648 227808 474700 227860
rect 486424 227808 486476 227860
rect 492312 227808 492364 227860
rect 530308 227808 530360 227860
rect 38108 227740 38160 227792
rect 44180 227740 44232 227792
rect 71872 227740 71924 227792
rect 110604 227740 110656 227792
rect 183928 227740 183980 227792
rect 222292 227740 222344 227792
rect 233976 227740 234028 227792
rect 240324 227740 240376 227792
rect 267832 227740 267884 227792
rect 306472 227740 306524 227792
rect 318064 227740 318116 227792
rect 324320 227740 324372 227792
rect 345664 227740 345716 227792
rect 362316 227740 362368 227792
rect 378876 227740 378928 227792
rect 390652 227740 390704 227792
rect 402244 227740 402296 227792
rect 408316 227740 408368 227792
rect 460204 227740 460256 227792
rect 464344 227740 464396 227792
rect 463976 227672 464028 227724
rect 502616 227740 502668 227792
rect 514024 227740 514076 227792
rect 520280 227740 520332 227792
rect 541624 227740 541676 227792
rect 558644 227740 558696 227792
rect 15200 227128 15252 227180
rect 16028 227128 16080 227180
rect 205088 225360 205140 225412
rect 345020 225224 345072 225276
rect 347044 225224 347096 225276
rect 205088 225156 205140 225208
rect 434628 225088 434680 225140
rect 487160 225088 487212 225140
rect 322848 225020 322900 225072
rect 375380 225020 375432 225072
rect 405648 225020 405700 225072
rect 458180 225020 458232 225072
rect 293868 224952 293920 225004
rect 346400 224952 346452 225004
rect 348424 224952 348476 225004
rect 352012 224952 352064 225004
rect 429108 224952 429160 225004
rect 429936 224952 429988 225004
rect 37280 222300 37332 222352
rect 38200 222300 38252 222352
rect 99380 222300 99432 222352
rect 99932 222300 99984 222352
rect 183560 222300 183612 222352
rect 184020 222300 184072 222352
rect 211160 222300 211212 222352
rect 211988 222300 212040 222352
rect 267740 222300 267792 222352
rect 267924 222300 267976 222352
rect 295340 222300 295392 222352
rect 295984 222300 296036 222352
rect 379520 222300 379572 222352
rect 379980 222300 380032 222352
rect 71780 221008 71832 221060
rect 71964 221008 72016 221060
rect 233240 220668 233292 220720
rect 234068 220668 234120 220720
rect 149244 220056 149296 220108
rect 149796 220056 149848 220108
rect 15292 202784 15344 202836
rect 36912 202784 36964 202836
rect 38200 202784 38252 202836
rect 64880 202784 64932 202836
rect 65064 202784 65116 202836
rect 92940 202784 92992 202836
rect 93032 202784 93084 202836
rect 120908 202784 120960 202836
rect 121092 202784 121144 202836
rect 148600 202784 148652 202836
rect 149796 202784 149848 202836
rect 176936 202784 176988 202836
rect 177028 202784 177080 202836
rect 204628 202784 204680 202836
rect 205180 202784 205232 202836
rect 232596 202784 232648 202836
rect 234068 202784 234120 202836
rect 260932 202784 260984 202836
rect 261024 202784 261076 202836
rect 288532 202784 288584 202836
rect 289084 202784 289136 202836
rect 316592 202784 316644 202836
rect 317052 202784 317104 202836
rect 344928 202784 344980 202836
rect 347044 202784 347096 202836
rect 372620 202784 372672 202836
rect 373080 202784 373132 202836
rect 400588 202784 400640 202836
rect 401048 202784 401100 202836
rect 428924 202784 428976 202836
rect 429936 202784 429988 202836
rect 456800 202784 456852 202836
rect 457076 202784 457128 202836
rect 484676 202784 484728 202836
rect 485044 202784 485096 202836
rect 512920 202784 512972 202836
rect 513104 202784 513156 202836
rect 540612 202784 540664 202836
rect 541072 202784 541124 202836
rect 568948 202784 569000 202836
rect 26608 202716 26660 202768
rect 38108 202716 38160 202768
rect 44640 202716 44692 202768
rect 65892 202716 65944 202768
rect 82636 202716 82688 202768
rect 99380 202716 99432 202768
rect 128636 202716 128688 202768
rect 149704 202716 149756 202768
rect 166632 202716 166684 202768
rect 183560 202716 183612 202768
rect 194968 202716 195020 202768
rect 211160 202716 211212 202768
rect 222936 202716 222988 202768
rect 233976 202716 234028 202768
rect 240324 202716 240376 202768
rect 261484 202716 261536 202768
rect 278504 202716 278556 202768
rect 295340 202716 295392 202768
rect 306932 202716 306984 202768
rect 318064 202716 318116 202768
rect 324320 202716 324372 202768
rect 345664 202716 345716 202768
rect 352656 202716 352708 202768
rect 378876 202716 378928 202768
rect 390928 202716 390980 202768
rect 402244 202716 402296 202768
rect 418620 202716 418672 202768
rect 429844 202716 429896 202768
rect 436652 202716 436704 202768
rect 458824 202716 458876 202768
rect 474464 202716 474516 202768
rect 486424 202716 486476 202768
rect 502616 202716 502668 202768
rect 514024 202716 514076 202768
rect 520648 202716 520700 202768
rect 541624 202716 541676 202768
rect 54852 202648 54904 202700
rect 71780 202648 71832 202700
rect 138940 202648 138992 202700
rect 149888 202648 149940 202700
rect 250628 202648 250680 202700
rect 267740 202648 267792 202700
rect 334624 202648 334676 202700
rect 348424 202648 348476 202700
rect 362868 202648 362920 202700
rect 379520 202648 379572 202700
rect 446956 202648 447008 202700
rect 460204 202648 460256 202700
rect 530952 202648 531004 202700
rect 547972 202648 548024 202700
rect 558644 202104 558696 202156
rect 568764 202104 568816 202156
rect 548340 200744 548392 200796
rect 569040 200744 569092 200796
rect 156328 200336 156380 200388
rect 177304 200336 177356 200388
rect 92756 200268 92808 200320
rect 110328 200268 110380 200320
rect 120724 200268 120776 200320
rect 138296 200268 138348 200320
rect 149704 200268 149756 200320
rect 165988 200268 166040 200320
rect 184020 200268 184072 200320
rect 204904 200268 204956 200320
rect 464344 200268 464396 200320
rect 485044 200268 485096 200320
rect 37004 200200 37056 200252
rect 54300 200200 54352 200252
rect 65892 200200 65944 200252
rect 81992 200200 82044 200252
rect 100024 200200 100076 200252
rect 120908 200200 120960 200252
rect 176752 200200 176804 200252
rect 194324 200200 194376 200252
rect 261484 200200 261536 200252
rect 278320 200200 278372 200252
rect 288900 200200 288952 200252
rect 306012 200200 306064 200252
rect 316776 200200 316828 200252
rect 334348 200200 334400 200252
rect 372896 200200 372948 200252
rect 390008 200200 390060 200252
rect 400772 200200 400824 200252
rect 418344 200200 418396 200252
rect 457444 200200 457496 200252
rect 474004 200200 474056 200252
rect 15200 200132 15252 200184
rect 26332 200132 26384 200184
rect 38108 200132 38160 200184
rect 64604 200132 64656 200184
rect 72332 200132 72384 200184
rect 93124 200132 93176 200184
rect 94504 200132 94556 200184
rect 120632 200132 120684 200184
rect 120816 200132 120868 200184
rect 148600 200132 148652 200184
rect 149796 200132 149848 200184
rect 176660 200132 176712 200184
rect 204812 200132 204864 200184
rect 222292 200132 222344 200184
rect 232780 200132 232832 200184
rect 250352 200132 250404 200184
rect 268016 200132 268068 200184
rect 289084 200132 289136 200184
rect 290464 200132 290516 200184
rect 316316 200132 316368 200184
rect 318064 200132 318116 200184
rect 344652 200132 344704 200184
rect 352012 200132 352064 200184
rect 373264 200132 373316 200184
rect 380348 200132 380400 200184
rect 400864 200132 400916 200184
rect 429844 200132 429896 200184
rect 456616 200132 456668 200184
rect 484860 200132 484912 200184
rect 502340 200132 502392 200184
rect 512736 200132 512788 200184
rect 530308 200132 530360 200184
rect 547144 200132 547196 200184
rect 558000 200132 558052 200184
rect 92756 198296 92808 198348
rect 232780 198296 232832 198348
rect 400772 198296 400824 198348
rect 400864 198296 400916 198348
rect 512736 198296 512788 198348
rect 568764 198296 568816 198348
rect 204720 198228 204772 198280
rect 204996 198228 205048 198280
rect 92756 198092 92808 198144
rect 232780 198092 232832 198144
rect 400772 198092 400824 198144
rect 400864 198092 400916 198144
rect 512736 198092 512788 198144
rect 568764 198092 568816 198144
rect 36820 195168 36872 195220
rect 37004 195168 37056 195220
rect 569316 191836 569368 191888
rect 580080 191836 580132 191888
rect 2780 187688 2832 187740
rect 5172 187688 5224 187740
rect 64880 185580 64932 185632
rect 65892 185580 65944 185632
rect 289084 182112 289136 182164
rect 295708 182112 295760 182164
rect 93124 181432 93176 181484
rect 99748 181432 99800 181484
rect 120908 181432 120960 181484
rect 127716 181432 127768 181484
rect 177304 181432 177356 181484
rect 183744 181432 183796 181484
rect 373264 181432 373316 181484
rect 379704 181432 379756 181484
rect 400864 181432 400916 181484
rect 407764 181432 407816 181484
rect 204904 180820 204956 180872
rect 211712 180820 211764 180872
rect 485044 180820 485096 180872
rect 491668 180820 491720 180872
rect 42708 179324 42760 179376
rect 95240 179324 95292 179376
rect 97908 179324 97960 179376
rect 150440 179324 150492 179376
rect 154488 179324 154540 179376
rect 207020 179324 207072 179376
rect 209688 179324 209740 179376
rect 262220 179324 262272 179376
rect 266268 179324 266320 179376
rect 318800 179324 318852 179376
rect 322848 179324 322900 179376
rect 375380 179324 375432 179376
rect 378048 179324 378100 179376
rect 430580 179324 430632 179376
rect 434628 179324 434680 179376
rect 487160 179324 487212 179376
rect 489828 179324 489880 179376
rect 542360 179324 542412 179376
rect 288808 178848 288860 178900
rect 288992 178848 289044 178900
rect 372804 178848 372856 178900
rect 372988 178848 373040 178900
rect 484768 178848 484820 178900
rect 484952 178848 485004 178900
rect 547880 178644 547932 178696
rect 548156 178644 548208 178696
rect 15384 176604 15436 176656
rect 43996 176604 44048 176656
rect 110328 176604 110380 176656
rect 120816 176604 120868 176656
rect 166632 176604 166684 176656
rect 204996 176604 205048 176656
rect 211252 176604 211304 176656
rect 240048 176604 240100 176656
rect 295432 176604 295484 176656
rect 324044 176604 324096 176656
rect 334348 176604 334400 176656
rect 372988 176604 373040 176656
rect 390468 176604 390520 176656
rect 428740 176604 428792 176656
rect 434812 176604 434864 176656
rect 26332 176536 26384 176588
rect 38108 176536 38160 176588
rect 42892 176536 42944 176588
rect 71780 176536 71832 176588
rect 82636 176536 82688 176588
rect 94504 176536 94556 176588
rect 138296 176536 138348 176588
rect 149796 176536 149848 176588
rect 194324 176536 194376 176588
rect 232872 176536 232924 176588
rect 238852 176536 238904 176588
rect 268016 176536 268068 176588
rect 278320 176536 278372 176588
rect 290464 176536 290516 176588
rect 306288 176536 306340 176588
rect 318064 176536 318116 176588
rect 323032 176536 323084 176588
rect 352012 176536 352064 176588
rect 362316 176536 362368 176588
rect 400956 176536 401008 176588
rect 407212 176536 407264 176588
rect 436008 176536 436060 176588
rect 491392 176604 491444 176656
rect 520004 176604 520056 176656
rect 530308 176604 530360 176656
rect 568856 176604 568908 176656
rect 463700 176536 463752 176588
rect 474648 176536 474700 176588
rect 512828 176536 512880 176588
rect 518992 176536 519044 176588
rect 547880 176536 547932 176588
rect 54300 176468 54352 176520
rect 92848 176468 92900 176520
rect 127072 176468 127124 176520
rect 156052 176468 156104 176520
rect 250352 176468 250404 176520
rect 288992 176468 289044 176520
rect 418344 176468 418396 176520
rect 429844 176468 429896 176520
rect 446312 176468 446364 176520
rect 484952 176468 485004 176520
rect 502340 176468 502392 176520
rect 540612 176468 540664 176520
rect 547144 176468 547196 176520
rect 548156 176468 548208 176520
rect 558000 176468 558052 176520
rect 540796 176400 540848 176452
rect 15200 175992 15252 176044
rect 16028 175992 16080 176044
rect 26608 174496 26660 174548
rect 36820 174496 36872 174548
rect 15384 174020 15436 174072
rect 54300 174020 54352 174072
rect 66904 174020 66956 174072
rect 82636 174020 82688 174072
rect 149704 174020 149756 174072
rect 166632 174020 166684 174072
rect 71872 173952 71924 174004
rect 110604 173952 110656 174004
rect 122104 173952 122156 174004
rect 128360 173952 128412 174004
rect 177304 173952 177356 174004
rect 194600 173952 194652 174004
rect 36912 173884 36964 173936
rect 43444 173884 43496 173936
rect 99380 173884 99432 173936
rect 138296 173884 138348 173936
rect 178684 173884 178736 173936
rect 184296 173884 184348 173936
rect 211252 174020 211304 174072
rect 183652 173816 183704 173868
rect 206284 173884 206336 173936
rect 209780 173884 209832 173936
rect 211988 173952 212040 174004
rect 374644 174020 374696 174072
rect 380348 174020 380400 174072
rect 407212 174020 407264 174072
rect 250628 173952 250680 174004
rect 262864 173952 262916 174004
rect 209964 173884 210016 173936
rect 222292 173884 222344 173936
rect 234068 173884 234120 173936
rect 240324 173884 240376 173936
rect 264244 173884 264296 173936
rect 267832 173952 267884 174004
rect 306472 173952 306524 174004
rect 318064 173952 318116 174004
rect 324320 173952 324372 174004
rect 345848 173952 345900 174004
rect 362316 173952 362368 174004
rect 373264 173952 373316 174004
rect 390652 173952 390704 174004
rect 402244 173952 402296 174004
rect 408316 173952 408368 174004
rect 491392 174020 491444 174072
rect 492404 174020 492456 174072
rect 446312 173952 446364 174004
rect 463792 173952 463844 174004
rect 502616 173952 502668 174004
rect 278596 173884 278648 173936
rect 295340 173884 295392 173936
rect 334624 173884 334676 173936
rect 345756 173884 345808 173936
rect 352012 173884 352064 173936
rect 379612 173884 379664 173936
rect 418620 173884 418672 173936
rect 429936 173884 429988 173936
rect 436100 173884 436152 173936
rect 457444 173884 457496 173936
rect 474648 173884 474700 173936
rect 486424 173884 486476 173936
rect 492312 173884 492364 173936
rect 492404 173884 492456 173936
rect 530308 174020 530360 174072
rect 541624 174020 541676 174072
rect 558644 174020 558696 174072
rect 514024 173884 514076 173936
rect 267924 173816 267976 173868
rect 520280 173884 520332 173936
rect 148968 172048 149020 172100
rect 153844 172048 153896 172100
rect 238668 171436 238720 171488
rect 291200 171436 291252 171488
rect 462228 171436 462280 171488
rect 514760 171436 514812 171488
rect 205088 171368 205140 171420
rect 209688 171368 209740 171420
rect 262220 171368 262272 171420
rect 434628 171368 434680 171420
rect 487160 171368 487212 171420
rect 541164 171232 541216 171284
rect 544384 171232 544436 171284
rect 40684 171164 40736 171216
rect 44180 171164 44232 171216
rect 71136 171164 71188 171216
rect 71964 171164 72016 171216
rect 205088 171164 205140 171216
rect 429108 171164 429160 171216
rect 429844 171164 429896 171216
rect 13544 171096 13596 171148
rect 66260 171096 66312 171148
rect 70308 171096 70360 171148
rect 122840 171096 122892 171148
rect 233240 166268 233292 166320
rect 233976 166268 234028 166320
rect 463700 166268 463752 166320
rect 464068 166268 464120 166320
rect 93124 153824 93176 153876
rect 99472 153824 99524 153876
rect 289176 153688 289228 153740
rect 295432 153688 295484 153740
rect 569408 151784 569460 151836
rect 580080 151784 580132 151836
rect 2780 149336 2832 149388
rect 5264 149336 5316 149388
rect 15292 148996 15344 149048
rect 36912 148996 36964 149048
rect 65064 148996 65116 149048
rect 92940 148996 92992 149048
rect 93032 148996 93084 149048
rect 120908 148996 120960 149048
rect 121092 148996 121144 149048
rect 148600 148996 148652 149048
rect 153844 148996 153896 149048
rect 176936 148996 176988 149048
rect 177028 148996 177080 149048
rect 204904 148996 204956 149048
rect 205180 148996 205232 149048
rect 232596 148996 232648 149048
rect 233976 148996 234028 149048
rect 260932 148996 260984 149048
rect 261024 148996 261076 149048
rect 288900 148996 288952 149048
rect 289084 148996 289136 149048
rect 316592 148996 316644 149048
rect 317052 148996 317104 149048
rect 344928 148996 344980 149048
rect 345664 148996 345716 149048
rect 372620 148996 372672 149048
rect 373080 148996 373132 149048
rect 400956 148996 401008 149048
rect 401048 148996 401100 149048
rect 428924 148996 428976 149048
rect 429844 148996 429896 149048
rect 456800 148996 456852 149048
rect 457076 148996 457128 149048
rect 484952 148996 485004 149048
rect 485044 148996 485096 149048
rect 512920 148996 512972 149048
rect 513104 148996 513156 149048
rect 540612 148996 540664 149048
rect 544384 148996 544436 149048
rect 568948 148996 569000 149048
rect 26608 148928 26660 148980
rect 40684 148928 40736 148980
rect 43444 148928 43496 148980
rect 64880 148928 64932 148980
rect 82636 148928 82688 148980
rect 93124 148928 93176 148980
rect 110604 148928 110656 148980
rect 122104 148928 122156 148980
rect 128636 148928 128688 148980
rect 149704 148928 149756 148980
rect 156328 148928 156380 148980
rect 177304 148928 177356 148980
rect 194600 148928 194652 148980
rect 206284 148928 206336 148980
rect 222936 148928 222988 148980
rect 234068 148928 234120 148980
rect 240324 148928 240376 148980
rect 262864 148928 262916 148980
rect 278596 148928 278648 148980
rect 289176 148928 289228 148980
rect 306932 148928 306984 148980
rect 318064 148928 318116 148980
rect 324320 148928 324372 148980
rect 345848 148928 345900 148980
rect 352656 148928 352708 148980
rect 373264 148928 373316 148980
rect 390652 148928 390704 148980
rect 402244 148928 402296 148980
rect 418620 148928 418672 148980
rect 429936 148928 429988 148980
rect 436652 148928 436704 148980
rect 457444 148928 457496 148980
rect 474648 148928 474700 148980
rect 486424 148928 486476 148980
rect 502616 148928 502668 148980
rect 514024 148928 514076 148980
rect 520648 148928 520700 148980
rect 541624 148928 541676 148980
rect 54852 148860 54904 148912
rect 71136 148860 71188 148912
rect 138940 148860 138992 148912
rect 155224 148860 155276 148912
rect 166632 148860 166684 148912
rect 178684 148860 178736 148912
rect 250628 148860 250680 148912
rect 264244 148860 264296 148912
rect 334624 148860 334676 148912
rect 345756 148860 345808 148912
rect 362868 148860 362920 148912
rect 374644 148860 374696 148912
rect 446956 148860 447008 148912
rect 463700 148860 463752 148912
rect 530952 148860 531004 148912
rect 547144 148860 547196 148912
rect 44640 148792 44692 148844
rect 66904 148792 66956 148844
rect 558644 148316 558696 148368
rect 568948 148316 569000 148368
rect 548340 146888 548392 146940
rect 569040 146888 569092 146940
rect 156328 146480 156380 146532
rect 180064 146480 180116 146532
rect 184020 146480 184072 146532
rect 204904 146480 204956 146532
rect 268016 146480 268068 146532
rect 289084 146480 289136 146532
rect 176844 146412 176896 146464
rect 194324 146412 194376 146464
rect 262864 146412 262916 146464
rect 278320 146412 278372 146464
rect 380348 146412 380400 146464
rect 401048 146412 401100 146464
rect 38200 146344 38252 146396
rect 54300 146344 54352 146396
rect 65892 146344 65944 146396
rect 81992 146344 82044 146396
rect 92940 146344 92992 146396
rect 110328 146344 110380 146396
rect 121000 146344 121052 146396
rect 138296 146344 138348 146396
rect 155224 146344 155276 146396
rect 165988 146344 166040 146396
rect 204812 146344 204864 146396
rect 222200 146344 222252 146396
rect 232780 146344 232832 146396
rect 250352 146344 250404 146396
rect 288808 146344 288860 146396
rect 306012 146344 306064 146396
rect 316776 146344 316828 146396
rect 334348 146344 334400 146396
rect 372896 146344 372948 146396
rect 390008 146344 390060 146396
rect 457444 146344 457496 146396
rect 474004 146344 474056 146396
rect 484860 146344 484912 146396
rect 502340 146344 502392 146396
rect 512736 146344 512788 146396
rect 530308 146344 530360 146396
rect 15292 146276 15344 146328
rect 26332 146276 26384 146328
rect 38108 146276 38160 146328
rect 64604 146276 64656 146328
rect 72332 146276 72384 146328
rect 93124 146276 93176 146328
rect 100024 146276 100076 146328
rect 121092 146276 121144 146328
rect 122104 146276 122156 146328
rect 148600 146276 148652 146328
rect 178684 146276 178736 146328
rect 204628 146276 204680 146328
rect 206284 146276 206336 146328
rect 232320 146276 232372 146328
rect 233976 146276 234028 146328
rect 260656 146276 260708 146328
rect 261484 146276 261536 146328
rect 288624 146276 288676 146328
rect 290464 146276 290516 146328
rect 316316 146276 316368 146328
rect 316868 146276 316920 146328
rect 344652 146276 344704 146328
rect 352012 146276 352064 146328
rect 373264 146276 373316 146328
rect 401140 146276 401192 146328
rect 418344 146276 418396 146328
rect 429844 146276 429896 146328
rect 456616 146276 456668 146328
rect 464344 146276 464396 146328
rect 485044 146276 485096 146328
rect 486424 146276 486476 146328
rect 512644 146276 512696 146328
rect 514024 146276 514076 146328
rect 540612 146276 540664 146328
rect 547144 146276 547196 146328
rect 558000 146276 558052 146328
rect 120724 144236 120776 144288
rect 121000 144236 121052 144288
rect 92756 144168 92808 144220
rect 92940 144168 92992 144220
rect 400772 144168 400824 144220
rect 401140 144168 401192 144220
rect 120816 144100 120868 144152
rect 121092 144100 121144 144152
rect 400864 144100 400916 144152
rect 401048 144100 401100 144152
rect 154488 143624 154540 143676
rect 207020 143624 207072 143676
rect 182088 143556 182140 143608
rect 234712 143556 234764 143608
rect 568764 142808 568816 142860
rect 568948 142808 569000 142860
rect 3332 136688 3384 136740
rect 7564 136688 7616 136740
rect 64880 128596 64932 128648
rect 65892 128596 65944 128648
rect 204904 128256 204956 128308
rect 211712 128256 211764 128308
rect 485044 128256 485096 128308
rect 491668 128256 491720 128308
rect 289084 127984 289136 128036
rect 295708 127984 295760 128036
rect 93124 127576 93176 127628
rect 99748 127576 99800 127628
rect 120816 127576 120868 127628
rect 127716 127576 127768 127628
rect 373264 127576 373316 127628
rect 379704 127576 379756 127628
rect 400864 127576 400916 127628
rect 407764 127576 407816 127628
rect 42708 125536 42760 125588
rect 95240 125536 95292 125588
rect 97908 125536 97960 125588
rect 150440 125536 150492 125588
rect 238668 125536 238720 125588
rect 291200 125536 291252 125588
rect 293868 125536 293920 125588
rect 346400 125536 346452 125588
rect 350448 125536 350500 125588
rect 402980 125536 403032 125588
rect 405648 125536 405700 125588
rect 458180 125536 458232 125588
rect 462228 125536 462280 125588
rect 514760 125536 514812 125588
rect 518808 125536 518860 125588
rect 571340 125536 571392 125588
rect 176752 124856 176804 124908
rect 372804 124856 372856 124908
rect 484768 124856 484820 124908
rect 15292 124652 15344 124704
rect 16120 124652 16172 124704
rect 36544 124652 36596 124704
rect 38200 124652 38252 124704
rect 176752 124652 176804 124704
rect 372804 124652 372856 124704
rect 484768 124652 484820 124704
rect 547880 124652 547932 124704
rect 548156 124652 548208 124704
rect 110328 122748 110380 122800
rect 122104 122748 122156 122800
rect 138296 122748 138348 122800
rect 176752 122748 176804 122800
rect 180064 122748 180116 122800
rect 184020 122748 184072 122800
rect 194324 122748 194376 122800
rect 206284 122748 206336 122800
rect 211252 122748 211304 122800
rect 240048 122748 240100 122800
rect 260656 122748 260708 122800
rect 262864 122748 262916 122800
rect 278320 122748 278372 122800
rect 290464 122748 290516 122800
rect 295432 122748 295484 122800
rect 324044 122748 324096 122800
rect 334348 122748 334400 122800
rect 372804 122748 372856 122800
rect 390468 122748 390520 122800
rect 428740 122748 428792 122800
rect 434812 122748 434864 122800
rect 26332 122680 26384 122732
rect 38108 122680 38160 122732
rect 42892 122680 42944 122732
rect 71780 122680 71832 122732
rect 82636 122680 82688 122732
rect 120908 122680 120960 122732
rect 127072 122680 127124 122732
rect 155960 122680 156012 122732
rect 166632 122680 166684 122732
rect 178684 122680 178736 122732
rect 222660 122680 222712 122732
rect 233976 122680 234028 122732
rect 250352 122680 250404 122732
rect 261484 122680 261536 122732
rect 306288 122680 306340 122732
rect 316868 122680 316920 122732
rect 323032 122680 323084 122732
rect 352012 122680 352064 122732
rect 362316 122680 362368 122732
rect 400956 122680 401008 122732
rect 407212 122680 407264 122732
rect 436008 122680 436060 122732
rect 491392 122748 491444 122800
rect 520004 122748 520056 122800
rect 530308 122748 530360 122800
rect 568856 122748 568908 122800
rect 463792 122680 463844 122732
rect 474648 122680 474700 122732
rect 486424 122680 486476 122732
rect 502340 122680 502392 122732
rect 514024 122680 514076 122732
rect 540612 122680 540664 122732
rect 547144 122680 547196 122732
rect 548156 122680 548208 122732
rect 558000 122680 558052 122732
rect 15384 122612 15436 122664
rect 43996 122612 44048 122664
rect 54300 122612 54352 122664
rect 92848 122612 92900 122664
rect 148600 122612 148652 122664
rect 155224 122612 155276 122664
rect 238852 122612 238904 122664
rect 268016 122612 268068 122664
rect 418344 122612 418396 122664
rect 429844 122612 429896 122664
rect 446312 122612 446364 122664
rect 484768 122612 484820 122664
rect 518992 122544 519044 122596
rect 547880 122544 547932 122596
rect 26608 120708 26660 120760
rect 36728 120708 36780 120760
rect 15568 120232 15620 120284
rect 54300 120232 54352 120284
rect 149704 120232 149756 120284
rect 166632 120232 166684 120284
rect 211160 120232 211212 120284
rect 250628 120232 250680 120284
rect 295432 120232 295484 120284
rect 71780 120164 71832 120216
rect 110604 120164 110656 120216
rect 122104 120164 122156 120216
rect 128360 120164 128412 120216
rect 149796 120164 149848 120216
rect 156328 120164 156380 120216
rect 183560 120164 183612 120216
rect 222292 120164 222344 120216
rect 262864 120164 262916 120216
rect 278228 120164 278280 120216
rect 290464 120164 290516 120216
rect 295984 120164 296036 120216
rect 407212 120232 407264 120284
rect 334624 120164 334676 120216
rect 378876 120164 378928 120216
rect 390744 120164 390796 120216
rect 402244 120164 402296 120216
rect 408316 120164 408368 120216
rect 429844 120232 429896 120284
rect 436100 120232 436152 120284
rect 491392 120232 491444 120284
rect 446312 120164 446364 120216
rect 457444 120164 457496 120216
rect 474372 120164 474424 120216
rect 486424 120164 486476 120216
rect 492312 120164 492364 120216
rect 541624 120232 541676 120284
rect 558644 120232 558696 120284
rect 530308 120164 530360 120216
rect 36912 120096 36964 120148
rect 43444 120096 43496 120148
rect 65892 120096 65944 120148
rect 82636 120096 82688 120148
rect 99380 120096 99432 120148
rect 138296 120096 138348 120148
rect 233976 120096 234028 120148
rect 240324 120096 240376 120148
rect 267832 120096 267884 120148
rect 306472 120096 306524 120148
rect 345664 120096 345716 120148
rect 362316 120096 362368 120148
rect 379520 120096 379572 120148
rect 418620 120096 418672 120148
rect 458824 120096 458876 120148
rect 464068 120096 464120 120148
rect 463792 120028 463844 120080
rect 502616 120096 502668 120148
rect 514024 120096 514076 120148
rect 520280 120096 520332 120148
rect 205088 117376 205140 117428
rect 293868 117376 293920 117428
rect 346400 117376 346452 117428
rect 40684 117240 40736 117292
rect 44088 117240 44140 117292
rect 238668 117308 238720 117360
rect 291200 117308 291252 117360
rect 322848 117308 322900 117360
rect 375380 117308 375432 117360
rect 434628 117308 434680 117360
rect 487160 117308 487212 117360
rect 264244 117240 264296 117292
rect 267924 117240 267976 117292
rect 345020 117240 345072 117292
rect 347044 117240 347096 117292
rect 348424 117240 348476 117292
rect 352012 117240 352064 117292
rect 429108 117240 429160 117292
rect 429936 117240 429988 117292
rect 541164 117240 541216 117292
rect 544384 117240 544436 117292
rect 205088 117172 205140 117224
rect 149244 115200 149296 115252
rect 149888 115200 149940 115252
rect 233240 114520 233292 114572
rect 234068 114520 234120 114572
rect 569500 111800 569552 111852
rect 580080 111800 580132 111852
rect 99380 100240 99432 100292
rect 99932 100240 99984 100292
rect 183560 100240 183612 100292
rect 184020 100240 184072 100292
rect 211160 100240 211212 100292
rect 211988 100240 212040 100292
rect 379520 100240 379572 100292
rect 379980 100240 380032 100292
rect 71780 97520 71832 97572
rect 72424 97520 72476 97572
rect 15200 95140 15252 95192
rect 36912 95140 36964 95192
rect 65064 95140 65116 95192
rect 92940 95140 92992 95192
rect 93032 95140 93084 95192
rect 120908 95140 120960 95192
rect 121092 95140 121144 95192
rect 148600 95140 148652 95192
rect 149888 95140 149940 95192
rect 176936 95140 176988 95192
rect 177028 95140 177080 95192
rect 204904 95140 204956 95192
rect 205180 95140 205232 95192
rect 232596 95140 232648 95192
rect 234068 95140 234120 95192
rect 260932 95140 260984 95192
rect 261024 95140 261076 95192
rect 288900 95140 288952 95192
rect 289084 95140 289136 95192
rect 316592 95140 316644 95192
rect 318064 95140 318116 95192
rect 344928 95140 344980 95192
rect 347044 95140 347096 95192
rect 372620 95140 372672 95192
rect 373080 95140 373132 95192
rect 400956 95140 401008 95192
rect 401048 95140 401100 95192
rect 428924 95140 428976 95192
rect 429936 95140 429988 95192
rect 456800 95140 456852 95192
rect 457076 95140 457128 95192
rect 484952 95140 485004 95192
rect 485044 95140 485096 95192
rect 512920 95140 512972 95192
rect 513104 95140 513156 95192
rect 540612 95140 540664 95192
rect 544384 95140 544436 95192
rect 568948 95140 569000 95192
rect 26608 95072 26660 95124
rect 40684 95072 40736 95124
rect 43444 95072 43496 95124
rect 64880 95072 64932 95124
rect 82636 95072 82688 95124
rect 99472 95072 99524 95124
rect 110604 95072 110656 95124
rect 122104 95072 122156 95124
rect 128636 95072 128688 95124
rect 149704 95072 149756 95124
rect 166632 95072 166684 95124
rect 183652 95072 183704 95124
rect 194600 95072 194652 95124
rect 211252 95072 211304 95124
rect 222936 95072 222988 95124
rect 233976 95072 234028 95124
rect 240324 95072 240376 95124
rect 262864 95072 262916 95124
rect 278596 95072 278648 95124
rect 290464 95072 290516 95124
rect 324320 95072 324372 95124
rect 345664 95072 345716 95124
rect 352656 95072 352708 95124
rect 378876 95072 378928 95124
rect 390652 95072 390704 95124
rect 402244 95072 402296 95124
rect 418620 95072 418672 95124
rect 429844 95072 429896 95124
rect 436652 95072 436704 95124
rect 457444 95072 457496 95124
rect 474648 95072 474700 95124
rect 486424 95072 486476 95124
rect 502616 95072 502668 95124
rect 514024 95072 514076 95124
rect 520648 95072 520700 95124
rect 541624 95072 541676 95124
rect 54944 95004 54996 95056
rect 72148 95004 72200 95056
rect 138940 95004 138992 95056
rect 149796 95004 149848 95056
rect 250628 95004 250680 95056
rect 264244 95004 264296 95056
rect 334624 95004 334676 95056
rect 348424 95004 348476 95056
rect 362868 95004 362920 95056
rect 379612 95004 379664 95056
rect 446956 95004 447008 95056
rect 458824 95004 458876 95056
rect 530952 95004 531004 95056
rect 547144 95004 547196 95056
rect 44640 94936 44692 94988
rect 65892 94936 65944 94988
rect 558644 94460 558696 94512
rect 568764 94460 568816 94512
rect 548340 93100 548392 93152
rect 569040 93100 569092 93152
rect 100024 92692 100076 92744
rect 120816 92692 120868 92744
rect 184020 92692 184072 92744
rect 204904 92692 204956 92744
rect 268016 92692 268068 92744
rect 289084 92692 289136 92744
rect 65892 92624 65944 92676
rect 81992 92624 82044 92676
rect 92756 92624 92808 92676
rect 110328 92624 110380 92676
rect 149796 92624 149848 92676
rect 165988 92624 166040 92676
rect 176752 92624 176804 92676
rect 194324 92624 194376 92676
rect 261576 92624 261628 92676
rect 278320 92624 278372 92676
rect 345756 92624 345808 92676
rect 362316 92624 362368 92676
rect 372804 92624 372856 92676
rect 390008 92624 390060 92676
rect 458824 92624 458876 92676
rect 474004 92624 474056 92676
rect 36912 92556 36964 92608
rect 54300 92556 54352 92608
rect 72332 92556 72384 92608
rect 93124 92556 93176 92608
rect 120724 92556 120776 92608
rect 138296 92556 138348 92608
rect 156328 92556 156380 92608
rect 180064 92556 180116 92608
rect 204812 92556 204864 92608
rect 222200 92556 222252 92608
rect 232780 92556 232832 92608
rect 250352 92556 250404 92608
rect 288808 92556 288860 92608
rect 306012 92556 306064 92608
rect 316776 92556 316828 92608
rect 334348 92556 334400 92608
rect 352012 92556 352064 92608
rect 376024 92556 376076 92608
rect 380348 92556 380400 92608
rect 400864 92556 400916 92608
rect 435364 92556 435416 92608
rect 446312 92556 446364 92608
rect 464344 92556 464396 92608
rect 485044 92556 485096 92608
rect 512920 92556 512972 92608
rect 530308 92556 530360 92608
rect 541716 92556 541768 92608
rect 558000 92556 558052 92608
rect 15200 92488 15252 92540
rect 26332 92488 26384 92540
rect 38108 92488 38160 92540
rect 64604 92488 64656 92540
rect 66904 92488 66956 92540
rect 92480 92488 92532 92540
rect 94504 92488 94556 92540
rect 120632 92488 120684 92540
rect 122104 92488 122156 92540
rect 148600 92488 148652 92540
rect 149704 92488 149756 92540
rect 176660 92488 176712 92540
rect 178684 92488 178736 92540
rect 204628 92488 204680 92540
rect 206284 92488 206336 92540
rect 232320 92488 232372 92540
rect 233976 92488 234028 92540
rect 260656 92488 260708 92540
rect 261484 92488 261536 92540
rect 288624 92488 288676 92540
rect 290464 92488 290516 92540
rect 316316 92488 316368 92540
rect 316868 92488 316920 92540
rect 344652 92488 344704 92540
rect 345664 92488 345716 92540
rect 372620 92488 372672 92540
rect 374644 92488 374696 92540
rect 400312 92488 400364 92540
rect 400772 92488 400824 92540
rect 418344 92488 418396 92540
rect 429844 92488 429896 92540
rect 456616 92488 456668 92540
rect 457444 92488 457496 92540
rect 484400 92488 484452 92540
rect 484768 92488 484820 92540
rect 502340 92488 502392 92540
rect 514024 92488 514076 92540
rect 540612 92488 540664 92540
rect 541624 92488 541676 92540
rect 568580 92488 568632 92540
rect 209688 89700 209740 89752
rect 262220 89700 262272 89752
rect 405648 89700 405700 89752
rect 458180 89700 458232 89752
rect 489828 89700 489880 89752
rect 542360 89700 542412 89752
rect 434720 87184 434772 87236
rect 435732 87184 435784 87236
rect 36820 85008 36872 85060
rect 37004 85008 37056 85060
rect 512828 85008 512880 85060
rect 513012 85008 513064 85060
rect 3332 84600 3384 84652
rect 9036 84600 9088 84652
rect 36820 77256 36872 77308
rect 37004 77256 37056 77308
rect 512828 77256 512880 77308
rect 513012 77256 513064 77308
rect 93124 73788 93176 73840
rect 99748 73788 99800 73840
rect 120816 73788 120868 73840
rect 127716 73788 127768 73840
rect 400864 73788 400916 73840
rect 407764 73788 407816 73840
rect 485044 73652 485096 73704
rect 491668 73652 491720 73704
rect 204904 73448 204956 73500
rect 211712 73448 211764 73500
rect 289084 73176 289136 73228
rect 295708 73176 295760 73228
rect 64880 72564 64932 72616
rect 65892 72564 65944 72616
rect 261024 72292 261076 72344
rect 261576 72292 261628 72344
rect 148968 71680 149020 71732
rect 149796 71680 149848 71732
rect 344928 71680 344980 71732
rect 345756 71680 345808 71732
rect 540888 71680 540940 71732
rect 541716 71680 541768 71732
rect 547880 70660 547932 70712
rect 548156 70660 548208 70712
rect 15200 69640 15252 69692
rect 16028 69640 16080 69692
rect 15384 68960 15436 69012
rect 43996 68960 44048 69012
rect 82636 68960 82688 69012
rect 94504 68960 94556 69012
rect 110328 68960 110380 69012
rect 122104 68960 122156 69012
rect 166632 68960 166684 69012
rect 178684 68960 178736 69012
rect 180064 68960 180116 69012
rect 184020 68960 184072 69012
rect 194324 68960 194376 69012
rect 206284 68960 206336 69012
rect 211252 68960 211304 69012
rect 240048 68960 240100 69012
rect 278320 68960 278372 69012
rect 290464 68960 290516 69012
rect 295432 68960 295484 69012
rect 324044 68960 324096 69012
rect 362316 68960 362368 69012
rect 374644 68960 374696 69012
rect 376024 68960 376076 69012
rect 379704 68960 379756 69012
rect 428648 68960 428700 69012
rect 435364 68960 435416 69012
rect 456616 68960 456668 69012
rect 458824 68960 458876 69012
rect 474648 68960 474700 69012
rect 512828 68960 512880 69012
rect 548156 68960 548208 69012
rect 558000 68960 558052 69012
rect 26332 68892 26384 68944
rect 38108 68892 38160 68944
rect 54300 68892 54352 68944
rect 66904 68892 66956 68944
rect 138296 68892 138348 68944
rect 149704 68892 149756 68944
rect 222660 68892 222712 68944
rect 233976 68892 234028 68944
rect 250352 68892 250404 68944
rect 261484 68892 261536 68944
rect 306288 68892 306340 68944
rect 316868 68892 316920 68944
rect 334348 68892 334400 68944
rect 345664 68892 345716 68944
rect 407212 68892 407264 68944
rect 436008 68892 436060 68944
rect 446312 68892 446364 68944
rect 457444 68892 457496 68944
rect 491392 68892 491444 68944
rect 520004 68892 520056 68944
rect 530308 68892 530360 68944
rect 541624 68892 541676 68944
rect 42892 68824 42944 68876
rect 71780 68824 71832 68876
rect 127072 68824 127124 68876
rect 156052 68824 156104 68876
rect 238852 68824 238904 68876
rect 268016 68824 268068 68876
rect 323032 68824 323084 68876
rect 352012 68824 352064 68876
rect 418344 68824 418396 68876
rect 429844 68824 429896 68876
rect 434720 68824 434772 68876
rect 463700 68824 463752 68876
rect 502340 68824 502392 68876
rect 514024 68824 514076 68876
rect 518900 68824 518952 68876
rect 547880 68824 547932 68876
rect 390468 68756 390520 68808
rect 428740 68756 428792 68808
rect 26608 66852 26660 66904
rect 36820 66852 36872 66904
rect 15384 66376 15436 66428
rect 54300 66376 54352 66428
rect 211252 66376 211304 66428
rect 250628 66376 250680 66428
rect 345664 66376 345716 66428
rect 362316 66376 362368 66428
rect 374644 66376 374696 66428
rect 380348 66376 380400 66428
rect 491392 66376 491444 66428
rect 65892 66308 65944 66360
rect 82636 66308 82688 66360
rect 99472 66308 99524 66360
rect 138296 66308 138348 66360
rect 149704 66308 149756 66360
rect 156328 66308 156380 66360
rect 183652 66308 183704 66360
rect 222384 66308 222436 66360
rect 267832 66308 267884 66360
rect 306380 66308 306432 66360
rect 318064 66308 318116 66360
rect 324320 66308 324372 66360
rect 373264 66308 373316 66360
rect 390652 66308 390704 66360
rect 407120 66308 407172 66360
rect 446312 66308 446364 66360
rect 457444 66308 457496 66360
rect 474648 66308 474700 66360
rect 486424 66308 486476 66360
rect 492312 66308 492364 66360
rect 530308 66308 530360 66360
rect 36912 66240 36964 66292
rect 43444 66240 43496 66292
rect 71872 66240 71924 66292
rect 110604 66240 110656 66292
rect 122104 66240 122156 66292
rect 128360 66240 128412 66292
rect 149888 66240 149940 66292
rect 166632 66240 166684 66292
rect 182824 66240 182876 66292
rect 194600 66240 194652 66292
rect 206284 66240 206336 66292
rect 211988 66240 212040 66292
rect 234068 66240 234120 66292
rect 240324 66240 240376 66292
rect 261484 66240 261536 66292
rect 278596 66240 278648 66292
rect 295432 66240 295484 66292
rect 334624 66240 334676 66292
rect 379612 66240 379664 66292
rect 418620 66240 418672 66292
rect 458824 66240 458876 66292
rect 464344 66240 464396 66292
rect 463792 66172 463844 66224
rect 502616 66240 502668 66292
rect 514024 66240 514076 66292
rect 520280 66240 520332 66292
rect 541624 66240 541676 66292
rect 558644 66240 558696 66292
rect 348424 63520 348476 63572
rect 352012 63520 352064 63572
rect 205088 63384 205140 63436
rect 40684 63248 40736 63300
rect 43996 63248 44048 63300
rect 345020 63248 345072 63300
rect 347044 63248 347096 63300
rect 429108 63248 429160 63300
rect 429844 63248 429896 63300
rect 205088 63180 205140 63232
rect 93124 61344 93176 61396
rect 99932 61344 99984 61396
rect 177304 61344 177356 61396
rect 184020 61344 184072 61396
rect 65984 60732 66036 60784
rect 71964 60732 72016 60784
rect 261576 60732 261628 60784
rect 267924 60732 267976 60784
rect 289176 60732 289228 60784
rect 295984 60732 296036 60784
rect 541716 60732 541768 60784
rect 548064 60732 548116 60784
rect 149244 59236 149296 59288
rect 149796 59236 149848 59288
rect 233240 59236 233292 59288
rect 233976 59236 234028 59288
rect 407120 50328 407172 50380
rect 407948 50328 408000 50380
rect 2964 44140 3016 44192
rect 11888 44140 11940 44192
rect 489828 44072 489880 44124
rect 542360 44072 542412 44124
rect 15292 41352 15344 41404
rect 36912 41352 36964 41404
rect 65064 41352 65116 41404
rect 92940 41352 92992 41404
rect 93032 41352 93084 41404
rect 120908 41352 120960 41404
rect 121092 41352 121144 41404
rect 148600 41352 148652 41404
rect 149796 41352 149848 41404
rect 176936 41352 176988 41404
rect 177028 41352 177080 41404
rect 204904 41352 204956 41404
rect 205180 41352 205232 41404
rect 232596 41352 232648 41404
rect 233976 41352 234028 41404
rect 260932 41352 260984 41404
rect 261024 41352 261076 41404
rect 288900 41352 288952 41404
rect 289084 41352 289136 41404
rect 316592 41352 316644 41404
rect 317052 41352 317104 41404
rect 344928 41352 344980 41404
rect 347044 41352 347096 41404
rect 372620 41352 372672 41404
rect 373080 41352 373132 41404
rect 400956 41352 401008 41404
rect 401048 41352 401100 41404
rect 428924 41352 428976 41404
rect 429844 41352 429896 41404
rect 456800 41352 456852 41404
rect 457076 41352 457128 41404
rect 484952 41352 485004 41404
rect 485044 41352 485096 41404
rect 512920 41352 512972 41404
rect 513104 41352 513156 41404
rect 540612 41352 540664 41404
rect 541072 41352 541124 41404
rect 568948 41352 569000 41404
rect 26608 41284 26660 41336
rect 40684 41284 40736 41336
rect 43444 41284 43496 41336
rect 64880 41284 64932 41336
rect 82636 41284 82688 41336
rect 93124 41284 93176 41336
rect 110604 41284 110656 41336
rect 122104 41284 122156 41336
rect 128636 41284 128688 41336
rect 149888 41284 149940 41336
rect 156328 41284 156380 41336
rect 182824 41284 182876 41336
rect 194600 41284 194652 41336
rect 206284 41284 206336 41336
rect 222936 41284 222988 41336
rect 234068 41284 234120 41336
rect 240324 41284 240376 41336
rect 261484 41284 261536 41336
rect 278596 41284 278648 41336
rect 289176 41284 289228 41336
rect 306932 41284 306984 41336
rect 318064 41284 318116 41336
rect 324320 41284 324372 41336
rect 345664 41284 345716 41336
rect 352656 41284 352708 41336
rect 373264 41284 373316 41336
rect 390652 41284 390704 41336
rect 407212 41284 407264 41336
rect 418620 41284 418672 41336
rect 436100 41284 436152 41336
rect 436652 41284 436704 41336
rect 457444 41284 457496 41336
rect 474648 41284 474700 41336
rect 486424 41284 486476 41336
rect 502616 41284 502668 41336
rect 514024 41284 514076 41336
rect 520648 41284 520700 41336
rect 541624 41284 541676 41336
rect 54944 41216 54996 41268
rect 65984 41216 66036 41268
rect 138940 41216 138992 41268
rect 149704 41216 149756 41268
rect 166632 41216 166684 41268
rect 177304 41216 177356 41268
rect 250628 41216 250680 41268
rect 261576 41216 261628 41268
rect 334624 41216 334676 41268
rect 348424 41216 348476 41268
rect 362868 41216 362920 41268
rect 374644 41216 374696 41268
rect 446956 41216 447008 41268
rect 458824 41216 458876 41268
rect 530952 41216 531004 41268
rect 541716 41216 541768 41268
rect 44640 41148 44692 41200
rect 65892 41148 65944 41200
rect 558644 40672 558696 40724
rect 568856 40672 568908 40724
rect 46940 39380 46992 39432
rect 205088 39380 205140 39432
rect 548340 39380 548392 39432
rect 569040 39380 569092 39432
rect 4988 39312 5040 39364
rect 41788 39312 41840 39364
rect 61108 39312 61160 39364
rect 569316 39312 569368 39364
rect 156328 38836 156380 38888
rect 180064 38836 180116 38888
rect 352012 38836 352064 38888
rect 373264 38836 373316 38888
rect 100024 38768 100076 38820
rect 121000 38768 121052 38820
rect 176844 38768 176896 38820
rect 194324 38768 194376 38820
rect 268016 38768 268068 38820
rect 289084 38768 289136 38820
rect 345664 38768 345716 38820
rect 362316 38768 362368 38820
rect 56600 38700 56652 38752
rect 92480 38700 92532 38752
rect 92756 38700 92808 38752
rect 110328 38700 110380 38752
rect 155224 38700 155276 38752
rect 165988 38700 166040 38752
rect 184020 38700 184072 38752
rect 204904 38700 204956 38752
rect 261484 38700 261536 38752
rect 278320 38700 278372 38752
rect 317144 38700 317196 38752
rect 334348 38700 334400 38752
rect 372804 38700 372856 38752
rect 390008 38700 390060 38752
rect 401048 38700 401100 38752
rect 418344 38700 418396 38752
rect 457444 38700 457496 38752
rect 474004 38700 474056 38752
rect 484860 38700 484912 38752
rect 502340 38700 502392 38752
rect 512736 38700 512788 38752
rect 530308 38700 530360 38752
rect 13728 38632 13780 38684
rect 81992 38632 82044 38684
rect 121092 38632 121144 38684
rect 138296 38632 138348 38684
rect 178684 38632 178736 38684
rect 204628 38632 204680 38684
rect 204812 38632 204864 38684
rect 222200 38632 222252 38684
rect 233976 38632 234028 38684
rect 260656 38632 260708 38684
rect 288900 38632 288952 38684
rect 306012 38632 306064 38684
rect 317052 38632 317104 38684
rect 344652 38632 344704 38684
rect 345756 38632 345808 38684
rect 372620 38632 372672 38684
rect 380348 38632 380400 38684
rect 401140 38632 401192 38684
rect 402244 38632 402296 38684
rect 428648 38632 428700 38684
rect 428740 38632 428792 38684
rect 446312 38632 446364 38684
rect 464344 38632 464396 38684
rect 485044 38632 485096 38684
rect 486424 38632 486476 38684
rect 512644 38632 512696 38684
rect 512828 38632 512880 38684
rect 540612 38632 540664 38684
rect 26976 38564 27028 38616
rect 37924 38564 37976 38616
rect 14464 38496 14516 38548
rect 38568 38496 38620 38548
rect 3976 38428 4028 38480
rect 33416 38428 33468 38480
rect 57888 38428 57940 38480
rect 65800 38428 65852 38480
rect 11704 38360 11756 38412
rect 22468 38360 22520 38412
rect 23756 38360 23808 38412
rect 152464 38360 152516 38412
rect 19248 38292 19300 38344
rect 234620 38292 234672 38344
rect 3424 38224 3476 38276
rect 54668 38224 54720 38276
rect 64604 38224 64656 38276
rect 569500 38224 569552 38276
rect 10324 38156 10376 38208
rect 30196 38156 30248 38208
rect 32128 38156 32180 38208
rect 545764 38156 545816 38208
rect 5172 38088 5224 38140
rect 45008 38088 45060 38140
rect 51448 38088 51500 38140
rect 569408 38088 569460 38140
rect 4804 38020 4856 38072
rect 20536 38020 20588 38072
rect 25688 38020 25740 38072
rect 580632 38020 580684 38072
rect 17316 37952 17368 38004
rect 580448 37952 580500 38004
rect 16028 37884 16080 37936
rect 580908 37884 580960 37936
rect 35348 37340 35400 37392
rect 38016 37340 38068 37392
rect 40040 37340 40092 37392
rect 48228 37340 48280 37392
rect 59820 37340 59872 37392
rect 65708 37340 65760 37392
rect 36636 37272 36688 37324
rect 95240 37272 95292 37324
rect 64512 36796 64564 36848
rect 95884 36796 95936 36848
rect 64236 36728 64288 36780
rect 569224 36728 569276 36780
rect 64420 36660 64472 36712
rect 580356 36660 580408 36712
rect 64328 36592 64380 36644
rect 580540 36592 580592 36644
rect 13544 36524 13596 36576
rect 580816 36524 580868 36576
rect 120724 36252 120776 36304
rect 121092 36252 121144 36304
rect 316868 36184 316920 36236
rect 317052 36184 317104 36236
rect 400772 36184 400824 36236
rect 401048 36184 401100 36236
rect 120816 36116 120868 36168
rect 121000 36116 121052 36168
rect 316776 36116 316828 36168
rect 317144 36116 317196 36168
rect 400864 36116 400916 36168
rect 401140 36116 401192 36168
rect 39856 36048 39908 36100
rect 61384 36048 61436 36100
rect 3424 35980 3476 36032
rect 43444 35980 43496 36032
rect 50528 35980 50580 36032
rect 61476 35980 61528 36032
rect 28724 35912 28776 35964
rect 580908 35912 580960 35964
rect 3792 35164 3844 35216
rect 61292 35164 61344 35216
rect 3332 31696 3384 31748
rect 12440 31696 12492 31748
rect 64328 31016 64380 31068
rect 64604 31016 64656 31068
rect 63500 27072 63552 27124
rect 65616 27072 65668 27124
rect 5080 23400 5132 23452
rect 12440 23400 12492 23452
rect 6184 22040 6236 22092
rect 12440 22040 12492 22092
rect 176752 21360 176804 21412
rect 176936 21360 176988 21412
rect 484768 21360 484820 21412
rect 484952 21360 485004 21412
rect 7564 20612 7616 20664
rect 12440 20612 12492 20664
rect 63500 19252 63552 19304
rect 69664 19252 69716 19304
rect 289084 18640 289136 18692
rect 295708 18640 295760 18692
rect 120816 18572 120868 18624
rect 127716 18572 127768 18624
rect 373264 18572 373316 18624
rect 379704 18572 379756 18624
rect 400864 18572 400916 18624
rect 407764 18572 407816 18624
rect 204904 17960 204956 18012
rect 211712 17960 211764 18012
rect 485044 17960 485096 18012
rect 491668 17960 491720 18012
rect 6276 17892 6328 17944
rect 12440 17892 12492 17944
rect 288532 16668 288584 16720
rect 288900 16668 288952 16720
rect 568488 16668 568540 16720
rect 569040 16668 569092 16720
rect 3792 16532 3844 16584
rect 63592 16532 63644 16584
rect 4896 15104 4948 15156
rect 35348 15104 35400 15156
rect 41788 15104 41840 15156
rect 429200 15104 429252 15156
rect 5264 15036 5316 15088
rect 22468 15036 22520 15088
rect 52736 15036 52788 15088
rect 233884 15036 233936 15088
rect 23756 14968 23808 15020
rect 65524 14968 65576 15020
rect 48228 14900 48280 14952
rect 71044 14900 71096 14952
rect 9036 13744 9088 13796
rect 16028 13744 16080 13796
rect 148600 13744 148652 13796
rect 155224 13744 155276 13796
rect 166632 13744 166684 13796
rect 178684 13744 178736 13796
rect 180064 13744 180116 13796
rect 184020 13744 184072 13796
rect 222660 13744 222712 13796
rect 233976 13744 234028 13796
rect 306288 13744 306340 13796
rect 316868 13744 316920 13796
rect 390468 13744 390520 13796
rect 402244 13744 402296 13796
rect 474648 13744 474700 13796
rect 486424 13744 486476 13796
rect 502340 13744 502392 13796
rect 512828 13744 512880 13796
rect 547880 13744 547932 13796
rect 558000 13744 558052 13796
rect 17316 13676 17368 13728
rect 574744 13676 574796 13728
rect 3516 13608 3568 13660
rect 28908 13608 28960 13660
rect 32128 13608 32180 13660
rect 580080 13608 580132 13660
rect 4068 13540 4120 13592
rect 25688 13540 25740 13592
rect 36636 13540 36688 13592
rect 580724 13540 580776 13592
rect 43076 13472 43128 13524
rect 580172 13472 580224 13524
rect 3700 13404 3752 13456
rect 57888 13404 57940 13456
rect 59820 13404 59872 13456
rect 580264 13404 580316 13456
rect 19248 13336 19300 13388
rect 518164 13336 518216 13388
rect 26976 13268 27028 13320
rect 378784 13268 378836 13320
rect 407212 13268 407264 13320
rect 436008 13268 436060 13320
rect 446312 13268 446364 13320
rect 484952 13268 485004 13320
rect 491392 13268 491444 13320
rect 520004 13336 520056 13388
rect 530308 13336 530360 13388
rect 568948 13336 569000 13388
rect 518992 13268 519044 13320
rect 547972 13268 548024 13320
rect 6920 13200 6972 13252
rect 55956 13200 56008 13252
rect 82636 13200 82688 13252
rect 120908 13200 120960 13252
rect 138296 13200 138348 13252
rect 176936 13200 176988 13252
rect 194324 13200 194376 13252
rect 232780 13200 232832 13252
rect 238852 13200 238904 13252
rect 11796 13132 11848 13184
rect 54668 13132 54720 13184
rect 71872 13132 71924 13184
rect 100024 13132 100076 13184
rect 110328 13132 110380 13184
rect 148784 13132 148836 13184
rect 211252 13132 211304 13184
rect 240048 13132 240100 13184
rect 250352 13200 250404 13252
rect 288808 13200 288860 13252
rect 295432 13200 295484 13252
rect 268016 13132 268068 13184
rect 278320 13132 278372 13184
rect 316960 13132 317012 13184
rect 323032 13200 323084 13252
rect 352012 13200 352064 13252
rect 362316 13200 362368 13252
rect 400956 13200 401008 13252
rect 434812 13200 434864 13252
rect 463700 13200 463752 13252
rect 324044 13132 324096 13184
rect 334348 13132 334400 13184
rect 345756 13132 345808 13184
rect 1400 13064 1452 13116
rect 33416 13064 33468 13116
rect 38568 13064 38620 13116
rect 72056 13064 72108 13116
rect 127072 13064 127124 13116
rect 156052 13064 156104 13116
rect 8944 12996 8996 13048
rect 30196 12996 30248 13048
rect 39856 12996 39908 13048
rect 68284 12996 68336 13048
rect 20536 12928 20588 12980
rect 578884 12928 578936 12980
rect 3608 12860 3660 12912
rect 46296 12860 46348 12912
rect 3884 12792 3936 12844
rect 51448 12792 51500 12844
rect 64236 3680 64288 3732
rect 125876 3680 125928 3732
rect 64144 3612 64196 3664
rect 126980 3612 127032 3664
rect 61476 3544 61528 3596
rect 132960 3544 133012 3596
rect 13728 3476 13780 3528
rect 129372 3476 129424 3528
rect 572 3408 624 3460
rect 48320 3408 48372 3460
rect 61384 3408 61436 3460
rect 136456 3408 136508 3460
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 2832 632088 2834 632097
rect 2778 632023 2834 632032
rect 2778 606112 2834 606121
rect 2778 606047 2834 606056
rect 2792 605946 2820 606047
rect 2780 605940 2832 605946
rect 2780 605882 2832 605888
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 2778 449576 2834 449585
rect 2778 449511 2834 449520
rect 2792 448866 2820 449511
rect 2780 448860 2832 448866
rect 2780 448802 2832 448808
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 410242 3188 410479
rect 3148 410236 3200 410242
rect 3148 410178 3200 410184
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 2778 345400 2834 345409
rect 2778 345335 2834 345344
rect 2792 345234 2820 345335
rect 2780 345228 2832 345234
rect 2780 345170 2832 345176
rect 3146 293176 3202 293185
rect 3146 293111 3202 293120
rect 3160 292738 3188 293111
rect 3148 292732 3200 292738
rect 3148 292674 3200 292680
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 3252 240174 3280 241023
rect 3240 240168 3292 240174
rect 3240 240110 3292 240116
rect 2778 188864 2834 188873
rect 2778 188799 2834 188808
rect 2792 187746 2820 188799
rect 2780 187740 2832 187746
rect 2780 187682 2832 187688
rect 2778 149832 2834 149841
rect 2778 149767 2834 149776
rect 2792 149394 2820 149767
rect 2780 149388 2832 149394
rect 2780 149330 2832 149336
rect 3330 136776 3386 136785
rect 3330 136711 3332 136720
rect 3384 136711 3386 136720
rect 3332 136682 3384 136688
rect 3330 84688 3386 84697
rect 3330 84623 3332 84632
rect 3384 84623 3386 84632
rect 3332 84594 3384 84600
rect 3330 58576 3386 58585
rect 3330 58511 3386 58520
rect 2962 45520 3018 45529
rect 2962 45455 3018 45464
rect 2976 44198 3004 45455
rect 2964 44192 3016 44198
rect 2964 44134 3016 44140
rect 3344 31754 3372 58511
rect 3436 38282 3464 684247
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 4804 632120 4856 632126
rect 4804 632062 4856 632068
rect 3514 580000 3570 580009
rect 3514 579935 3570 579944
rect 3424 38276 3476 38282
rect 3424 38218 3476 38224
rect 3424 36032 3476 36038
rect 3424 35974 3476 35980
rect 3332 31748 3384 31754
rect 3332 31690 3384 31696
rect 1400 13116 1452 13122
rect 1400 13058 1452 13064
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 542 -960 654 480
rect 1412 354 1440 13058
rect 3436 6497 3464 35974
rect 3528 13666 3556 579935
rect 3606 553888 3662 553897
rect 3606 553823 3662 553832
rect 3620 553450 3648 553823
rect 3608 553444 3660 553450
rect 3608 553386 3660 553392
rect 3606 501800 3662 501809
rect 3606 501735 3662 501744
rect 3516 13660 3568 13666
rect 3516 13602 3568 13608
rect 3620 12918 3648 501735
rect 3698 475688 3754 475697
rect 3698 475623 3754 475632
rect 3712 13462 3740 475623
rect 3790 358456 3846 358465
rect 3790 358391 3846 358400
rect 3804 35222 3832 358391
rect 3882 306232 3938 306241
rect 3882 306167 3938 306176
rect 3792 35216 3844 35222
rect 3792 35158 3844 35164
rect 3790 19408 3846 19417
rect 3790 19343 3846 19352
rect 3804 16590 3832 19343
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3700 13456 3752 13462
rect 3700 13398 3752 13404
rect 3608 12912 3660 12918
rect 3608 12854 3660 12860
rect 3896 12850 3924 306167
rect 3974 254144 4030 254153
rect 3974 254079 4030 254088
rect 3988 38486 4016 254079
rect 4066 97608 4122 97617
rect 4066 97543 4122 97552
rect 3976 38480 4028 38486
rect 3976 38422 4028 38428
rect 4080 13598 4108 97543
rect 4816 38078 4844 632062
rect 4896 605940 4948 605946
rect 4896 605882 4948 605888
rect 4804 38072 4856 38078
rect 4804 38014 4856 38020
rect 4908 15162 4936 605882
rect 6184 527196 6236 527202
rect 6184 527138 6236 527144
rect 4988 448860 5040 448866
rect 4988 448802 5040 448808
rect 5000 39370 5028 448802
rect 5080 345228 5132 345234
rect 5080 345170 5132 345176
rect 4988 39364 5040 39370
rect 4988 39306 5040 39312
rect 5092 23458 5120 345170
rect 5172 187740 5224 187746
rect 5172 187682 5224 187688
rect 5184 38146 5212 187682
rect 5264 149388 5316 149394
rect 5264 149330 5316 149336
rect 5172 38140 5224 38146
rect 5172 38082 5224 38088
rect 5080 23452 5132 23458
rect 5080 23394 5132 23400
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 5276 15094 5304 149330
rect 6196 22098 6224 527138
rect 6276 292732 6328 292738
rect 6276 292674 6328 292680
rect 6184 22092 6236 22098
rect 6184 22034 6236 22040
rect 6288 17950 6316 292674
rect 6276 17944 6328 17950
rect 6276 17886 6328 17892
rect 5264 15088 5316 15094
rect 5264 15030 5316 15036
rect 4068 13592 4120 13598
rect 4068 13534 4120 13540
rect 6932 13258 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 37924 700800 37976 700806
rect 37924 700742 37976 700748
rect 13452 700528 13504 700534
rect 13452 700470 13504 700476
rect 11704 656940 11756 656946
rect 11704 656882 11756 656888
rect 10324 553444 10376 553450
rect 10324 553386 10376 553392
rect 8944 410236 8996 410242
rect 8944 410178 8996 410184
rect 7564 136740 7616 136746
rect 7564 136682 7616 136688
rect 7576 20670 7604 136682
rect 7564 20664 7616 20670
rect 7564 20606 7616 20612
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 8956 13054 8984 410178
rect 9036 84652 9088 84658
rect 9036 84594 9088 84600
rect 9048 13802 9076 84594
rect 10336 38214 10364 553386
rect 11716 38418 11744 656882
rect 11796 397520 11848 397526
rect 11796 397462 11848 397468
rect 11704 38412 11756 38418
rect 11704 38354 11756 38360
rect 10324 38208 10376 38214
rect 10324 38150 10376 38156
rect 9036 13796 9088 13802
rect 9036 13738 9088 13744
rect 11808 13190 11836 397462
rect 11888 44192 11940 44198
rect 11888 44134 11940 44140
rect 11900 34513 11928 44134
rect 11886 34504 11942 34513
rect 11886 34439 11942 34448
rect 13464 33153 13492 700470
rect 36912 687336 36964 687342
rect 36912 687278 36964 687284
rect 15292 687268 15344 687274
rect 15292 687210 15344 687216
rect 26332 687268 26384 687274
rect 26332 687210 26384 687216
rect 13634 674248 13690 674257
rect 13634 674183 13690 674192
rect 13648 665961 13676 674183
rect 13634 665952 13690 665961
rect 13634 665887 13690 665896
rect 15304 664766 15332 687210
rect 26344 684964 26372 687210
rect 15396 684270 16054 684298
rect 36662 684270 36768 684298
rect 15292 664760 15344 664766
rect 15292 664702 15344 664708
rect 15396 662386 15424 684270
rect 36740 680218 36768 684270
rect 36740 680190 36860 680218
rect 36832 676214 36860 680190
rect 36740 676186 36860 676214
rect 36740 673454 36768 676186
rect 36740 673426 36860 673454
rect 36832 668642 36860 673426
rect 36820 668636 36872 668642
rect 36820 668578 36872 668584
rect 36924 664766 36952 687278
rect 37004 668636 37056 668642
rect 37004 668578 37056 668584
rect 16120 664760 16172 664766
rect 16120 664702 16172 664708
rect 36544 664760 36596 664766
rect 36912 664760 36964 664766
rect 36596 664708 36662 664714
rect 36544 664702 36662 664708
rect 36912 664702 36964 664708
rect 15488 664006 16054 664034
rect 15384 662380 15436 662386
rect 15384 662322 15436 662328
rect 13636 661700 13688 661706
rect 13636 661642 13688 661648
rect 13542 620256 13598 620265
rect 13542 620191 13598 620200
rect 13556 611969 13584 620191
rect 13542 611960 13598 611969
rect 13542 611895 13598 611904
rect 13542 602032 13598 602041
rect 13542 601967 13598 601976
rect 13556 593745 13584 601967
rect 13542 593736 13598 593745
rect 13542 593671 13598 593680
rect 13542 574696 13598 574705
rect 13542 574631 13598 574640
rect 13556 566273 13584 574631
rect 13542 566264 13598 566273
rect 13542 566199 13598 566208
rect 13542 548040 13598 548049
rect 13542 547975 13598 547984
rect 13556 539753 13584 547975
rect 13542 539744 13598 539753
rect 13542 539679 13598 539688
rect 13542 485752 13598 485761
rect 13542 485687 13598 485696
rect 13556 477329 13584 485687
rect 13542 477320 13598 477329
rect 13542 477255 13598 477264
rect 13542 466712 13598 466721
rect 13542 466647 13598 466656
rect 13556 458289 13584 466647
rect 13542 458280 13598 458289
rect 13542 458215 13598 458224
rect 13542 404288 13598 404297
rect 13542 404223 13598 404232
rect 13556 396001 13584 404223
rect 13542 395992 13598 396001
rect 13542 395927 13598 395936
rect 13542 377768 13598 377777
rect 13542 377703 13598 377712
rect 13556 369345 13584 377703
rect 13542 369336 13598 369345
rect 13542 369271 13598 369280
rect 13542 350296 13598 350305
rect 13542 350231 13598 350240
rect 13556 342009 13584 350231
rect 13542 342000 13598 342009
rect 13542 341935 13598 341944
rect 13542 323776 13598 323785
rect 13542 323711 13598 323720
rect 13556 315353 13584 323711
rect 13542 315344 13598 315353
rect 13542 315279 13598 315288
rect 13542 278080 13598 278089
rect 13542 278015 13598 278024
rect 13556 269793 13584 278015
rect 13542 269784 13598 269793
rect 13542 269719 13598 269728
rect 13542 242312 13598 242321
rect 13542 242247 13598 242256
rect 13556 234025 13584 242247
rect 13542 234016 13598 234025
rect 13542 233951 13598 233960
rect 13542 224088 13598 224097
rect 13542 224023 13598 224032
rect 13556 215801 13584 224023
rect 13542 215792 13598 215801
rect 13542 215727 13598 215736
rect 13542 196752 13598 196761
rect 13542 196687 13598 196696
rect 13556 188329 13584 196687
rect 13542 188320 13598 188329
rect 13542 188255 13598 188264
rect 13544 171148 13596 171154
rect 13544 171090 13596 171096
rect 13556 161809 13584 171090
rect 13542 161800 13598 161809
rect 13542 161735 13598 161744
rect 13542 142760 13598 142769
rect 13542 142695 13598 142704
rect 13556 134337 13584 142695
rect 13542 134328 13598 134337
rect 13542 134263 13598 134272
rect 13542 116104 13598 116113
rect 13542 116039 13598 116048
rect 13556 107817 13584 116039
rect 13542 107808 13598 107817
rect 13542 107743 13598 107752
rect 13542 88768 13598 88777
rect 13542 88703 13598 88712
rect 13556 80345 13584 88703
rect 13542 80336 13598 80345
rect 13542 80271 13598 80280
rect 13542 53816 13598 53825
rect 13542 53751 13598 53760
rect 13556 45393 13584 53751
rect 13542 45384 13598 45393
rect 13542 45319 13598 45328
rect 13544 36576 13596 36582
rect 13544 36518 13596 36524
rect 13450 33144 13506 33153
rect 13450 33079 13506 33088
rect 12440 31748 12492 31754
rect 12440 31690 12492 31696
rect 12452 31113 12480 31690
rect 12438 31104 12494 31113
rect 12438 31039 12494 31048
rect 13556 29753 13584 36518
rect 13542 29744 13598 29753
rect 13542 29679 13598 29688
rect 13648 27713 13676 661642
rect 15488 659002 15516 664006
rect 15568 659728 15620 659734
rect 15568 659670 15620 659676
rect 15212 658974 15516 659002
rect 13726 656024 13782 656033
rect 13726 655959 13782 655968
rect 13740 647737 13768 655959
rect 13726 647728 13782 647737
rect 13726 647663 13782 647672
rect 15212 634778 15240 658974
rect 15580 654134 15608 659670
rect 16132 657914 16160 664702
rect 36556 664686 36662 664702
rect 26344 662318 26372 664020
rect 37016 663794 37044 668578
rect 36832 663766 37044 663794
rect 26332 662312 26384 662318
rect 26332 662254 26384 662260
rect 36832 660346 36860 663766
rect 26608 660340 26660 660346
rect 26608 660282 26660 660288
rect 36820 660340 36872 660346
rect 36820 660282 36872 660288
rect 16132 657886 16330 657914
rect 26620 657900 26648 660282
rect 36938 657206 37136 657234
rect 15580 654106 15976 654134
rect 15948 637786 15976 654106
rect 15948 637758 16330 637786
rect 15200 634772 15252 634778
rect 15200 634714 15252 634720
rect 26620 634710 26648 637092
rect 36924 634778 36952 637092
rect 37108 634778 37136 657206
rect 36912 634772 36964 634778
rect 36912 634714 36964 634720
rect 37096 634772 37148 634778
rect 37096 634714 37148 634720
rect 26608 634704 26660 634710
rect 26608 634646 26660 634652
rect 37096 632188 37148 632194
rect 37096 632130 37148 632136
rect 15292 632120 15344 632126
rect 15292 632062 15344 632068
rect 26332 632120 26384 632126
rect 26332 632062 26384 632068
rect 15304 610162 15332 632062
rect 26344 630972 26372 632062
rect 36662 630414 37044 630442
rect 15396 630278 16054 630306
rect 36728 630284 36780 630290
rect 15292 610156 15344 610162
rect 15292 610098 15344 610104
rect 15396 608598 15424 630278
rect 36728 630226 36780 630232
rect 36740 610722 36768 630226
rect 37016 621058 37044 630414
rect 37108 630290 37136 632130
rect 37096 630284 37148 630290
rect 37096 630226 37148 630232
rect 36662 610694 36768 610722
rect 36832 621030 37044 621058
rect 15488 610014 16054 610042
rect 15384 608592 15436 608598
rect 15384 608534 15436 608540
rect 15488 608002 15516 610014
rect 15936 609952 15988 609958
rect 15936 609894 15988 609900
rect 15212 607974 15516 608002
rect 15212 580990 15240 607974
rect 15384 606008 15436 606014
rect 15384 605950 15436 605956
rect 15396 596174 15424 605950
rect 15948 603922 15976 609894
rect 26344 608530 26372 610028
rect 26332 608524 26384 608530
rect 26332 608466 26384 608472
rect 36832 606490 36860 621030
rect 26608 606484 26660 606490
rect 26608 606426 26660 606432
rect 36820 606484 36872 606490
rect 36820 606426 36872 606432
rect 15948 603894 16330 603922
rect 26620 603908 26648 606426
rect 36938 603214 37320 603242
rect 37292 599758 37320 603214
rect 37280 599752 37332 599758
rect 37280 599694 37332 599700
rect 15396 596146 15976 596174
rect 15948 583794 15976 596146
rect 15948 583766 16330 583794
rect 15200 580984 15252 580990
rect 15200 580926 15252 580932
rect 26620 580922 26648 583100
rect 36924 580990 36952 583100
rect 36912 580984 36964 580990
rect 36912 580926 36964 580932
rect 26608 580916 26660 580922
rect 26608 580858 26660 580864
rect 36912 578332 36964 578338
rect 36912 578274 36964 578280
rect 15292 578264 15344 578270
rect 15292 578206 15344 578212
rect 26332 578264 26384 578270
rect 26332 578206 26384 578212
rect 15304 553382 15332 578206
rect 26344 576980 26372 578206
rect 15396 576286 16054 576314
rect 36662 576286 36860 576314
rect 15396 554742 15424 576286
rect 36832 571266 36860 576286
rect 36820 571260 36872 571266
rect 36820 571202 36872 571208
rect 36924 569954 36952 578274
rect 37004 571260 37056 571266
rect 37004 571202 37056 571208
rect 36740 569926 36952 569954
rect 36740 556730 36768 569926
rect 37016 567202 37044 571202
rect 36662 556702 36768 556730
rect 36832 567174 37044 567202
rect 15488 556022 16054 556050
rect 15384 554736 15436 554742
rect 15384 554678 15436 554684
rect 15292 553376 15344 553382
rect 15292 553318 15344 553324
rect 15488 551970 15516 556022
rect 26344 554674 26372 556036
rect 26332 554668 26384 554674
rect 26332 554610 26384 554616
rect 16028 553376 16080 553382
rect 16028 553318 16080 553324
rect 15568 552220 15620 552226
rect 15568 552162 15620 552168
rect 15212 551942 15516 551970
rect 15212 527134 15240 551942
rect 15580 547874 15608 552162
rect 16040 549930 16068 553318
rect 36832 552702 36860 567174
rect 26608 552696 26660 552702
rect 26608 552638 26660 552644
rect 36820 552696 36872 552702
rect 36820 552638 36872 552644
rect 16040 549902 16330 549930
rect 26620 549916 26648 552638
rect 36938 549358 37320 549386
rect 37292 548554 37320 549358
rect 37280 548548 37332 548554
rect 37280 548490 37332 548496
rect 15396 547846 15608 547874
rect 15396 538214 15424 547846
rect 15396 538186 15976 538214
rect 15948 529666 15976 538186
rect 15948 529638 16330 529666
rect 15200 527128 15252 527134
rect 15200 527070 15252 527076
rect 26620 527066 26648 529108
rect 36924 527134 36952 529108
rect 36912 527128 36964 527134
rect 36912 527070 36964 527076
rect 26608 527060 26660 527066
rect 26608 527002 26660 527008
rect 37096 524544 37148 524550
rect 37096 524486 37148 524492
rect 15292 524476 15344 524482
rect 15292 524418 15344 524424
rect 26332 524476 26384 524482
rect 26332 524418 26384 524424
rect 13726 520704 13782 520713
rect 13726 520639 13782 520648
rect 13740 512281 13768 520639
rect 13726 512272 13782 512281
rect 13726 512207 13782 512216
rect 15304 497418 15332 524418
rect 26344 522852 26372 524418
rect 36662 522430 37044 522458
rect 15396 522294 16054 522322
rect 36728 522300 36780 522306
rect 15396 500954 15424 522294
rect 36728 522242 36780 522248
rect 36740 502738 36768 522242
rect 37016 518514 37044 522430
rect 37108 522306 37136 524486
rect 37096 522300 37148 522306
rect 37096 522242 37148 522248
rect 36662 502710 36768 502738
rect 36832 518486 37044 518514
rect 15488 502030 16054 502058
rect 15384 500948 15436 500954
rect 15384 500890 15436 500896
rect 15292 497412 15344 497418
rect 15292 497354 15344 497360
rect 15488 489914 15516 502030
rect 26344 500886 26372 502044
rect 26332 500880 26384 500886
rect 26332 500822 26384 500828
rect 36832 498846 36860 518486
rect 26608 498840 26660 498846
rect 26608 498782 26660 498788
rect 36820 498840 36872 498846
rect 36820 498782 36872 498788
rect 15936 498364 15988 498370
rect 15936 498306 15988 498312
rect 15212 489886 15516 489914
rect 15212 473346 15240 489886
rect 15948 475674 15976 498306
rect 16028 497412 16080 497418
rect 16028 497354 16080 497360
rect 16040 495938 16068 497354
rect 16040 495910 16330 495938
rect 26620 495924 26648 498782
rect 36938 495502 37320 495530
rect 37292 492590 37320 495502
rect 37280 492584 37332 492590
rect 37280 492526 37332 492532
rect 15948 475646 16330 475674
rect 15200 473340 15252 473346
rect 15200 473282 15252 473288
rect 26620 473278 26648 475116
rect 36924 473346 36952 475116
rect 36912 473340 36964 473346
rect 36912 473282 36964 473288
rect 26608 473272 26660 473278
rect 26608 473214 26660 473220
rect 15292 470620 15344 470626
rect 15292 470562 15344 470568
rect 26332 470620 26384 470626
rect 26332 470562 26384 470568
rect 36728 470620 36780 470626
rect 36728 470562 36780 470568
rect 15304 448186 15332 470562
rect 26344 468860 26372 470562
rect 36740 468450 36768 470562
rect 36728 468444 36780 468450
rect 36728 468386 36780 468392
rect 15488 468302 16054 468330
rect 36662 468302 36860 468330
rect 15292 448180 15344 448186
rect 15292 448122 15344 448128
rect 15488 445738 15516 468302
rect 36728 468240 36780 468246
rect 36728 468182 36780 468188
rect 36740 448746 36768 468182
rect 36662 448718 36768 448746
rect 16120 448180 16172 448186
rect 16120 448122 16172 448128
rect 15580 448038 16054 448066
rect 15476 445732 15528 445738
rect 15476 445674 15528 445680
rect 15580 444802 15608 448038
rect 15212 444774 15608 444802
rect 13726 431760 13782 431769
rect 13726 431695 13782 431704
rect 13740 423337 13768 431695
rect 13726 423328 13782 423337
rect 13726 423263 13782 423272
rect 15212 419490 15240 444774
rect 15384 444508 15436 444514
rect 15384 444450 15436 444456
rect 15396 441614 15424 444450
rect 16132 441946 16160 448122
rect 26344 445670 26372 448052
rect 26332 445664 26384 445670
rect 26332 445606 26384 445612
rect 36832 445058 36860 468302
rect 26608 445052 26660 445058
rect 26608 444994 26660 445000
rect 36820 445052 36872 445058
rect 36820 444994 36872 445000
rect 16132 441918 16330 441946
rect 26620 441932 26648 444994
rect 15396 441586 15976 441614
rect 15948 421682 15976 441586
rect 36938 441238 37320 441266
rect 37096 438932 37148 438938
rect 37096 438874 37148 438880
rect 15948 421654 16330 421682
rect 15200 419484 15252 419490
rect 15200 419426 15252 419432
rect 26620 419422 26648 421124
rect 36924 419490 36952 421124
rect 36912 419484 36964 419490
rect 36912 419426 36964 419432
rect 37108 419422 37136 438874
rect 37292 436626 37320 441238
rect 37280 436620 37332 436626
rect 37280 436562 37332 436568
rect 26608 419416 26660 419422
rect 26608 419358 26660 419364
rect 37096 419416 37148 419422
rect 37096 419358 37148 419364
rect 15292 416832 15344 416838
rect 15292 416774 15344 416780
rect 26332 416832 26384 416838
rect 26332 416774 26384 416780
rect 36912 416832 36964 416838
rect 36912 416774 36964 416780
rect 15304 394738 15332 416774
rect 26344 414868 26372 416774
rect 15396 414310 16054 414338
rect 36662 414310 36860 414338
rect 15292 394732 15344 394738
rect 15292 394674 15344 394680
rect 15396 391950 15424 414310
rect 36728 414248 36780 414254
rect 36728 414190 36780 414196
rect 36740 394754 36768 414190
rect 36832 412826 36860 414310
rect 36924 414254 36952 416774
rect 36912 414248 36964 414254
rect 36912 414190 36964 414196
rect 36820 412820 36872 412826
rect 36820 412762 36872 412768
rect 36820 412616 36872 412622
rect 36820 412558 36872 412564
rect 16120 394732 16172 394738
rect 36662 394726 36768 394754
rect 16120 394674 16172 394680
rect 15488 394046 16054 394074
rect 15384 391944 15436 391950
rect 15384 391886 15436 391892
rect 15488 389450 15516 394046
rect 15212 389422 15516 389450
rect 15212 365702 15240 389422
rect 15384 389360 15436 389366
rect 15384 389302 15436 389308
rect 15396 383654 15424 389302
rect 16132 387954 16160 394674
rect 26344 391882 26372 394060
rect 26332 391876 26384 391882
rect 26332 391818 26384 391824
rect 36832 389842 36860 412558
rect 26608 389836 26660 389842
rect 26608 389778 26660 389784
rect 36820 389836 36872 389842
rect 36820 389778 36872 389784
rect 16132 387926 16330 387954
rect 26620 387940 26648 389778
rect 36938 387246 37320 387274
rect 37292 385490 37320 387246
rect 37280 385484 37332 385490
rect 37280 385426 37332 385432
rect 15396 383626 15976 383654
rect 15948 367690 15976 383626
rect 15948 367662 16330 367690
rect 15200 365696 15252 365702
rect 15200 365638 15252 365644
rect 26620 365634 26648 367132
rect 36924 365702 36952 367132
rect 36912 365696 36964 365702
rect 36912 365638 36964 365644
rect 26608 365628 26660 365634
rect 26608 365570 26660 365576
rect 36912 363044 36964 363050
rect 36912 362986 36964 362992
rect 15292 362976 15344 362982
rect 15292 362918 15344 362924
rect 26332 362976 26384 362982
rect 26332 362918 26384 362924
rect 15304 340202 15332 362918
rect 26344 360876 26372 362918
rect 36662 360590 36860 360618
rect 15396 360318 16054 360346
rect 15292 340196 15344 340202
rect 15292 340138 15344 340144
rect 15396 338094 15424 360318
rect 36832 355434 36860 360590
rect 36820 355428 36872 355434
rect 36820 355370 36872 355376
rect 36924 352594 36952 362986
rect 37004 355428 37056 355434
rect 37004 355370 37056 355376
rect 36740 352566 36952 352594
rect 36740 340762 36768 352566
rect 37016 347818 37044 355370
rect 36820 347812 36872 347818
rect 36820 347754 36872 347760
rect 37004 347812 37056 347818
rect 37004 347754 37056 347760
rect 36662 340734 36768 340762
rect 15488 340054 16054 340082
rect 15384 338088 15436 338094
rect 15384 338030 15436 338036
rect 15488 337770 15516 340054
rect 15936 339992 15988 339998
rect 15936 339934 15988 339940
rect 15212 337742 15516 337770
rect 15212 311846 15240 337742
rect 15384 335504 15436 335510
rect 15384 335446 15436 335452
rect 15396 325694 15424 335446
rect 15948 333962 15976 339934
rect 26344 338026 26372 340068
rect 26332 338020 26384 338026
rect 26332 337962 26384 337968
rect 36832 336054 36860 347754
rect 26608 336048 26660 336054
rect 26608 335990 26660 335996
rect 36820 336048 36872 336054
rect 36820 335990 36872 335996
rect 15948 333934 16330 333962
rect 26620 333948 26648 335990
rect 36938 333254 37320 333282
rect 37292 329526 37320 333254
rect 37280 329520 37332 329526
rect 37280 329462 37332 329468
rect 15396 325666 15976 325694
rect 15948 313698 15976 325666
rect 15948 313670 16330 313698
rect 15200 311840 15252 311846
rect 15200 311782 15252 311788
rect 26620 311778 26648 313140
rect 36924 311846 36952 313140
rect 36912 311840 36964 311846
rect 36912 311782 36964 311788
rect 26608 311772 26660 311778
rect 26608 311714 26660 311720
rect 36912 309256 36964 309262
rect 36912 309198 36964 309204
rect 15200 309188 15252 309194
rect 15200 309130 15252 309136
rect 26332 309188 26384 309194
rect 26332 309130 26384 309136
rect 13726 296304 13782 296313
rect 13726 296239 13782 296248
rect 13740 288017 13768 296239
rect 13726 288008 13782 288017
rect 13726 287943 13782 287952
rect 15212 283218 15240 309130
rect 26344 306884 26372 309130
rect 15580 306326 16054 306354
rect 36662 306326 36860 306354
rect 15580 296714 15608 306326
rect 36728 306264 36780 306270
rect 36728 306206 36780 306212
rect 15396 296686 15608 296714
rect 15396 284306 15424 296686
rect 36740 286770 36768 306206
rect 36832 305794 36860 306326
rect 36924 306270 36952 309198
rect 36912 306264 36964 306270
rect 36912 306206 36964 306212
rect 36820 305788 36872 305794
rect 36820 305730 36872 305736
rect 36820 305584 36872 305590
rect 36820 305526 36872 305532
rect 36662 286742 36768 286770
rect 15488 286062 16054 286090
rect 15384 284300 15436 284306
rect 15384 284242 15436 284248
rect 15200 283212 15252 283218
rect 15200 283154 15252 283160
rect 15488 281738 15516 286062
rect 26344 284238 26372 286076
rect 26332 284232 26384 284238
rect 26332 284174 26384 284180
rect 16028 283212 16080 283218
rect 16028 283154 16080 283160
rect 15304 281710 15516 281738
rect 15304 256698 15332 281710
rect 15384 281580 15436 281586
rect 15384 281522 15436 281528
rect 15396 267734 15424 281522
rect 16040 279970 16068 283154
rect 36832 282198 36860 305526
rect 26608 282192 26660 282198
rect 26608 282134 26660 282140
rect 36820 282192 36872 282198
rect 36820 282134 36872 282140
rect 16040 279942 16330 279970
rect 26620 279956 26648 282134
rect 36938 279262 37136 279290
rect 15396 267706 15976 267734
rect 15948 259706 15976 267706
rect 15948 259678 16330 259706
rect 15292 256692 15344 256698
rect 15292 256634 15344 256640
rect 26620 256630 26648 259148
rect 36924 256698 36952 259148
rect 37108 256698 37136 279262
rect 36912 256692 36964 256698
rect 36912 256634 36964 256640
rect 37096 256692 37148 256698
rect 37096 256634 37148 256640
rect 26608 256624 26660 256630
rect 26608 256566 26660 256572
rect 37648 255400 37700 255406
rect 37648 255342 37700 255348
rect 15200 255332 15252 255338
rect 15200 255274 15252 255280
rect 26332 255332 26384 255338
rect 26332 255274 26384 255280
rect 14464 240168 14516 240174
rect 14464 240110 14516 240116
rect 13728 38684 13780 38690
rect 13728 38626 13780 38632
rect 13634 27704 13690 27713
rect 13634 27639 13690 27648
rect 13740 26353 13768 38626
rect 14476 38554 14504 240110
rect 15212 227186 15240 255274
rect 26344 252892 26372 255274
rect 36662 252470 37044 252498
rect 15396 252334 16054 252362
rect 36728 252340 36780 252346
rect 15396 230450 15424 252334
rect 36728 252282 36780 252288
rect 36740 232778 36768 252282
rect 37016 248282 37044 252470
rect 37660 252346 37688 255342
rect 37648 252340 37700 252346
rect 37648 252282 37700 252288
rect 36662 232750 36768 232778
rect 36832 248254 37044 248282
rect 15580 232070 16054 232098
rect 15384 230444 15436 230450
rect 15384 230386 15436 230392
rect 15200 227180 15252 227186
rect 15200 227122 15252 227128
rect 15580 219434 15608 232070
rect 26344 230382 26372 232084
rect 26332 230376 26384 230382
rect 26332 230318 26384 230324
rect 36832 228410 36860 248254
rect 26608 228404 26660 228410
rect 26608 228346 26660 228352
rect 36820 228404 36872 228410
rect 36820 228346 36872 228352
rect 15936 227928 15988 227934
rect 15936 227870 15988 227876
rect 15304 219406 15608 219434
rect 15304 202842 15332 219406
rect 15948 205714 15976 227870
rect 16028 227180 16080 227186
rect 16028 227122 16080 227128
rect 16040 225978 16068 227122
rect 16040 225950 16330 225978
rect 26620 225964 26648 228346
rect 36938 225270 37320 225298
rect 37292 222358 37320 225270
rect 37280 222352 37332 222358
rect 37280 222294 37332 222300
rect 15948 205686 16330 205714
rect 15292 202836 15344 202842
rect 15292 202778 15344 202784
rect 26620 202774 26648 205020
rect 36924 202842 36952 205020
rect 36912 202836 36964 202842
rect 36912 202778 36964 202784
rect 26608 202768 26660 202774
rect 26608 202710 26660 202716
rect 37004 200252 37056 200258
rect 37004 200194 37056 200200
rect 15200 200184 15252 200190
rect 15200 200126 15252 200132
rect 26332 200184 26384 200190
rect 26332 200126 26384 200132
rect 15212 176050 15240 200126
rect 26344 198900 26372 200126
rect 36662 198478 36860 198506
rect 15396 198206 16054 198234
rect 15396 176662 15424 198206
rect 36832 195378 36860 198478
rect 36832 195350 36952 195378
rect 36820 195220 36872 195226
rect 36820 195162 36872 195168
rect 36832 195106 36860 195162
rect 36740 195078 36860 195106
rect 36740 178786 36768 195078
rect 36924 193214 36952 195350
rect 37016 195226 37044 200194
rect 37004 195220 37056 195226
rect 37004 195162 37056 195168
rect 36662 178758 36768 178786
rect 36832 193186 36952 193214
rect 15488 178078 16054 178106
rect 15384 176656 15436 176662
rect 15384 176598 15436 176604
rect 15200 176044 15252 176050
rect 15200 175986 15252 175992
rect 15488 174570 15516 178078
rect 26344 176594 26372 178092
rect 26332 176588 26384 176594
rect 26332 176530 26384 176536
rect 16028 176044 16080 176050
rect 16028 175986 16080 175992
rect 15304 174542 15516 174570
rect 15304 149054 15332 174542
rect 15384 174072 15436 174078
rect 15384 174014 15436 174020
rect 15396 171134 15424 174014
rect 16040 171986 16068 175986
rect 36832 174554 36860 193186
rect 26608 174548 26660 174554
rect 26608 174490 26660 174496
rect 36820 174548 36872 174554
rect 36820 174490 36872 174496
rect 16040 171958 16330 171986
rect 26620 171972 26648 174490
rect 36912 173936 36964 173942
rect 36912 173878 36964 173884
rect 36924 171972 36952 173878
rect 15396 171106 15976 171134
rect 15948 151722 15976 171106
rect 15948 151694 16330 151722
rect 15292 149048 15344 149054
rect 15292 148990 15344 148996
rect 26620 148986 26648 151028
rect 36924 149054 36952 151028
rect 36912 149048 36964 149054
rect 36912 148990 36964 148996
rect 26608 148980 26660 148986
rect 26608 148922 26660 148928
rect 15292 146328 15344 146334
rect 15292 146270 15344 146276
rect 26332 146328 26384 146334
rect 26332 146270 26384 146276
rect 15304 124710 15332 146270
rect 26344 144908 26372 146270
rect 15396 144214 16054 144242
rect 36662 144214 36768 144242
rect 15292 124704 15344 124710
rect 15292 124646 15344 124652
rect 15396 122670 15424 144214
rect 16120 124704 16172 124710
rect 16120 124646 16172 124652
rect 36544 124704 36596 124710
rect 36596 124652 36662 124658
rect 36544 124646 36662 124652
rect 15488 124086 16054 124114
rect 15384 122664 15436 122670
rect 15384 122606 15436 122612
rect 15488 117994 15516 124086
rect 15568 120284 15620 120290
rect 15568 120226 15620 120232
rect 15212 117966 15516 117994
rect 15212 95198 15240 117966
rect 15580 113174 15608 120226
rect 16132 117994 16160 124646
rect 36556 124630 36662 124646
rect 26344 122738 26372 124100
rect 26332 122732 26384 122738
rect 26332 122674 26384 122680
rect 36740 120766 36768 144214
rect 26608 120760 26660 120766
rect 26608 120702 26660 120708
rect 36728 120760 36780 120766
rect 36728 120702 36780 120708
rect 16132 117966 16330 117994
rect 26620 117980 26648 120702
rect 36912 120148 36964 120154
rect 36912 120090 36964 120096
rect 36924 117980 36952 120090
rect 15580 113146 15976 113174
rect 15948 97730 15976 113146
rect 15948 97702 16330 97730
rect 15200 95192 15252 95198
rect 15200 95134 15252 95140
rect 26620 95130 26648 97036
rect 36924 95198 36952 97036
rect 36912 95192 36964 95198
rect 36912 95134 36964 95140
rect 26608 95124 26660 95130
rect 26608 95066 26660 95072
rect 36912 92608 36964 92614
rect 36912 92550 36964 92556
rect 15200 92540 15252 92546
rect 15200 92482 15252 92488
rect 26332 92540 26384 92546
rect 26332 92482 26384 92488
rect 15212 69698 15240 92482
rect 26344 90916 26372 92482
rect 36662 90494 36860 90522
rect 15396 90222 16054 90250
rect 15200 69692 15252 69698
rect 15200 69634 15252 69640
rect 15396 69018 15424 90222
rect 36832 85066 36860 90494
rect 36820 85060 36872 85066
rect 36820 85002 36872 85008
rect 36924 82090 36952 92550
rect 37004 85060 37056 85066
rect 37004 85002 37056 85008
rect 36740 82062 36952 82090
rect 36740 70666 36768 82062
rect 37016 77314 37044 85002
rect 36820 77308 36872 77314
rect 36820 77250 36872 77256
rect 37004 77308 37056 77314
rect 37004 77250 37056 77256
rect 36662 70638 36768 70666
rect 15488 70094 16054 70122
rect 15384 69012 15436 69018
rect 15384 68954 15436 68960
rect 15488 67538 15516 70094
rect 16028 69692 16080 69698
rect 16028 69634 16080 69640
rect 15304 67510 15516 67538
rect 15304 41410 15332 67510
rect 15384 66428 15436 66434
rect 15384 66370 15436 66376
rect 15396 55214 15424 66370
rect 16040 63866 16068 69634
rect 26344 68950 26372 70108
rect 26332 68944 26384 68950
rect 26332 68886 26384 68892
rect 36832 66910 36860 77250
rect 26608 66904 26660 66910
rect 26608 66846 26660 66852
rect 36820 66904 36872 66910
rect 36820 66846 36872 66852
rect 16040 63838 16330 63866
rect 26620 63852 26648 66846
rect 36912 66292 36964 66298
rect 36912 66234 36964 66240
rect 36924 63852 36952 66234
rect 15396 55186 15976 55214
rect 15948 43738 15976 55186
rect 15948 43710 16330 43738
rect 15292 41404 15344 41410
rect 15292 41346 15344 41352
rect 26620 41342 26648 43044
rect 36924 41410 36952 43044
rect 36912 41404 36964 41410
rect 36912 41346 36964 41352
rect 26608 41336 26660 41342
rect 26608 41278 26660 41284
rect 37936 38622 37964 700742
rect 39304 687268 39356 687274
rect 39304 687210 39356 687216
rect 38658 674248 38714 674257
rect 38658 674183 38714 674192
rect 38016 659796 38068 659802
rect 38016 659738 38068 659744
rect 38028 634710 38056 659738
rect 38672 647737 38700 674183
rect 39316 662318 39344 687210
rect 39304 662312 39356 662318
rect 39304 662254 39356 662260
rect 38658 647728 38714 647737
rect 38658 647663 38714 647672
rect 38016 634704 38068 634710
rect 38016 634646 38068 634652
rect 39304 632120 39356 632126
rect 39304 632062 39356 632068
rect 38658 620256 38714 620265
rect 38658 620191 38714 620200
rect 38108 605872 38160 605878
rect 38108 605814 38160 605820
rect 38016 599752 38068 599758
rect 38016 599694 38068 599700
rect 38028 580990 38056 599694
rect 38016 580984 38068 580990
rect 38016 580926 38068 580932
rect 38120 580922 38148 605814
rect 38672 593745 38700 620191
rect 39316 608530 39344 632062
rect 39304 608524 39356 608530
rect 39304 608466 39356 608472
rect 38658 593736 38714 593745
rect 38658 593671 38714 593680
rect 38108 580916 38160 580922
rect 38108 580858 38160 580864
rect 39304 578264 39356 578270
rect 39304 578206 39356 578212
rect 38658 566264 38714 566273
rect 38658 566199 38714 566208
rect 38016 552084 38068 552090
rect 38016 552026 38068 552032
rect 38028 527066 38056 552026
rect 38108 548548 38160 548554
rect 38108 548490 38160 548496
rect 38120 527134 38148 548490
rect 38672 539753 38700 566199
rect 39316 554674 39344 578206
rect 39304 554668 39356 554674
rect 39304 554610 39356 554616
rect 38658 539744 38714 539753
rect 38658 539679 38714 539688
rect 38108 527128 38160 527134
rect 38108 527070 38160 527076
rect 38016 527060 38068 527066
rect 38016 527002 38068 527008
rect 38016 524476 38068 524482
rect 38016 524418 38068 524424
rect 38028 500886 38056 524418
rect 38658 512272 38714 512281
rect 38658 512207 38714 512216
rect 38016 500880 38068 500886
rect 38016 500822 38068 500828
rect 38108 498228 38160 498234
rect 38108 498170 38160 498176
rect 38016 492584 38068 492590
rect 38016 492526 38068 492532
rect 38028 473346 38056 492526
rect 38016 473340 38068 473346
rect 38016 473282 38068 473288
rect 38120 473278 38148 498170
rect 38672 485761 38700 512207
rect 38658 485752 38714 485761
rect 38658 485687 38714 485696
rect 38108 473272 38160 473278
rect 38108 473214 38160 473220
rect 38658 458280 38714 458289
rect 38658 458215 38714 458224
rect 38016 436620 38068 436626
rect 38016 436562 38068 436568
rect 38028 419490 38056 436562
rect 38672 431769 38700 458215
rect 38658 431760 38714 431769
rect 38658 431695 38714 431704
rect 38016 419484 38068 419490
rect 38016 419426 38068 419432
rect 38658 404288 38714 404297
rect 38658 404223 38714 404232
rect 38016 389224 38068 389230
rect 38016 389166 38068 389172
rect 38028 365634 38056 389166
rect 38108 385484 38160 385490
rect 38108 385426 38160 385432
rect 38120 365702 38148 385426
rect 38672 377777 38700 404223
rect 38658 377768 38714 377777
rect 38658 377703 38714 377712
rect 38108 365696 38160 365702
rect 38108 365638 38160 365644
rect 38016 365628 38068 365634
rect 38016 365570 38068 365576
rect 38016 362976 38068 362982
rect 38016 362918 38068 362924
rect 38028 338026 38056 362918
rect 38658 350296 38714 350305
rect 38658 350231 38714 350240
rect 38016 338020 38068 338026
rect 38016 337962 38068 337968
rect 38016 335368 38068 335374
rect 38016 335310 38068 335316
rect 38028 311778 38056 335310
rect 38108 329520 38160 329526
rect 38108 329462 38160 329468
rect 38120 311846 38148 329462
rect 38672 323785 38700 350231
rect 38658 323776 38714 323785
rect 38658 323711 38714 323720
rect 38108 311840 38160 311846
rect 38108 311782 38160 311788
rect 38016 311772 38068 311778
rect 38016 311714 38068 311720
rect 38016 309188 38068 309194
rect 38016 309130 38068 309136
rect 38028 284238 38056 309130
rect 38658 296304 38714 296313
rect 38658 296239 38714 296248
rect 38016 284232 38068 284238
rect 38016 284174 38068 284180
rect 38016 281648 38068 281654
rect 38016 281590 38068 281596
rect 38028 256630 38056 281590
rect 38672 269793 38700 296239
rect 38658 269784 38714 269793
rect 38658 269719 38714 269728
rect 38016 256624 38068 256630
rect 38016 256566 38068 256572
rect 38108 255332 38160 255338
rect 38108 255274 38160 255280
rect 38016 231872 38068 231878
rect 38016 231814 38068 231820
rect 26976 38616 27028 38622
rect 26976 38558 27028 38564
rect 37924 38616 37976 38622
rect 37924 38558 37976 38564
rect 14464 38548 14516 38554
rect 14464 38490 14516 38496
rect 22468 38412 22520 38418
rect 22468 38354 22520 38360
rect 23756 38412 23808 38418
rect 23756 38354 23808 38360
rect 19248 38344 19300 38350
rect 19248 38286 19300 38292
rect 17316 38004 17368 38010
rect 17316 37946 17368 37952
rect 16028 37936 16080 37942
rect 16028 37878 16080 37884
rect 16040 35972 16068 37878
rect 17328 35972 17356 37946
rect 19260 35972 19288 38286
rect 20536 38072 20588 38078
rect 20536 38014 20588 38020
rect 20548 35972 20576 38014
rect 22480 35972 22508 38354
rect 23768 35972 23796 38354
rect 25688 38072 25740 38078
rect 25688 38014 25740 38020
rect 25700 35972 25728 38014
rect 26988 35972 27016 38558
rect 33416 38480 33468 38486
rect 33416 38422 33468 38428
rect 30196 38208 30248 38214
rect 30196 38150 30248 38156
rect 32128 38208 32180 38214
rect 32128 38150 32180 38156
rect 28736 35970 28934 35986
rect 30208 35972 30236 38150
rect 32140 35972 32168 38150
rect 33428 35972 33456 38422
rect 38028 37398 38056 231814
rect 38120 230382 38148 255274
rect 38658 242312 38714 242321
rect 38658 242247 38714 242256
rect 38108 230376 38160 230382
rect 38108 230318 38160 230324
rect 38108 227792 38160 227798
rect 38108 227734 38160 227740
rect 38120 202774 38148 227734
rect 38200 222352 38252 222358
rect 38200 222294 38252 222300
rect 38212 202842 38240 222294
rect 38672 215801 38700 242247
rect 38658 215792 38714 215801
rect 38658 215727 38714 215736
rect 38200 202836 38252 202842
rect 38200 202778 38252 202784
rect 38108 202768 38160 202774
rect 38108 202710 38160 202716
rect 38108 200184 38160 200190
rect 38108 200126 38160 200132
rect 38120 176594 38148 200126
rect 38658 188320 38714 188329
rect 38658 188255 38714 188264
rect 38108 176588 38160 176594
rect 38108 176530 38160 176536
rect 38672 161809 38700 188255
rect 38658 161800 38714 161809
rect 38658 161735 38714 161744
rect 38200 146396 38252 146402
rect 38200 146338 38252 146344
rect 38108 146328 38160 146334
rect 38108 146270 38160 146276
rect 38120 122738 38148 146270
rect 38212 124710 38240 146338
rect 38658 134328 38714 134337
rect 38658 134263 38714 134272
rect 38200 124704 38252 124710
rect 38200 124646 38252 124652
rect 38108 122732 38160 122738
rect 38108 122674 38160 122680
rect 38672 107817 38700 134263
rect 38658 107808 38714 107817
rect 38658 107743 38714 107752
rect 38108 92540 38160 92546
rect 38108 92482 38160 92488
rect 38120 68950 38148 92482
rect 38658 80336 38714 80345
rect 38658 80271 38714 80280
rect 38108 68944 38160 68950
rect 38108 68886 38160 68892
rect 38672 53825 38700 80271
rect 38658 53816 38714 53825
rect 38658 53751 38714 53760
rect 38568 38548 38620 38554
rect 38568 38490 38620 38496
rect 35348 37392 35400 37398
rect 35348 37334 35400 37340
rect 38016 37392 38068 37398
rect 38016 37334 38068 37340
rect 35360 35972 35388 37334
rect 36636 37324 36688 37330
rect 36636 37266 36688 37272
rect 36648 35972 36676 37266
rect 38580 35972 38608 38490
rect 40052 37398 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 65616 700732 65668 700738
rect 65616 700674 65668 700680
rect 65524 700392 65576 700398
rect 65524 700334 65576 700340
rect 54300 687336 54352 687342
rect 54300 687278 54352 687284
rect 54312 684964 54340 687278
rect 64604 687268 64656 687274
rect 64604 687210 64656 687216
rect 64616 684964 64644 687210
rect 42904 684270 44022 684298
rect 42706 674248 42762 674257
rect 42706 674183 42762 674192
rect 42720 665174 42748 674183
rect 42708 665168 42760 665174
rect 42708 665110 42760 665116
rect 42904 662318 42932 684270
rect 64880 669112 64932 669118
rect 64880 669054 64932 669060
rect 64892 664714 64920 669054
rect 64630 664686 64920 664714
rect 43640 664006 44022 664034
rect 54326 664006 54616 664034
rect 43640 662386 43668 664006
rect 43628 662380 43680 662386
rect 43628 662322 43680 662328
rect 42892 662312 42944 662318
rect 42892 662254 42944 662260
rect 54588 662250 54616 664006
rect 54576 662244 54628 662250
rect 54576 662186 54628 662192
rect 44180 659796 44232 659802
rect 44180 659738 44232 659744
rect 44192 657914 44220 659738
rect 54300 659728 54352 659734
rect 54300 659670 54352 659676
rect 54312 657914 54340 659670
rect 44192 657886 44344 657914
rect 54312 657886 54648 657914
rect 64952 657206 65104 657234
rect 42708 656940 42760 656946
rect 42708 656882 42760 656888
rect 42720 647737 42748 656882
rect 42706 647728 42762 647737
rect 42706 647663 42762 647672
rect 44344 637078 44680 637106
rect 54648 637078 54984 637106
rect 44652 634817 44680 637078
rect 44638 634808 44694 634817
rect 44638 634743 44694 634752
rect 54956 634710 54984 637078
rect 64938 636834 64966 637092
rect 64892 636806 64966 636834
rect 64892 634778 64920 636806
rect 65076 634778 65104 657206
rect 64880 634772 64932 634778
rect 64880 634714 64932 634720
rect 65064 634772 65116 634778
rect 65064 634714 65116 634720
rect 54944 634704 54996 634710
rect 54944 634646 54996 634652
rect 54300 632188 54352 632194
rect 54300 632130 54352 632136
rect 54312 630972 54340 632130
rect 64604 632120 64656 632126
rect 64604 632062 64656 632068
rect 64616 630972 64644 632062
rect 42904 630278 44022 630306
rect 42706 620256 42762 620265
rect 42706 620191 42762 620200
rect 42720 611318 42748 620191
rect 42708 611312 42760 611318
rect 42708 611254 42760 611260
rect 42904 608530 42932 630278
rect 64880 613148 64932 613154
rect 64880 613090 64932 613096
rect 64892 610722 64920 613090
rect 64630 610694 64920 610722
rect 44008 608598 44036 610028
rect 43996 608592 44048 608598
rect 43996 608534 44048 608540
rect 42892 608524 42944 608530
rect 42892 608466 42944 608472
rect 54312 608394 54340 610028
rect 54300 608388 54352 608394
rect 54300 608330 54352 608336
rect 54300 606008 54352 606014
rect 54300 605950 54352 605956
rect 44180 605872 44232 605878
rect 44180 605814 44232 605820
rect 44192 603922 44220 605814
rect 54312 603922 54340 605950
rect 44192 603894 44344 603922
rect 54312 603894 54648 603922
rect 64952 603214 65104 603242
rect 42706 602168 42762 602177
rect 42706 602103 42762 602112
rect 42720 593745 42748 602103
rect 42706 593736 42762 593745
rect 42706 593671 42762 593680
rect 44344 583086 44680 583114
rect 54648 583086 54892 583114
rect 44652 580922 44680 583086
rect 44640 580916 44692 580922
rect 44640 580858 44692 580864
rect 54864 580854 54892 583086
rect 64938 582842 64966 583100
rect 64892 582814 64966 582842
rect 64892 580990 64920 582814
rect 65076 580990 65104 603214
rect 64880 580984 64932 580990
rect 64880 580926 64932 580932
rect 65064 580984 65116 580990
rect 65064 580926 65116 580932
rect 54852 580848 54904 580854
rect 54852 580790 54904 580796
rect 53932 578332 53984 578338
rect 53932 578274 53984 578280
rect 53944 576994 53972 578274
rect 64236 578264 64288 578270
rect 64236 578206 64288 578212
rect 64248 576994 64276 578206
rect 53944 576966 54326 576994
rect 64248 576966 64630 576994
rect 42904 576286 44022 576314
rect 42706 566264 42762 566273
rect 42706 566199 42762 566208
rect 42720 557530 42748 566199
rect 42708 557524 42760 557530
rect 42708 557466 42760 557472
rect 42904 554674 42932 576286
rect 64880 562352 64932 562358
rect 64880 562294 64932 562300
rect 64892 556730 64920 562294
rect 64630 556702 64920 556730
rect 44008 554742 44036 556036
rect 43996 554736 44048 554742
rect 43996 554678 44048 554684
rect 42892 554668 42944 554674
rect 42892 554610 42944 554616
rect 54312 554538 54340 556036
rect 54300 554532 54352 554538
rect 54300 554474 54352 554480
rect 54300 552220 54352 552226
rect 54300 552162 54352 552168
rect 44180 552084 44232 552090
rect 44180 552026 44232 552032
rect 44192 549930 44220 552026
rect 54312 549930 54340 552162
rect 44192 549902 44344 549930
rect 54312 549902 54648 549930
rect 64952 549222 65104 549250
rect 42706 548176 42762 548185
rect 42706 548111 42762 548120
rect 42720 539753 42748 548111
rect 42706 539744 42762 539753
rect 42706 539679 42762 539688
rect 44344 529094 44680 529122
rect 54648 529094 54984 529122
rect 44652 527066 44680 529094
rect 44640 527060 44692 527066
rect 44640 527002 44692 527008
rect 54956 526998 54984 529094
rect 64938 528850 64966 529108
rect 64892 528822 64966 528850
rect 64892 527134 64920 528822
rect 65076 527134 65104 549222
rect 64880 527128 64932 527134
rect 64880 527070 64932 527076
rect 65064 527128 65116 527134
rect 65064 527070 65116 527076
rect 54944 526992 54996 526998
rect 54944 526934 54996 526940
rect 54300 524544 54352 524550
rect 54300 524486 54352 524492
rect 54312 522852 54340 524486
rect 64604 524476 64656 524482
rect 64604 524418 64656 524424
rect 64616 522852 64644 524418
rect 42904 522294 44022 522322
rect 42904 500886 42932 522294
rect 64880 503260 64932 503266
rect 64880 503202 64932 503208
rect 64892 502330 64920 503202
rect 64630 502302 64920 502330
rect 44008 500954 44036 502044
rect 43996 500948 44048 500954
rect 43996 500890 44048 500896
rect 42892 500880 42944 500886
rect 42892 500822 42944 500828
rect 54312 500750 54340 502044
rect 54300 500744 54352 500750
rect 54300 500686 54352 500692
rect 54300 498364 54352 498370
rect 54300 498306 54352 498312
rect 44180 498228 44232 498234
rect 44180 498170 44232 498176
rect 44192 495938 44220 498170
rect 54312 495938 54340 498306
rect 44192 495910 44344 495938
rect 54312 495910 54648 495938
rect 64952 495230 65104 495258
rect 42706 485752 42762 485761
rect 42706 485687 42762 485696
rect 42720 477193 42748 485687
rect 42706 477184 42762 477193
rect 42706 477119 42762 477128
rect 44344 475102 44680 475130
rect 54648 475102 54984 475130
rect 44652 473278 44680 475102
rect 44640 473272 44692 473278
rect 44640 473214 44692 473220
rect 54956 473210 54984 475102
rect 64938 474858 64966 475116
rect 64892 474830 64966 474858
rect 64892 473346 64920 474830
rect 65076 473346 65104 495230
rect 64880 473340 64932 473346
rect 64880 473282 64932 473288
rect 65064 473340 65116 473346
rect 65064 473282 65116 473288
rect 54944 473204 54996 473210
rect 54944 473146 54996 473152
rect 54300 470620 54352 470626
rect 54300 470562 54352 470568
rect 54312 468860 54340 470562
rect 42904 468302 44022 468330
rect 64630 468302 64828 468330
rect 42904 445602 42932 468302
rect 44008 445738 44036 448052
rect 54312 445738 54340 448052
rect 43996 445732 44048 445738
rect 43996 445674 44048 445680
rect 54300 445732 54352 445738
rect 54300 445674 54352 445680
rect 64616 445641 64644 448052
rect 64800 445670 64828 468302
rect 64788 445664 64840 445670
rect 64602 445632 64658 445641
rect 42892 445596 42944 445602
rect 64788 445606 64840 445612
rect 64602 445567 64658 445576
rect 42892 445538 42944 445544
rect 54300 444508 54352 444514
rect 54300 444450 54352 444456
rect 54312 441946 54340 444450
rect 54312 441918 54648 441946
rect 44192 441238 44344 441266
rect 64952 441238 65104 441266
rect 44192 438938 44220 441238
rect 44180 438932 44232 438938
rect 44180 438874 44232 438880
rect 42706 431760 42762 431769
rect 42706 431695 42762 431704
rect 42720 423201 42748 431695
rect 42706 423192 42762 423201
rect 42706 423127 42762 423136
rect 44344 421110 44680 421138
rect 54648 421110 54984 421138
rect 44652 419422 44680 421110
rect 44640 419416 44692 419422
rect 44640 419358 44692 419364
rect 54956 419354 54984 421110
rect 64938 420866 64966 421124
rect 64892 420838 64966 420866
rect 64892 419490 64920 420838
rect 65076 419490 65104 441238
rect 64880 419484 64932 419490
rect 64880 419426 64932 419432
rect 65064 419484 65116 419490
rect 65064 419426 65116 419432
rect 54944 419348 54996 419354
rect 54944 419290 54996 419296
rect 54300 416832 54352 416838
rect 54300 416774 54352 416780
rect 54312 414868 54340 416774
rect 42904 414310 44022 414338
rect 64630 414310 64828 414338
rect 42904 391814 42932 414310
rect 44008 391950 44036 394060
rect 54312 391950 54340 394060
rect 43996 391944 44048 391950
rect 43996 391886 44048 391892
rect 54300 391944 54352 391950
rect 64616 391921 64644 394060
rect 54300 391886 54352 391892
rect 64602 391912 64658 391921
rect 64800 391882 64828 414310
rect 64602 391847 64658 391856
rect 64788 391876 64840 391882
rect 64788 391818 64840 391824
rect 42892 391808 42944 391814
rect 42892 391750 42944 391756
rect 54300 389360 54352 389366
rect 54300 389302 54352 389308
rect 44180 389224 44232 389230
rect 44180 389166 44232 389172
rect 44192 387954 44220 389166
rect 54312 387954 54340 389302
rect 44192 387926 44344 387954
rect 54312 387926 54648 387954
rect 64952 387246 65104 387274
rect 42706 377768 42762 377777
rect 42706 377703 42762 377712
rect 42720 368490 42748 377703
rect 42708 368484 42760 368490
rect 42708 368426 42760 368432
rect 44344 367118 44680 367146
rect 54648 367118 54984 367146
rect 44652 365634 44680 367118
rect 44640 365628 44692 365634
rect 44640 365570 44692 365576
rect 54956 365566 54984 367118
rect 64938 366874 64966 367132
rect 64892 366846 64966 366874
rect 64892 365702 64920 366846
rect 65076 365702 65104 387246
rect 64880 365696 64932 365702
rect 64880 365638 64932 365644
rect 65064 365696 65116 365702
rect 65064 365638 65116 365644
rect 54944 365560 54996 365566
rect 54944 365502 54996 365508
rect 54300 363044 54352 363050
rect 54300 362986 54352 362992
rect 54312 360876 54340 362986
rect 64604 362976 64656 362982
rect 64604 362918 64656 362924
rect 64616 360876 64644 362918
rect 42904 360318 44022 360346
rect 42904 338026 42932 360318
rect 64880 342916 64932 342922
rect 64880 342858 64932 342864
rect 64892 340762 64920 342858
rect 64630 340734 64920 340762
rect 44008 338094 44036 340068
rect 43996 338088 44048 338094
rect 43996 338030 44048 338036
rect 42892 338020 42944 338026
rect 42892 337962 42944 337968
rect 54312 337890 54340 340068
rect 54300 337884 54352 337890
rect 54300 337826 54352 337832
rect 54300 335504 54352 335510
rect 54300 335446 54352 335452
rect 44180 335368 44232 335374
rect 44180 335310 44232 335316
rect 44192 333962 44220 335310
rect 54312 333962 54340 335446
rect 44192 333934 44344 333962
rect 54312 333934 54648 333962
rect 64952 333254 65104 333282
rect 42708 332648 42760 332654
rect 42708 332590 42760 332596
rect 42720 323785 42748 332590
rect 42706 323776 42762 323785
rect 42706 323711 42762 323720
rect 44344 313126 44680 313154
rect 54648 313126 54984 313154
rect 44652 311778 44680 313126
rect 44640 311772 44692 311778
rect 44640 311714 44692 311720
rect 54956 311710 54984 313126
rect 64938 312882 64966 313140
rect 64892 312854 64966 312882
rect 64892 311846 64920 312854
rect 65076 311846 65104 333254
rect 64880 311840 64932 311846
rect 64880 311782 64932 311788
rect 65064 311840 65116 311846
rect 65064 311782 65116 311788
rect 54944 311704 54996 311710
rect 54944 311646 54996 311652
rect 54300 309256 54352 309262
rect 54300 309198 54352 309204
rect 54312 306884 54340 309198
rect 64604 309188 64656 309194
rect 64604 309130 64656 309136
rect 64616 306884 64644 309130
rect 43548 306326 44022 306354
rect 43548 296714 43576 306326
rect 42904 296686 43576 296714
rect 42904 284238 42932 296686
rect 64880 291916 64932 291922
rect 64880 291858 64932 291864
rect 64892 286770 64920 291858
rect 64630 286742 64920 286770
rect 44008 284306 44036 286076
rect 43996 284300 44048 284306
rect 43996 284242 44048 284248
rect 42892 284232 42944 284238
rect 42892 284174 42944 284180
rect 54312 284102 54340 286076
rect 54300 284096 54352 284102
rect 54300 284038 54352 284044
rect 44180 281648 44232 281654
rect 44180 281590 44232 281596
rect 44192 279970 44220 281590
rect 54300 281580 54352 281586
rect 54300 281522 54352 281528
rect 54312 279970 54340 281522
rect 44192 279942 44344 279970
rect 54312 279942 54648 279970
rect 64952 279262 65104 279290
rect 42708 278792 42760 278798
rect 42708 278734 42760 278740
rect 42720 269793 42748 278734
rect 42706 269784 42762 269793
rect 42706 269719 42762 269728
rect 44344 259134 44680 259162
rect 54648 259134 54984 259162
rect 44652 256601 44680 259134
rect 54956 256630 54984 259134
rect 64938 258890 64966 259148
rect 64892 258862 64966 258890
rect 64892 256698 64920 258862
rect 65076 256698 65104 279262
rect 64880 256692 64932 256698
rect 64880 256634 64932 256640
rect 65064 256692 65116 256698
rect 65064 256634 65116 256640
rect 54944 256624 54996 256630
rect 44638 256592 44694 256601
rect 54944 256566 54996 256572
rect 44638 256527 44694 256536
rect 54300 255400 54352 255406
rect 54300 255342 54352 255348
rect 54312 252892 54340 255342
rect 64604 255332 64656 255338
rect 64604 255274 64656 255280
rect 64616 252892 64644 255274
rect 42904 252334 44022 252362
rect 42706 242312 42762 242321
rect 42706 242247 42762 242256
rect 42720 233238 42748 242247
rect 42708 233232 42760 233238
rect 42708 233174 42760 233180
rect 42904 230382 42932 252334
rect 64880 235748 64932 235754
rect 64880 235690 64932 235696
rect 64892 232778 64920 235690
rect 64630 232750 64920 232778
rect 44008 230450 44036 232084
rect 43996 230444 44048 230450
rect 43996 230386 44048 230392
rect 42892 230376 42944 230382
rect 42892 230318 42944 230324
rect 54312 230246 54340 232084
rect 54300 230240 54352 230246
rect 54300 230182 54352 230188
rect 54300 227928 54352 227934
rect 54300 227870 54352 227876
rect 44180 227792 44232 227798
rect 44180 227734 44232 227740
rect 44192 225978 44220 227734
rect 54312 225978 54340 227870
rect 44192 225950 44344 225978
rect 54312 225950 54648 225978
rect 64952 225270 65104 225298
rect 42706 224224 42762 224233
rect 42706 224159 42762 224168
rect 42720 215801 42748 224159
rect 42706 215792 42762 215801
rect 42706 215727 42762 215736
rect 44344 205006 44680 205034
rect 54648 205006 54892 205034
rect 44652 202774 44680 205006
rect 44640 202768 44692 202774
rect 44640 202710 44692 202716
rect 54864 202706 54892 205006
rect 64938 204762 64966 205020
rect 64892 204734 64966 204762
rect 64892 202842 64920 204734
rect 65076 202842 65104 225270
rect 64880 202836 64932 202842
rect 64880 202778 64932 202784
rect 65064 202836 65116 202842
rect 65064 202778 65116 202784
rect 54852 202700 54904 202706
rect 54852 202642 54904 202648
rect 54300 200252 54352 200258
rect 54300 200194 54352 200200
rect 54312 198900 54340 200194
rect 64604 200184 64656 200190
rect 64604 200126 64656 200132
rect 64616 198900 64644 200126
rect 42904 198206 44022 198234
rect 42706 188320 42762 188329
rect 42706 188255 42762 188264
rect 42720 179382 42748 188255
rect 42708 179376 42760 179382
rect 42708 179318 42760 179324
rect 42904 176594 42932 198206
rect 64880 185632 64932 185638
rect 64880 185574 64932 185580
rect 64892 178786 64920 185574
rect 64630 178758 64920 178786
rect 44008 176662 44036 178092
rect 43996 176656 44048 176662
rect 43996 176598 44048 176604
rect 42892 176588 42944 176594
rect 42892 176530 42944 176536
rect 54312 176526 54340 178092
rect 54300 176520 54352 176526
rect 54300 176462 54352 176468
rect 54300 174072 54352 174078
rect 54300 174014 54352 174020
rect 43444 173936 43496 173942
rect 43444 173878 43496 173884
rect 40684 171216 40736 171222
rect 40684 171158 40736 171164
rect 40696 148986 40724 171158
rect 42706 170096 42762 170105
rect 42706 170031 42762 170040
rect 42720 161809 42748 170031
rect 42706 161800 42762 161809
rect 42706 161735 42762 161744
rect 43456 148986 43484 173878
rect 54312 171986 54340 174014
rect 54312 171958 54648 171986
rect 44192 171278 44344 171306
rect 64952 171278 65104 171306
rect 44192 171222 44220 171278
rect 44180 171216 44232 171222
rect 44180 171158 44232 171164
rect 44344 151014 44680 151042
rect 54648 151014 54892 151042
rect 40684 148980 40736 148986
rect 40684 148922 40736 148928
rect 43444 148980 43496 148986
rect 43444 148922 43496 148928
rect 44652 148850 44680 151014
rect 54864 148918 54892 151014
rect 64938 150770 64966 151028
rect 64892 150742 64966 150770
rect 64892 148986 64920 150742
rect 65076 149054 65104 171278
rect 65064 149048 65116 149054
rect 65064 148990 65116 148996
rect 64880 148980 64932 148986
rect 64880 148922 64932 148928
rect 54852 148912 54904 148918
rect 54852 148854 54904 148860
rect 44640 148844 44692 148850
rect 44640 148786 44692 148792
rect 54300 146396 54352 146402
rect 54300 146338 54352 146344
rect 54312 144908 54340 146338
rect 64604 146328 64656 146334
rect 64604 146270 64656 146276
rect 64616 144908 64644 146270
rect 42904 144214 44022 144242
rect 42706 134328 42762 134337
rect 42706 134263 42762 134272
rect 42720 125594 42748 134263
rect 42708 125588 42760 125594
rect 42708 125530 42760 125536
rect 42904 122738 42932 144214
rect 64880 128648 64932 128654
rect 64880 128590 64932 128596
rect 64892 124794 64920 128590
rect 64630 124766 64920 124794
rect 42892 122732 42944 122738
rect 42892 122674 42944 122680
rect 44008 122670 44036 124100
rect 54312 122670 54340 124100
rect 43996 122664 44048 122670
rect 43996 122606 44048 122612
rect 54300 122664 54352 122670
rect 54300 122606 54352 122612
rect 54300 120284 54352 120290
rect 54300 120226 54352 120232
rect 43444 120148 43496 120154
rect 43444 120090 43496 120096
rect 40684 117292 40736 117298
rect 40684 117234 40736 117240
rect 40696 95130 40724 117234
rect 42706 116240 42762 116249
rect 42706 116175 42762 116184
rect 42720 107817 42748 116175
rect 42706 107808 42762 107817
rect 42706 107743 42762 107752
rect 43456 95130 43484 120090
rect 54312 117994 54340 120226
rect 54312 117966 54648 117994
rect 44100 117298 44344 117314
rect 44088 117292 44344 117298
rect 44140 117286 44344 117292
rect 64952 117286 65104 117314
rect 44088 117234 44140 117240
rect 44344 97022 44680 97050
rect 54648 97022 54984 97050
rect 40684 95124 40736 95130
rect 40684 95066 40736 95072
rect 43444 95124 43496 95130
rect 43444 95066 43496 95072
rect 44652 94994 44680 97022
rect 54956 95062 54984 97022
rect 64938 96778 64966 97036
rect 64892 96750 64966 96778
rect 64892 95130 64920 96750
rect 65076 95198 65104 117286
rect 65064 95192 65116 95198
rect 65064 95134 65116 95140
rect 64880 95124 64932 95130
rect 64880 95066 64932 95072
rect 54944 95056 54996 95062
rect 54944 94998 54996 95004
rect 44640 94988 44692 94994
rect 44640 94930 44692 94936
rect 54300 92608 54352 92614
rect 54300 92550 54352 92556
rect 54312 90916 54340 92550
rect 64604 92540 64656 92546
rect 64604 92482 64656 92488
rect 64616 90916 64644 92482
rect 42904 90222 44022 90250
rect 42904 68882 42932 90222
rect 64880 72616 64932 72622
rect 64880 72558 64932 72564
rect 64892 70666 64920 72558
rect 64630 70638 64920 70666
rect 44008 69018 44036 70108
rect 43996 69012 44048 69018
rect 43996 68954 44048 68960
rect 54312 68950 54340 70108
rect 54300 68944 54352 68950
rect 54300 68886 54352 68892
rect 42892 68876 42944 68882
rect 42892 68818 42944 68824
rect 54300 66428 54352 66434
rect 54300 66370 54352 66376
rect 43444 66292 43496 66298
rect 43444 66234 43496 66240
rect 40684 63300 40736 63306
rect 40684 63242 40736 63248
rect 40696 41342 40724 63242
rect 42706 53816 42762 53825
rect 42706 53751 42762 53760
rect 42720 45257 42748 53751
rect 42706 45248 42762 45257
rect 42706 45183 42762 45192
rect 43456 41342 43484 66234
rect 54312 63866 54340 66370
rect 54312 63838 54648 63866
rect 44008 63306 44344 63322
rect 43996 63300 44344 63306
rect 44048 63294 44344 63300
rect 64952 63294 65104 63322
rect 43996 63242 44048 63248
rect 44344 43030 44680 43058
rect 54648 43030 54984 43058
rect 40684 41336 40736 41342
rect 40684 41278 40736 41284
rect 43444 41336 43496 41342
rect 43444 41278 43496 41284
rect 44652 41206 44680 43030
rect 54956 41274 54984 43030
rect 64938 42786 64966 43044
rect 64892 42758 64966 42786
rect 64892 41342 64920 42758
rect 65076 41410 65104 63294
rect 65064 41404 65116 41410
rect 65064 41346 65116 41352
rect 64880 41336 64932 41342
rect 64880 41278 64932 41284
rect 54944 41268 54996 41274
rect 54944 41210 54996 41216
rect 44640 41200 44692 41206
rect 44640 41142 44692 41148
rect 46940 39432 46992 39438
rect 46940 39374 46992 39380
rect 41788 39364 41840 39370
rect 41788 39306 41840 39312
rect 40040 37392 40092 37398
rect 40040 37334 40092 37340
rect 39856 36100 39908 36106
rect 39856 36042 39908 36048
rect 39868 35972 39896 36042
rect 41800 35972 41828 39306
rect 45008 38140 45060 38146
rect 45008 38082 45060 38088
rect 43444 36032 43496 36038
rect 43496 35980 43746 35986
rect 43444 35974 43746 35980
rect 28724 35964 28934 35970
rect 28776 35958 28934 35964
rect 43456 35958 43746 35974
rect 45020 35972 45048 38082
rect 46952 35972 46980 39374
rect 61108 39364 61160 39370
rect 61108 39306 61160 39312
rect 56600 38752 56652 38758
rect 56600 38694 56652 38700
rect 54668 38276 54720 38282
rect 54668 38218 54720 38224
rect 51448 38140 51500 38146
rect 51448 38082 51500 38088
rect 48228 37392 48280 37398
rect 48228 37334 48280 37340
rect 48240 35972 48268 37334
rect 50528 36032 50580 36038
rect 50186 35980 50528 35986
rect 50186 35974 50580 35980
rect 50186 35958 50568 35974
rect 51460 35972 51488 38082
rect 53378 37904 53434 37913
rect 53378 37839 53434 37848
rect 53392 35972 53420 37839
rect 54680 35972 54708 38218
rect 56612 35972 56640 38694
rect 57888 38480 57940 38486
rect 57888 38422 57940 38428
rect 57900 35972 57928 38422
rect 59820 37392 59872 37398
rect 59820 37334 59872 37340
rect 59832 35972 59860 37334
rect 61120 35972 61148 39306
rect 64604 38276 64656 38282
rect 64604 38218 64656 38224
rect 64512 36848 64564 36854
rect 64512 36790 64564 36796
rect 64236 36780 64288 36786
rect 64236 36722 64288 36728
rect 61384 36100 61436 36106
rect 61384 36042 61436 36048
rect 28724 35906 28776 35912
rect 61292 35216 61344 35222
rect 61292 35158 61344 35164
rect 61304 34377 61332 35158
rect 61290 34368 61346 34377
rect 61290 34303 61346 34312
rect 13726 26344 13782 26353
rect 13726 26279 13782 26288
rect 13726 24168 13782 24177
rect 13726 24103 13782 24112
rect 12440 23452 12492 23458
rect 12440 23394 12492 23400
rect 12452 22953 12480 23394
rect 12438 22944 12494 22953
rect 12438 22879 12494 22888
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 12452 20913 12480 22034
rect 12438 20904 12494 20913
rect 12438 20839 12494 20848
rect 12440 20664 12492 20670
rect 12440 20606 12492 20612
rect 12452 19553 12480 20606
rect 12438 19544 12494 19553
rect 12438 19479 12494 19488
rect 12440 17944 12492 17950
rect 12440 17886 12492 17892
rect 12452 17513 12480 17886
rect 12438 17504 12494 17513
rect 12438 17439 12494 17448
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 8944 13048 8996 13054
rect 8944 12990 8996 12996
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 13740 3534 13768 24103
rect 16040 13802 16068 16116
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 17328 13734 17356 16116
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 19260 13394 19288 16116
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 20548 12986 20576 16116
rect 22480 15094 22508 16116
rect 22468 15088 22520 15094
rect 22468 15030 22520 15036
rect 23768 15026 23796 16116
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 25700 13598 25728 16116
rect 25688 13592 25740 13598
rect 25688 13534 25740 13540
rect 26988 13326 27016 16116
rect 28920 13666 28948 16116
rect 28908 13660 28960 13666
rect 28908 13602 28960 13608
rect 26976 13320 27028 13326
rect 26976 13262 27028 13268
rect 30208 13054 30236 16116
rect 32140 13666 32168 16116
rect 32128 13660 32180 13666
rect 32128 13602 32180 13608
rect 33428 13122 33456 16116
rect 35360 15162 35388 16116
rect 35348 15156 35400 15162
rect 35348 15098 35400 15104
rect 36648 13598 36676 16116
rect 36636 13592 36688 13598
rect 36636 13534 36688 13540
rect 38580 13122 38608 16116
rect 33416 13116 33468 13122
rect 33416 13058 33468 13064
rect 38568 13116 38620 13122
rect 38568 13058 38620 13064
rect 39868 13054 39896 16116
rect 41800 15162 41828 16116
rect 41788 15156 41840 15162
rect 41788 15098 41840 15104
rect 43088 13530 43116 16116
rect 45020 13705 45048 16116
rect 45006 13696 45062 13705
rect 45006 13631 45062 13640
rect 43076 13524 43128 13530
rect 43076 13466 43128 13472
rect 30196 13048 30248 13054
rect 30196 12990 30248 12996
rect 39856 13048 39908 13054
rect 39856 12990 39908 12996
rect 20536 12980 20588 12986
rect 20536 12922 20588 12928
rect 46308 12918 46336 16116
rect 48240 14958 48268 16116
rect 48332 16102 49542 16130
rect 48228 14952 48280 14958
rect 48228 14894 48280 14900
rect 46296 12912 46348 12918
rect 46296 12854 46348 12860
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 48332 3466 48360 16102
rect 51460 12850 51488 16116
rect 52748 15094 52776 16116
rect 52736 15088 52788 15094
rect 52736 15030 52788 15036
rect 54680 13190 54708 16116
rect 55968 13258 55996 16116
rect 57900 13462 57928 16116
rect 59832 13462 59860 16116
rect 61120 13569 61148 16116
rect 61106 13560 61162 13569
rect 61106 13495 61162 13504
rect 57888 13456 57940 13462
rect 57888 13398 57940 13404
rect 59820 13456 59872 13462
rect 59820 13398 59872 13404
rect 55956 13252 56008 13258
rect 55956 13194 56008 13200
rect 54668 13184 54720 13190
rect 54668 13126 54720 13132
rect 51448 12844 51500 12850
rect 51448 12786 51500 12792
rect 61396 3466 61424 36042
rect 61476 36032 61528 36038
rect 61476 35974 61528 35980
rect 61488 3602 61516 35974
rect 64248 35193 64276 36722
rect 64420 36712 64472 36718
rect 64420 36654 64472 36660
rect 64328 36644 64380 36650
rect 64328 36586 64380 36592
rect 64234 35184 64290 35193
rect 64234 35119 64290 35128
rect 64340 31226 64368 36586
rect 64432 31657 64460 36654
rect 64418 31648 64474 31657
rect 64418 31583 64474 31592
rect 64248 31198 64368 31226
rect 64142 30288 64198 30297
rect 64142 30223 64198 30232
rect 63500 27124 63552 27130
rect 63500 27066 63552 27072
rect 63512 27033 63540 27066
rect 63498 27024 63554 27033
rect 63498 26959 63554 26968
rect 63590 21448 63646 21457
rect 63590 21383 63646 21392
rect 63500 19304 63552 19310
rect 63500 19246 63552 19252
rect 63512 18193 63540 19246
rect 63498 18184 63554 18193
rect 63498 18119 63554 18128
rect 63604 16590 63632 21383
rect 63592 16584 63644 16590
rect 63592 16526 63644 16532
rect 64156 3670 64184 30223
rect 64248 28393 64276 31198
rect 64328 31068 64380 31074
rect 64328 31010 64380 31016
rect 64234 28384 64290 28393
rect 64234 28319 64290 28328
rect 64234 24984 64290 24993
rect 64234 24919 64290 24928
rect 64248 3738 64276 24919
rect 64340 16833 64368 31010
rect 64524 26234 64552 36790
rect 64616 31074 64644 38218
rect 64604 31068 64656 31074
rect 64604 31010 64656 31016
rect 64432 26206 64552 26234
rect 64432 23633 64460 26206
rect 64418 23624 64474 23633
rect 64418 23559 64474 23568
rect 64326 16824 64382 16833
rect 64326 16759 64382 16768
rect 65536 15026 65564 700334
rect 65628 27130 65656 700674
rect 65708 700664 65760 700670
rect 65708 700606 65760 700612
rect 65720 37398 65748 700606
rect 71044 700460 71096 700466
rect 71044 700402 71096 700408
rect 65800 700324 65852 700330
rect 65800 700266 65852 700272
rect 65812 38486 65840 700266
rect 68284 699712 68336 699718
rect 68284 699654 68336 699660
rect 65892 687336 65944 687342
rect 65892 687278 65944 687284
rect 65904 669118 65932 687278
rect 66258 674248 66314 674257
rect 66258 674183 66314 674192
rect 65892 669112 65944 669118
rect 65892 669054 65944 669060
rect 66272 665961 66300 674183
rect 66258 665952 66314 665961
rect 66258 665887 66314 665896
rect 66258 656024 66314 656033
rect 66258 655959 66314 655968
rect 66272 647737 66300 655959
rect 66258 647728 66314 647737
rect 66258 647663 66314 647672
rect 65892 632188 65944 632194
rect 65892 632130 65944 632136
rect 65904 613154 65932 632130
rect 66258 620256 66314 620265
rect 66258 620191 66314 620200
rect 65892 613148 65944 613154
rect 65892 613090 65944 613096
rect 66272 611969 66300 620191
rect 66258 611960 66314 611969
rect 66258 611895 66314 611904
rect 65892 605872 65944 605878
rect 65892 605814 65944 605820
rect 65904 580922 65932 605814
rect 65892 580916 65944 580922
rect 65892 580858 65944 580864
rect 65892 578332 65944 578338
rect 65892 578274 65944 578280
rect 65904 562358 65932 578274
rect 66258 574696 66314 574705
rect 66258 574631 66314 574640
rect 66272 566273 66300 574631
rect 66258 566264 66314 566273
rect 66258 566199 66314 566208
rect 65892 562352 65944 562358
rect 65892 562294 65944 562300
rect 65892 552084 65944 552090
rect 65892 552026 65944 552032
rect 65904 527066 65932 552026
rect 65892 527060 65944 527066
rect 65892 527002 65944 527008
rect 65892 524544 65944 524550
rect 65892 524486 65944 524492
rect 65904 503266 65932 524486
rect 66258 520704 66314 520713
rect 66258 520639 66314 520648
rect 66272 512281 66300 520639
rect 66258 512272 66314 512281
rect 66258 512207 66314 512216
rect 65892 503260 65944 503266
rect 65892 503202 65944 503208
rect 65892 498296 65944 498302
rect 65892 498238 65944 498244
rect 65904 473278 65932 498238
rect 65892 473272 65944 473278
rect 65892 473214 65944 473220
rect 66258 466712 66314 466721
rect 66258 466647 66314 466656
rect 66272 458289 66300 466647
rect 66258 458280 66314 458289
rect 66258 458215 66314 458224
rect 65892 444508 65944 444514
rect 65892 444450 65944 444456
rect 65904 419422 65932 444450
rect 65984 438932 66036 438938
rect 65984 438874 66036 438880
rect 65892 419416 65944 419422
rect 65892 419358 65944 419364
rect 65996 419354 66024 438874
rect 65984 419348 66036 419354
rect 65984 419290 66036 419296
rect 66258 404288 66314 404297
rect 66258 404223 66314 404232
rect 66272 396001 66300 404223
rect 66258 395992 66314 396001
rect 66258 395927 66314 395936
rect 65892 389292 65944 389298
rect 65892 389234 65944 389240
rect 65904 365634 65932 389234
rect 66258 377768 66314 377777
rect 66258 377703 66314 377712
rect 66272 369345 66300 377703
rect 66258 369336 66314 369345
rect 66258 369271 66314 369280
rect 65892 365628 65944 365634
rect 65892 365570 65944 365576
rect 65892 363044 65944 363050
rect 65892 362986 65944 362992
rect 65904 342922 65932 362986
rect 66258 350296 66314 350305
rect 66258 350231 66314 350240
rect 65892 342916 65944 342922
rect 65892 342858 65944 342864
rect 66272 342009 66300 350231
rect 66258 342000 66314 342009
rect 66258 341935 66314 341944
rect 65892 335368 65944 335374
rect 65892 335310 65944 335316
rect 65904 311778 65932 335310
rect 66258 323776 66314 323785
rect 66258 323711 66314 323720
rect 66272 315353 66300 323711
rect 66258 315344 66314 315353
rect 66258 315279 66314 315288
rect 65892 311772 65944 311778
rect 65892 311714 65944 311720
rect 65892 309256 65944 309262
rect 65892 309198 65944 309204
rect 65904 291922 65932 309198
rect 66258 296304 66314 296313
rect 66258 296239 66314 296248
rect 65892 291916 65944 291922
rect 65892 291858 65944 291864
rect 66272 288017 66300 296239
rect 66258 288008 66314 288017
rect 66258 287943 66314 287952
rect 66258 278080 66314 278089
rect 66258 278015 66314 278024
rect 66272 269793 66300 278015
rect 66258 269784 66314 269793
rect 66258 269719 66314 269728
rect 65892 255400 65944 255406
rect 65892 255342 65944 255348
rect 65904 235754 65932 255342
rect 66258 242312 66314 242321
rect 66258 242247 66314 242256
rect 65892 235748 65944 235754
rect 65892 235690 65944 235696
rect 66272 234025 66300 242247
rect 66258 234016 66314 234025
rect 66258 233951 66314 233960
rect 65892 227860 65944 227866
rect 65892 227802 65944 227808
rect 65904 202774 65932 227802
rect 65892 202768 65944 202774
rect 65892 202710 65944 202716
rect 65892 200252 65944 200258
rect 65892 200194 65944 200200
rect 65904 185638 65932 200194
rect 66258 196752 66314 196761
rect 66258 196687 66314 196696
rect 66272 188329 66300 196687
rect 66258 188320 66314 188329
rect 66258 188255 66314 188264
rect 65892 185632 65944 185638
rect 65892 185574 65944 185580
rect 66904 174072 66956 174078
rect 66904 174014 66956 174020
rect 66260 171148 66312 171154
rect 66260 171090 66312 171096
rect 66272 161809 66300 171090
rect 66258 161800 66314 161809
rect 66258 161735 66314 161744
rect 66916 148850 66944 174014
rect 66904 148844 66956 148850
rect 66904 148786 66956 148792
rect 65892 146396 65944 146402
rect 65892 146338 65944 146344
rect 65904 128654 65932 146338
rect 66258 142760 66314 142769
rect 66258 142695 66314 142704
rect 66272 134337 66300 142695
rect 66258 134328 66314 134337
rect 66258 134263 66314 134272
rect 65892 128648 65944 128654
rect 65892 128590 65944 128596
rect 65892 120148 65944 120154
rect 65892 120090 65944 120096
rect 65904 94994 65932 120090
rect 65892 94988 65944 94994
rect 65892 94930 65944 94936
rect 65892 92676 65944 92682
rect 65892 92618 65944 92624
rect 65904 72622 65932 92618
rect 66904 92540 66956 92546
rect 66904 92482 66956 92488
rect 66258 88768 66314 88777
rect 66258 88703 66314 88712
rect 66272 80345 66300 88703
rect 66258 80336 66314 80345
rect 66258 80271 66314 80280
rect 65892 72616 65944 72622
rect 65892 72558 65944 72564
rect 66916 68950 66944 92482
rect 66904 68944 66956 68950
rect 66904 68886 66956 68892
rect 65892 66360 65944 66366
rect 65892 66302 65944 66308
rect 65904 41206 65932 66302
rect 65984 60784 66036 60790
rect 65984 60726 66036 60732
rect 65996 41274 66024 60726
rect 65984 41268 66036 41274
rect 65984 41210 66036 41216
rect 65892 41200 65944 41206
rect 65892 41142 65944 41148
rect 65800 38480 65852 38486
rect 65800 38422 65852 38428
rect 65708 37392 65760 37398
rect 65708 37334 65760 37340
rect 65616 27124 65668 27130
rect 65616 27066 65668 27072
rect 65524 15020 65576 15026
rect 65524 14962 65576 14968
rect 68296 13054 68324 699654
rect 70306 673840 70362 673849
rect 70306 673775 70362 673784
rect 70320 665961 70348 673775
rect 70306 665952 70362 665961
rect 70306 665887 70362 665896
rect 70306 656024 70362 656033
rect 70306 655959 70362 655968
rect 70320 647737 70348 655959
rect 70306 647728 70362 647737
rect 70306 647663 70362 647672
rect 70306 620256 70362 620265
rect 70306 620191 70362 620200
rect 70320 611969 70348 620191
rect 70306 611960 70362 611969
rect 70306 611895 70362 611904
rect 70306 602032 70362 602041
rect 70306 601967 70362 601976
rect 70320 593745 70348 601967
rect 70306 593736 70362 593745
rect 70306 593671 70362 593680
rect 70306 574696 70362 574705
rect 70306 574631 70362 574640
rect 70320 566273 70348 574631
rect 70306 566264 70362 566273
rect 70306 566199 70362 566208
rect 70306 548040 70362 548049
rect 70306 547975 70362 547984
rect 70320 539753 70348 547975
rect 70306 539744 70362 539753
rect 70306 539679 70362 539688
rect 70306 520840 70362 520849
rect 70306 520775 70362 520784
rect 70320 512281 70348 520775
rect 70306 512272 70362 512281
rect 70306 512207 70362 512216
rect 70306 485752 70362 485761
rect 70306 485687 70362 485696
rect 70320 477329 70348 485687
rect 70306 477320 70362 477329
rect 70306 477255 70362 477264
rect 69664 470620 69716 470626
rect 69664 470562 69716 470568
rect 69676 19310 69704 470562
rect 70306 466712 70362 466721
rect 70306 466647 70362 466656
rect 70320 458289 70348 466647
rect 70306 458280 70362 458289
rect 70306 458215 70362 458224
rect 70306 431760 70362 431769
rect 70306 431695 70362 431704
rect 70320 423337 70348 431695
rect 70306 423328 70362 423337
rect 70306 423263 70362 423272
rect 70306 404288 70362 404297
rect 70306 404223 70362 404232
rect 70320 396001 70348 404223
rect 70306 395992 70362 396001
rect 70306 395927 70362 395936
rect 70306 377768 70362 377777
rect 70306 377703 70362 377712
rect 70320 369345 70348 377703
rect 70306 369336 70362 369345
rect 70306 369271 70362 369280
rect 70306 350296 70362 350305
rect 70306 350231 70362 350240
rect 70320 341873 70348 350231
rect 70306 341864 70362 341873
rect 70306 341799 70362 341808
rect 70306 323776 70362 323785
rect 70306 323711 70362 323720
rect 70320 315353 70348 323711
rect 70306 315344 70362 315353
rect 70306 315279 70362 315288
rect 70306 296304 70362 296313
rect 70306 296239 70362 296248
rect 70320 288017 70348 296239
rect 70306 288008 70362 288017
rect 70306 287943 70362 287952
rect 70306 278080 70362 278089
rect 70306 278015 70362 278024
rect 70320 269793 70348 278015
rect 70306 269784 70362 269793
rect 70306 269719 70362 269728
rect 70306 242312 70362 242321
rect 70306 242247 70362 242256
rect 70320 234025 70348 242247
rect 70306 234016 70362 234025
rect 70306 233951 70362 233960
rect 70306 224088 70362 224097
rect 70306 224023 70362 224032
rect 70320 215801 70348 224023
rect 70306 215792 70362 215801
rect 70306 215727 70362 215736
rect 70306 196752 70362 196761
rect 70306 196687 70362 196696
rect 70320 188329 70348 196687
rect 70306 188320 70362 188329
rect 70306 188255 70362 188264
rect 70308 171148 70360 171154
rect 70308 171090 70360 171096
rect 70320 161809 70348 171090
rect 70306 161800 70362 161809
rect 70306 161735 70362 161744
rect 70306 142760 70362 142769
rect 70306 142695 70362 142704
rect 70320 134337 70348 142695
rect 70306 134328 70362 134337
rect 70306 134263 70362 134272
rect 70306 116104 70362 116113
rect 70306 116039 70362 116048
rect 70320 108361 70348 116039
rect 70306 108352 70362 108361
rect 70306 108287 70362 108296
rect 70306 88768 70362 88777
rect 70306 88703 70362 88712
rect 70320 80345 70348 88703
rect 70306 80336 70362 80345
rect 70306 80271 70362 80280
rect 70306 53272 70362 53281
rect 70306 53207 70362 53216
rect 70320 45393 70348 53207
rect 70306 45384 70362 45393
rect 70306 45319 70362 45328
rect 70306 34912 70362 34921
rect 70306 34847 70362 34856
rect 70320 26897 70348 34847
rect 70306 26888 70362 26897
rect 70306 26823 70362 26832
rect 69664 19304 69716 19310
rect 69664 19246 69716 19252
rect 71056 14958 71084 700402
rect 72988 699718 73016 703520
rect 105464 700806 105492 703520
rect 105452 700800 105504 700806
rect 105452 700742 105504 700748
rect 95884 700596 95936 700602
rect 95884 700538 95936 700544
rect 72976 699712 73028 699718
rect 72976 699654 73028 699660
rect 81992 687336 82044 687342
rect 81992 687278 82044 687284
rect 92940 687336 92992 687342
rect 92940 687278 92992 687284
rect 72332 687268 72384 687274
rect 72332 687210 72384 687216
rect 72344 684978 72372 687210
rect 72036 684950 72372 684978
rect 82004 684978 82032 687278
rect 82004 684950 82340 684978
rect 92644 684542 92888 684570
rect 92756 684276 92808 684282
rect 92756 684218 92808 684224
rect 92768 664714 92796 684218
rect 92644 664686 92796 664714
rect 71792 664006 72036 664034
rect 82340 664006 82676 664034
rect 71792 662318 71820 664006
rect 82648 662318 82676 664006
rect 71780 662312 71832 662318
rect 71780 662254 71832 662260
rect 82636 662312 82688 662318
rect 82636 662254 82688 662260
rect 92860 662250 92888 684542
rect 92952 684282 92980 687278
rect 93124 687268 93176 687274
rect 93124 687210 93176 687216
rect 92940 684276 92992 684282
rect 92940 684218 92992 684224
rect 93136 667214 93164 687210
rect 95238 674248 95294 674257
rect 95238 674183 95294 674192
rect 93124 667208 93176 667214
rect 93124 667150 93176 667156
rect 95252 665174 95280 674183
rect 95240 665168 95292 665174
rect 95240 665110 95292 665116
rect 92848 662244 92900 662250
rect 92848 662186 92900 662192
rect 71872 659796 71924 659802
rect 71872 659738 71924 659744
rect 71780 655716 71832 655722
rect 71780 655658 71832 655664
rect 71792 634710 71820 655658
rect 71884 637786 71912 659738
rect 82266 657384 82322 657393
rect 82322 657342 82662 657370
rect 82266 657319 82322 657328
rect 71976 657206 72358 657234
rect 92966 657206 93072 657234
rect 71976 655722 72004 657206
rect 71964 655716 72016 655722
rect 71964 655658 72016 655664
rect 71884 637758 72358 637786
rect 82648 634710 82676 637092
rect 92952 634778 92980 637092
rect 93044 634778 93072 657206
rect 95240 656940 95292 656946
rect 95240 656882 95292 656888
rect 95252 647737 95280 656882
rect 95238 647728 95294 647737
rect 95238 647663 95294 647672
rect 92940 634772 92992 634778
rect 92940 634714 92992 634720
rect 93032 634772 93084 634778
rect 93032 634714 93084 634720
rect 71780 634704 71832 634710
rect 71780 634646 71832 634652
rect 82636 634704 82688 634710
rect 82636 634646 82688 634652
rect 81992 632188 82044 632194
rect 81992 632130 82044 632136
rect 92848 632188 92900 632194
rect 92848 632130 92900 632136
rect 72332 632120 72384 632126
rect 72332 632062 72384 632068
rect 72344 630986 72372 632062
rect 72036 630958 72372 630986
rect 82004 630986 82032 632130
rect 82004 630958 82340 630986
rect 92644 630278 92796 630306
rect 92768 614038 92796 630278
rect 92756 614032 92808 614038
rect 92756 613974 92808 613980
rect 92860 610994 92888 632130
rect 93124 632120 93176 632126
rect 93124 632062 93176 632068
rect 92940 614032 92992 614038
rect 92940 613974 92992 613980
rect 92768 610966 92888 610994
rect 92768 610722 92796 610966
rect 92644 610694 92796 610722
rect 71792 610014 72036 610042
rect 82340 610014 82676 610042
rect 71792 608530 71820 610014
rect 71780 608524 71832 608530
rect 71780 608466 71832 608472
rect 82648 608462 82676 610014
rect 82636 608456 82688 608462
rect 82636 608398 82688 608404
rect 92952 608394 92980 613974
rect 93136 613426 93164 632062
rect 95238 620256 95294 620265
rect 95238 620191 95294 620200
rect 93124 613420 93176 613426
rect 93124 613362 93176 613368
rect 95252 611318 95280 620191
rect 95240 611312 95292 611318
rect 95240 611254 95292 611260
rect 92940 608388 92992 608394
rect 92940 608330 92992 608336
rect 71872 605940 71924 605946
rect 71872 605882 71924 605888
rect 71780 599752 71832 599758
rect 71780 599694 71832 599700
rect 71792 580854 71820 599694
rect 71884 583794 71912 605882
rect 82636 605872 82688 605878
rect 82636 605814 82688 605820
rect 82648 603908 82676 605814
rect 71976 603214 72358 603242
rect 92966 603214 93072 603242
rect 71976 599758 72004 603214
rect 71964 599752 72016 599758
rect 71964 599694 72016 599700
rect 71884 583766 72358 583794
rect 82648 580922 82676 583100
rect 92952 580990 92980 583100
rect 93044 580990 93072 603214
rect 93124 585812 93176 585818
rect 93124 585754 93176 585760
rect 92940 580984 92992 580990
rect 92940 580926 92992 580932
rect 93032 580984 93084 580990
rect 93032 580926 93084 580932
rect 93136 580922 93164 585754
rect 82636 580916 82688 580922
rect 82636 580858 82688 580864
rect 93124 580916 93176 580922
rect 93124 580858 93176 580864
rect 71780 580848 71832 580854
rect 71780 580790 71832 580796
rect 81992 578332 82044 578338
rect 81992 578274 82044 578280
rect 92848 578332 92900 578338
rect 92848 578274 92900 578280
rect 72332 578264 72384 578270
rect 72332 578206 72384 578212
rect 72344 576994 72372 578206
rect 72036 576966 72372 576994
rect 82004 576994 82032 578274
rect 82004 576966 82340 576994
rect 92644 576286 92796 576314
rect 92768 556646 92796 576286
rect 92860 560294 92888 578274
rect 93124 578264 93176 578270
rect 93124 578206 93176 578212
rect 92860 560266 92980 560294
rect 87420 556640 87472 556646
rect 87420 556582 87472 556588
rect 92756 556640 92808 556646
rect 92756 556582 92808 556588
rect 71792 556022 72036 556050
rect 82340 556022 82676 556050
rect 71792 554674 71820 556022
rect 71780 554668 71832 554674
rect 71780 554610 71832 554616
rect 82648 554606 82676 556022
rect 82636 554600 82688 554606
rect 82636 554542 82688 554548
rect 87432 554538 87460 556582
rect 92952 556458 92980 560266
rect 93136 559570 93164 578206
rect 95238 566264 95294 566273
rect 95238 566199 95294 566208
rect 93124 559564 93176 559570
rect 93124 559506 93176 559512
rect 95252 557530 95280 566199
rect 95240 557524 95292 557530
rect 95240 557466 95292 557472
rect 92644 556430 92980 556458
rect 87420 554532 87472 554538
rect 87420 554474 87472 554480
rect 71780 552152 71832 552158
rect 71780 552094 71832 552100
rect 71792 533662 71820 552094
rect 82636 552084 82688 552090
rect 82636 552026 82688 552032
rect 82648 549916 82676 552026
rect 71884 549222 72358 549250
rect 92966 549222 93072 549250
rect 71780 533656 71832 533662
rect 71780 533598 71832 533604
rect 71884 530482 71912 549222
rect 72056 533656 72108 533662
rect 72056 533598 72108 533604
rect 71792 530454 71912 530482
rect 71792 528554 71820 530454
rect 72068 529666 72096 533598
rect 72068 529638 72358 529666
rect 71792 528526 71912 528554
rect 71884 526998 71912 528526
rect 82648 527066 82676 529108
rect 92952 527134 92980 529108
rect 93044 527134 93072 549222
rect 92940 527128 92992 527134
rect 92940 527070 92992 527076
rect 93032 527128 93084 527134
rect 93032 527070 93084 527076
rect 82636 527060 82688 527066
rect 82636 527002 82688 527008
rect 71872 526992 71924 526998
rect 71872 526934 71924 526940
rect 81992 524544 82044 524550
rect 81992 524486 82044 524492
rect 92848 524544 92900 524550
rect 92848 524486 92900 524492
rect 72332 524476 72384 524482
rect 72332 524418 72384 524424
rect 72344 522866 72372 524418
rect 72036 522838 72372 522866
rect 82004 522866 82032 524486
rect 82004 522838 82340 522866
rect 92644 522294 92796 522322
rect 92768 507210 92796 522294
rect 92756 507204 92808 507210
rect 92756 507146 92808 507152
rect 92860 503010 92888 524486
rect 93124 524476 93176 524482
rect 93124 524418 93176 524424
rect 92940 507204 92992 507210
rect 92940 507146 92992 507152
rect 92768 502982 92888 503010
rect 92768 502738 92796 502982
rect 92644 502710 92796 502738
rect 71792 502030 72036 502058
rect 82340 502030 82676 502058
rect 71792 500886 71820 502030
rect 71780 500880 71832 500886
rect 71780 500822 71832 500828
rect 82648 500818 82676 502030
rect 82636 500812 82688 500818
rect 82636 500754 82688 500760
rect 92952 500750 92980 507146
rect 93136 505782 93164 524418
rect 95238 520976 95294 520985
rect 95238 520911 95294 520920
rect 95252 512281 95280 520911
rect 95238 512272 95294 512281
rect 95238 512207 95294 512216
rect 93124 505776 93176 505782
rect 93124 505718 93176 505724
rect 92940 500744 92992 500750
rect 92940 500686 92992 500692
rect 82636 498296 82688 498302
rect 82636 498238 82688 498244
rect 71780 498228 71832 498234
rect 71780 498170 71832 498176
rect 71792 475726 71820 498170
rect 82648 495924 82676 498238
rect 71884 495230 72358 495258
rect 92966 495230 93072 495258
rect 71780 475720 71832 475726
rect 71780 475662 71832 475668
rect 71884 473210 71912 495230
rect 72056 475720 72108 475726
rect 72108 475668 72358 475674
rect 72056 475662 72358 475668
rect 72068 475646 72358 475662
rect 82648 473278 82676 475116
rect 92952 473346 92980 475116
rect 93044 473346 93072 495230
rect 92940 473340 92992 473346
rect 92940 473282 92992 473288
rect 93032 473340 93084 473346
rect 93032 473282 93084 473288
rect 82636 473272 82688 473278
rect 82636 473214 82688 473220
rect 71872 473204 71924 473210
rect 71872 473146 71924 473152
rect 92848 470756 92900 470762
rect 92848 470698 92900 470704
rect 72332 470688 72384 470694
rect 72332 470630 72384 470636
rect 72344 468874 72372 470630
rect 72036 468846 72372 468874
rect 81990 468480 82046 468489
rect 82046 468438 82340 468466
rect 81990 468415 82046 468424
rect 92644 468302 92796 468330
rect 92768 451994 92796 468302
rect 92756 451988 92808 451994
rect 92756 451930 92808 451936
rect 92860 448746 92888 470698
rect 93124 470688 93176 470694
rect 93124 470630 93176 470636
rect 92940 451988 92992 451994
rect 92940 451930 92992 451936
rect 92644 448718 92888 448746
rect 71792 448038 72036 448066
rect 82340 448038 82676 448066
rect 71792 445602 71820 448038
rect 82648 445670 82676 448038
rect 92952 445738 92980 451930
rect 93136 451926 93164 470630
rect 95238 466848 95294 466857
rect 95238 466783 95294 466792
rect 95252 458289 95280 466783
rect 95238 458280 95294 458289
rect 95238 458215 95294 458224
rect 93124 451920 93176 451926
rect 93124 451862 93176 451868
rect 92940 445732 92992 445738
rect 92940 445674 92992 445680
rect 82636 445664 82688 445670
rect 82636 445606 82688 445612
rect 71780 445596 71832 445602
rect 71780 445538 71832 445544
rect 82636 444508 82688 444514
rect 82636 444450 82688 444456
rect 71872 444440 71924 444446
rect 71872 444382 71924 444388
rect 71884 421682 71912 444382
rect 82648 441932 82676 444450
rect 71976 441238 72358 441266
rect 92966 441238 93072 441266
rect 71976 438938 72004 441238
rect 71964 438932 72016 438938
rect 71964 438874 72016 438880
rect 71884 421654 72358 421682
rect 82648 419422 82676 421124
rect 92952 419490 92980 421124
rect 93044 419490 93072 441238
rect 93124 439544 93176 439550
rect 93124 439486 93176 439492
rect 92940 419484 92992 419490
rect 92940 419426 92992 419432
rect 93032 419484 93084 419490
rect 93032 419426 93084 419432
rect 93136 419422 93164 439486
rect 82636 419416 82688 419422
rect 82636 419358 82688 419364
rect 93124 419416 93176 419422
rect 93124 419358 93176 419364
rect 92848 416900 92900 416906
rect 92848 416842 92900 416848
rect 72332 416832 72384 416838
rect 72332 416774 72384 416780
rect 72344 414882 72372 416774
rect 72036 414854 72372 414882
rect 81990 414488 82046 414497
rect 82046 414446 82340 414474
rect 81990 414423 82046 414432
rect 92644 414310 92796 414338
rect 92768 394874 92796 414310
rect 92756 394868 92808 394874
rect 92756 394810 92808 394816
rect 92860 394754 92888 416842
rect 93124 416832 93176 416838
rect 93124 416774 93176 416780
rect 93136 396778 93164 416774
rect 95238 404288 95294 404297
rect 95238 404223 95294 404232
rect 93124 396772 93176 396778
rect 93124 396714 93176 396720
rect 95252 395865 95280 404223
rect 95238 395856 95294 395865
rect 95238 395791 95294 395800
rect 92644 394726 92888 394754
rect 92756 394664 92808 394670
rect 92756 394606 92808 394612
rect 71792 394046 72036 394074
rect 82340 394046 82676 394074
rect 71792 391814 71820 394046
rect 82648 391882 82676 394046
rect 92768 391950 92796 394606
rect 92756 391944 92808 391950
rect 92756 391886 92808 391892
rect 82636 391876 82688 391882
rect 82636 391818 82688 391824
rect 71780 391808 71832 391814
rect 71780 391750 71832 391756
rect 82636 389292 82688 389298
rect 82636 389234 82688 389240
rect 71780 389224 71832 389230
rect 71780 389166 71832 389172
rect 71792 367742 71820 389166
rect 82648 387940 82676 389234
rect 71884 387246 72358 387274
rect 92966 387246 93072 387274
rect 71884 383654 71912 387246
rect 71884 383626 72096 383654
rect 72068 376754 72096 383626
rect 71884 376726 72096 376754
rect 71780 367736 71832 367742
rect 71780 367678 71832 367684
rect 71884 365566 71912 376726
rect 72056 367736 72108 367742
rect 72108 367684 72358 367690
rect 72056 367678 72358 367684
rect 72068 367662 72358 367678
rect 82648 365634 82676 367132
rect 92952 365702 92980 367132
rect 93044 365702 93072 387246
rect 95238 377768 95294 377777
rect 95238 377703 95294 377712
rect 95252 368490 95280 377703
rect 95240 368484 95292 368490
rect 95240 368426 95292 368432
rect 92940 365696 92992 365702
rect 92940 365638 92992 365644
rect 93032 365696 93084 365702
rect 93032 365638 93084 365644
rect 82636 365628 82688 365634
rect 82636 365570 82688 365576
rect 71872 365560 71924 365566
rect 71872 365502 71924 365508
rect 81992 363044 82044 363050
rect 81992 362986 82044 362992
rect 92848 363044 92900 363050
rect 92848 362986 92900 362992
rect 72332 362976 72384 362982
rect 72332 362918 72384 362924
rect 72344 360890 72372 362918
rect 72036 360862 72372 360890
rect 82004 360890 82032 362986
rect 82004 360862 82340 360890
rect 92644 360318 92796 360346
rect 92768 345710 92796 360318
rect 92756 345704 92808 345710
rect 92756 345646 92808 345652
rect 92860 340490 92888 362986
rect 93124 362976 93176 362982
rect 93124 362918 93176 362924
rect 92940 345704 92992 345710
rect 92940 345646 92992 345652
rect 92644 340462 92888 340490
rect 71792 340054 72036 340082
rect 82340 340054 82676 340082
rect 71792 338026 71820 340054
rect 71780 338020 71832 338026
rect 71780 337962 71832 337968
rect 82648 337958 82676 340054
rect 82636 337952 82688 337958
rect 82636 337894 82688 337900
rect 92952 337890 92980 345646
rect 93136 342922 93164 362918
rect 95238 350296 95294 350305
rect 95238 350231 95294 350240
rect 93124 342916 93176 342922
rect 93124 342858 93176 342864
rect 95252 341737 95280 350231
rect 95238 341728 95294 341737
rect 95238 341663 95294 341672
rect 92940 337884 92992 337890
rect 92940 337826 92992 337832
rect 71780 335436 71832 335442
rect 71780 335378 71832 335384
rect 71792 313478 71820 335378
rect 82636 335368 82688 335374
rect 82636 335310 82688 335316
rect 82648 333948 82676 335310
rect 71884 333254 72358 333282
rect 92966 333254 93072 333282
rect 71884 325694 71912 333254
rect 71884 325666 72096 325694
rect 72068 321554 72096 325666
rect 71976 321526 72096 321554
rect 71780 313472 71832 313478
rect 71780 313414 71832 313420
rect 71976 311894 72004 321526
rect 72056 313472 72108 313478
rect 72108 313420 72358 313426
rect 72056 313414 72358 313420
rect 72068 313398 72358 313414
rect 71976 311866 72096 311894
rect 72068 311710 72096 311866
rect 82648 311778 82676 313140
rect 92952 311846 92980 313140
rect 93044 311846 93072 333254
rect 95240 332648 95292 332654
rect 95240 332590 95292 332596
rect 95252 323785 95280 332590
rect 95238 323776 95294 323785
rect 95238 323711 95294 323720
rect 92940 311840 92992 311846
rect 92940 311782 92992 311788
rect 93032 311840 93084 311846
rect 93032 311782 93084 311788
rect 82636 311772 82688 311778
rect 82636 311714 82688 311720
rect 72056 311704 72108 311710
rect 72056 311646 72108 311652
rect 81992 309256 82044 309262
rect 81992 309198 82044 309204
rect 92940 309256 92992 309262
rect 92940 309198 92992 309204
rect 72332 309188 72384 309194
rect 72332 309130 72384 309136
rect 72344 306898 72372 309130
rect 72036 306870 72372 306898
rect 82004 306898 82032 309198
rect 82004 306870 82340 306898
rect 92644 306326 92888 306354
rect 92756 301572 92808 301578
rect 92756 301514 92808 301520
rect 92768 286770 92796 301514
rect 92644 286742 92796 286770
rect 71792 286062 72036 286090
rect 82340 286062 82676 286090
rect 71792 284238 71820 286062
rect 71780 284232 71832 284238
rect 71780 284174 71832 284180
rect 82648 284170 82676 286062
rect 82636 284164 82688 284170
rect 82636 284106 82688 284112
rect 92860 284102 92888 306326
rect 92952 301578 92980 309198
rect 93124 309188 93176 309194
rect 93124 309130 93176 309136
rect 92940 301572 92992 301578
rect 92940 301514 92992 301520
rect 93136 289134 93164 309130
rect 95238 296304 95294 296313
rect 95238 296239 95294 296248
rect 93124 289128 93176 289134
rect 93124 289070 93176 289076
rect 95252 287881 95280 296239
rect 95238 287872 95294 287881
rect 95238 287807 95294 287816
rect 92848 284096 92900 284102
rect 92848 284038 92900 284044
rect 71872 281648 71924 281654
rect 71872 281590 71924 281596
rect 71780 272604 71832 272610
rect 71780 272546 71832 272552
rect 71792 256630 71820 272546
rect 71884 259706 71912 281590
rect 82266 279304 82322 279313
rect 71976 279262 72358 279290
rect 71976 272610 72004 279262
rect 82322 279262 82662 279290
rect 92966 279262 93072 279290
rect 82266 279239 82322 279248
rect 71964 272604 72016 272610
rect 71964 272546 72016 272552
rect 71884 259678 72358 259706
rect 82648 256630 82676 259148
rect 92952 256698 92980 259148
rect 93044 256698 93072 279262
rect 95240 278792 95292 278798
rect 95240 278734 95292 278740
rect 95252 269793 95280 278734
rect 95238 269784 95294 269793
rect 95238 269719 95294 269728
rect 92940 256692 92992 256698
rect 92940 256634 92992 256640
rect 93032 256692 93084 256698
rect 93032 256634 93084 256640
rect 71780 256624 71832 256630
rect 71780 256566 71832 256572
rect 82636 256624 82688 256630
rect 82636 256566 82688 256572
rect 81992 255400 82044 255406
rect 81992 255342 82044 255348
rect 92940 255400 92992 255406
rect 92940 255342 92992 255348
rect 72332 255332 72384 255338
rect 72332 255274 72384 255280
rect 72344 252906 72372 255274
rect 72036 252878 72372 252906
rect 82004 252906 82032 255342
rect 82004 252878 82340 252906
rect 92644 252606 92888 252634
rect 92756 251796 92808 251802
rect 92756 251738 92808 251744
rect 92768 232778 92796 251738
rect 92644 232750 92796 232778
rect 71792 232070 72036 232098
rect 82340 232070 82676 232098
rect 71792 230382 71820 232070
rect 71780 230376 71832 230382
rect 71780 230318 71832 230324
rect 82648 230314 82676 232070
rect 82636 230308 82688 230314
rect 82636 230250 82688 230256
rect 92860 230246 92888 252606
rect 92952 251802 92980 255342
rect 93124 255332 93176 255338
rect 93124 255274 93176 255280
rect 92940 251796 92992 251802
rect 92940 251738 92992 251744
rect 93136 235278 93164 255274
rect 95238 242312 95294 242321
rect 95238 242247 95294 242256
rect 93124 235272 93176 235278
rect 93124 235214 93176 235220
rect 95252 233238 95280 242247
rect 95240 233232 95292 233238
rect 95240 233174 95292 233180
rect 92848 230240 92900 230246
rect 92848 230182 92900 230188
rect 82636 227860 82688 227866
rect 82636 227802 82688 227808
rect 71872 227792 71924 227798
rect 71872 227734 71924 227740
rect 71780 221060 71832 221066
rect 71780 221002 71832 221008
rect 71792 202706 71820 221002
rect 71884 205714 71912 227734
rect 82648 225964 82676 227802
rect 71976 225270 72358 225298
rect 92966 225270 93072 225298
rect 71976 221066 72004 225270
rect 71964 221060 72016 221066
rect 71964 221002 72016 221008
rect 71884 205686 72358 205714
rect 82648 202774 82676 205020
rect 92952 202842 92980 205020
rect 93044 202842 93072 225270
rect 92940 202836 92992 202842
rect 92940 202778 92992 202784
rect 93032 202836 93084 202842
rect 93032 202778 93084 202784
rect 82636 202768 82688 202774
rect 82636 202710 82688 202716
rect 71780 202700 71832 202706
rect 71780 202642 71832 202648
rect 92756 200320 92808 200326
rect 92756 200262 92808 200268
rect 81992 200252 82044 200258
rect 81992 200194 82044 200200
rect 72332 200184 72384 200190
rect 72332 200126 72384 200132
rect 72344 198914 72372 200126
rect 72036 198886 72372 198914
rect 82004 198914 82032 200194
rect 82004 198886 82340 198914
rect 92768 198354 92796 200262
rect 93124 200184 93176 200190
rect 93124 200126 93176 200132
rect 94504 200184 94556 200190
rect 94504 200126 94556 200132
rect 92756 198348 92808 198354
rect 92756 198290 92808 198296
rect 92644 198206 92888 198234
rect 92756 198144 92808 198150
rect 92756 198086 92808 198092
rect 92768 178786 92796 198086
rect 92644 178758 92796 178786
rect 71792 178078 72036 178106
rect 82340 178078 82676 178106
rect 71792 176594 71820 178078
rect 82648 176594 82676 178078
rect 71780 176588 71832 176594
rect 71780 176530 71832 176536
rect 82636 176588 82688 176594
rect 82636 176530 82688 176536
rect 92860 176526 92888 198206
rect 93136 181490 93164 200126
rect 93124 181484 93176 181490
rect 93124 181426 93176 181432
rect 94516 176594 94544 200126
rect 95238 188320 95294 188329
rect 95238 188255 95294 188264
rect 95252 179382 95280 188255
rect 95240 179376 95292 179382
rect 95240 179318 95292 179324
rect 94504 176588 94556 176594
rect 94504 176530 94556 176536
rect 92848 176520 92900 176526
rect 92848 176462 92900 176468
rect 82636 174072 82688 174078
rect 82636 174014 82688 174020
rect 71872 174004 71924 174010
rect 71872 173946 71924 173952
rect 71136 171216 71188 171222
rect 71136 171158 71188 171164
rect 71148 148918 71176 171158
rect 71884 151722 71912 173946
rect 82648 171972 82676 174014
rect 71976 171278 72358 171306
rect 92966 171278 93072 171306
rect 71976 171222 72004 171278
rect 71964 171216 72016 171222
rect 71964 171158 72016 171164
rect 71884 151694 72358 151722
rect 82648 148986 82676 151028
rect 92952 149054 92980 151028
rect 93044 149054 93072 171278
rect 95238 170096 95294 170105
rect 95238 170031 95294 170040
rect 95252 161809 95280 170031
rect 95238 161800 95294 161809
rect 95238 161735 95294 161744
rect 93124 153876 93176 153882
rect 93124 153818 93176 153824
rect 92940 149048 92992 149054
rect 92940 148990 92992 148996
rect 93032 149048 93084 149054
rect 93032 148990 93084 148996
rect 93136 148986 93164 153818
rect 82636 148980 82688 148986
rect 82636 148922 82688 148928
rect 93124 148980 93176 148986
rect 93124 148922 93176 148928
rect 71136 148912 71188 148918
rect 71136 148854 71188 148860
rect 81992 146396 82044 146402
rect 81992 146338 82044 146344
rect 92940 146396 92992 146402
rect 92940 146338 92992 146344
rect 72332 146328 72384 146334
rect 72332 146270 72384 146276
rect 72344 144922 72372 146270
rect 72036 144894 72372 144922
rect 82004 144922 82032 146338
rect 82004 144894 82340 144922
rect 92644 144486 92888 144514
rect 92756 144220 92808 144226
rect 92756 144162 92808 144168
rect 92768 124794 92796 144162
rect 92644 124766 92796 124794
rect 71792 124086 72036 124114
rect 82340 124086 82676 124114
rect 71792 122738 71820 124086
rect 82648 122738 82676 124086
rect 71780 122732 71832 122738
rect 71780 122674 71832 122680
rect 82636 122732 82688 122738
rect 82636 122674 82688 122680
rect 92860 122670 92888 144486
rect 92952 144226 92980 146338
rect 93124 146328 93176 146334
rect 93124 146270 93176 146276
rect 92940 144220 92992 144226
rect 92940 144162 92992 144168
rect 93136 127634 93164 146270
rect 95238 134328 95294 134337
rect 95238 134263 95294 134272
rect 93124 127628 93176 127634
rect 93124 127570 93176 127576
rect 95252 125594 95280 134263
rect 95240 125588 95292 125594
rect 95240 125530 95292 125536
rect 92848 122664 92900 122670
rect 92848 122606 92900 122612
rect 71780 120216 71832 120222
rect 71780 120158 71832 120164
rect 71792 97578 71820 120158
rect 82636 120148 82688 120154
rect 82636 120090 82688 120096
rect 82648 117980 82676 120090
rect 71884 117286 72358 117314
rect 92966 117286 93072 117314
rect 71884 113174 71912 117286
rect 71884 113146 72096 113174
rect 71780 97572 71832 97578
rect 71780 97514 71832 97520
rect 72068 96614 72096 113146
rect 72358 97578 72464 97594
rect 72358 97572 72476 97578
rect 72358 97566 72424 97572
rect 72424 97514 72476 97520
rect 72068 96586 72188 96614
rect 72160 95062 72188 96586
rect 82648 95130 82676 97036
rect 92952 95198 92980 97036
rect 93044 95198 93072 117286
rect 92940 95192 92992 95198
rect 92940 95134 92992 95140
rect 93032 95192 93084 95198
rect 93032 95134 93084 95140
rect 82636 95124 82688 95130
rect 82636 95066 82688 95072
rect 72148 95056 72200 95062
rect 72148 94998 72200 95004
rect 81992 92676 82044 92682
rect 81992 92618 82044 92624
rect 92756 92676 92808 92682
rect 92756 92618 92808 92624
rect 72332 92608 72384 92614
rect 72332 92550 72384 92556
rect 72344 90930 72372 92550
rect 72036 90902 72372 90930
rect 82004 90930 82032 92618
rect 92480 92540 92532 92546
rect 92480 92482 92532 92488
rect 92492 90930 92520 92482
rect 82004 90902 82340 90930
rect 92492 90902 92644 90930
rect 92768 70666 92796 92618
rect 93124 92608 93176 92614
rect 93124 92550 93176 92556
rect 93136 73846 93164 92550
rect 94504 92540 94556 92546
rect 94504 92482 94556 92488
rect 93124 73840 93176 73846
rect 93124 73782 93176 73788
rect 92644 70638 92796 70666
rect 71792 70094 72036 70122
rect 82340 70094 82676 70122
rect 71792 68882 71820 70094
rect 82648 69018 82676 70094
rect 94516 69018 94544 92482
rect 95238 88904 95294 88913
rect 95238 88839 95294 88848
rect 95252 80345 95280 88839
rect 95238 80336 95294 80345
rect 95238 80271 95294 80280
rect 82636 69012 82688 69018
rect 82636 68954 82688 68960
rect 94504 69012 94556 69018
rect 94504 68954 94556 68960
rect 71780 68876 71832 68882
rect 71780 68818 71832 68824
rect 82636 66360 82688 66366
rect 82636 66302 82688 66308
rect 71872 66292 71924 66298
rect 71872 66234 71924 66240
rect 71884 43738 71912 66234
rect 82648 63852 82676 66302
rect 71976 63294 72358 63322
rect 92966 63294 93072 63322
rect 71976 60790 72004 63294
rect 71964 60784 72016 60790
rect 71964 60726 72016 60732
rect 71884 43710 72358 43738
rect 82648 41342 82676 43044
rect 92952 41410 92980 43044
rect 93044 41410 93072 63294
rect 93124 61396 93176 61402
rect 93124 61338 93176 61344
rect 92940 41404 92992 41410
rect 92940 41346 92992 41352
rect 93032 41404 93084 41410
rect 93032 41346 93084 41352
rect 93136 41342 93164 61338
rect 82636 41336 82688 41342
rect 82636 41278 82688 41284
rect 93124 41336 93176 41342
rect 93124 41278 93176 41284
rect 92480 38752 92532 38758
rect 92480 38694 92532 38700
rect 92756 38752 92808 38758
rect 92756 38694 92808 38700
rect 81992 38684 82044 38690
rect 81992 38626 82044 38632
rect 82004 36938 82032 38626
rect 92492 36938 92520 38694
rect 82004 36910 82340 36938
rect 92492 36910 92644 36938
rect 71792 36230 72036 36258
rect 71792 35894 71820 36230
rect 71792 35866 71912 35894
rect 71044 14952 71096 14958
rect 71044 14894 71096 14900
rect 71884 13190 71912 35866
rect 92768 16674 92796 38694
rect 95240 37324 95292 37330
rect 95240 37266 95292 37272
rect 95252 26353 95280 37266
rect 95896 36854 95924 700538
rect 137848 700398 137876 703520
rect 170324 700466 170352 703520
rect 170312 700460 170364 700466
rect 170312 700402 170364 700408
rect 137836 700392 137888 700398
rect 137836 700334 137888 700340
rect 152464 700392 152516 700398
rect 152464 700334 152516 700340
rect 100024 687404 100076 687410
rect 100024 687346 100076 687352
rect 121092 687404 121144 687410
rect 121092 687346 121144 687352
rect 100036 684964 100064 687346
rect 110328 687336 110380 687342
rect 110328 687278 110380 687284
rect 110340 684964 110368 687278
rect 121000 687268 121052 687274
rect 121000 687210 121052 687216
rect 120658 684542 120948 684570
rect 120724 684276 120776 684282
rect 120724 684218 120776 684224
rect 97906 674248 97962 674257
rect 97906 674183 97962 674192
rect 97920 665174 97948 674183
rect 99748 667208 99800 667214
rect 99748 667150 99800 667156
rect 97908 665168 97960 665174
rect 97908 665110 97960 665116
rect 99760 664714 99788 667150
rect 120736 664714 120764 684218
rect 120816 684208 120868 684214
rect 120816 684150 120868 684156
rect 120828 667214 120856 684150
rect 120816 667208 120868 667214
rect 120816 667150 120868 667156
rect 99760 664686 100050 664714
rect 120658 664686 120764 664714
rect 110340 662250 110368 664020
rect 120920 662318 120948 684542
rect 121012 684282 121040 687210
rect 121000 684276 121052 684282
rect 121000 684218 121052 684224
rect 121104 684214 121132 687346
rect 138296 687268 138348 687274
rect 138296 687210 138348 687216
rect 138308 684964 138336 687210
rect 127084 684270 128018 684298
rect 148626 684270 148824 684298
rect 121092 684208 121144 684214
rect 121092 684150 121144 684156
rect 122838 674248 122894 674257
rect 122838 674183 122894 674192
rect 126886 674248 126942 674257
rect 126886 674183 126942 674192
rect 122852 665961 122880 674183
rect 126900 665961 126928 674183
rect 122838 665952 122894 665961
rect 122838 665887 122894 665896
rect 126886 665952 126942 665961
rect 126886 665887 126942 665896
rect 127084 662318 127112 684270
rect 127716 667208 127768 667214
rect 127716 667150 127768 667156
rect 127728 664714 127756 667150
rect 127728 664686 128018 664714
rect 138322 664006 138704 664034
rect 138676 662386 138704 664006
rect 148520 664006 148626 664034
rect 148520 663794 148548 664006
rect 148520 663766 148732 663794
rect 148704 662425 148732 663766
rect 148690 662416 148746 662425
rect 138664 662380 138716 662386
rect 148690 662351 148746 662360
rect 138664 662322 138716 662328
rect 120908 662312 120960 662318
rect 120908 662254 120960 662260
rect 127072 662312 127124 662318
rect 127072 662254 127124 662260
rect 148796 662250 148824 684270
rect 150438 674248 150494 674257
rect 150438 674183 150494 674192
rect 150452 665174 150480 674183
rect 150440 665168 150492 665174
rect 150440 665110 150492 665116
rect 110328 662244 110380 662250
rect 110328 662186 110380 662192
rect 148784 662244 148836 662250
rect 148784 662186 148836 662192
rect 110604 659796 110656 659802
rect 110604 659738 110656 659744
rect 99472 659728 99524 659734
rect 99472 659670 99524 659676
rect 97908 656940 97960 656946
rect 97908 656882 97960 656888
rect 97920 647737 97948 656882
rect 99380 655716 99432 655722
rect 99380 655658 99432 655664
rect 97906 647728 97962 647737
rect 97906 647663 97962 647672
rect 99392 634710 99420 655658
rect 99484 654134 99512 659670
rect 110616 657900 110644 659738
rect 138296 659728 138348 659734
rect 138296 659670 138348 659676
rect 149796 659728 149848 659734
rect 149796 659670 149848 659676
rect 138308 657914 138336 659670
rect 138308 657886 138644 657914
rect 128450 657384 128506 657393
rect 128340 657342 128450 657370
rect 128450 657319 128506 657328
rect 99944 657206 100326 657234
rect 120934 657206 121132 657234
rect 148948 657206 149744 657234
rect 99944 655722 99972 657206
rect 99932 655716 99984 655722
rect 99932 655658 99984 655664
rect 99484 654106 99880 654134
rect 99852 637786 99880 654106
rect 99852 637758 100326 637786
rect 110616 634817 110644 637092
rect 110602 634808 110658 634817
rect 120920 634778 120948 637092
rect 121104 634778 121132 657206
rect 122838 656024 122894 656033
rect 122838 655959 122894 655968
rect 126886 656024 126942 656033
rect 126886 655959 126942 655968
rect 122852 647737 122880 655959
rect 126900 647737 126928 655959
rect 122838 647728 122894 647737
rect 122838 647663 122894 647672
rect 126886 647728 126942 647737
rect 126886 647663 126942 647672
rect 128340 637078 128676 637106
rect 138644 637078 138980 637106
rect 110602 634743 110658 634752
rect 120908 634772 120960 634778
rect 120908 634714 120960 634720
rect 121092 634772 121144 634778
rect 121092 634714 121144 634720
rect 128648 634710 128676 637078
rect 99380 634704 99432 634710
rect 99380 634646 99432 634652
rect 128636 634704 128688 634710
rect 128636 634646 128688 634652
rect 138952 634642 138980 637078
rect 148612 637078 148948 637106
rect 148612 634778 148640 637078
rect 149716 634778 149744 657206
rect 148600 634772 148652 634778
rect 148600 634714 148652 634720
rect 149704 634772 149756 634778
rect 149704 634714 149756 634720
rect 149808 634710 149836 659670
rect 150440 656940 150492 656946
rect 150440 656882 150492 656888
rect 150452 647737 150480 656882
rect 150438 647728 150494 647737
rect 150438 647663 150494 647672
rect 149796 634704 149848 634710
rect 149796 634646 149848 634652
rect 138940 634636 138992 634642
rect 138940 634578 138992 634584
rect 100024 632256 100076 632262
rect 100024 632198 100076 632204
rect 121092 632256 121144 632262
rect 121092 632198 121144 632204
rect 100036 630972 100064 632198
rect 110328 632188 110380 632194
rect 110328 632130 110380 632136
rect 110340 630972 110368 632130
rect 121000 632120 121052 632126
rect 121000 632062 121052 632068
rect 120658 630550 120948 630578
rect 120724 630284 120776 630290
rect 120724 630226 120776 630232
rect 97906 620256 97962 620265
rect 97906 620191 97962 620200
rect 97920 611318 97948 620191
rect 99748 613420 99800 613426
rect 99748 613362 99800 613368
rect 97908 611312 97960 611318
rect 97908 611254 97960 611260
rect 99760 610722 99788 613362
rect 120736 610722 120764 630226
rect 120816 630216 120868 630222
rect 120816 630158 120868 630164
rect 120828 613426 120856 630158
rect 120816 613420 120868 613426
rect 120816 613362 120868 613368
rect 99760 610694 100050 610722
rect 120658 610694 120764 610722
rect 110340 608530 110368 610028
rect 110328 608524 110380 608530
rect 110328 608466 110380 608472
rect 120920 608462 120948 630550
rect 121012 630290 121040 632062
rect 121000 630284 121052 630290
rect 121000 630226 121052 630232
rect 121104 630222 121132 632198
rect 138296 632120 138348 632126
rect 138296 632062 138348 632068
rect 138308 630972 138336 632062
rect 127084 630278 128018 630306
rect 148626 630278 148824 630306
rect 121092 630216 121144 630222
rect 121092 630158 121144 630164
rect 122838 620256 122894 620265
rect 122838 620191 122894 620200
rect 126886 620256 126942 620265
rect 126886 620191 126942 620200
rect 122852 611969 122880 620191
rect 126900 611969 126928 620191
rect 122838 611960 122894 611969
rect 122838 611895 122894 611904
rect 126886 611960 126942 611969
rect 126886 611895 126942 611904
rect 127084 608462 127112 630278
rect 127716 613420 127768 613426
rect 127716 613362 127768 613368
rect 127728 610722 127756 613362
rect 127728 610694 128018 610722
rect 138308 608598 138336 610028
rect 138296 608592 138348 608598
rect 148612 608569 148640 610028
rect 138296 608534 138348 608540
rect 148598 608560 148654 608569
rect 148796 608530 148824 630278
rect 150438 620256 150494 620265
rect 150438 620191 150494 620200
rect 150452 611318 150480 620191
rect 150440 611312 150492 611318
rect 150440 611254 150492 611260
rect 148598 608495 148654 608504
rect 148784 608524 148836 608530
rect 148784 608466 148836 608472
rect 120908 608456 120960 608462
rect 120908 608398 120960 608404
rect 127072 608456 127124 608462
rect 127072 608398 127124 608404
rect 110604 605940 110656 605946
rect 110604 605882 110656 605888
rect 149888 605940 149940 605946
rect 149888 605882 149940 605888
rect 99380 605872 99432 605878
rect 99380 605814 99432 605820
rect 97906 602168 97962 602177
rect 97906 602103 97962 602112
rect 97920 593745 97948 602103
rect 97906 593736 97962 593745
rect 97906 593671 97962 593680
rect 99392 583930 99420 605814
rect 110616 603908 110644 605882
rect 138296 605872 138348 605878
rect 138296 605814 138348 605820
rect 149796 605872 149848 605878
rect 149796 605814 149848 605820
rect 138308 603922 138336 605814
rect 138308 603894 138644 603922
rect 128450 603392 128506 603401
rect 128340 603350 128450 603378
rect 128450 603327 128506 603336
rect 99484 603214 100326 603242
rect 120934 603214 121132 603242
rect 148948 603214 149744 603242
rect 99484 585818 99512 603214
rect 99472 585812 99524 585818
rect 99472 585754 99524 585760
rect 99392 583902 99880 583930
rect 99852 583794 99880 583902
rect 99852 583766 100326 583794
rect 110616 580961 110644 583100
rect 120920 580990 120948 583100
rect 121104 580990 121132 603214
rect 122838 602032 122894 602041
rect 122838 601967 122894 601976
rect 126886 602032 126942 602041
rect 126886 601967 126942 601976
rect 122852 593745 122880 601967
rect 126900 593745 126928 601967
rect 122838 593736 122894 593745
rect 122838 593671 122894 593680
rect 126886 593736 126942 593745
rect 126886 593671 126942 593680
rect 128340 583086 128676 583114
rect 138644 583086 138980 583114
rect 120908 580984 120960 580990
rect 110602 580952 110658 580961
rect 120908 580926 120960 580932
rect 121092 580984 121144 580990
rect 121092 580926 121144 580932
rect 128648 580922 128676 583086
rect 110602 580887 110658 580896
rect 128636 580916 128688 580922
rect 128636 580858 128688 580864
rect 138952 580854 138980 583086
rect 148612 583086 148948 583114
rect 148612 580990 148640 583086
rect 149716 580990 149744 603214
rect 148600 580984 148652 580990
rect 148600 580926 148652 580932
rect 149704 580984 149756 580990
rect 149704 580926 149756 580932
rect 149808 580922 149836 605814
rect 149796 580916 149848 580922
rect 149796 580858 149848 580864
rect 149900 580854 149928 605882
rect 138940 580848 138992 580854
rect 138940 580790 138992 580796
rect 149888 580848 149940 580854
rect 149888 580790 149940 580796
rect 100024 578400 100076 578406
rect 100024 578342 100076 578348
rect 121000 578400 121052 578406
rect 121000 578342 121052 578348
rect 100036 576980 100064 578342
rect 110328 578332 110380 578338
rect 110328 578274 110380 578280
rect 110340 576980 110368 578274
rect 120658 576558 120948 576586
rect 120724 576292 120776 576298
rect 120724 576234 120776 576240
rect 97906 566264 97962 566273
rect 97906 566199 97962 566208
rect 97920 557530 97948 566199
rect 99748 559564 99800 559570
rect 99748 559506 99800 559512
rect 97908 557524 97960 557530
rect 97908 557466 97960 557472
rect 99760 556730 99788 559506
rect 120736 556730 120764 576234
rect 120920 568002 120948 576558
rect 120908 567996 120960 568002
rect 120908 567938 120960 567944
rect 120908 567792 120960 567798
rect 120908 567734 120960 567740
rect 120816 565140 120868 565146
rect 120816 565082 120868 565088
rect 120828 559570 120856 565082
rect 120816 559564 120868 559570
rect 120816 559506 120868 559512
rect 99760 556702 100050 556730
rect 120658 556702 120764 556730
rect 110340 554674 110368 556036
rect 110328 554668 110380 554674
rect 110328 554610 110380 554616
rect 120920 554606 120948 567734
rect 121012 565146 121040 578342
rect 121092 578264 121144 578270
rect 121092 578206 121144 578212
rect 138020 578264 138072 578270
rect 138020 578206 138072 578212
rect 121104 576298 121132 578206
rect 138032 576994 138060 578206
rect 138032 576966 138322 576994
rect 121092 576292 121144 576298
rect 121092 576234 121144 576240
rect 127084 576286 128018 576314
rect 148626 576286 148824 576314
rect 122838 574696 122894 574705
rect 122838 574631 122894 574640
rect 126886 574696 126942 574705
rect 126886 574631 126942 574640
rect 122852 566273 122880 574631
rect 126900 566273 126928 574631
rect 122838 566264 122894 566273
rect 122838 566199 122894 566208
rect 126886 566264 126942 566273
rect 126886 566199 126942 566208
rect 121000 565140 121052 565146
rect 121000 565082 121052 565088
rect 127084 554606 127112 576286
rect 127716 559564 127768 559570
rect 127716 559506 127768 559512
rect 127728 556730 127756 559506
rect 127728 556702 128018 556730
rect 138308 554742 138336 556036
rect 138296 554736 138348 554742
rect 148612 554713 148640 556036
rect 138296 554678 138348 554684
rect 148598 554704 148654 554713
rect 148796 554674 148824 576286
rect 150438 566264 150494 566273
rect 150438 566199 150494 566208
rect 150452 557530 150480 566199
rect 150440 557524 150492 557530
rect 150440 557466 150492 557472
rect 148598 554639 148654 554648
rect 148784 554668 148836 554674
rect 148784 554610 148836 554616
rect 120908 554600 120960 554606
rect 120908 554542 120960 554548
rect 127072 554600 127124 554606
rect 127072 554542 127124 554548
rect 110604 552152 110656 552158
rect 110604 552094 110656 552100
rect 149888 552152 149940 552158
rect 149888 552094 149940 552100
rect 99380 552084 99432 552090
rect 99380 552026 99432 552032
rect 97906 548176 97962 548185
rect 97906 548111 97962 548120
rect 97920 539753 97948 548111
rect 97906 539744 97962 539753
rect 97906 539679 97962 539688
rect 99392 533662 99420 552026
rect 110616 549916 110644 552094
rect 138296 552084 138348 552090
rect 138296 552026 138348 552032
rect 149796 552084 149848 552090
rect 149796 552026 149848 552032
rect 138308 549930 138336 552026
rect 138308 549902 138644 549930
rect 128450 549400 128506 549409
rect 128340 549358 128450 549386
rect 128450 549335 128506 549344
rect 99484 549222 100326 549250
rect 120934 549222 121132 549250
rect 148948 549222 149744 549250
rect 99380 533656 99432 533662
rect 99380 533598 99432 533604
rect 99484 527066 99512 549222
rect 99932 533656 99984 533662
rect 99932 533598 99984 533604
rect 99944 529666 99972 533598
rect 99944 529638 100326 529666
rect 110616 527105 110644 529108
rect 120920 527134 120948 529108
rect 121104 527134 121132 549222
rect 122838 548040 122894 548049
rect 122838 547975 122894 547984
rect 126886 548040 126942 548049
rect 126886 547975 126942 547984
rect 122852 539753 122880 547975
rect 126900 539753 126928 547975
rect 122838 539744 122894 539753
rect 122838 539679 122894 539688
rect 126886 539744 126942 539753
rect 126886 539679 126942 539688
rect 128340 529094 128676 529122
rect 138644 529094 138980 529122
rect 120908 527128 120960 527134
rect 110602 527096 110658 527105
rect 99472 527060 99524 527066
rect 120908 527070 120960 527076
rect 121092 527128 121144 527134
rect 121092 527070 121144 527076
rect 128648 527066 128676 529094
rect 110602 527031 110658 527040
rect 128636 527060 128688 527066
rect 99472 527002 99524 527008
rect 128636 527002 128688 527008
rect 138952 526998 138980 529094
rect 148612 529094 148948 529122
rect 148612 527134 148640 529094
rect 149716 527134 149744 549222
rect 148600 527128 148652 527134
rect 148600 527070 148652 527076
rect 149704 527128 149756 527134
rect 149704 527070 149756 527076
rect 149808 527066 149836 552026
rect 149796 527060 149848 527066
rect 149796 527002 149848 527008
rect 149900 526998 149928 552094
rect 138940 526992 138992 526998
rect 138940 526934 138992 526940
rect 149888 526992 149940 526998
rect 149888 526934 149940 526940
rect 110328 524544 110380 524550
rect 110328 524486 110380 524492
rect 121000 524544 121052 524550
rect 121000 524486 121052 524492
rect 138296 524544 138348 524550
rect 138296 524486 138348 524492
rect 100024 524476 100076 524482
rect 100024 524418 100076 524424
rect 100036 522852 100064 524418
rect 110340 522852 110368 524486
rect 120658 522566 120948 522594
rect 120724 522300 120776 522306
rect 120724 522242 120776 522248
rect 97906 520704 97962 520713
rect 97906 520639 97962 520648
rect 97920 512281 97948 520639
rect 97906 512272 97962 512281
rect 97906 512207 97962 512216
rect 99748 505776 99800 505782
rect 99748 505718 99800 505724
rect 99760 502738 99788 505718
rect 120736 502738 120764 522242
rect 120816 522232 120868 522238
rect 120816 522174 120868 522180
rect 120828 505782 120856 522174
rect 120816 505776 120868 505782
rect 120816 505718 120868 505724
rect 99760 502710 100050 502738
rect 120658 502710 120764 502738
rect 110340 500886 110368 502044
rect 110328 500880 110380 500886
rect 110328 500822 110380 500828
rect 120920 500818 120948 522566
rect 121012 522306 121040 524486
rect 121092 524476 121144 524482
rect 121092 524418 121144 524424
rect 121000 522300 121052 522306
rect 121000 522242 121052 522248
rect 121104 522238 121132 524418
rect 138308 522852 138336 524486
rect 127084 522294 128018 522322
rect 148626 522294 148824 522322
rect 121092 522232 121144 522238
rect 121092 522174 121144 522180
rect 126886 520976 126942 520985
rect 126886 520911 126942 520920
rect 122838 520840 122894 520849
rect 122838 520775 122894 520784
rect 122852 512281 122880 520775
rect 126900 512281 126928 520911
rect 122838 512272 122894 512281
rect 122838 512207 122894 512216
rect 126886 512272 126942 512281
rect 126886 512207 126942 512216
rect 127084 500818 127112 522294
rect 127716 505776 127768 505782
rect 127716 505718 127768 505724
rect 127728 502738 127756 505718
rect 127728 502710 128018 502738
rect 138308 500954 138336 502044
rect 138296 500948 138348 500954
rect 138296 500890 138348 500896
rect 148612 500857 148640 502044
rect 148796 500886 148824 522294
rect 150438 520704 150494 520713
rect 150438 520639 150494 520648
rect 150452 512281 150480 520639
rect 150438 512272 150494 512281
rect 150438 512207 150494 512216
rect 148784 500880 148836 500886
rect 148598 500848 148654 500857
rect 120908 500812 120960 500818
rect 120908 500754 120960 500760
rect 127072 500812 127124 500818
rect 148784 500822 148836 500828
rect 148598 500783 148654 500792
rect 127072 500754 127124 500760
rect 99380 498296 99432 498302
rect 99380 498238 99432 498244
rect 138296 498296 138348 498302
rect 138296 498238 138348 498244
rect 149704 498296 149756 498302
rect 149704 498238 149756 498244
rect 97906 485752 97962 485761
rect 97906 485687 97962 485696
rect 97920 477193 97948 485687
rect 99392 477698 99420 498238
rect 110604 498228 110656 498234
rect 110604 498170 110656 498176
rect 110616 495924 110644 498170
rect 138308 495938 138336 498238
rect 138308 495910 138644 495938
rect 128174 495272 128230 495281
rect 99484 495230 100326 495258
rect 120934 495230 121132 495258
rect 99380 477692 99432 477698
rect 99380 477634 99432 477640
rect 97906 477184 97962 477193
rect 97906 477119 97962 477128
rect 99484 473278 99512 495230
rect 99932 477692 99984 477698
rect 99932 477634 99984 477640
rect 99944 475674 99972 477634
rect 99944 475646 100326 475674
rect 99472 473272 99524 473278
rect 110616 473249 110644 475116
rect 120920 473346 120948 475116
rect 121104 473346 121132 495230
rect 128230 495230 128340 495258
rect 148948 495230 149284 495258
rect 128174 495207 128230 495216
rect 149256 492590 149284 495230
rect 149244 492584 149296 492590
rect 149244 492526 149296 492532
rect 122838 485752 122894 485761
rect 122838 485687 122894 485696
rect 126886 485752 126942 485761
rect 126886 485687 126942 485696
rect 122852 477329 122880 485687
rect 126900 477329 126928 485687
rect 122838 477320 122894 477329
rect 122838 477255 122894 477264
rect 126886 477320 126942 477329
rect 126886 477255 126942 477264
rect 128340 475102 128676 475130
rect 138644 475102 138980 475130
rect 120908 473340 120960 473346
rect 120908 473282 120960 473288
rect 121092 473340 121144 473346
rect 121092 473282 121144 473288
rect 128648 473278 128676 475102
rect 128636 473272 128688 473278
rect 99472 473214 99524 473220
rect 110602 473240 110658 473249
rect 128636 473214 128688 473220
rect 138952 473210 138980 475102
rect 148612 475102 148948 475130
rect 148612 473346 148640 475102
rect 148600 473340 148652 473346
rect 148600 473282 148652 473288
rect 149716 473210 149744 498238
rect 149888 498228 149940 498234
rect 149888 498170 149940 498176
rect 149796 492584 149848 492590
rect 149796 492526 149848 492532
rect 149808 473346 149836 492526
rect 149796 473340 149848 473346
rect 149796 473282 149848 473288
rect 149900 473278 149928 498170
rect 149888 473272 149940 473278
rect 149888 473214 149940 473220
rect 110602 473175 110658 473184
rect 138940 473204 138992 473210
rect 138940 473146 138992 473152
rect 149704 473204 149756 473210
rect 149704 473146 149756 473152
rect 100024 470824 100076 470830
rect 100024 470766 100076 470772
rect 120816 470824 120868 470830
rect 120816 470766 120868 470772
rect 100036 468860 100064 470766
rect 110328 470756 110380 470762
rect 110328 470698 110380 470704
rect 110340 468860 110368 470698
rect 120724 470688 120776 470694
rect 120724 470630 120776 470636
rect 120736 468450 120764 470630
rect 120828 468450 120856 470766
rect 138296 470688 138348 470694
rect 138296 470630 138348 470636
rect 138308 468860 138336 470630
rect 120724 468444 120776 468450
rect 120724 468386 120776 468392
rect 120816 468444 120868 468450
rect 120816 468386 120868 468392
rect 120658 468302 120948 468330
rect 120724 468240 120776 468246
rect 120724 468182 120776 468188
rect 120816 468240 120868 468246
rect 120816 468182 120868 468188
rect 97906 466848 97962 466857
rect 97906 466783 97962 466792
rect 97920 458289 97948 466783
rect 97906 458280 97962 458289
rect 97906 458215 97962 458224
rect 99748 451920 99800 451926
rect 99748 451862 99800 451868
rect 99760 448746 99788 451862
rect 120736 448746 120764 468182
rect 120828 451926 120856 468182
rect 120816 451920 120868 451926
rect 120816 451862 120868 451868
rect 99760 448718 100050 448746
rect 120658 448718 120764 448746
rect 110340 445738 110368 448052
rect 110328 445732 110380 445738
rect 110328 445674 110380 445680
rect 120920 445670 120948 468302
rect 127084 468302 128018 468330
rect 148626 468302 148824 468330
rect 122838 466712 122894 466721
rect 122838 466647 122894 466656
rect 122852 458289 122880 466647
rect 122838 458280 122894 458289
rect 122838 458215 122894 458224
rect 120908 445664 120960 445670
rect 120908 445606 120960 445612
rect 127084 445602 127112 468302
rect 127716 451920 127768 451926
rect 127716 451862 127768 451868
rect 127728 448746 127756 451862
rect 127728 448718 128018 448746
rect 138308 445670 138336 448052
rect 138296 445664 138348 445670
rect 148612 445641 148640 448052
rect 148796 445738 148824 468302
rect 150438 466848 150494 466857
rect 150438 466783 150494 466792
rect 150452 458289 150480 466783
rect 150438 458280 150494 458289
rect 150438 458215 150494 458224
rect 148784 445732 148836 445738
rect 148784 445674 148836 445680
rect 138296 445606 138348 445612
rect 148598 445632 148654 445641
rect 127072 445596 127124 445602
rect 148598 445567 148654 445576
rect 127072 445538 127124 445544
rect 99472 444508 99524 444514
rect 99472 444450 99524 444456
rect 138296 444508 138348 444514
rect 138296 444450 138348 444456
rect 149888 444508 149940 444514
rect 149888 444450 149940 444456
rect 99484 441614 99512 444450
rect 110604 444440 110656 444446
rect 110604 444382 110656 444388
rect 110616 441932 110644 444382
rect 138308 441946 138336 444450
rect 149796 444440 149848 444446
rect 149796 444382 149848 444388
rect 138308 441918 138644 441946
rect 128450 441688 128506 441697
rect 128340 441646 128450 441674
rect 128450 441623 128506 441632
rect 99484 441586 99880 441614
rect 97906 431760 97962 431769
rect 97906 431695 97962 431704
rect 97920 423201 97948 431695
rect 97906 423192 97962 423201
rect 97906 423127 97962 423136
rect 99852 421682 99880 441586
rect 99944 441238 100326 441266
rect 120934 441238 121132 441266
rect 148948 441238 149744 441266
rect 99944 439550 99972 441238
rect 99932 439544 99984 439550
rect 99932 439486 99984 439492
rect 99852 421654 100326 421682
rect 110616 419529 110644 421124
rect 110602 419520 110658 419529
rect 120920 419490 120948 421124
rect 121104 419490 121132 441238
rect 122838 431760 122894 431769
rect 122838 431695 122894 431704
rect 126886 431760 126942 431769
rect 126886 431695 126942 431704
rect 122852 423337 122880 431695
rect 126900 423337 126928 431695
rect 122838 423328 122894 423337
rect 122838 423263 122894 423272
rect 126886 423328 126942 423337
rect 126886 423263 126942 423272
rect 128340 421110 128676 421138
rect 138644 421110 138980 421138
rect 110602 419455 110658 419464
rect 120908 419484 120960 419490
rect 120908 419426 120960 419432
rect 121092 419484 121144 419490
rect 121092 419426 121144 419432
rect 128648 419422 128676 421110
rect 128636 419416 128688 419422
rect 128636 419358 128688 419364
rect 138952 419354 138980 421110
rect 148612 421110 148948 421138
rect 148612 419490 148640 421110
rect 149716 419490 149744 441238
rect 148600 419484 148652 419490
rect 148600 419426 148652 419432
rect 149704 419484 149756 419490
rect 149704 419426 149756 419432
rect 149808 419422 149836 444382
rect 149796 419416 149848 419422
rect 149796 419358 149848 419364
rect 149900 419354 149928 444450
rect 138940 419348 138992 419354
rect 138940 419290 138992 419296
rect 149888 419348 149940 419354
rect 149888 419290 149940 419296
rect 100024 416968 100076 416974
rect 100024 416910 100076 416916
rect 121092 416968 121144 416974
rect 121092 416910 121144 416916
rect 100036 414868 100064 416910
rect 110328 416900 110380 416906
rect 110328 416842 110380 416848
rect 110340 414868 110368 416842
rect 121000 416832 121052 416838
rect 121000 416774 121052 416780
rect 120658 414582 120948 414610
rect 120724 414316 120776 414322
rect 120724 414258 120776 414264
rect 97906 404288 97962 404297
rect 97906 404223 97962 404232
rect 97920 395865 97948 404223
rect 99748 396772 99800 396778
rect 99748 396714 99800 396720
rect 97906 395856 97962 395865
rect 97906 395791 97962 395800
rect 99760 394754 99788 396714
rect 120736 394754 120764 414258
rect 120816 414248 120868 414254
rect 120816 414190 120868 414196
rect 120828 396778 120856 414190
rect 120816 396772 120868 396778
rect 120816 396714 120868 396720
rect 99760 394726 100050 394754
rect 120658 394726 120764 394754
rect 110340 391814 110368 394060
rect 120920 391882 120948 414582
rect 121012 414322 121040 416774
rect 121000 414316 121052 414322
rect 121000 414258 121052 414264
rect 121104 414254 121132 416910
rect 138296 416832 138348 416838
rect 138296 416774 138348 416780
rect 138308 414868 138336 416774
rect 127084 414310 128018 414338
rect 148626 414310 148824 414338
rect 121092 414248 121144 414254
rect 121092 414190 121144 414196
rect 122838 404288 122894 404297
rect 122838 404223 122894 404232
rect 122852 396001 122880 404223
rect 122838 395992 122894 396001
rect 122838 395927 122894 395936
rect 127084 391882 127112 414310
rect 127716 396772 127768 396778
rect 127716 396714 127768 396720
rect 127728 394754 127756 396714
rect 127728 394726 128018 394754
rect 138308 391950 138336 394060
rect 138296 391944 138348 391950
rect 148612 391921 148640 394060
rect 138296 391886 138348 391892
rect 148598 391912 148654 391921
rect 120908 391876 120960 391882
rect 120908 391818 120960 391824
rect 127072 391876 127124 391882
rect 148598 391847 148654 391856
rect 127072 391818 127124 391824
rect 148796 391814 148824 414310
rect 150438 404288 150494 404297
rect 150438 404223 150494 404232
rect 150452 395865 150480 404223
rect 150438 395856 150494 395865
rect 150438 395791 150494 395800
rect 110328 391808 110380 391814
rect 110328 391750 110380 391756
rect 148784 391808 148836 391814
rect 148784 391750 148836 391756
rect 99472 389292 99524 389298
rect 99472 389234 99524 389240
rect 138296 389292 138348 389298
rect 138296 389234 138348 389240
rect 149704 389292 149756 389298
rect 149704 389234 149756 389240
rect 99380 385484 99432 385490
rect 99380 385426 99432 385432
rect 97906 377768 97962 377777
rect 97906 377703 97962 377712
rect 97920 368490 97948 377703
rect 97908 368484 97960 368490
rect 97908 368426 97960 368432
rect 99392 365634 99420 385426
rect 99484 383654 99512 389234
rect 110604 389224 110656 389230
rect 110604 389166 110656 389172
rect 110616 387940 110644 389166
rect 138308 387954 138336 389234
rect 138308 387926 138644 387954
rect 128450 387424 128506 387433
rect 128340 387382 128450 387410
rect 128450 387359 128506 387368
rect 99944 387246 100326 387274
rect 120934 387246 121132 387274
rect 148948 387246 149284 387274
rect 99944 385490 99972 387246
rect 99932 385484 99984 385490
rect 99932 385426 99984 385432
rect 99484 383626 99880 383654
rect 99852 367690 99880 383626
rect 99852 367662 100326 367690
rect 110616 365673 110644 367132
rect 120920 365702 120948 367132
rect 121104 365702 121132 387246
rect 149256 385490 149284 387246
rect 149244 385484 149296 385490
rect 149244 385426 149296 385432
rect 122838 377768 122894 377777
rect 122838 377703 122894 377712
rect 126886 377768 126942 377777
rect 126886 377703 126942 377712
rect 122852 369345 122880 377703
rect 126900 369345 126928 377703
rect 122838 369336 122894 369345
rect 122838 369271 122894 369280
rect 126886 369336 126942 369345
rect 126886 369271 126942 369280
rect 128340 367118 128676 367146
rect 138644 367118 138980 367146
rect 120908 365696 120960 365702
rect 110602 365664 110658 365673
rect 99380 365628 99432 365634
rect 120908 365638 120960 365644
rect 121092 365696 121144 365702
rect 121092 365638 121144 365644
rect 128648 365634 128676 367118
rect 110602 365599 110658 365608
rect 128636 365628 128688 365634
rect 99380 365570 99432 365576
rect 128636 365570 128688 365576
rect 138952 365566 138980 367118
rect 148612 367118 148948 367146
rect 148612 365702 148640 367118
rect 148600 365696 148652 365702
rect 148600 365638 148652 365644
rect 149716 365566 149744 389234
rect 149796 389224 149848 389230
rect 149796 389166 149848 389172
rect 149808 365634 149836 389166
rect 149888 385484 149940 385490
rect 149888 385426 149940 385432
rect 149900 365702 149928 385426
rect 150438 377768 150494 377777
rect 150438 377703 150494 377712
rect 150452 368490 150480 377703
rect 150440 368484 150492 368490
rect 150440 368426 150492 368432
rect 149888 365696 149940 365702
rect 149888 365638 149940 365644
rect 149796 365628 149848 365634
rect 149796 365570 149848 365576
rect 138940 365560 138992 365566
rect 138940 365502 138992 365508
rect 149704 365560 149756 365566
rect 149704 365502 149756 365508
rect 100024 363112 100076 363118
rect 100024 363054 100076 363060
rect 121092 363112 121144 363118
rect 121092 363054 121144 363060
rect 100036 360876 100064 363054
rect 110328 363044 110380 363050
rect 110328 362986 110380 362992
rect 110340 360876 110368 362986
rect 121000 362976 121052 362982
rect 121000 362918 121052 362924
rect 120658 360590 120948 360618
rect 120724 360256 120776 360262
rect 120724 360198 120776 360204
rect 97906 350296 97962 350305
rect 97906 350231 97962 350240
rect 97920 342009 97948 350231
rect 99748 342916 99800 342922
rect 99748 342858 99800 342864
rect 97906 342000 97962 342009
rect 97906 341935 97962 341944
rect 99760 340762 99788 342858
rect 120736 340762 120764 360198
rect 120816 360188 120868 360194
rect 120816 360130 120868 360136
rect 120828 342922 120856 360130
rect 120816 342916 120868 342922
rect 120816 342858 120868 342864
rect 99760 340734 100050 340762
rect 120658 340734 120764 340762
rect 110340 338026 110368 340068
rect 110328 338020 110380 338026
rect 110328 337962 110380 337968
rect 120920 337958 120948 360590
rect 121012 360262 121040 362918
rect 121000 360256 121052 360262
rect 121000 360198 121052 360204
rect 121104 360194 121132 363054
rect 138296 362976 138348 362982
rect 138296 362918 138348 362924
rect 138308 360876 138336 362918
rect 127084 360318 128018 360346
rect 148626 360318 148824 360346
rect 121092 360188 121144 360194
rect 121092 360130 121144 360136
rect 122838 350296 122894 350305
rect 122838 350231 122894 350240
rect 122852 341873 122880 350231
rect 122838 341864 122894 341873
rect 122838 341799 122894 341808
rect 127084 337958 127112 360318
rect 127716 342916 127768 342922
rect 127716 342858 127768 342864
rect 127728 340762 127756 342858
rect 127728 340734 128018 340762
rect 138308 338094 138336 340068
rect 138296 338088 138348 338094
rect 148612 338065 148640 340068
rect 138296 338030 138348 338036
rect 148598 338056 148654 338065
rect 148796 338026 148824 360318
rect 150438 350296 150494 350305
rect 150438 350231 150494 350240
rect 150452 342009 150480 350231
rect 150438 342000 150494 342009
rect 150438 341935 150494 341944
rect 148598 337991 148654 338000
rect 148784 338020 148836 338026
rect 148784 337962 148836 337968
rect 120908 337952 120960 337958
rect 120908 337894 120960 337900
rect 127072 337952 127124 337958
rect 127072 337894 127124 337900
rect 110604 335436 110656 335442
rect 110604 335378 110656 335384
rect 149704 335436 149756 335442
rect 149704 335378 149756 335384
rect 99380 335368 99432 335374
rect 99380 335310 99432 335316
rect 97908 332648 97960 332654
rect 97908 332590 97960 332596
rect 97920 323785 97948 332590
rect 97906 323776 97962 323785
rect 97906 323711 97962 323720
rect 99392 314634 99420 335310
rect 110616 333948 110644 335378
rect 138296 335368 138348 335374
rect 138296 335310 138348 335316
rect 138308 333962 138336 335310
rect 138308 333934 138644 333962
rect 128450 333296 128506 333305
rect 99484 333254 100326 333282
rect 120934 333254 121132 333282
rect 128340 333254 128450 333282
rect 99380 314628 99432 314634
rect 99380 314570 99432 314576
rect 99484 311778 99512 333254
rect 99932 314628 99984 314634
rect 99932 314570 99984 314576
rect 99944 313698 99972 314570
rect 99944 313670 100326 313698
rect 110616 311817 110644 313140
rect 120920 311846 120948 313140
rect 121104 311846 121132 333254
rect 148948 333254 149284 333282
rect 128450 333231 128506 333240
rect 149256 329526 149284 333254
rect 149244 329520 149296 329526
rect 149244 329462 149296 329468
rect 122838 323776 122894 323785
rect 122838 323711 122894 323720
rect 126886 323776 126942 323785
rect 126886 323711 126942 323720
rect 122852 315353 122880 323711
rect 126900 315353 126928 323711
rect 122838 315344 122894 315353
rect 122838 315279 122894 315288
rect 126886 315344 126942 315353
rect 126886 315279 126942 315288
rect 128340 313126 128676 313154
rect 138644 313126 138980 313154
rect 120908 311840 120960 311846
rect 110602 311808 110658 311817
rect 99472 311772 99524 311778
rect 120908 311782 120960 311788
rect 121092 311840 121144 311846
rect 121092 311782 121144 311788
rect 128648 311778 128676 313126
rect 110602 311743 110658 311752
rect 128636 311772 128688 311778
rect 99472 311714 99524 311720
rect 128636 311714 128688 311720
rect 138952 311710 138980 313126
rect 148612 313126 148948 313154
rect 148612 311846 148640 313126
rect 148600 311840 148652 311846
rect 148600 311782 148652 311788
rect 149716 311710 149744 335378
rect 149888 335368 149940 335374
rect 149888 335310 149940 335316
rect 149796 329520 149848 329526
rect 149796 329462 149848 329468
rect 149808 311846 149836 329462
rect 149796 311840 149848 311846
rect 149796 311782 149848 311788
rect 149900 311778 149928 335310
rect 150440 332648 150492 332654
rect 150440 332590 150492 332596
rect 150452 323785 150480 332590
rect 150438 323776 150494 323785
rect 150438 323711 150494 323720
rect 149888 311772 149940 311778
rect 149888 311714 149940 311720
rect 138940 311704 138992 311710
rect 138940 311646 138992 311652
rect 149704 311704 149756 311710
rect 149704 311646 149756 311652
rect 100024 309324 100076 309330
rect 100024 309266 100076 309272
rect 121000 309324 121052 309330
rect 121000 309266 121052 309272
rect 100036 306884 100064 309266
rect 110328 309256 110380 309262
rect 110328 309198 110380 309204
rect 110340 306884 110368 309198
rect 120658 306598 120948 306626
rect 120724 306332 120776 306338
rect 120724 306274 120776 306280
rect 97906 296304 97962 296313
rect 97906 296239 97962 296248
rect 97920 287881 97948 296239
rect 99748 289128 99800 289134
rect 99748 289070 99800 289076
rect 97906 287872 97962 287881
rect 97906 287807 97962 287816
rect 99760 286770 99788 289070
rect 120736 286770 120764 306274
rect 120816 306264 120868 306270
rect 120816 306206 120868 306212
rect 120828 289134 120856 306206
rect 120816 289128 120868 289134
rect 120816 289070 120868 289076
rect 99760 286742 100050 286770
rect 120658 286742 120764 286770
rect 110340 284238 110368 286076
rect 110328 284232 110380 284238
rect 110328 284174 110380 284180
rect 120920 284170 120948 306598
rect 121012 306270 121040 309266
rect 121092 309188 121144 309194
rect 121092 309130 121144 309136
rect 138296 309188 138348 309194
rect 138296 309130 138348 309136
rect 121104 306338 121132 309130
rect 138308 306884 138336 309130
rect 121092 306332 121144 306338
rect 121092 306274 121144 306280
rect 127084 306326 128018 306354
rect 148626 306326 148824 306354
rect 121000 306264 121052 306270
rect 121000 306206 121052 306212
rect 122838 296304 122894 296313
rect 122838 296239 122894 296248
rect 126886 296304 126942 296313
rect 126886 296239 126942 296248
rect 122852 288017 122880 296239
rect 126900 288017 126928 296239
rect 122838 288008 122894 288017
rect 122838 287943 122894 287952
rect 126886 288008 126942 288017
rect 126886 287943 126942 287952
rect 127084 284170 127112 306326
rect 127716 289128 127768 289134
rect 127716 289070 127768 289076
rect 127728 286770 127756 289070
rect 127728 286742 128018 286770
rect 138308 284306 138336 286076
rect 138296 284300 138348 284306
rect 138296 284242 138348 284248
rect 148612 284209 148640 286076
rect 148796 284238 148824 306326
rect 150438 296304 150494 296313
rect 150438 296239 150494 296248
rect 150452 287881 150480 296239
rect 150438 287872 150494 287881
rect 150438 287807 150494 287816
rect 148784 284232 148836 284238
rect 148598 284200 148654 284209
rect 120908 284164 120960 284170
rect 120908 284106 120960 284112
rect 127072 284164 127124 284170
rect 148784 284174 148836 284180
rect 148598 284135 148654 284144
rect 127072 284106 127124 284112
rect 110604 281648 110656 281654
rect 110604 281590 110656 281596
rect 99472 281580 99524 281586
rect 99472 281522 99524 281528
rect 97908 278792 97960 278798
rect 97908 278734 97960 278740
rect 97920 269793 97948 278734
rect 99380 272604 99432 272610
rect 99380 272546 99432 272552
rect 97906 269784 97962 269793
rect 97906 269719 97962 269728
rect 99392 256630 99420 272546
rect 99484 267734 99512 281522
rect 110616 279956 110644 281590
rect 138296 281580 138348 281586
rect 138296 281522 138348 281528
rect 149704 281580 149756 281586
rect 149704 281522 149756 281528
rect 138308 279970 138336 281522
rect 138308 279942 138644 279970
rect 128450 279304 128506 279313
rect 99944 279262 100326 279290
rect 120934 279262 121132 279290
rect 128340 279262 128450 279290
rect 99944 272610 99972 279262
rect 99932 272604 99984 272610
rect 99932 272546 99984 272552
rect 99484 267706 99880 267734
rect 99852 259706 99880 267706
rect 99852 259678 100326 259706
rect 99380 256624 99432 256630
rect 110616 256601 110644 259148
rect 120920 256698 120948 259148
rect 121104 256698 121132 279262
rect 148948 279262 149284 279290
rect 128450 279239 128506 279248
rect 149256 278390 149284 279262
rect 149244 278384 149296 278390
rect 149244 278326 149296 278332
rect 122838 278080 122894 278089
rect 122838 278015 122894 278024
rect 126886 278080 126942 278089
rect 126886 278015 126942 278024
rect 122852 269793 122880 278015
rect 126900 269793 126928 278015
rect 122838 269784 122894 269793
rect 122838 269719 122894 269728
rect 126886 269784 126942 269793
rect 126886 269719 126942 269728
rect 128340 259134 128676 259162
rect 138644 259134 138980 259162
rect 120908 256692 120960 256698
rect 120908 256634 120960 256640
rect 121092 256692 121144 256698
rect 121092 256634 121144 256640
rect 128648 256630 128676 259134
rect 128636 256624 128688 256630
rect 99380 256566 99432 256572
rect 110602 256592 110658 256601
rect 128636 256566 128688 256572
rect 138952 256562 138980 259134
rect 148612 259134 148948 259162
rect 148612 256698 148640 259134
rect 148600 256692 148652 256698
rect 148600 256634 148652 256640
rect 149716 256630 149744 281522
rect 150440 278792 150492 278798
rect 150440 278734 150492 278740
rect 149796 278384 149848 278390
rect 149796 278326 149848 278332
rect 149808 256698 149836 278326
rect 150452 269793 150480 278734
rect 150438 269784 150494 269793
rect 150438 269719 150494 269728
rect 149796 256692 149848 256698
rect 149796 256634 149848 256640
rect 149704 256624 149756 256630
rect 149704 256566 149756 256572
rect 110602 256527 110658 256536
rect 138940 256556 138992 256562
rect 138940 256498 138992 256504
rect 100024 255468 100076 255474
rect 100024 255410 100076 255416
rect 121092 255468 121144 255474
rect 121092 255410 121144 255416
rect 100036 252892 100064 255410
rect 110328 255400 110380 255406
rect 110328 255342 110380 255348
rect 110340 252892 110368 255342
rect 121000 255332 121052 255338
rect 121000 255274 121052 255280
rect 120658 252606 120948 252634
rect 120724 252272 120776 252278
rect 120724 252214 120776 252220
rect 97906 242312 97962 242321
rect 97906 242247 97962 242256
rect 97920 233238 97948 242247
rect 99748 235272 99800 235278
rect 99748 235214 99800 235220
rect 97908 233232 97960 233238
rect 97908 233174 97960 233180
rect 99760 232778 99788 235214
rect 120736 232778 120764 252214
rect 120816 252204 120868 252210
rect 120816 252146 120868 252152
rect 120828 235278 120856 252146
rect 120816 235272 120868 235278
rect 120816 235214 120868 235220
rect 99760 232750 100050 232778
rect 120658 232750 120764 232778
rect 110340 230382 110368 232084
rect 110328 230376 110380 230382
rect 110328 230318 110380 230324
rect 120920 230314 120948 252606
rect 121012 252278 121040 255274
rect 121000 252272 121052 252278
rect 121000 252214 121052 252220
rect 121104 252210 121132 255410
rect 138296 255332 138348 255338
rect 138296 255274 138348 255280
rect 138308 252892 138336 255274
rect 127084 252334 128018 252362
rect 148626 252334 148824 252362
rect 121092 252204 121144 252210
rect 121092 252146 121144 252152
rect 122838 242312 122894 242321
rect 122838 242247 122894 242256
rect 126886 242312 126942 242321
rect 126886 242247 126942 242256
rect 122852 234025 122880 242247
rect 126900 234025 126928 242247
rect 122838 234016 122894 234025
rect 122838 233951 122894 233960
rect 126886 234016 126942 234025
rect 126886 233951 126942 233960
rect 127084 230314 127112 252334
rect 127716 235272 127768 235278
rect 127716 235214 127768 235220
rect 127728 232778 127756 235214
rect 127728 232750 128018 232778
rect 138308 230450 138336 232084
rect 148612 230489 148640 232084
rect 148598 230480 148654 230489
rect 138296 230444 138348 230450
rect 148598 230415 148654 230424
rect 138296 230386 138348 230392
rect 148796 230382 148824 252334
rect 150438 242312 150494 242321
rect 150438 242247 150494 242256
rect 150452 233238 150480 242247
rect 150440 233232 150492 233238
rect 150440 233174 150492 233180
rect 148784 230376 148836 230382
rect 148784 230318 148836 230324
rect 120908 230308 120960 230314
rect 120908 230250 120960 230256
rect 127072 230308 127124 230314
rect 127072 230250 127124 230256
rect 149704 227928 149756 227934
rect 149704 227870 149756 227876
rect 99840 227860 99892 227866
rect 99840 227802 99892 227808
rect 138296 227860 138348 227866
rect 138296 227802 138348 227808
rect 97906 224224 97962 224233
rect 97906 224159 97962 224168
rect 97920 215801 97948 224159
rect 99380 222352 99432 222358
rect 99380 222294 99432 222300
rect 97906 215792 97962 215801
rect 97906 215727 97962 215736
rect 99392 202774 99420 222294
rect 99852 205714 99880 227802
rect 110604 227792 110656 227798
rect 110604 227734 110656 227740
rect 110616 225964 110644 227734
rect 138308 225978 138336 227802
rect 138308 225950 138644 225978
rect 128450 225312 128506 225321
rect 99944 225270 100326 225298
rect 120934 225270 121132 225298
rect 128340 225270 128450 225298
rect 99944 222358 99972 225270
rect 99932 222352 99984 222358
rect 99932 222294 99984 222300
rect 99852 205686 100326 205714
rect 110616 202881 110644 205020
rect 110602 202872 110658 202881
rect 120920 202842 120948 205020
rect 121104 202842 121132 225270
rect 148948 225270 149284 225298
rect 128450 225247 128506 225256
rect 122838 224088 122894 224097
rect 122838 224023 122894 224032
rect 126886 224088 126942 224097
rect 126886 224023 126942 224032
rect 122852 215801 122880 224023
rect 126900 215801 126928 224023
rect 149256 220114 149284 225270
rect 149244 220108 149296 220114
rect 149244 220050 149296 220056
rect 122838 215792 122894 215801
rect 122838 215727 122894 215736
rect 126886 215792 126942 215801
rect 126886 215727 126942 215736
rect 128340 205006 128676 205034
rect 138644 205006 138980 205034
rect 110602 202807 110658 202816
rect 120908 202836 120960 202842
rect 120908 202778 120960 202784
rect 121092 202836 121144 202842
rect 121092 202778 121144 202784
rect 128648 202774 128676 205006
rect 99380 202768 99432 202774
rect 99380 202710 99432 202716
rect 128636 202768 128688 202774
rect 128636 202710 128688 202716
rect 138952 202706 138980 205006
rect 148612 205006 148948 205034
rect 148612 202842 148640 205006
rect 148600 202836 148652 202842
rect 148600 202778 148652 202784
rect 149716 202774 149744 227870
rect 149888 227860 149940 227866
rect 149888 227802 149940 227808
rect 149796 220108 149848 220114
rect 149796 220050 149848 220056
rect 149808 202842 149836 220050
rect 149796 202836 149848 202842
rect 149796 202778 149848 202784
rect 149704 202768 149756 202774
rect 149704 202710 149756 202716
rect 149900 202706 149928 227802
rect 138940 202700 138992 202706
rect 138940 202642 138992 202648
rect 149888 202700 149940 202706
rect 149888 202642 149940 202648
rect 110328 200320 110380 200326
rect 110328 200262 110380 200268
rect 120724 200320 120776 200326
rect 120724 200262 120776 200268
rect 138296 200320 138348 200326
rect 138296 200262 138348 200268
rect 149704 200320 149756 200326
rect 149704 200262 149756 200268
rect 100024 200252 100076 200258
rect 100024 200194 100076 200200
rect 100036 198900 100064 200194
rect 110340 198900 110368 200262
rect 120632 200184 120684 200190
rect 120632 200126 120684 200132
rect 120644 198900 120672 200126
rect 97906 188320 97962 188329
rect 97906 188255 97962 188264
rect 97920 179382 97948 188255
rect 99748 181484 99800 181490
rect 99748 181426 99800 181432
rect 97908 179376 97960 179382
rect 97908 179318 97960 179324
rect 99760 178786 99788 181426
rect 120736 178786 120764 200262
rect 120908 200252 120960 200258
rect 120908 200194 120960 200200
rect 120816 200184 120868 200190
rect 120816 200126 120868 200132
rect 99760 178758 100050 178786
rect 120658 178758 120764 178786
rect 110340 176662 110368 178092
rect 120828 176662 120856 200126
rect 120920 181490 120948 200194
rect 138308 198900 138336 200262
rect 148600 200184 148652 200190
rect 148600 200126 148652 200132
rect 148612 198900 148640 200126
rect 127084 198206 128018 198234
rect 122838 196752 122894 196761
rect 122838 196687 122894 196696
rect 126886 196752 126942 196761
rect 126886 196687 126942 196696
rect 122852 188329 122880 196687
rect 126900 188329 126928 196687
rect 122838 188320 122894 188329
rect 122838 188255 122894 188264
rect 126886 188320 126942 188329
rect 126886 188255 126942 188264
rect 120908 181484 120960 181490
rect 120908 181426 120960 181432
rect 110328 176656 110380 176662
rect 110328 176598 110380 176604
rect 120816 176656 120868 176662
rect 120816 176598 120868 176604
rect 127084 176526 127112 198206
rect 127716 181484 127768 181490
rect 127716 181426 127768 181432
rect 127728 178786 127756 181426
rect 149716 180794 149744 200262
rect 149796 200184 149848 200190
rect 149796 200126 149848 200132
rect 149072 180766 149744 180794
rect 149072 178786 149100 180766
rect 127728 178758 128018 178786
rect 148626 178758 149100 178786
rect 138308 176594 138336 178092
rect 149808 176594 149836 200126
rect 150438 188320 150494 188329
rect 150438 188255 150494 188264
rect 150452 179382 150480 188255
rect 150440 179376 150492 179382
rect 150440 179318 150492 179324
rect 138296 176588 138348 176594
rect 138296 176530 138348 176536
rect 149796 176588 149848 176594
rect 149796 176530 149848 176536
rect 127072 176520 127124 176526
rect 127072 176462 127124 176468
rect 149704 174072 149756 174078
rect 149704 174014 149756 174020
rect 110604 174004 110656 174010
rect 110604 173946 110656 173952
rect 122104 174004 122156 174010
rect 122104 173946 122156 173952
rect 128360 174004 128412 174010
rect 128360 173946 128412 173952
rect 99380 173936 99432 173942
rect 99380 173878 99432 173884
rect 97906 170640 97962 170649
rect 97906 170575 97962 170584
rect 97920 161809 97948 170575
rect 97906 161800 97962 161809
rect 97906 161735 97962 161744
rect 99392 151814 99420 173878
rect 110616 171972 110644 173946
rect 99484 171278 100326 171306
rect 120934 171278 121132 171306
rect 99484 153882 99512 171278
rect 99472 153876 99524 153882
rect 99472 153818 99524 153824
rect 99392 151786 99880 151814
rect 99852 151722 99880 151786
rect 99852 151694 100326 151722
rect 110616 148986 110644 151028
rect 120920 149054 120948 151028
rect 121104 149054 121132 171278
rect 120908 149048 120960 149054
rect 120908 148990 120960 148996
rect 121092 149048 121144 149054
rect 121092 148990 121144 148996
rect 122116 148986 122144 173946
rect 128372 171986 128400 173946
rect 138296 173936 138348 173942
rect 138296 173878 138348 173884
rect 128340 171958 128400 171986
rect 138308 171986 138336 173878
rect 148968 172100 149020 172106
rect 148968 172042 149020 172048
rect 148980 171986 149008 172042
rect 138308 171958 138644 171986
rect 148948 171958 149008 171986
rect 122840 171148 122892 171154
rect 122840 171090 122892 171096
rect 122852 161809 122880 171090
rect 122838 161800 122894 161809
rect 122838 161735 122894 161744
rect 128340 151014 128676 151042
rect 138644 151014 138980 151042
rect 128648 148986 128676 151014
rect 110604 148980 110656 148986
rect 110604 148922 110656 148928
rect 122104 148980 122156 148986
rect 122104 148922 122156 148928
rect 128636 148980 128688 148986
rect 128636 148922 128688 148928
rect 138952 148918 138980 151014
rect 148612 151014 148948 151042
rect 148612 149054 148640 151014
rect 148600 149048 148652 149054
rect 148600 148990 148652 148996
rect 149716 148986 149744 174014
rect 149704 148980 149756 148986
rect 149704 148922 149756 148928
rect 138940 148912 138992 148918
rect 138940 148854 138992 148860
rect 110328 146396 110380 146402
rect 110328 146338 110380 146344
rect 121000 146396 121052 146402
rect 121000 146338 121052 146344
rect 138296 146396 138348 146402
rect 138296 146338 138348 146344
rect 100024 146328 100076 146334
rect 100024 146270 100076 146276
rect 100036 144908 100064 146270
rect 110340 144908 110368 146338
rect 120658 144486 120948 144514
rect 120724 144288 120776 144294
rect 120724 144230 120776 144236
rect 97906 134328 97962 134337
rect 97906 134263 97962 134272
rect 97920 125594 97948 134263
rect 99748 127628 99800 127634
rect 99748 127570 99800 127576
rect 97908 125588 97960 125594
rect 97908 125530 97960 125536
rect 99760 124794 99788 127570
rect 120736 124794 120764 144230
rect 120816 144152 120868 144158
rect 120816 144094 120868 144100
rect 120828 127634 120856 144094
rect 120816 127628 120868 127634
rect 120816 127570 120868 127576
rect 99760 124766 100050 124794
rect 120658 124766 120764 124794
rect 110340 122806 110368 124100
rect 110328 122800 110380 122806
rect 110328 122742 110380 122748
rect 120920 122738 120948 144486
rect 121012 144294 121040 146338
rect 121092 146328 121144 146334
rect 121092 146270 121144 146276
rect 122104 146328 122156 146334
rect 122104 146270 122156 146276
rect 121000 144288 121052 144294
rect 121000 144230 121052 144236
rect 121104 144158 121132 146270
rect 121092 144152 121144 144158
rect 121092 144094 121144 144100
rect 122116 122806 122144 146270
rect 138308 144908 138336 146338
rect 148600 146328 148652 146334
rect 148600 146270 148652 146276
rect 148612 144908 148640 146270
rect 127084 144214 128018 144242
rect 122838 142760 122894 142769
rect 122838 142695 122894 142704
rect 126886 142760 126942 142769
rect 126886 142695 126942 142704
rect 122852 134337 122880 142695
rect 126900 134337 126928 142695
rect 122838 134328 122894 134337
rect 122838 134263 122894 134272
rect 126886 134328 126942 134337
rect 126886 134263 126942 134272
rect 122104 122800 122156 122806
rect 122104 122742 122156 122748
rect 127084 122738 127112 144214
rect 150438 134328 150494 134337
rect 150438 134263 150494 134272
rect 127716 127628 127768 127634
rect 127716 127570 127768 127576
rect 127728 124794 127756 127570
rect 150452 125594 150480 134263
rect 150440 125588 150492 125594
rect 150440 125530 150492 125536
rect 127728 124766 128018 124794
rect 138308 122806 138336 124100
rect 138296 122800 138348 122806
rect 138296 122742 138348 122748
rect 120908 122732 120960 122738
rect 120908 122674 120960 122680
rect 127072 122732 127124 122738
rect 127072 122674 127124 122680
rect 148612 122670 148640 124100
rect 148600 122664 148652 122670
rect 148600 122606 148652 122612
rect 149704 120284 149756 120290
rect 149704 120226 149756 120232
rect 110604 120216 110656 120222
rect 110604 120158 110656 120164
rect 122104 120216 122156 120222
rect 122104 120158 122156 120164
rect 128360 120216 128412 120222
rect 128360 120158 128412 120164
rect 99380 120148 99432 120154
rect 99380 120090 99432 120096
rect 97906 116240 97962 116249
rect 97906 116175 97962 116184
rect 97920 107817 97948 116175
rect 97906 107808 97962 107817
rect 97906 107743 97962 107752
rect 99392 100298 99420 120090
rect 110616 117980 110644 120158
rect 99484 117286 100326 117314
rect 120934 117286 121132 117314
rect 99380 100292 99432 100298
rect 99380 100234 99432 100240
rect 99484 95130 99512 117286
rect 99932 100292 99984 100298
rect 99932 100234 99984 100240
rect 99944 97730 99972 100234
rect 99944 97702 100326 97730
rect 110616 95130 110644 97036
rect 120920 95198 120948 97036
rect 121104 95198 121132 117286
rect 120908 95192 120960 95198
rect 120908 95134 120960 95140
rect 121092 95192 121144 95198
rect 121092 95134 121144 95140
rect 122116 95130 122144 120158
rect 128372 117994 128400 120158
rect 138296 120148 138348 120154
rect 138296 120090 138348 120096
rect 128340 117966 128400 117994
rect 138308 117994 138336 120090
rect 138308 117966 138644 117994
rect 148948 117286 149284 117314
rect 126886 116376 126942 116385
rect 126886 116311 126942 116320
rect 122838 116104 122894 116113
rect 122838 116039 122894 116048
rect 122852 107817 122880 116039
rect 126900 107817 126928 116311
rect 149256 115258 149284 117286
rect 149244 115252 149296 115258
rect 149244 115194 149296 115200
rect 122838 107808 122894 107817
rect 122838 107743 122894 107752
rect 126886 107808 126942 107817
rect 126886 107743 126942 107752
rect 128340 97022 128676 97050
rect 138644 97022 138980 97050
rect 128648 95130 128676 97022
rect 99472 95124 99524 95130
rect 99472 95066 99524 95072
rect 110604 95124 110656 95130
rect 110604 95066 110656 95072
rect 122104 95124 122156 95130
rect 122104 95066 122156 95072
rect 128636 95124 128688 95130
rect 128636 95066 128688 95072
rect 138952 95062 138980 97022
rect 148612 97022 148948 97050
rect 148612 95198 148640 97022
rect 148600 95192 148652 95198
rect 148600 95134 148652 95140
rect 149716 95130 149744 120226
rect 149796 120216 149848 120222
rect 149796 120158 149848 120164
rect 149704 95124 149756 95130
rect 149704 95066 149756 95072
rect 149808 95062 149836 120158
rect 149888 115252 149940 115258
rect 149888 115194 149940 115200
rect 149900 95198 149928 115194
rect 149888 95192 149940 95198
rect 149888 95134 149940 95140
rect 138940 95056 138992 95062
rect 138940 94998 138992 95004
rect 149796 95056 149848 95062
rect 149796 94998 149848 95004
rect 100024 92744 100076 92750
rect 100024 92686 100076 92692
rect 120816 92744 120868 92750
rect 120816 92686 120868 92692
rect 100036 90916 100064 92686
rect 110328 92676 110380 92682
rect 110328 92618 110380 92624
rect 110340 90916 110368 92618
rect 120724 92608 120776 92614
rect 120724 92550 120776 92556
rect 120632 92540 120684 92546
rect 120632 92482 120684 92488
rect 120644 90916 120672 92482
rect 97906 88904 97962 88913
rect 97906 88839 97962 88848
rect 97920 80345 97948 88839
rect 97906 80336 97962 80345
rect 97906 80271 97962 80280
rect 99748 73840 99800 73846
rect 99748 73782 99800 73788
rect 99760 70666 99788 73782
rect 120736 70666 120764 92550
rect 120828 73846 120856 92686
rect 149796 92676 149848 92682
rect 149796 92618 149848 92624
rect 138296 92608 138348 92614
rect 138296 92550 138348 92556
rect 122104 92540 122156 92546
rect 122104 92482 122156 92488
rect 120816 73840 120868 73846
rect 120816 73782 120868 73788
rect 99760 70638 100050 70666
rect 120658 70638 120764 70666
rect 110340 69018 110368 70108
rect 122116 69018 122144 92482
rect 138308 90916 138336 92550
rect 148600 92540 148652 92546
rect 148600 92482 148652 92488
rect 149704 92540 149756 92546
rect 149704 92482 149756 92488
rect 148612 90916 148640 92482
rect 127084 90222 128018 90250
rect 122838 88768 122894 88777
rect 122838 88703 122894 88712
rect 126886 88768 126942 88777
rect 126886 88703 126942 88712
rect 122852 80345 122880 88703
rect 126900 80345 126928 88703
rect 122838 80336 122894 80345
rect 122838 80271 122894 80280
rect 126886 80336 126942 80345
rect 126886 80271 126942 80280
rect 110328 69012 110380 69018
rect 110328 68954 110380 68960
rect 122104 69012 122156 69018
rect 122104 68954 122156 68960
rect 127084 68882 127112 90222
rect 127716 73840 127768 73846
rect 127716 73782 127768 73788
rect 127728 70666 127756 73782
rect 148968 71732 149020 71738
rect 148968 71674 149020 71680
rect 148980 70666 149008 71674
rect 127728 70638 128018 70666
rect 148626 70638 149008 70666
rect 138308 68950 138336 70108
rect 149716 68950 149744 92482
rect 149808 71738 149836 92618
rect 150438 88904 150494 88913
rect 150438 88839 150494 88848
rect 150452 80345 150480 88839
rect 150438 80336 150494 80345
rect 150438 80271 150494 80280
rect 149796 71732 149848 71738
rect 149796 71674 149848 71680
rect 138296 68944 138348 68950
rect 138296 68886 138348 68892
rect 149704 68944 149756 68950
rect 149704 68886 149756 68892
rect 127072 68876 127124 68882
rect 127072 68818 127124 68824
rect 99472 66360 99524 66366
rect 99472 66302 99524 66308
rect 138296 66360 138348 66366
rect 138296 66302 138348 66308
rect 149704 66360 149756 66366
rect 149704 66302 149756 66308
rect 99484 55214 99512 66302
rect 110604 66292 110656 66298
rect 110604 66234 110656 66240
rect 122104 66292 122156 66298
rect 122104 66234 122156 66240
rect 128360 66292 128412 66298
rect 128360 66234 128412 66240
rect 110616 63852 110644 66234
rect 99944 63294 100326 63322
rect 120934 63294 121132 63322
rect 99944 61402 99972 63294
rect 99932 61396 99984 61402
rect 99932 61338 99984 61344
rect 99484 55186 99880 55214
rect 97906 53816 97962 53825
rect 97906 53751 97962 53760
rect 97920 45257 97948 53751
rect 97906 45248 97962 45257
rect 97906 45183 97962 45192
rect 99852 43738 99880 55186
rect 99852 43710 100326 43738
rect 110616 41342 110644 43044
rect 120920 41410 120948 43044
rect 121104 41410 121132 63294
rect 120908 41404 120960 41410
rect 120908 41346 120960 41352
rect 121092 41404 121144 41410
rect 121092 41346 121144 41352
rect 122116 41342 122144 66234
rect 128372 63866 128400 66234
rect 128340 63838 128400 63866
rect 138308 63866 138336 66302
rect 138308 63838 138644 63866
rect 148948 63294 149284 63322
rect 149256 59294 149284 63294
rect 149244 59288 149296 59294
rect 149244 59230 149296 59236
rect 122838 53816 122894 53825
rect 122838 53751 122894 53760
rect 126886 53816 126942 53825
rect 126886 53751 126942 53760
rect 122852 45393 122880 53751
rect 126900 45393 126928 53751
rect 122838 45384 122894 45393
rect 122838 45319 122894 45328
rect 126886 45384 126942 45393
rect 126886 45319 126942 45328
rect 128340 43030 128676 43058
rect 138644 43030 138980 43058
rect 128648 41342 128676 43030
rect 110604 41336 110656 41342
rect 110604 41278 110656 41284
rect 122104 41336 122156 41342
rect 122104 41278 122156 41284
rect 128636 41336 128688 41342
rect 128636 41278 128688 41284
rect 138952 41274 138980 43030
rect 148612 43030 148948 43058
rect 148612 41410 148640 43030
rect 148600 41404 148652 41410
rect 148600 41346 148652 41352
rect 149716 41274 149744 66302
rect 149888 66292 149940 66298
rect 149888 66234 149940 66240
rect 149796 59288 149848 59294
rect 149796 59230 149848 59236
rect 149808 41410 149836 59230
rect 149796 41404 149848 41410
rect 149796 41346 149848 41352
rect 149900 41342 149928 66234
rect 149888 41336 149940 41342
rect 149888 41278 149940 41284
rect 138940 41268 138992 41274
rect 138940 41210 138992 41216
rect 149704 41268 149756 41274
rect 149704 41210 149756 41216
rect 100024 38820 100076 38826
rect 100024 38762 100076 38768
rect 121000 38820 121052 38826
rect 121000 38762 121052 38768
rect 100036 36924 100064 38762
rect 110328 38752 110380 38758
rect 110328 38694 110380 38700
rect 110340 36924 110368 38694
rect 95884 36848 95936 36854
rect 95884 36790 95936 36796
rect 120658 36502 120948 36530
rect 120724 36304 120776 36310
rect 120724 36246 120776 36252
rect 97906 34776 97962 34785
rect 97906 34711 97962 34720
rect 97920 26353 97948 34711
rect 95238 26344 95294 26353
rect 95238 26279 95294 26288
rect 97906 26344 97962 26353
rect 97906 26279 97962 26288
rect 120736 16674 120764 36246
rect 120816 36168 120868 36174
rect 120816 36110 120868 36116
rect 120828 18630 120856 36110
rect 120816 18624 120868 18630
rect 120816 18566 120868 18572
rect 92644 16646 92796 16674
rect 120658 16646 120764 16674
rect 72036 16102 72096 16130
rect 82340 16102 82676 16130
rect 71872 13184 71924 13190
rect 71872 13126 71924 13132
rect 72068 13122 72096 16102
rect 82648 13258 82676 16102
rect 82636 13252 82688 13258
rect 82636 13194 82688 13200
rect 100036 13190 100064 16116
rect 110340 13190 110368 16116
rect 120920 13258 120948 36502
rect 121012 36174 121040 38762
rect 121092 38684 121144 38690
rect 121092 38626 121144 38632
rect 138296 38684 138348 38690
rect 138296 38626 138348 38632
rect 121104 36310 121132 38626
rect 138308 36924 138336 38626
rect 152476 38418 152504 700334
rect 202800 700330 202828 703520
rect 205088 700460 205140 700466
rect 205088 700402 205140 700408
rect 202788 700324 202840 700330
rect 202788 700266 202840 700272
rect 176936 687336 176988 687342
rect 176936 687278 176988 687284
rect 194324 687336 194376 687342
rect 194324 687278 194376 687284
rect 156328 687268 156380 687274
rect 156328 687210 156380 687216
rect 156340 684978 156368 687210
rect 156032 684950 156368 684978
rect 165986 684584 166042 684593
rect 166042 684542 166336 684570
rect 165986 684519 166042 684528
rect 176640 684270 176792 684298
rect 176764 683330 176792 684270
rect 176752 683324 176804 683330
rect 176752 683266 176804 683272
rect 176844 683120 176896 683126
rect 176844 683062 176896 683068
rect 176752 679516 176804 679522
rect 176752 679458 176804 679464
rect 154486 674248 154542 674257
rect 154486 674183 154542 674192
rect 154500 665174 154528 674183
rect 154488 665168 154540 665174
rect 154488 665110 154540 665116
rect 176764 664714 176792 679458
rect 176640 664686 176792 664714
rect 156018 663794 156046 664020
rect 166336 664006 166672 664034
rect 155972 663766 156046 663794
rect 155972 662318 156000 663766
rect 166644 662318 166672 664006
rect 176856 662386 176884 683062
rect 176948 679522 176976 687278
rect 177304 687268 177356 687274
rect 177304 687210 177356 687216
rect 184020 687268 184072 687274
rect 184020 687210 184072 687216
rect 176936 679516 176988 679522
rect 176936 679458 176988 679464
rect 177316 667214 177344 687210
rect 184032 684964 184060 687210
rect 194336 684964 194364 687278
rect 204720 687268 204772 687274
rect 204720 687210 204772 687216
rect 204732 684434 204760 687210
rect 204732 684406 204852 684434
rect 204654 684282 204760 684298
rect 204654 684276 204772 684282
rect 204654 684270 204720 684276
rect 204720 684218 204772 684224
rect 204824 683114 204852 684406
rect 204996 684276 205048 684282
rect 204996 684218 205048 684224
rect 204824 683086 204944 683114
rect 204812 681760 204864 681766
rect 204812 681702 204864 681708
rect 178038 674248 178094 674257
rect 178038 674183 178094 674192
rect 182086 674248 182142 674257
rect 182086 674183 182142 674192
rect 177304 667208 177356 667214
rect 177304 667150 177356 667156
rect 178052 665961 178080 674183
rect 182100 665961 182128 674183
rect 183652 667208 183704 667214
rect 183652 667150 183704 667156
rect 178038 665952 178094 665961
rect 178038 665887 178094 665896
rect 182086 665952 182142 665961
rect 182086 665887 182142 665896
rect 183664 664714 183692 667150
rect 204824 664714 204852 681702
rect 204916 667894 204944 683086
rect 204904 667888 204956 667894
rect 204904 667830 204956 667836
rect 183664 664686 184046 664714
rect 204654 664686 204852 664714
rect 194336 662386 194364 664020
rect 176844 662380 176896 662386
rect 176844 662322 176896 662328
rect 194324 662380 194376 662386
rect 194324 662322 194376 662328
rect 205008 662318 205036 684218
rect 155960 662312 156012 662318
rect 155960 662254 156012 662260
rect 166632 662312 166684 662318
rect 166632 662254 166684 662260
rect 204996 662312 205048 662318
rect 204996 662254 205048 662260
rect 166632 659728 166684 659734
rect 166632 659670 166684 659676
rect 183652 659728 183704 659734
rect 183652 659670 183704 659676
rect 166644 657900 166672 659670
rect 155972 657206 156354 657234
rect 176962 657206 177068 657234
rect 154488 656940 154540 656946
rect 154488 656882 154540 656888
rect 154500 647737 154528 656882
rect 154486 647728 154542 647737
rect 154486 647663 154542 647672
rect 155972 634642 156000 657206
rect 156340 634817 156368 637092
rect 156326 634808 156382 634817
rect 156326 634743 156382 634752
rect 166644 634710 166672 637092
rect 176948 634778 176976 637092
rect 177040 634778 177068 657206
rect 183560 655716 183612 655722
rect 183560 655658 183612 655664
rect 176936 634772 176988 634778
rect 176936 634714 176988 634720
rect 177028 634772 177080 634778
rect 177028 634714 177080 634720
rect 183572 634710 183600 655658
rect 183664 654134 183692 659670
rect 194782 657384 194838 657393
rect 194626 657342 194782 657370
rect 205100 657354 205128 700402
rect 233884 700324 233936 700330
rect 233884 700266 233936 700272
rect 209044 687268 209096 687274
rect 209044 687210 209096 687216
rect 222200 687268 222252 687274
rect 222200 687210 222252 687216
rect 232964 687268 233016 687274
rect 232964 687210 233016 687216
rect 209056 681766 209084 687210
rect 222212 684978 222240 687210
rect 222212 684950 222364 684978
rect 232668 684542 232912 684570
rect 211264 684270 212060 684298
rect 232780 684276 232832 684282
rect 209044 681760 209096 681766
rect 209044 681702 209096 681708
rect 207018 674248 207074 674257
rect 207018 674183 207074 674192
rect 209686 674248 209742 674257
rect 209686 674183 209742 674192
rect 207032 665174 207060 674183
rect 209700 665174 209728 674183
rect 207020 665168 207072 665174
rect 207020 665110 207072 665116
rect 209688 665168 209740 665174
rect 209688 665110 209740 665116
rect 211264 662318 211292 684270
rect 232780 684218 232832 684224
rect 211712 667888 211764 667894
rect 211712 667830 211764 667836
rect 211724 664714 211752 667830
rect 232792 664714 232820 684218
rect 211724 664686 212060 664714
rect 232668 664686 232820 664714
rect 222364 664006 222700 664034
rect 222672 662425 222700 664006
rect 222658 662416 222714 662425
rect 232884 662386 232912 684542
rect 232976 684282 233004 687210
rect 232964 684276 233016 684282
rect 232964 684218 233016 684224
rect 222658 662351 222714 662360
rect 232872 662380 232924 662386
rect 232872 662322 232924 662328
rect 211252 662312 211304 662318
rect 211252 662254 211304 662260
rect 211252 659796 211304 659802
rect 211252 659738 211304 659744
rect 194782 657319 194838 657328
rect 205088 657348 205140 657354
rect 205088 657290 205140 657296
rect 184032 657206 184322 657234
rect 204930 657206 205220 657234
rect 184032 655722 184060 657206
rect 205088 657144 205140 657150
rect 205088 657086 205140 657092
rect 184202 656024 184258 656033
rect 184202 655959 184258 655968
rect 184020 655716 184072 655722
rect 184020 655658 184072 655664
rect 183664 654106 183968 654134
rect 183940 637786 183968 654106
rect 184216 648281 184244 655959
rect 184202 648272 184258 648281
rect 184202 648207 184258 648216
rect 183940 637758 184322 637786
rect 194612 634710 194640 637092
rect 204916 634778 204944 637092
rect 204904 634772 204956 634778
rect 204904 634714 204956 634720
rect 166632 634704 166684 634710
rect 166632 634646 166684 634652
rect 183560 634704 183612 634710
rect 183560 634646 183612 634652
rect 194600 634704 194652 634710
rect 194600 634646 194652 634652
rect 155960 634636 156012 634642
rect 155960 634578 156012 634584
rect 184020 632256 184072 632262
rect 184020 632198 184072 632204
rect 204904 632256 204956 632262
rect 204904 632198 204956 632204
rect 176844 632188 176896 632194
rect 176844 632130 176896 632136
rect 156328 632120 156380 632126
rect 156328 632062 156380 632068
rect 156340 630986 156368 632062
rect 156032 630958 156368 630986
rect 165986 630456 166042 630465
rect 166042 630414 166336 630442
rect 165986 630391 166042 630400
rect 176640 630278 176792 630306
rect 154486 620256 154542 620265
rect 154486 620191 154542 620200
rect 154500 611318 154528 620191
rect 154488 611312 154540 611318
rect 154488 611254 154540 611260
rect 176764 610842 176792 630278
rect 176752 610836 176804 610842
rect 176752 610778 176804 610784
rect 176856 610450 176884 632130
rect 177304 632120 177356 632126
rect 177304 632062 177356 632068
rect 177316 613426 177344 632062
rect 184032 630972 184060 632198
rect 194324 632188 194376 632194
rect 194324 632130 194376 632136
rect 194336 630972 194364 632130
rect 204812 632120 204864 632126
rect 204812 632062 204864 632068
rect 204654 630290 204760 630306
rect 204654 630284 204772 630290
rect 204654 630278 204720 630284
rect 204720 630226 204772 630232
rect 178038 620256 178094 620265
rect 178038 620191 178094 620200
rect 182086 620256 182142 620265
rect 182086 620191 182142 620200
rect 177304 613420 177356 613426
rect 177304 613362 177356 613368
rect 178052 611969 178080 620191
rect 182100 611969 182128 620191
rect 183652 613420 183704 613426
rect 183652 613362 183704 613368
rect 178038 611960 178094 611969
rect 178038 611895 178094 611904
rect 182086 611960 182142 611969
rect 182086 611895 182142 611904
rect 176936 610836 176988 610842
rect 176936 610778 176988 610784
rect 176640 610422 176884 610450
rect 156032 610014 156092 610042
rect 166336 610014 166672 610042
rect 156064 608462 156092 610014
rect 166644 608530 166672 610014
rect 176948 608598 176976 610778
rect 183664 610722 183692 613362
rect 204824 610722 204852 632062
rect 204916 613154 204944 632198
rect 204996 630284 205048 630290
rect 204996 630226 205048 630232
rect 204904 613148 204956 613154
rect 204904 613090 204956 613096
rect 183664 610694 184046 610722
rect 204654 610694 204852 610722
rect 194336 608598 194364 610028
rect 176936 608592 176988 608598
rect 176936 608534 176988 608540
rect 194324 608592 194376 608598
rect 194324 608534 194376 608540
rect 205008 608530 205036 630226
rect 166632 608524 166684 608530
rect 166632 608466 166684 608472
rect 204996 608524 205048 608530
rect 204996 608466 205048 608472
rect 156052 608456 156104 608462
rect 156052 608398 156104 608404
rect 156328 605940 156380 605946
rect 156328 605882 156380 605888
rect 156340 603908 156368 605882
rect 166632 605872 166684 605878
rect 166632 605814 166684 605820
rect 183560 605872 183612 605878
rect 183560 605814 183612 605820
rect 166644 603908 166672 605814
rect 176962 603214 177068 603242
rect 154486 602168 154542 602177
rect 154486 602103 154542 602112
rect 154500 593745 154528 602103
rect 154486 593736 154542 593745
rect 154486 593671 154542 593680
rect 156340 580961 156368 583100
rect 156326 580952 156382 580961
rect 166644 580922 166672 583100
rect 176948 580990 176976 583100
rect 177040 580990 177068 603214
rect 182086 602032 182142 602041
rect 182086 601967 182142 601976
rect 182100 593745 182128 601967
rect 182086 593736 182142 593745
rect 182086 593671 182142 593680
rect 177120 585812 177172 585818
rect 177120 585754 177172 585760
rect 176936 580984 176988 580990
rect 176936 580926 176988 580932
rect 177028 580984 177080 580990
rect 177028 580926 177080 580932
rect 177132 580922 177160 585754
rect 183572 583930 183600 605814
rect 194782 603392 194838 603401
rect 194626 603350 194782 603378
rect 205100 603362 205128 657086
rect 205192 634778 205220 657206
rect 207020 656940 207072 656946
rect 207020 656882 207072 656888
rect 209688 656940 209740 656946
rect 209688 656882 209740 656888
rect 207032 647737 207060 656882
rect 209700 647737 209728 656882
rect 211160 655716 211212 655722
rect 211160 655658 211212 655664
rect 207018 647728 207074 647737
rect 207018 647663 207074 647672
rect 209686 647728 209742 647737
rect 209686 647663 209742 647672
rect 205180 634772 205232 634778
rect 205180 634714 205232 634720
rect 211172 634710 211200 655658
rect 211264 654134 211292 659738
rect 222292 659728 222344 659734
rect 222292 659670 222344 659676
rect 222304 657914 222332 659670
rect 222304 657886 222640 657914
rect 212000 657206 212336 657234
rect 232944 657206 233096 657234
rect 212000 655722 212028 657206
rect 211988 655716 212040 655722
rect 211988 655658 212040 655664
rect 211264 654106 211936 654134
rect 211908 637786 211936 654106
rect 211908 637758 212336 637786
rect 222640 637078 222976 637106
rect 222948 634710 222976 637078
rect 232608 637078 232944 637106
rect 232608 634778 232636 637078
rect 233068 634778 233096 657206
rect 232596 634772 232648 634778
rect 232596 634714 232648 634720
rect 233056 634772 233108 634778
rect 233056 634714 233108 634720
rect 211160 634704 211212 634710
rect 211160 634646 211212 634652
rect 222936 634704 222988 634710
rect 222936 634646 222988 634652
rect 222200 632120 222252 632126
rect 222200 632062 222252 632068
rect 232964 632120 233016 632126
rect 232964 632062 233016 632068
rect 222212 630986 222240 632062
rect 222212 630958 222364 630986
rect 232668 630550 232912 630578
rect 211264 630278 212060 630306
rect 207018 620256 207074 620265
rect 207018 620191 207074 620200
rect 209686 620256 209742 620265
rect 209686 620191 209742 620200
rect 207032 611318 207060 620191
rect 209700 611318 209728 620191
rect 207020 611312 207072 611318
rect 207020 611254 207072 611260
rect 209688 611312 209740 611318
rect 209688 611254 209740 611260
rect 211264 608530 211292 630278
rect 232780 628652 232832 628658
rect 232780 628594 232832 628600
rect 211712 613148 211764 613154
rect 211712 613090 211764 613096
rect 211724 610722 211752 613090
rect 232792 610722 232820 628594
rect 211724 610694 212060 610722
rect 232668 610694 232820 610722
rect 222364 610014 222700 610042
rect 222672 608569 222700 610014
rect 232884 608598 232912 630550
rect 232976 628658 233004 632062
rect 232964 628652 233016 628658
rect 232964 628594 233016 628600
rect 232872 608592 232924 608598
rect 222658 608560 222714 608569
rect 211252 608524 211304 608530
rect 232872 608534 232924 608540
rect 222658 608495 222714 608504
rect 211252 608466 211304 608472
rect 211252 605940 211304 605946
rect 211252 605882 211304 605888
rect 194782 603327 194838 603336
rect 205088 603356 205140 603362
rect 205088 603298 205140 603304
rect 183664 603214 184322 603242
rect 204930 603214 205220 603242
rect 183664 585818 183692 603214
rect 205088 603152 205140 603158
rect 205088 603094 205140 603100
rect 183652 585812 183704 585818
rect 183652 585754 183704 585760
rect 183572 583902 183968 583930
rect 183940 583794 183968 583902
rect 183940 583766 184322 583794
rect 194612 580922 194640 583100
rect 204916 580990 204944 583100
rect 204904 580984 204956 580990
rect 204904 580926 204956 580932
rect 156326 580887 156382 580896
rect 166632 580916 166684 580922
rect 166632 580858 166684 580864
rect 177120 580916 177172 580922
rect 177120 580858 177172 580864
rect 194600 580916 194652 580922
rect 194600 580858 194652 580864
rect 184020 578400 184072 578406
rect 184020 578342 184072 578348
rect 204904 578400 204956 578406
rect 204904 578342 204956 578348
rect 176752 578332 176804 578338
rect 176752 578274 176804 578280
rect 156328 578264 156380 578270
rect 156328 578206 156380 578212
rect 156340 576994 156368 578206
rect 156032 576966 156368 576994
rect 165986 576464 166042 576473
rect 166042 576422 166336 576450
rect 176764 576434 176792 578274
rect 177304 578264 177356 578270
rect 177304 578206 177356 578212
rect 176752 576428 176804 576434
rect 165986 576399 166042 576408
rect 176752 576370 176804 576376
rect 176640 576286 176884 576314
rect 176752 576224 176804 576230
rect 176752 576166 176804 576172
rect 154486 566264 154542 566273
rect 154486 566199 154542 566208
rect 154500 557530 154528 566199
rect 154488 557524 154540 557530
rect 154488 557466 154540 557472
rect 176764 556730 176792 576166
rect 176640 556702 176792 556730
rect 156032 556022 156092 556050
rect 166336 556022 166672 556050
rect 156064 554606 156092 556022
rect 166644 554674 166672 556022
rect 176856 554742 176884 576286
rect 177316 559570 177344 578206
rect 184032 576980 184060 578342
rect 194324 578332 194376 578338
rect 194324 578274 194376 578280
rect 194336 576980 194364 578274
rect 204812 578264 204864 578270
rect 204812 578206 204864 578212
rect 204654 576298 204760 576314
rect 204654 576292 204772 576298
rect 204654 576286 204720 576292
rect 204720 576234 204772 576240
rect 178038 574696 178094 574705
rect 178038 574631 178094 574640
rect 182086 574696 182142 574705
rect 182086 574631 182142 574640
rect 178052 566273 178080 574631
rect 182100 566273 182128 574631
rect 178038 566264 178094 566273
rect 178038 566199 178094 566208
rect 182086 566264 182142 566273
rect 182086 566199 182142 566208
rect 177304 559564 177356 559570
rect 177304 559506 177356 559512
rect 183744 559564 183796 559570
rect 183744 559506 183796 559512
rect 183756 556730 183784 559506
rect 204824 556730 204852 578206
rect 204916 558958 204944 578342
rect 204996 576292 205048 576298
rect 204996 576234 205048 576240
rect 204904 558952 204956 558958
rect 204904 558894 204956 558900
rect 183756 556702 184046 556730
rect 204654 556702 204852 556730
rect 194336 554742 194364 556036
rect 176844 554736 176896 554742
rect 176844 554678 176896 554684
rect 194324 554736 194376 554742
rect 194324 554678 194376 554684
rect 205008 554674 205036 576234
rect 166632 554668 166684 554674
rect 166632 554610 166684 554616
rect 204996 554668 205048 554674
rect 204996 554610 205048 554616
rect 156052 554600 156104 554606
rect 156052 554542 156104 554548
rect 156328 552152 156380 552158
rect 156328 552094 156380 552100
rect 156340 549916 156368 552094
rect 166632 552084 166684 552090
rect 166632 552026 166684 552032
rect 183560 552084 183612 552090
rect 183560 552026 183612 552032
rect 166644 549916 166672 552026
rect 176962 549222 177068 549250
rect 154486 548176 154542 548185
rect 154486 548111 154542 548120
rect 154500 539753 154528 548111
rect 154486 539744 154542 539753
rect 154486 539679 154542 539688
rect 156340 527105 156368 529108
rect 156326 527096 156382 527105
rect 166644 527066 166672 529108
rect 176948 527134 176976 529108
rect 177040 527134 177068 549222
rect 182086 548040 182142 548049
rect 182086 547975 182142 547984
rect 182100 539753 182128 547975
rect 182086 539744 182142 539753
rect 182086 539679 182142 539688
rect 183572 533662 183600 552026
rect 194782 549400 194838 549409
rect 194626 549358 194782 549386
rect 205100 549370 205128 603094
rect 205192 580990 205220 603214
rect 207018 602168 207074 602177
rect 207018 602103 207074 602112
rect 209686 602168 209742 602177
rect 209686 602103 209742 602112
rect 207032 593745 207060 602103
rect 209700 593745 209728 602103
rect 211160 599752 211212 599758
rect 211160 599694 211212 599700
rect 207018 593736 207074 593745
rect 207018 593671 207074 593680
rect 209686 593736 209742 593745
rect 209686 593671 209742 593680
rect 205180 580984 205232 580990
rect 205180 580926 205232 580932
rect 211172 580922 211200 599694
rect 211264 596174 211292 605882
rect 222384 605872 222436 605878
rect 222384 605814 222436 605820
rect 222396 603922 222424 605814
rect 222396 603894 222640 603922
rect 212000 603214 212336 603242
rect 232944 603214 233280 603242
rect 212000 599758 212028 603214
rect 233252 599758 233280 603214
rect 211988 599752 212040 599758
rect 211988 599694 212040 599700
rect 233240 599752 233292 599758
rect 233240 599694 233292 599700
rect 211264 596146 211936 596174
rect 211908 583794 211936 596146
rect 211908 583766 212336 583794
rect 222640 583086 222976 583114
rect 222948 580922 222976 583086
rect 232608 583086 232944 583114
rect 232608 580990 232636 583086
rect 232596 580984 232648 580990
rect 232596 580926 232648 580932
rect 211160 580916 211212 580922
rect 211160 580858 211212 580864
rect 222936 580916 222988 580922
rect 222936 580858 222988 580864
rect 222200 578264 222252 578270
rect 222200 578206 222252 578212
rect 232780 578264 232832 578270
rect 232780 578206 232832 578212
rect 222212 576994 222240 578206
rect 222212 576966 222364 576994
rect 232792 576434 232820 578206
rect 232780 576428 232832 576434
rect 232780 576370 232832 576376
rect 211264 576286 212060 576314
rect 232668 576286 232912 576314
rect 207018 566264 207074 566273
rect 207018 566199 207074 566208
rect 209686 566264 209742 566273
rect 209686 566199 209742 566208
rect 207032 557530 207060 566199
rect 209700 557530 209728 566199
rect 207020 557524 207072 557530
rect 207020 557466 207072 557472
rect 209688 557524 209740 557530
rect 209688 557466 209740 557472
rect 211264 554674 211292 576286
rect 232780 576224 232832 576230
rect 232780 576166 232832 576172
rect 211712 558952 211764 558958
rect 211712 558894 211764 558900
rect 211724 556730 211752 558894
rect 232792 556730 232820 576166
rect 211724 556702 212060 556730
rect 232668 556702 232820 556730
rect 222364 556022 222700 556050
rect 222672 554713 222700 556022
rect 232884 554742 232912 576286
rect 232872 554736 232924 554742
rect 222658 554704 222714 554713
rect 211252 554668 211304 554674
rect 232872 554678 232924 554684
rect 222658 554639 222714 554648
rect 211252 554610 211304 554616
rect 211160 552152 211212 552158
rect 211160 552094 211212 552100
rect 194782 549335 194838 549344
rect 205088 549364 205140 549370
rect 205088 549306 205140 549312
rect 183664 549222 184322 549250
rect 204930 549222 205220 549250
rect 183560 533656 183612 533662
rect 183560 533598 183612 533604
rect 176936 527128 176988 527134
rect 176936 527070 176988 527076
rect 177028 527128 177080 527134
rect 177028 527070 177080 527076
rect 183664 527066 183692 549222
rect 205088 549160 205140 549166
rect 205088 549102 205140 549108
rect 184020 533656 184072 533662
rect 184020 533598 184072 533604
rect 184032 529666 184060 533598
rect 184032 529638 184322 529666
rect 194612 527066 194640 529108
rect 204916 527134 204944 529108
rect 204904 527128 204956 527134
rect 204904 527070 204956 527076
rect 156326 527031 156382 527040
rect 166632 527060 166684 527066
rect 166632 527002 166684 527008
rect 183652 527060 183704 527066
rect 183652 527002 183704 527008
rect 194600 527060 194652 527066
rect 194600 527002 194652 527008
rect 184020 524612 184072 524618
rect 184020 524554 184072 524560
rect 204904 524612 204956 524618
rect 204904 524554 204956 524560
rect 177028 524544 177080 524550
rect 177028 524486 177080 524492
rect 156328 524476 156380 524482
rect 156328 524418 156380 524424
rect 156340 522866 156368 524418
rect 156032 522838 156368 522866
rect 165986 522472 166042 522481
rect 166042 522430 166336 522458
rect 165986 522407 166042 522416
rect 177040 522322 177068 524486
rect 177304 524476 177356 524482
rect 177304 524418 177356 524424
rect 176640 522294 176884 522322
rect 176856 522034 176884 522294
rect 176948 522294 177068 522322
rect 176844 522028 176896 522034
rect 176844 521970 176896 521976
rect 155866 520840 155922 520849
rect 155866 520775 155922 520784
rect 155880 518906 155908 520775
rect 176948 519602 176976 522294
rect 177028 522028 177080 522034
rect 177028 521970 177080 521976
rect 176764 519574 176976 519602
rect 154488 518900 154540 518906
rect 154488 518842 154540 518848
rect 155868 518900 155920 518906
rect 155868 518842 155920 518848
rect 154500 512281 154528 518842
rect 154486 512272 154542 512281
rect 154486 512207 154542 512216
rect 176764 502738 176792 519574
rect 177040 514842 177068 521970
rect 176640 502710 176792 502738
rect 176856 514814 177068 514842
rect 156032 502030 156092 502058
rect 166336 502030 166672 502058
rect 156064 500818 156092 502030
rect 166644 500886 166672 502030
rect 176856 500954 176884 514814
rect 177316 505782 177344 524418
rect 184032 522852 184060 524554
rect 194324 524544 194376 524550
rect 194324 524486 194376 524492
rect 194336 522852 194364 524486
rect 204812 524476 204864 524482
rect 204812 524418 204864 524424
rect 204654 522306 204760 522322
rect 204654 522300 204772 522306
rect 204654 522294 204720 522300
rect 204720 522242 204772 522248
rect 182086 520704 182142 520713
rect 182086 520639 182142 520648
rect 182100 512281 182128 520639
rect 182086 512272 182142 512281
rect 182086 512207 182142 512216
rect 177304 505776 177356 505782
rect 177304 505718 177356 505724
rect 183652 505776 183704 505782
rect 183652 505718 183704 505724
rect 183664 502738 183692 505718
rect 204824 502738 204852 524418
rect 204916 505986 204944 524554
rect 204996 522300 205048 522306
rect 204996 522242 205048 522248
rect 204904 505980 204956 505986
rect 204904 505922 204956 505928
rect 183664 502710 184046 502738
rect 204654 502710 204852 502738
rect 194336 500954 194364 502044
rect 176844 500948 176896 500954
rect 176844 500890 176896 500896
rect 194324 500948 194376 500954
rect 194324 500890 194376 500896
rect 205008 500886 205036 522242
rect 166632 500880 166684 500886
rect 166632 500822 166684 500828
rect 204996 500880 205048 500886
rect 204996 500822 205048 500828
rect 156052 500812 156104 500818
rect 156052 500754 156104 500760
rect 156328 498296 156380 498302
rect 156328 498238 156380 498244
rect 156340 495924 156368 498238
rect 166632 498228 166684 498234
rect 166632 498170 166684 498176
rect 183560 498228 183612 498234
rect 183560 498170 183612 498176
rect 166644 495924 166672 498170
rect 176962 495230 177068 495258
rect 154486 485752 154542 485761
rect 154486 485687 154542 485696
rect 154500 477193 154528 485687
rect 154486 477184 154542 477193
rect 154486 477119 154542 477128
rect 156340 473249 156368 475116
rect 166644 473278 166672 475116
rect 176948 473346 176976 475116
rect 177040 473346 177068 495230
rect 182086 485752 182142 485761
rect 182086 485687 182142 485696
rect 182100 477329 182128 485687
rect 183572 477698 183600 498170
rect 194782 495544 194838 495553
rect 194626 495502 194782 495530
rect 194782 495479 194838 495488
rect 205100 495378 205128 549102
rect 205192 527134 205220 549222
rect 207018 548176 207074 548185
rect 207018 548111 207074 548120
rect 207032 539753 207060 548111
rect 207018 539744 207074 539753
rect 207018 539679 207074 539688
rect 211172 533662 211200 552094
rect 222292 552084 222344 552090
rect 222292 552026 222344 552032
rect 222304 549930 222332 552026
rect 222304 549902 222640 549930
rect 232944 549358 233280 549386
rect 211264 549222 212336 549250
rect 211160 533656 211212 533662
rect 211160 533598 211212 533604
rect 205180 527128 205232 527134
rect 205180 527070 205232 527076
rect 211264 527066 211292 549222
rect 233252 548554 233280 549358
rect 233240 548548 233292 548554
rect 233240 548490 233292 548496
rect 211988 533656 212040 533662
rect 211988 533598 212040 533604
rect 212000 529666 212028 533598
rect 212000 529638 212336 529666
rect 222640 529094 222976 529122
rect 222948 527066 222976 529094
rect 232608 529094 232944 529122
rect 232608 527134 232636 529094
rect 232596 527128 232648 527134
rect 232596 527070 232648 527076
rect 211252 527060 211304 527066
rect 211252 527002 211304 527008
rect 222936 527060 222988 527066
rect 222936 527002 222988 527008
rect 222200 524476 222252 524482
rect 222200 524418 222252 524424
rect 232964 524476 233016 524482
rect 232964 524418 233016 524424
rect 222212 522866 222240 524418
rect 222212 522838 222364 522866
rect 232668 522566 232912 522594
rect 211264 522294 212060 522322
rect 207018 520840 207074 520849
rect 207018 520775 207074 520784
rect 207032 512281 207060 520775
rect 207018 512272 207074 512281
rect 207018 512207 207074 512216
rect 211264 500886 211292 522294
rect 232780 521688 232832 521694
rect 232780 521630 232832 521636
rect 211712 505980 211764 505986
rect 211712 505922 211764 505928
rect 211724 502738 211752 505922
rect 232792 502738 232820 521630
rect 211724 502710 212060 502738
rect 232668 502710 232820 502738
rect 222364 502030 222700 502058
rect 211252 500880 211304 500886
rect 222672 500857 222700 502030
rect 232884 500954 232912 522566
rect 232976 521694 233004 524418
rect 232964 521688 233016 521694
rect 232964 521630 233016 521636
rect 232872 500948 232924 500954
rect 232872 500890 232924 500896
rect 211252 500822 211304 500828
rect 222658 500848 222714 500857
rect 222658 500783 222714 500792
rect 211160 498296 211212 498302
rect 211160 498238 211212 498244
rect 205088 495372 205140 495378
rect 205088 495314 205140 495320
rect 183664 495230 184322 495258
rect 204930 495230 205220 495258
rect 183560 477692 183612 477698
rect 183560 477634 183612 477640
rect 182086 477320 182142 477329
rect 182086 477255 182142 477264
rect 176936 473340 176988 473346
rect 176936 473282 176988 473288
rect 177028 473340 177080 473346
rect 177028 473282 177080 473288
rect 183664 473278 183692 495230
rect 205088 495168 205140 495174
rect 205088 495110 205140 495116
rect 184020 477692 184072 477698
rect 184020 477634 184072 477640
rect 184032 475674 184060 477634
rect 184032 475646 184322 475674
rect 194612 473278 194640 475116
rect 204916 473346 204944 475116
rect 204904 473340 204956 473346
rect 204904 473282 204956 473288
rect 166632 473272 166684 473278
rect 156326 473240 156382 473249
rect 166632 473214 166684 473220
rect 183652 473272 183704 473278
rect 183652 473214 183704 473220
rect 194600 473272 194652 473278
rect 194600 473214 194652 473220
rect 156326 473175 156382 473184
rect 184020 470824 184072 470830
rect 184020 470766 184072 470772
rect 204904 470824 204956 470830
rect 204904 470766 204956 470772
rect 176844 470756 176896 470762
rect 176844 470698 176896 470704
rect 156328 470688 156380 470694
rect 156328 470630 156380 470636
rect 156340 468874 156368 470630
rect 156032 468846 156368 468874
rect 165986 468480 166042 468489
rect 166042 468438 166336 468466
rect 165986 468415 166042 468424
rect 176640 468302 176792 468330
rect 154486 466848 154542 466857
rect 154486 466783 154542 466792
rect 154500 458289 154528 466783
rect 154486 458280 154542 458289
rect 154486 458215 154542 458224
rect 176764 448866 176792 468302
rect 176752 448860 176804 448866
rect 176752 448802 176804 448808
rect 176856 448474 176884 470698
rect 177304 470688 177356 470694
rect 177304 470630 177356 470636
rect 177316 451926 177344 470630
rect 184032 468860 184060 470766
rect 194324 470756 194376 470762
rect 194324 470698 194376 470704
rect 194336 468860 194364 470698
rect 204812 470688 204864 470694
rect 204812 470630 204864 470636
rect 204654 468314 204760 468330
rect 204654 468308 204772 468314
rect 204654 468302 204720 468308
rect 204720 468250 204772 468256
rect 178038 466712 178094 466721
rect 178038 466647 178094 466656
rect 182086 466712 182142 466721
rect 182086 466647 182142 466656
rect 178052 458289 178080 466647
rect 182100 458289 182128 466647
rect 178038 458280 178094 458289
rect 178038 458215 178094 458224
rect 182086 458280 182142 458289
rect 182086 458215 182142 458224
rect 177304 451920 177356 451926
rect 177304 451862 177356 451868
rect 183744 451920 183796 451926
rect 183744 451862 183796 451868
rect 176936 448860 176988 448866
rect 176936 448802 176988 448808
rect 176640 448446 176884 448474
rect 156032 448038 156092 448066
rect 166336 448038 166672 448066
rect 156064 445602 156092 448038
rect 166644 445602 166672 448038
rect 176948 445670 176976 448802
rect 183756 448746 183784 451862
rect 204824 448746 204852 470630
rect 204916 451314 204944 470766
rect 204996 468308 205048 468314
rect 204996 468250 205048 468256
rect 204904 451308 204956 451314
rect 204904 451250 204956 451256
rect 183756 448718 184046 448746
rect 204654 448718 204852 448746
rect 194336 445738 194364 448052
rect 194324 445732 194376 445738
rect 194324 445674 194376 445680
rect 176936 445664 176988 445670
rect 176936 445606 176988 445612
rect 205008 445602 205036 468250
rect 156052 445596 156104 445602
rect 156052 445538 156104 445544
rect 166632 445596 166684 445602
rect 166632 445538 166684 445544
rect 204996 445596 205048 445602
rect 204996 445538 205048 445544
rect 156328 444508 156380 444514
rect 156328 444450 156380 444456
rect 156340 441932 156368 444450
rect 166632 444440 166684 444446
rect 166632 444382 166684 444388
rect 183652 444440 183704 444446
rect 183652 444382 183704 444388
rect 166644 441932 166672 444382
rect 183664 441614 183692 444382
rect 194782 441688 194838 441697
rect 194626 441646 194782 441674
rect 194782 441623 194838 441632
rect 183664 441586 183968 441614
rect 176962 441238 177068 441266
rect 154486 431760 154542 431769
rect 154486 431695 154542 431704
rect 154500 423201 154528 431695
rect 154486 423192 154542 423201
rect 154486 423127 154542 423136
rect 156340 419529 156368 421124
rect 156326 419520 156382 419529
rect 156326 419455 156382 419464
rect 166644 419422 166672 421124
rect 176948 419490 176976 421124
rect 177040 419490 177068 441238
rect 177304 439544 177356 439550
rect 177304 439486 177356 439492
rect 176936 419484 176988 419490
rect 176936 419426 176988 419432
rect 177028 419484 177080 419490
rect 177028 419426 177080 419432
rect 177316 419422 177344 439486
rect 182086 431760 182142 431769
rect 182086 431695 182142 431704
rect 182100 423337 182128 431695
rect 182086 423328 182142 423337
rect 182086 423263 182142 423272
rect 183940 421682 183968 441586
rect 205100 441386 205128 495110
rect 205192 473346 205220 495230
rect 207018 485752 207074 485761
rect 207018 485687 207074 485696
rect 207032 477193 207060 485687
rect 211172 477698 211200 498238
rect 222292 498228 222344 498234
rect 222292 498170 222344 498176
rect 222304 495938 222332 498170
rect 222304 495910 222640 495938
rect 211264 495230 212336 495258
rect 232944 495230 233280 495258
rect 211160 477692 211212 477698
rect 211160 477634 211212 477640
rect 207018 477184 207074 477193
rect 207018 477119 207074 477128
rect 205180 473340 205232 473346
rect 205180 473282 205232 473288
rect 211264 473278 211292 495230
rect 233252 492590 233280 495230
rect 233240 492584 233292 492590
rect 233240 492526 233292 492532
rect 211988 477692 212040 477698
rect 211988 477634 212040 477640
rect 212000 475674 212028 477634
rect 212000 475646 212336 475674
rect 222640 475102 222976 475130
rect 222948 473278 222976 475102
rect 232608 475102 232944 475130
rect 232608 473346 232636 475102
rect 232596 473340 232648 473346
rect 232596 473282 232648 473288
rect 211252 473272 211304 473278
rect 211252 473214 211304 473220
rect 222936 473272 222988 473278
rect 222936 473214 222988 473220
rect 222292 470688 222344 470694
rect 222292 470630 222344 470636
rect 232780 470688 232832 470694
rect 232780 470630 232832 470636
rect 222304 468874 222332 470630
rect 222304 468846 222364 468874
rect 232792 468450 232820 470630
rect 232780 468444 232832 468450
rect 232780 468386 232832 468392
rect 211264 468302 212060 468330
rect 232668 468302 232912 468330
rect 207018 466848 207074 466857
rect 207018 466783 207074 466792
rect 207032 458289 207060 466783
rect 207018 458280 207074 458289
rect 207018 458215 207074 458224
rect 211264 445670 211292 468302
rect 232780 468240 232832 468246
rect 232780 468182 232832 468188
rect 211712 451308 211764 451314
rect 211712 451250 211764 451256
rect 211724 448746 211752 451250
rect 232792 448746 232820 468182
rect 211724 448718 212060 448746
rect 232668 448718 232820 448746
rect 222364 448038 222700 448066
rect 211252 445664 211304 445670
rect 222672 445641 222700 448038
rect 232884 445738 232912 468302
rect 232872 445732 232924 445738
rect 232872 445674 232924 445680
rect 211252 445606 211304 445612
rect 222658 445632 222714 445641
rect 222658 445567 222714 445576
rect 211160 444508 211212 444514
rect 211160 444450 211212 444456
rect 205088 441380 205140 441386
rect 205088 441322 205140 441328
rect 184032 441238 184322 441266
rect 204930 441238 205220 441266
rect 184032 439550 184060 441238
rect 205088 441176 205140 441182
rect 205088 441118 205140 441124
rect 184020 439544 184072 439550
rect 184020 439486 184072 439492
rect 183940 421654 184322 421682
rect 194612 419422 194640 421124
rect 204916 419490 204944 421124
rect 204904 419484 204956 419490
rect 204904 419426 204956 419432
rect 166632 419416 166684 419422
rect 166632 419358 166684 419364
rect 177304 419416 177356 419422
rect 177304 419358 177356 419364
rect 194600 419416 194652 419422
rect 194600 419358 194652 419364
rect 176844 416900 176896 416906
rect 176844 416842 176896 416848
rect 194324 416900 194376 416906
rect 194324 416842 194376 416848
rect 204812 416900 204864 416906
rect 204812 416842 204864 416848
rect 156328 416832 156380 416838
rect 156328 416774 156380 416780
rect 156340 414882 156368 416774
rect 156032 414854 156368 414882
rect 165986 414488 166042 414497
rect 166042 414446 166336 414474
rect 165986 414423 166042 414432
rect 176640 414310 176792 414338
rect 154486 404288 154542 404297
rect 154486 404223 154542 404232
rect 154500 395865 154528 404223
rect 154486 395856 154542 395865
rect 154486 395791 154542 395800
rect 176764 394874 176792 414310
rect 176752 394868 176804 394874
rect 176752 394810 176804 394816
rect 176856 394754 176884 416842
rect 177304 416832 177356 416838
rect 177304 416774 177356 416780
rect 184020 416832 184072 416838
rect 184020 416774 184072 416780
rect 177316 396778 177344 416774
rect 184032 414868 184060 416774
rect 194336 414868 194364 416842
rect 204654 414310 204760 414338
rect 204732 414254 204760 414310
rect 204720 414248 204772 414254
rect 204720 414190 204772 414196
rect 178038 404288 178094 404297
rect 178038 404223 178094 404232
rect 182086 404288 182142 404297
rect 182086 404223 182142 404232
rect 177304 396772 177356 396778
rect 177304 396714 177356 396720
rect 178052 396001 178080 404223
rect 182100 396001 182128 404223
rect 183652 396772 183704 396778
rect 183652 396714 183704 396720
rect 178038 395992 178094 396001
rect 178038 395927 178094 395936
rect 182086 395992 182142 396001
rect 182086 395927 182142 395936
rect 176640 394726 176884 394754
rect 183664 394754 183692 396714
rect 204824 394754 204852 416842
rect 204904 416832 204956 416838
rect 204904 416774 204956 416780
rect 204916 397458 204944 416774
rect 204996 414248 205048 414254
rect 204996 414190 205048 414196
rect 204904 397452 204956 397458
rect 204904 397394 204956 397400
rect 183664 394726 184046 394754
rect 204654 394726 204852 394754
rect 176752 394664 176804 394670
rect 176752 394606 176804 394612
rect 156018 393802 156046 394060
rect 166336 394046 166672 394074
rect 155972 393774 156046 393802
rect 155972 391882 156000 393774
rect 166644 391882 166672 394046
rect 176764 391950 176792 394606
rect 194336 391950 194364 394060
rect 176752 391944 176804 391950
rect 176752 391886 176804 391892
rect 194324 391944 194376 391950
rect 194324 391886 194376 391892
rect 205008 391882 205036 414190
rect 155960 391876 156012 391882
rect 155960 391818 156012 391824
rect 166632 391876 166684 391882
rect 166632 391818 166684 391824
rect 204996 391876 205048 391882
rect 204996 391818 205048 391824
rect 156328 389292 156380 389298
rect 156328 389234 156380 389240
rect 156340 387940 156368 389234
rect 166632 389224 166684 389230
rect 166632 389166 166684 389172
rect 183560 389224 183612 389230
rect 183560 389166 183612 389172
rect 166644 387940 166672 389166
rect 176962 387246 177068 387274
rect 154486 377768 154542 377777
rect 154486 377703 154542 377712
rect 154500 368490 154528 377703
rect 154488 368484 154540 368490
rect 154488 368426 154540 368432
rect 156340 365673 156368 367132
rect 156326 365664 156382 365673
rect 166644 365634 166672 367132
rect 176948 365702 176976 367132
rect 177040 365702 177068 387246
rect 182086 377768 182142 377777
rect 182086 377703 182142 377712
rect 182100 369345 182128 377703
rect 183572 370598 183600 389166
rect 194782 387424 194838 387433
rect 194626 387382 194782 387410
rect 205100 387394 205128 441118
rect 205192 419490 205220 441238
rect 207018 431760 207074 431769
rect 207018 431695 207074 431704
rect 209686 431760 209742 431769
rect 209686 431695 209742 431704
rect 207032 423201 207060 431695
rect 209700 423201 209728 431695
rect 211172 427174 211200 444450
rect 222292 444440 222344 444446
rect 222292 444382 222344 444388
rect 222304 441946 222332 444382
rect 222304 441918 222640 441946
rect 211264 441238 212336 441266
rect 232944 441238 233280 441266
rect 211160 427168 211212 427174
rect 211160 427110 211212 427116
rect 207018 423192 207074 423201
rect 207018 423127 207074 423136
rect 209686 423192 209742 423201
rect 209686 423127 209742 423136
rect 205180 419484 205232 419490
rect 205180 419426 205232 419432
rect 211264 419422 211292 441238
rect 233252 436626 233280 441238
rect 233240 436620 233292 436626
rect 233240 436562 233292 436568
rect 211988 427168 212040 427174
rect 211988 427110 212040 427116
rect 212000 421682 212028 427110
rect 212000 421654 212336 421682
rect 222640 421110 222976 421138
rect 222948 419422 222976 421110
rect 232608 421110 232944 421138
rect 232608 419490 232636 421110
rect 232596 419484 232648 419490
rect 232596 419426 232648 419432
rect 211252 419416 211304 419422
rect 211252 419358 211304 419364
rect 222936 419416 222988 419422
rect 222936 419358 222988 419364
rect 222200 416900 222252 416906
rect 222200 416842 222252 416848
rect 222212 414882 222240 416842
rect 232964 416832 233016 416838
rect 232964 416774 233016 416780
rect 222212 414854 222364 414882
rect 232668 414582 232912 414610
rect 211264 414310 212060 414338
rect 232780 414316 232832 414322
rect 207018 404288 207074 404297
rect 207018 404223 207074 404232
rect 207032 395865 207060 404223
rect 207018 395856 207074 395865
rect 207018 395791 207074 395800
rect 211264 391882 211292 414310
rect 232780 414258 232832 414264
rect 211712 397452 211764 397458
rect 211712 397394 211764 397400
rect 211724 394754 211752 397394
rect 232792 394754 232820 414258
rect 211724 394726 212060 394754
rect 232668 394726 232820 394754
rect 222364 394046 222700 394074
rect 222672 391921 222700 394046
rect 232884 391950 232912 414582
rect 232976 414322 233004 416774
rect 232964 414316 233016 414322
rect 232964 414258 233016 414264
rect 232872 391944 232924 391950
rect 222658 391912 222714 391921
rect 211252 391876 211304 391882
rect 232872 391886 232924 391892
rect 222658 391847 222714 391856
rect 211252 391818 211304 391824
rect 211252 389292 211304 389298
rect 211252 389234 211304 389240
rect 194782 387359 194838 387368
rect 205088 387388 205140 387394
rect 205088 387330 205140 387336
rect 183664 387246 184322 387274
rect 204930 387246 205220 387274
rect 183560 370592 183612 370598
rect 183560 370534 183612 370540
rect 182086 369336 182142 369345
rect 182086 369271 182142 369280
rect 176936 365696 176988 365702
rect 176936 365638 176988 365644
rect 177028 365696 177080 365702
rect 177028 365638 177080 365644
rect 183664 365634 183692 387246
rect 205088 387184 205140 387190
rect 205088 387126 205140 387132
rect 184020 370592 184072 370598
rect 184020 370534 184072 370540
rect 184032 367690 184060 370534
rect 184032 367662 184322 367690
rect 194612 365634 194640 367132
rect 204916 365702 204944 367132
rect 204904 365696 204956 365702
rect 204904 365638 204956 365644
rect 156326 365599 156382 365608
rect 166632 365628 166684 365634
rect 166632 365570 166684 365576
rect 183652 365628 183704 365634
rect 183652 365570 183704 365576
rect 194600 365628 194652 365634
rect 194600 365570 194652 365576
rect 184020 363112 184072 363118
rect 184020 363054 184072 363060
rect 204904 363112 204956 363118
rect 204904 363054 204956 363060
rect 176844 363044 176896 363050
rect 176844 362986 176896 362992
rect 156328 362976 156380 362982
rect 156328 362918 156380 362924
rect 156340 360890 156368 362918
rect 156032 360862 156368 360890
rect 165986 360496 166042 360505
rect 166042 360454 166336 360482
rect 165986 360431 166042 360440
rect 176640 360318 176792 360346
rect 154486 350296 154542 350305
rect 154486 350231 154542 350240
rect 154500 341873 154528 350231
rect 154486 341864 154542 341873
rect 154486 341799 154542 341808
rect 176764 340882 176792 360318
rect 176752 340876 176804 340882
rect 176752 340818 176804 340824
rect 176856 340490 176884 362986
rect 177304 362976 177356 362982
rect 177304 362918 177356 362924
rect 177316 342922 177344 362918
rect 184032 360876 184060 363054
rect 194324 363044 194376 363050
rect 194324 362986 194376 362992
rect 194336 360876 194364 362986
rect 204812 362976 204864 362982
rect 204812 362918 204864 362924
rect 204654 360318 204760 360346
rect 204732 360262 204760 360318
rect 204720 360256 204772 360262
rect 204720 360198 204772 360204
rect 178038 350296 178094 350305
rect 178038 350231 178094 350240
rect 182086 350296 182142 350305
rect 182086 350231 182142 350240
rect 177304 342916 177356 342922
rect 177304 342858 177356 342864
rect 178052 341737 178080 350231
rect 182100 342009 182128 350231
rect 183652 342916 183704 342922
rect 183652 342858 183704 342864
rect 182086 342000 182142 342009
rect 182086 341935 182142 341944
rect 178038 341728 178094 341737
rect 178038 341663 178094 341672
rect 176936 340876 176988 340882
rect 176936 340818 176988 340824
rect 176640 340462 176884 340490
rect 156032 340054 156092 340082
rect 166336 340054 166672 340082
rect 156064 337958 156092 340054
rect 166644 338026 166672 340054
rect 176948 338094 176976 340818
rect 183664 340762 183692 342858
rect 204824 340762 204852 362918
rect 204916 342650 204944 363054
rect 204996 360256 205048 360262
rect 204996 360198 205048 360204
rect 204904 342644 204956 342650
rect 204904 342586 204956 342592
rect 183664 340734 184046 340762
rect 204654 340734 204852 340762
rect 194336 338094 194364 340068
rect 176936 338088 176988 338094
rect 176936 338030 176988 338036
rect 194324 338088 194376 338094
rect 194324 338030 194376 338036
rect 205008 338026 205036 360198
rect 166632 338020 166684 338026
rect 166632 337962 166684 337968
rect 204996 338020 205048 338026
rect 204996 337962 205048 337968
rect 156052 337952 156104 337958
rect 156052 337894 156104 337900
rect 156328 335436 156380 335442
rect 156328 335378 156380 335384
rect 156340 333948 156368 335378
rect 166632 335368 166684 335374
rect 166632 335310 166684 335316
rect 183560 335368 183612 335374
rect 183560 335310 183612 335316
rect 166644 333948 166672 335310
rect 176962 333254 177068 333282
rect 154488 332648 154540 332654
rect 154488 332590 154540 332596
rect 154500 323785 154528 332590
rect 154486 323776 154542 323785
rect 154486 323711 154542 323720
rect 156340 311817 156368 313140
rect 156326 311808 156382 311817
rect 166644 311778 166672 313140
rect 176948 311846 176976 313140
rect 177040 311846 177068 333254
rect 182086 323776 182142 323785
rect 182086 323711 182142 323720
rect 182100 315353 182128 323711
rect 182086 315344 182142 315353
rect 182086 315279 182142 315288
rect 183572 314634 183600 335310
rect 205100 333402 205128 387126
rect 205192 365702 205220 387246
rect 211160 385484 211212 385490
rect 211160 385426 211212 385432
rect 207018 377768 207074 377777
rect 207018 377703 207074 377712
rect 209686 377768 209742 377777
rect 209686 377703 209742 377712
rect 207032 368490 207060 377703
rect 209700 368490 209728 377703
rect 207020 368484 207072 368490
rect 207020 368426 207072 368432
rect 209688 368484 209740 368490
rect 209688 368426 209740 368432
rect 205180 365696 205232 365702
rect 205180 365638 205232 365644
rect 211172 365634 211200 385426
rect 211264 383654 211292 389234
rect 222292 389224 222344 389230
rect 222292 389166 222344 389172
rect 222304 387954 222332 389166
rect 222304 387926 222640 387954
rect 212000 387246 212336 387274
rect 232944 387246 233280 387274
rect 212000 385490 212028 387246
rect 233252 385490 233280 387246
rect 211988 385484 212040 385490
rect 211988 385426 212040 385432
rect 233240 385484 233292 385490
rect 233240 385426 233292 385432
rect 211264 383626 211936 383654
rect 211908 367690 211936 383626
rect 211908 367662 212336 367690
rect 222640 367118 222976 367146
rect 222948 365634 222976 367118
rect 232608 367118 232944 367146
rect 232608 365702 232636 367118
rect 232596 365696 232648 365702
rect 232596 365638 232648 365644
rect 211160 365628 211212 365634
rect 211160 365570 211212 365576
rect 222936 365628 222988 365634
rect 222936 365570 222988 365576
rect 222200 362976 222252 362982
rect 222200 362918 222252 362924
rect 232964 362976 233016 362982
rect 232964 362918 233016 362924
rect 222212 360890 222240 362918
rect 222212 360862 222364 360890
rect 232668 360590 232912 360618
rect 211264 360318 212060 360346
rect 207018 350296 207074 350305
rect 207018 350231 207074 350240
rect 207032 341873 207060 350231
rect 207018 341864 207074 341873
rect 207018 341799 207074 341808
rect 211264 338026 211292 360318
rect 232780 358828 232832 358834
rect 232780 358770 232832 358776
rect 211712 342644 211764 342650
rect 211712 342586 211764 342592
rect 211724 340762 211752 342586
rect 232792 340762 232820 358770
rect 211724 340734 212060 340762
rect 232668 340734 232820 340762
rect 222364 340054 222700 340082
rect 222672 338065 222700 340054
rect 232884 338094 232912 360590
rect 232976 358834 233004 362918
rect 232964 358828 233016 358834
rect 232964 358770 233016 358776
rect 232872 338088 232924 338094
rect 222658 338056 222714 338065
rect 211252 338020 211304 338026
rect 232872 338030 232924 338036
rect 222658 337991 222714 338000
rect 211252 337962 211304 337968
rect 211160 335436 211212 335442
rect 211160 335378 211212 335384
rect 205088 333396 205140 333402
rect 205088 333338 205140 333344
rect 194782 333296 194838 333305
rect 183664 333254 184322 333282
rect 194626 333254 194782 333282
rect 183560 314628 183612 314634
rect 183560 314570 183612 314576
rect 176936 311840 176988 311846
rect 176936 311782 176988 311788
rect 177028 311840 177080 311846
rect 177028 311782 177080 311788
rect 183664 311778 183692 333254
rect 204930 333254 205220 333282
rect 194782 333231 194838 333240
rect 205088 333192 205140 333198
rect 205088 333134 205140 333140
rect 184020 314628 184072 314634
rect 184020 314570 184072 314576
rect 184032 313698 184060 314570
rect 184032 313670 184322 313698
rect 194612 311778 194640 313140
rect 204916 311846 204944 313140
rect 204904 311840 204956 311846
rect 204904 311782 204956 311788
rect 156326 311743 156382 311752
rect 166632 311772 166684 311778
rect 166632 311714 166684 311720
rect 183652 311772 183704 311778
rect 183652 311714 183704 311720
rect 194600 311772 194652 311778
rect 194600 311714 194652 311720
rect 176936 309256 176988 309262
rect 176936 309198 176988 309204
rect 194324 309256 194376 309262
rect 194324 309198 194376 309204
rect 156328 309188 156380 309194
rect 156328 309130 156380 309136
rect 156340 306898 156368 309130
rect 156032 306870 156368 306898
rect 165986 306504 166042 306513
rect 166042 306462 166336 306490
rect 165986 306439 166042 306448
rect 176640 306326 176884 306354
rect 176856 297498 176884 306326
rect 176844 297492 176896 297498
rect 176844 297434 176896 297440
rect 176844 297288 176896 297294
rect 176844 297230 176896 297236
rect 154486 296304 154542 296313
rect 154486 296239 154542 296248
rect 154500 287881 154528 296239
rect 176752 292528 176804 292534
rect 176752 292470 176804 292476
rect 154486 287872 154542 287881
rect 154486 287807 154542 287816
rect 176764 286770 176792 292470
rect 176640 286742 176792 286770
rect 156032 286062 156092 286090
rect 166336 286062 166672 286090
rect 156064 284170 156092 286062
rect 166644 284238 166672 286062
rect 176856 284306 176884 297230
rect 176948 292534 176976 309198
rect 177304 309188 177356 309194
rect 177304 309130 177356 309136
rect 184020 309188 184072 309194
rect 184020 309130 184072 309136
rect 176936 292528 176988 292534
rect 176936 292470 176988 292476
rect 177316 289134 177344 309130
rect 184032 306884 184060 309130
rect 194336 306884 194364 309198
rect 204904 309188 204956 309194
rect 204904 309130 204956 309136
rect 204654 306326 204852 306354
rect 204824 303822 204852 306326
rect 204812 303816 204864 303822
rect 204812 303758 204864 303764
rect 204812 303680 204864 303686
rect 204812 303622 204864 303628
rect 182086 296304 182142 296313
rect 182086 296239 182142 296248
rect 177304 289128 177356 289134
rect 177304 289070 177356 289076
rect 182100 288017 182128 296239
rect 183744 289128 183796 289134
rect 183744 289070 183796 289076
rect 182086 288008 182142 288017
rect 182086 287943 182142 287952
rect 183756 286770 183784 289070
rect 204824 286770 204852 303622
rect 204916 288454 204944 309130
rect 204996 303816 205048 303822
rect 204996 303758 205048 303764
rect 204904 288448 204956 288454
rect 204904 288390 204956 288396
rect 183756 286742 184046 286770
rect 204654 286742 204852 286770
rect 194336 284306 194364 286076
rect 176844 284300 176896 284306
rect 176844 284242 176896 284248
rect 194324 284300 194376 284306
rect 194324 284242 194376 284248
rect 205008 284238 205036 303758
rect 166632 284232 166684 284238
rect 166632 284174 166684 284180
rect 204996 284232 205048 284238
rect 204996 284174 205048 284180
rect 156052 284164 156104 284170
rect 156052 284106 156104 284112
rect 166632 281580 166684 281586
rect 166632 281522 166684 281528
rect 183652 281580 183704 281586
rect 183652 281522 183704 281528
rect 166644 279956 166672 281522
rect 155972 279262 156354 279290
rect 176962 279262 177068 279290
rect 154488 278792 154540 278798
rect 154488 278734 154540 278740
rect 154500 269793 154528 278734
rect 154486 269784 154542 269793
rect 154486 269719 154542 269728
rect 155972 256562 156000 279262
rect 156340 256601 156368 259148
rect 166644 256630 166672 259148
rect 176948 256698 176976 259148
rect 177040 256698 177068 279262
rect 182086 278080 182142 278089
rect 182086 278015 182142 278024
rect 182100 269793 182128 278015
rect 183560 272604 183612 272610
rect 183560 272546 183612 272552
rect 182086 269784 182142 269793
rect 182086 269719 182142 269728
rect 176936 256692 176988 256698
rect 176936 256634 176988 256640
rect 177028 256692 177080 256698
rect 177028 256634 177080 256640
rect 183572 256630 183600 272546
rect 183664 267734 183692 281522
rect 205100 279410 205128 333134
rect 205192 311846 205220 333254
rect 207020 332648 207072 332654
rect 207020 332590 207072 332596
rect 209688 332648 209740 332654
rect 209688 332590 209740 332596
rect 207032 323785 207060 332590
rect 209700 323785 209728 332590
rect 207018 323776 207074 323785
rect 207018 323711 207074 323720
rect 209686 323776 209742 323785
rect 209686 323711 209742 323720
rect 211172 314634 211200 335378
rect 222384 335368 222436 335374
rect 222384 335310 222436 335316
rect 222396 333962 222424 335310
rect 222396 333934 222640 333962
rect 211264 333254 212336 333282
rect 232944 333254 233280 333282
rect 211160 314628 211212 314634
rect 211160 314570 211212 314576
rect 205180 311840 205232 311846
rect 205180 311782 205232 311788
rect 211264 311778 211292 333254
rect 233252 329526 233280 333254
rect 233240 329520 233292 329526
rect 233240 329462 233292 329468
rect 211988 314628 212040 314634
rect 211988 314570 212040 314576
rect 212000 313698 212028 314570
rect 212000 313670 212336 313698
rect 222640 313126 222976 313154
rect 222948 311778 222976 313126
rect 232608 313126 232944 313154
rect 232608 311846 232636 313126
rect 232596 311840 232648 311846
rect 232596 311782 232648 311788
rect 211252 311772 211304 311778
rect 211252 311714 211304 311720
rect 222936 311772 222988 311778
rect 222936 311714 222988 311720
rect 209044 309188 209096 309194
rect 209044 309130 209096 309136
rect 222200 309188 222252 309194
rect 222200 309130 222252 309136
rect 232964 309188 233016 309194
rect 232964 309130 233016 309136
rect 209056 303686 209084 309130
rect 222212 306898 222240 309130
rect 222212 306870 222364 306898
rect 211264 306326 212060 306354
rect 232668 306326 232912 306354
rect 209044 303680 209096 303686
rect 209044 303622 209096 303628
rect 207018 296304 207074 296313
rect 207018 296239 207074 296248
rect 207032 287881 207060 296239
rect 207018 287872 207074 287881
rect 207018 287807 207074 287816
rect 211264 284238 211292 306326
rect 232780 301572 232832 301578
rect 232780 301514 232832 301520
rect 211712 288448 211764 288454
rect 211712 288390 211764 288396
rect 211724 286770 211752 288390
rect 232792 286770 232820 301514
rect 211724 286742 212060 286770
rect 232668 286742 232820 286770
rect 222364 286062 222700 286090
rect 211252 284232 211304 284238
rect 222672 284209 222700 286062
rect 232884 284306 232912 306326
rect 232976 301578 233004 309130
rect 232964 301572 233016 301578
rect 232964 301514 233016 301520
rect 232872 284300 232924 284306
rect 232872 284242 232924 284248
rect 211252 284174 211304 284180
rect 222658 284200 222714 284209
rect 222658 284135 222714 284144
rect 211252 281648 211304 281654
rect 211252 281590 211304 281596
rect 205088 279404 205140 279410
rect 205088 279346 205140 279352
rect 194782 279304 194838 279313
rect 184032 279262 184322 279290
rect 194626 279262 194782 279290
rect 184032 272610 184060 279262
rect 204930 279262 205220 279290
rect 194782 279239 194838 279248
rect 205088 279200 205140 279206
rect 205088 279142 205140 279148
rect 184020 272604 184072 272610
rect 184020 272546 184072 272552
rect 183664 267706 183968 267734
rect 183940 259706 183968 267706
rect 183940 259678 184322 259706
rect 194612 256630 194640 259148
rect 204916 256698 204944 259148
rect 204904 256692 204956 256698
rect 204904 256634 204956 256640
rect 166632 256624 166684 256630
rect 156326 256592 156382 256601
rect 155960 256556 156012 256562
rect 166632 256566 166684 256572
rect 183560 256624 183612 256630
rect 183560 256566 183612 256572
rect 194600 256624 194652 256630
rect 194600 256566 194652 256572
rect 156326 256527 156382 256536
rect 155960 256498 156012 256504
rect 177028 255400 177080 255406
rect 177028 255342 177080 255348
rect 194324 255400 194376 255406
rect 194324 255342 194376 255348
rect 156328 255332 156380 255338
rect 156328 255274 156380 255280
rect 156340 252906 156368 255274
rect 156032 252878 156368 252906
rect 165986 252648 166042 252657
rect 166042 252606 166336 252634
rect 165986 252583 166042 252592
rect 177040 252362 177068 255342
rect 177304 255332 177356 255338
rect 177304 255274 177356 255280
rect 184020 255332 184072 255338
rect 184020 255274 184072 255280
rect 176640 252334 176792 252362
rect 176764 251394 176792 252334
rect 176948 252334 177068 252362
rect 176752 251388 176804 251394
rect 176752 251330 176804 251336
rect 176948 249098 176976 252334
rect 177028 251388 177080 251394
rect 177028 251330 177080 251336
rect 176764 249070 176976 249098
rect 154486 242312 154542 242321
rect 154486 242247 154542 242256
rect 154500 233238 154528 242247
rect 154488 233232 154540 233238
rect 154488 233174 154540 233180
rect 176764 232778 176792 249070
rect 177040 244338 177068 251330
rect 176640 232750 176792 232778
rect 176856 244310 177068 244338
rect 156032 232070 156092 232098
rect 166336 232070 166672 232098
rect 156064 230314 156092 232070
rect 166644 230382 166672 232070
rect 176856 230450 176884 244310
rect 177316 235278 177344 255274
rect 184032 252892 184060 255274
rect 194336 252892 194364 255342
rect 204996 255332 205048 255338
rect 204996 255274 205048 255280
rect 205008 252362 205036 255274
rect 204654 252334 204760 252362
rect 204732 252278 204760 252334
rect 204916 252334 205036 252362
rect 204720 252272 204772 252278
rect 204720 252214 204772 252220
rect 204812 250572 204864 250578
rect 204812 250514 204864 250520
rect 178038 242312 178094 242321
rect 178038 242247 178094 242256
rect 182086 242312 182142 242321
rect 182086 242247 182142 242256
rect 177304 235272 177356 235278
rect 177304 235214 177356 235220
rect 178052 234025 178080 242247
rect 182100 234025 182128 242247
rect 183652 235272 183704 235278
rect 183652 235214 183704 235220
rect 178038 234016 178094 234025
rect 178038 233951 178094 233960
rect 182086 234016 182142 234025
rect 182086 233951 182142 233960
rect 183664 232778 183692 235214
rect 204824 232778 204852 250514
rect 204916 235482 204944 252334
rect 204996 252272 205048 252278
rect 204996 252214 205048 252220
rect 204904 235476 204956 235482
rect 204904 235418 204956 235424
rect 183664 232750 184046 232778
rect 204654 232750 204852 232778
rect 194336 230450 194364 232084
rect 176844 230444 176896 230450
rect 176844 230386 176896 230392
rect 194324 230444 194376 230450
rect 194324 230386 194376 230392
rect 205008 230382 205036 252214
rect 166632 230376 166684 230382
rect 166632 230318 166684 230324
rect 204996 230376 205048 230382
rect 204996 230318 205048 230324
rect 156052 230308 156104 230314
rect 156052 230250 156104 230256
rect 166632 227928 166684 227934
rect 166632 227870 166684 227876
rect 156328 227860 156380 227866
rect 156328 227802 156380 227808
rect 156340 225964 156368 227802
rect 166644 225964 166672 227870
rect 183928 227792 183980 227798
rect 183928 227734 183980 227740
rect 176962 225270 177068 225298
rect 154486 224224 154542 224233
rect 154486 224159 154542 224168
rect 154500 215801 154528 224159
rect 154486 215792 154542 215801
rect 154486 215727 154542 215736
rect 156340 202881 156368 205020
rect 156326 202872 156382 202881
rect 156326 202807 156382 202816
rect 166644 202774 166672 205020
rect 176948 202842 176976 205020
rect 177040 202842 177068 225270
rect 182086 224088 182142 224097
rect 182086 224023 182142 224032
rect 182100 215801 182128 224023
rect 183560 222352 183612 222358
rect 183560 222294 183612 222300
rect 182086 215792 182142 215801
rect 182086 215727 182142 215736
rect 176936 202836 176988 202842
rect 176936 202778 176988 202784
rect 177028 202836 177080 202842
rect 177028 202778 177080 202784
rect 183572 202774 183600 222294
rect 183940 205714 183968 227734
rect 205100 225418 205128 279142
rect 205192 256698 205220 279262
rect 207020 278792 207072 278798
rect 207020 278734 207072 278740
rect 209688 278792 209740 278798
rect 209688 278734 209740 278740
rect 207032 269793 207060 278734
rect 209700 269793 209728 278734
rect 211160 272604 211212 272610
rect 211160 272546 211212 272552
rect 207018 269784 207074 269793
rect 207018 269719 207074 269728
rect 209686 269784 209742 269793
rect 209686 269719 209742 269728
rect 205180 256692 205232 256698
rect 205180 256634 205232 256640
rect 211172 256630 211200 272546
rect 211264 267734 211292 281590
rect 222292 281580 222344 281586
rect 222292 281522 222344 281528
rect 222304 279970 222332 281522
rect 222304 279942 222640 279970
rect 212000 279262 212336 279290
rect 232944 279262 233096 279290
rect 212000 272610 212028 279262
rect 211988 272604 212040 272610
rect 211988 272546 212040 272552
rect 211264 267706 211936 267734
rect 211908 259706 211936 267706
rect 211908 259678 212336 259706
rect 222640 259134 222976 259162
rect 222948 256630 222976 259134
rect 232608 259134 232944 259162
rect 232608 256698 232636 259134
rect 233068 256698 233096 279262
rect 232596 256692 232648 256698
rect 232596 256634 232648 256640
rect 233056 256692 233108 256698
rect 233056 256634 233108 256640
rect 211160 256624 211212 256630
rect 211160 256566 211212 256572
rect 222936 256624 222988 256630
rect 222936 256566 222988 256572
rect 208400 255332 208452 255338
rect 208400 255274 208452 255280
rect 222200 255332 222252 255338
rect 222200 255274 222252 255280
rect 232964 255332 233016 255338
rect 232964 255274 233016 255280
rect 208412 250578 208440 255274
rect 222212 252906 222240 255274
rect 222212 252878 222364 252906
rect 232668 252606 232912 252634
rect 211264 252334 212060 252362
rect 208400 250572 208452 250578
rect 208400 250514 208452 250520
rect 207018 242312 207074 242321
rect 207018 242247 207074 242256
rect 209686 242312 209742 242321
rect 209686 242247 209742 242256
rect 207032 233238 207060 242247
rect 209700 233238 209728 242247
rect 207020 233232 207072 233238
rect 207020 233174 207072 233180
rect 209688 233232 209740 233238
rect 209688 233174 209740 233180
rect 211264 230382 211292 252334
rect 232780 251864 232832 251870
rect 232780 251806 232832 251812
rect 211712 235476 211764 235482
rect 211712 235418 211764 235424
rect 211724 232778 211752 235418
rect 232792 232778 232820 251806
rect 211724 232750 212060 232778
rect 232668 232750 232820 232778
rect 222364 232070 222700 232098
rect 222672 230489 222700 232070
rect 222658 230480 222714 230489
rect 232884 230450 232912 252606
rect 232976 251870 233004 255274
rect 232964 251864 233016 251870
rect 232964 251806 233016 251812
rect 222658 230415 222714 230424
rect 232872 230444 232924 230450
rect 232872 230386 232924 230392
rect 211252 230376 211304 230382
rect 211252 230318 211304 230324
rect 211896 227860 211948 227866
rect 211896 227802 211948 227808
rect 205088 225412 205140 225418
rect 205088 225354 205140 225360
rect 194782 225312 194838 225321
rect 184032 225270 184322 225298
rect 194626 225270 194782 225298
rect 184032 222358 184060 225270
rect 204930 225270 205220 225298
rect 194782 225247 194838 225256
rect 205088 225208 205140 225214
rect 205088 225150 205140 225156
rect 184020 222352 184072 222358
rect 184020 222294 184072 222300
rect 183940 205686 184322 205714
rect 194626 205006 195008 205034
rect 194980 202774 195008 205006
rect 204640 205006 204930 205034
rect 204640 202842 204668 205006
rect 204628 202836 204680 202842
rect 204628 202778 204680 202784
rect 166632 202768 166684 202774
rect 166632 202710 166684 202716
rect 183560 202768 183612 202774
rect 183560 202710 183612 202716
rect 194968 202768 195020 202774
rect 194968 202710 195020 202716
rect 156328 200388 156380 200394
rect 156328 200330 156380 200336
rect 177304 200388 177356 200394
rect 177304 200330 177356 200336
rect 156340 198914 156368 200330
rect 165988 200320 166040 200326
rect 165988 200262 166040 200268
rect 156032 198886 156368 198914
rect 166000 198914 166028 200262
rect 176752 200252 176804 200258
rect 176752 200194 176804 200200
rect 176660 200184 176712 200190
rect 176660 200126 176712 200132
rect 176672 198914 176700 200126
rect 166000 198886 166336 198914
rect 176640 198886 176700 198914
rect 154486 188320 154542 188329
rect 154486 188255 154542 188264
rect 154500 179382 154528 188255
rect 154488 179376 154540 179382
rect 154488 179318 154540 179324
rect 176764 178786 176792 200194
rect 177316 181490 177344 200330
rect 184020 200320 184072 200326
rect 184020 200262 184072 200268
rect 204904 200320 204956 200326
rect 204904 200262 204956 200268
rect 184032 198900 184060 200262
rect 194324 200252 194376 200258
rect 194324 200194 194376 200200
rect 194336 198900 194364 200194
rect 204812 200184 204864 200190
rect 204812 200126 204864 200132
rect 204720 198280 204772 198286
rect 204654 198228 204720 198234
rect 204654 198222 204772 198228
rect 204654 198206 204760 198222
rect 178038 196752 178094 196761
rect 178038 196687 178094 196696
rect 182086 196752 182142 196761
rect 182086 196687 182142 196696
rect 178052 188329 178080 196687
rect 182100 188329 182128 196687
rect 178038 188320 178094 188329
rect 178038 188255 178094 188264
rect 182086 188320 182142 188329
rect 182086 188255 182142 188264
rect 177304 181484 177356 181490
rect 177304 181426 177356 181432
rect 183744 181484 183796 181490
rect 183744 181426 183796 181432
rect 176640 178758 176792 178786
rect 183756 178786 183784 181426
rect 204824 178786 204852 200126
rect 204916 180878 204944 200262
rect 204996 198280 205048 198286
rect 204996 198222 205048 198228
rect 204904 180872 204956 180878
rect 204904 180814 204956 180820
rect 183756 178758 184046 178786
rect 204654 178758 204852 178786
rect 156032 178078 156092 178106
rect 166336 178078 166672 178106
rect 156064 176526 156092 178078
rect 166644 176662 166672 178078
rect 166632 176656 166684 176662
rect 166632 176598 166684 176604
rect 194336 176594 194364 178092
rect 205008 176662 205036 198222
rect 204996 176656 205048 176662
rect 204996 176598 205048 176604
rect 194324 176588 194376 176594
rect 194324 176530 194376 176536
rect 156052 176520 156104 176526
rect 156052 176462 156104 176468
rect 166632 174072 166684 174078
rect 166632 174014 166684 174020
rect 153844 172100 153896 172106
rect 153844 172042 153896 172048
rect 153856 149054 153884 172042
rect 166644 171972 166672 174014
rect 177304 174004 177356 174010
rect 177304 173946 177356 173952
rect 194600 174004 194652 174010
rect 194600 173946 194652 173952
rect 155880 171278 156354 171306
rect 176962 171278 177068 171306
rect 154486 170232 154542 170241
rect 154486 170167 154542 170176
rect 154500 161809 154528 170167
rect 154486 161800 154542 161809
rect 154486 161735 154542 161744
rect 155880 161474 155908 171278
rect 155236 161446 155908 161474
rect 153844 149048 153896 149054
rect 153844 148990 153896 148996
rect 155236 148918 155264 161446
rect 156340 148986 156368 151028
rect 156328 148980 156380 148986
rect 156328 148922 156380 148928
rect 166644 148918 166672 151028
rect 176948 149054 176976 151028
rect 177040 149054 177068 171278
rect 176936 149048 176988 149054
rect 176936 148990 176988 148996
rect 177028 149048 177080 149054
rect 177028 148990 177080 148996
rect 177316 148986 177344 173946
rect 178684 173936 178736 173942
rect 178684 173878 178736 173884
rect 184296 173936 184348 173942
rect 184296 173878 184348 173884
rect 178038 170368 178094 170377
rect 178038 170303 178094 170312
rect 178052 161809 178080 170303
rect 178038 161800 178094 161809
rect 178038 161735 178094 161744
rect 177304 148980 177356 148986
rect 177304 148922 177356 148928
rect 178696 148918 178724 173878
rect 183652 173868 183704 173874
rect 183652 173810 183704 173816
rect 183664 171134 183692 173810
rect 184308 171972 184336 173878
rect 194612 171972 194640 173946
rect 205100 171426 205128 225150
rect 205192 202842 205220 225270
rect 207018 224224 207074 224233
rect 207018 224159 207074 224168
rect 209686 224224 209742 224233
rect 209686 224159 209742 224168
rect 207032 215801 207060 224159
rect 209700 215801 209728 224159
rect 211160 222352 211212 222358
rect 211160 222294 211212 222300
rect 207018 215792 207074 215801
rect 207018 215727 207074 215736
rect 209686 215792 209742 215801
rect 209686 215727 209742 215736
rect 205180 202836 205232 202842
rect 205180 202778 205232 202784
rect 211172 202774 211200 222294
rect 211908 205714 211936 227802
rect 222292 227792 222344 227798
rect 222292 227734 222344 227740
rect 222304 225978 222332 227734
rect 222304 225950 222640 225978
rect 212000 225270 212336 225298
rect 232944 225270 233280 225298
rect 212000 222358 212028 225270
rect 211988 222352 212040 222358
rect 211988 222294 212040 222300
rect 233252 220726 233280 225270
rect 233240 220720 233292 220726
rect 233240 220662 233292 220668
rect 211908 205686 212336 205714
rect 222640 205006 222976 205034
rect 222948 202774 222976 205006
rect 232608 205006 232944 205034
rect 232608 202842 232636 205006
rect 232596 202836 232648 202842
rect 232596 202778 232648 202784
rect 211160 202768 211212 202774
rect 211160 202710 211212 202716
rect 222936 202768 222988 202774
rect 222936 202710 222988 202716
rect 222292 200184 222344 200190
rect 222292 200126 222344 200132
rect 232780 200184 232832 200190
rect 232780 200126 232832 200132
rect 222304 198914 222332 200126
rect 222304 198886 222364 198914
rect 232792 198354 232820 200126
rect 232780 198348 232832 198354
rect 232780 198290 232832 198296
rect 211264 198206 212060 198234
rect 232668 198206 232912 198234
rect 207018 188320 207074 188329
rect 207018 188255 207074 188264
rect 209686 188320 209742 188329
rect 209686 188255 209742 188264
rect 207032 179382 207060 188255
rect 209700 179382 209728 188255
rect 207020 179376 207072 179382
rect 207020 179318 207072 179324
rect 209688 179376 209740 179382
rect 209688 179318 209740 179324
rect 211264 176662 211292 198206
rect 232780 198144 232832 198150
rect 232780 198086 232832 198092
rect 211712 180872 211764 180878
rect 211712 180814 211764 180820
rect 211724 178786 211752 180814
rect 232792 178786 232820 198086
rect 211724 178758 212060 178786
rect 232668 178758 232820 178786
rect 222364 178078 222700 178106
rect 211252 176656 211304 176662
rect 222672 176633 222700 178078
rect 211252 176598 211304 176604
rect 222658 176624 222714 176633
rect 232884 176594 232912 198206
rect 222658 176559 222714 176568
rect 232872 176588 232924 176594
rect 232872 176530 232924 176536
rect 211252 174072 211304 174078
rect 211252 174014 211304 174020
rect 206284 173936 206336 173942
rect 206284 173878 206336 173884
rect 209780 173936 209832 173942
rect 209964 173936 210016 173942
rect 209832 173884 209964 173890
rect 209780 173878 210016 173884
rect 205088 171420 205140 171426
rect 205088 171362 205140 171368
rect 204930 171278 205220 171306
rect 205088 171216 205140 171222
rect 205088 171158 205140 171164
rect 183664 171106 183968 171134
rect 182086 170096 182142 170105
rect 182086 170031 182142 170040
rect 182100 161809 182128 170031
rect 182086 161800 182142 161809
rect 182086 161735 182142 161744
rect 183940 151722 183968 171106
rect 183940 151694 184322 151722
rect 194612 148986 194640 151028
rect 204916 149054 204944 151028
rect 204904 149048 204956 149054
rect 204904 148990 204956 148996
rect 194600 148980 194652 148986
rect 194600 148922 194652 148928
rect 155224 148912 155276 148918
rect 155224 148854 155276 148860
rect 166632 148912 166684 148918
rect 166632 148854 166684 148860
rect 178684 148912 178736 148918
rect 178684 148854 178736 148860
rect 156328 146532 156380 146538
rect 156328 146474 156380 146480
rect 180064 146532 180116 146538
rect 180064 146474 180116 146480
rect 184020 146532 184072 146538
rect 184020 146474 184072 146480
rect 204904 146532 204956 146538
rect 204904 146474 204956 146480
rect 155224 146396 155276 146402
rect 155224 146338 155276 146344
rect 154488 143676 154540 143682
rect 154488 143618 154540 143624
rect 154500 134337 154528 143618
rect 154486 134328 154542 134337
rect 154486 134263 154542 134272
rect 155236 122670 155264 146338
rect 156340 144922 156368 146474
rect 176844 146464 176896 146470
rect 176844 146406 176896 146412
rect 165988 146396 166040 146402
rect 165988 146338 166040 146344
rect 156032 144894 156368 144922
rect 166000 144922 166028 146338
rect 166000 144894 166336 144922
rect 176640 144214 176792 144242
rect 176764 124914 176792 144214
rect 176752 124908 176804 124914
rect 176752 124850 176804 124856
rect 176856 124794 176884 146406
rect 178684 146328 178736 146334
rect 178684 146270 178736 146276
rect 178038 142760 178094 142769
rect 178038 142695 178094 142704
rect 178052 134337 178080 142695
rect 178038 134328 178094 134337
rect 178038 134263 178094 134272
rect 176640 124766 176884 124794
rect 176752 124704 176804 124710
rect 176752 124646 176804 124652
rect 156018 123842 156046 124100
rect 166336 124086 166672 124114
rect 155972 123814 156046 123842
rect 155972 122738 156000 123814
rect 166644 122738 166672 124086
rect 176764 122806 176792 124646
rect 176752 122800 176804 122806
rect 176752 122742 176804 122748
rect 178696 122738 178724 146270
rect 180076 122806 180104 146474
rect 184032 144908 184060 146474
rect 194324 146464 194376 146470
rect 194324 146406 194376 146412
rect 194336 144908 194364 146406
rect 204812 146396 204864 146402
rect 204812 146338 204864 146344
rect 204628 146328 204680 146334
rect 204628 146270 204680 146276
rect 204640 144908 204668 146270
rect 182088 143608 182140 143614
rect 182088 143550 182140 143556
rect 182100 134337 182128 143550
rect 182086 134328 182142 134337
rect 182086 134263 182142 134272
rect 204824 124794 204852 146338
rect 204916 128314 204944 146474
rect 204904 128308 204956 128314
rect 204904 128250 204956 128256
rect 204654 124766 204852 124794
rect 184032 122806 184060 124100
rect 194336 122806 194364 124100
rect 180064 122800 180116 122806
rect 180064 122742 180116 122748
rect 184020 122800 184072 122806
rect 184020 122742 184072 122748
rect 194324 122800 194376 122806
rect 194324 122742 194376 122748
rect 155960 122732 156012 122738
rect 155960 122674 156012 122680
rect 166632 122732 166684 122738
rect 166632 122674 166684 122680
rect 178684 122732 178736 122738
rect 178684 122674 178736 122680
rect 155224 122664 155276 122670
rect 155224 122606 155276 122612
rect 166632 120284 166684 120290
rect 166632 120226 166684 120232
rect 156328 120216 156380 120222
rect 156328 120158 156380 120164
rect 156340 117980 156368 120158
rect 166644 117980 166672 120226
rect 183560 120216 183612 120222
rect 183560 120158 183612 120164
rect 176962 117286 177068 117314
rect 154486 116104 154542 116113
rect 154486 116039 154542 116048
rect 154500 107817 154528 116039
rect 154486 107808 154542 107817
rect 154486 107743 154542 107752
rect 156340 95169 156368 97036
rect 156326 95160 156382 95169
rect 166644 95130 166672 97036
rect 176948 95198 176976 97036
rect 177040 95198 177068 117286
rect 182086 116376 182142 116385
rect 182086 116311 182142 116320
rect 182100 107817 182128 116311
rect 182086 107808 182142 107817
rect 182086 107743 182142 107752
rect 183572 100298 183600 120158
rect 205100 117434 205128 171158
rect 205192 149054 205220 171278
rect 205180 149048 205232 149054
rect 205180 148990 205232 148996
rect 206296 148986 206324 173878
rect 209792 173862 210004 173878
rect 209688 171420 209740 171426
rect 209688 171362 209740 171368
rect 207018 170232 207074 170241
rect 207018 170167 207074 170176
rect 207032 161809 207060 170167
rect 209700 161809 209728 171362
rect 211264 171134 211292 174014
rect 211988 174004 212040 174010
rect 211988 173946 212040 173952
rect 212000 171986 212028 173946
rect 222292 173936 222344 173942
rect 222292 173878 222344 173884
rect 222304 171986 222332 173878
rect 212000 171958 212336 171986
rect 222304 171958 222640 171986
rect 232944 171278 233280 171306
rect 211264 171106 211936 171134
rect 207018 161800 207074 161809
rect 207018 161735 207074 161744
rect 209686 161800 209742 161809
rect 209686 161735 209742 161744
rect 211908 151722 211936 171106
rect 233252 166326 233280 171278
rect 233240 166320 233292 166326
rect 233240 166262 233292 166268
rect 211908 151694 212336 151722
rect 222640 151014 222976 151042
rect 222948 148986 222976 151014
rect 232608 151014 232944 151042
rect 232608 149054 232636 151014
rect 232596 149048 232648 149054
rect 232596 148990 232648 148996
rect 206284 148980 206336 148986
rect 206284 148922 206336 148928
rect 222936 148980 222988 148986
rect 222936 148922 222988 148928
rect 222200 146396 222252 146402
rect 222200 146338 222252 146344
rect 232780 146396 232832 146402
rect 232780 146338 232832 146344
rect 206284 146328 206336 146334
rect 206284 146270 206336 146276
rect 206296 122806 206324 146270
rect 222212 144922 222240 146338
rect 232320 146328 232372 146334
rect 232320 146270 232372 146276
rect 232332 144922 232360 146270
rect 222212 144894 222364 144922
rect 232332 144894 232668 144922
rect 211264 144214 212060 144242
rect 207020 143676 207072 143682
rect 207020 143618 207072 143624
rect 207032 134337 207060 143618
rect 209686 142760 209742 142769
rect 209686 142695 209742 142704
rect 209700 134337 209728 142695
rect 207018 134328 207074 134337
rect 207018 134263 207074 134272
rect 209686 134328 209742 134337
rect 209686 134263 209742 134272
rect 211264 122806 211292 144214
rect 211712 128308 211764 128314
rect 211712 128250 211764 128256
rect 211724 124794 211752 128250
rect 232792 124794 232820 146338
rect 211724 124766 212060 124794
rect 232668 124766 232820 124794
rect 222364 124086 222700 124114
rect 206284 122800 206336 122806
rect 206284 122742 206336 122748
rect 211252 122800 211304 122806
rect 211252 122742 211304 122748
rect 222672 122738 222700 124086
rect 222660 122732 222712 122738
rect 222660 122674 222712 122680
rect 211160 120284 211212 120290
rect 211160 120226 211212 120232
rect 205088 117428 205140 117434
rect 205088 117370 205140 117376
rect 194782 117328 194838 117337
rect 183664 117286 184322 117314
rect 194626 117286 194782 117314
rect 183560 100292 183612 100298
rect 183560 100234 183612 100240
rect 176936 95192 176988 95198
rect 176936 95134 176988 95140
rect 177028 95192 177080 95198
rect 177028 95134 177080 95140
rect 183664 95130 183692 117286
rect 204930 117286 205220 117314
rect 194782 117263 194838 117272
rect 205088 117224 205140 117230
rect 205088 117166 205140 117172
rect 184020 100292 184072 100298
rect 184020 100234 184072 100240
rect 184032 97730 184060 100234
rect 184032 97702 184322 97730
rect 194612 95130 194640 97036
rect 204916 95198 204944 97036
rect 204904 95192 204956 95198
rect 204904 95134 204956 95140
rect 156326 95095 156382 95104
rect 166632 95124 166684 95130
rect 166632 95066 166684 95072
rect 183652 95124 183704 95130
rect 183652 95066 183704 95072
rect 194600 95124 194652 95130
rect 194600 95066 194652 95072
rect 184020 92744 184072 92750
rect 184020 92686 184072 92692
rect 204904 92744 204956 92750
rect 204904 92686 204956 92692
rect 165988 92676 166040 92682
rect 165988 92618 166040 92624
rect 176752 92676 176804 92682
rect 176752 92618 176804 92624
rect 156328 92608 156380 92614
rect 156328 92550 156380 92556
rect 156340 90930 156368 92550
rect 156032 90902 156368 90930
rect 166000 90930 166028 92618
rect 176660 92540 176712 92546
rect 176660 92482 176712 92488
rect 176672 90930 176700 92482
rect 166000 90902 166336 90930
rect 176640 90902 176700 90930
rect 154486 88904 154542 88913
rect 154486 88839 154542 88848
rect 154500 80345 154528 88839
rect 154486 80336 154542 80345
rect 154486 80271 154542 80280
rect 176764 70666 176792 92618
rect 180064 92608 180116 92614
rect 180064 92550 180116 92556
rect 178684 92540 178736 92546
rect 178684 92482 178736 92488
rect 176640 70638 176792 70666
rect 156032 70094 156092 70122
rect 166336 70094 166672 70122
rect 156064 68882 156092 70094
rect 166644 69018 166672 70094
rect 178696 69018 178724 92482
rect 180076 69018 180104 92550
rect 184032 90916 184060 92686
rect 194324 92676 194376 92682
rect 194324 92618 194376 92624
rect 194336 90916 194364 92618
rect 204812 92608 204864 92614
rect 204812 92550 204864 92556
rect 204628 92540 204680 92546
rect 204628 92482 204680 92488
rect 204640 90916 204668 92482
rect 182086 88768 182142 88777
rect 182086 88703 182142 88712
rect 182100 80345 182128 88703
rect 182086 80336 182142 80345
rect 182086 80271 182142 80280
rect 204824 70666 204852 92550
rect 204916 73506 204944 92686
rect 204904 73500 204956 73506
rect 204904 73442 204956 73448
rect 204654 70638 204852 70666
rect 184032 69018 184060 70108
rect 194336 69018 194364 70108
rect 166632 69012 166684 69018
rect 166632 68954 166684 68960
rect 178684 69012 178736 69018
rect 178684 68954 178736 68960
rect 180064 69012 180116 69018
rect 180064 68954 180116 68960
rect 184020 69012 184072 69018
rect 184020 68954 184072 68960
rect 194324 69012 194376 69018
rect 194324 68954 194376 68960
rect 156052 68876 156104 68882
rect 156052 68818 156104 68824
rect 156328 66360 156380 66366
rect 156328 66302 156380 66308
rect 183652 66360 183704 66366
rect 183652 66302 183704 66308
rect 156340 63852 156368 66302
rect 166632 66292 166684 66298
rect 166632 66234 166684 66240
rect 182824 66292 182876 66298
rect 182824 66234 182876 66240
rect 166644 63852 166672 66234
rect 176962 63294 177068 63322
rect 154486 53816 154542 53825
rect 154486 53751 154542 53760
rect 154500 45257 154528 53751
rect 154486 45248 154542 45257
rect 154486 45183 154542 45192
rect 156340 41342 156368 43044
rect 156328 41336 156380 41342
rect 156328 41278 156380 41284
rect 166644 41274 166672 43044
rect 176948 41410 176976 43044
rect 177040 41410 177068 63294
rect 177304 61396 177356 61402
rect 177304 61338 177356 61344
rect 176936 41404 176988 41410
rect 176936 41346 176988 41352
rect 177028 41404 177080 41410
rect 177028 41346 177080 41352
rect 177316 41274 177344 61338
rect 182086 53816 182142 53825
rect 182086 53751 182142 53760
rect 182100 45393 182128 53751
rect 182086 45384 182142 45393
rect 182086 45319 182142 45328
rect 182836 41342 182864 66234
rect 183664 55214 183692 66302
rect 194600 66292 194652 66298
rect 194600 66234 194652 66240
rect 194612 63852 194640 66234
rect 205100 63442 205128 117166
rect 205192 95198 205220 117286
rect 209686 116512 209742 116521
rect 209686 116447 209742 116456
rect 207018 116104 207074 116113
rect 207018 116039 207074 116048
rect 207032 107817 207060 116039
rect 209700 107817 209728 116447
rect 207018 107808 207074 107817
rect 207018 107743 207074 107752
rect 209686 107808 209742 107817
rect 209686 107743 209742 107752
rect 211172 100298 211200 120226
rect 222292 120216 222344 120222
rect 222292 120158 222344 120164
rect 222304 117994 222332 120158
rect 222304 117966 222640 117994
rect 211264 117286 212336 117314
rect 232944 117286 233280 117314
rect 211160 100292 211212 100298
rect 211160 100234 211212 100240
rect 205180 95192 205232 95198
rect 205180 95134 205232 95140
rect 211264 95130 211292 117286
rect 233252 114578 233280 117286
rect 233240 114572 233292 114578
rect 233240 114514 233292 114520
rect 211988 100292 212040 100298
rect 211988 100234 212040 100240
rect 212000 97730 212028 100234
rect 212000 97702 212336 97730
rect 222640 97022 222976 97050
rect 222948 95130 222976 97022
rect 232608 97022 232944 97050
rect 232608 95198 232636 97022
rect 232596 95192 232648 95198
rect 232596 95134 232648 95140
rect 211252 95124 211304 95130
rect 211252 95066 211304 95072
rect 222936 95124 222988 95130
rect 222936 95066 222988 95072
rect 222200 92608 222252 92614
rect 222200 92550 222252 92556
rect 232780 92608 232832 92614
rect 232780 92550 232832 92556
rect 206284 92540 206336 92546
rect 206284 92482 206336 92488
rect 206296 69018 206324 92482
rect 222212 90930 222240 92550
rect 232320 92540 232372 92546
rect 232320 92482 232372 92488
rect 232332 90930 232360 92482
rect 222212 90902 222364 90930
rect 232332 90902 232668 90930
rect 211264 90222 212060 90250
rect 209688 89752 209740 89758
rect 209688 89694 209740 89700
rect 207018 88904 207074 88913
rect 207018 88839 207074 88848
rect 207032 80345 207060 88839
rect 209700 80345 209728 89694
rect 207018 80336 207074 80345
rect 207018 80271 207074 80280
rect 209686 80336 209742 80345
rect 209686 80271 209742 80280
rect 211264 69018 211292 90222
rect 211712 73500 211764 73506
rect 211712 73442 211764 73448
rect 211724 70666 211752 73442
rect 232792 70666 232820 92550
rect 211724 70638 212060 70666
rect 232668 70638 232820 70666
rect 222364 70094 222700 70122
rect 206284 69012 206336 69018
rect 206284 68954 206336 68960
rect 211252 69012 211304 69018
rect 211252 68954 211304 68960
rect 222672 68950 222700 70094
rect 222660 68944 222712 68950
rect 222660 68886 222712 68892
rect 211252 66428 211304 66434
rect 211252 66370 211304 66376
rect 206284 66292 206336 66298
rect 206284 66234 206336 66240
rect 205088 63436 205140 63442
rect 205088 63378 205140 63384
rect 184032 63294 184322 63322
rect 204930 63294 205220 63322
rect 184032 61402 184060 63294
rect 205088 63232 205140 63238
rect 205088 63174 205140 63180
rect 184020 61396 184072 61402
rect 184020 61338 184072 61344
rect 183664 55186 183968 55214
rect 183940 43738 183968 55186
rect 183940 43710 184322 43738
rect 194612 41342 194640 43044
rect 204916 41410 204944 43044
rect 204904 41404 204956 41410
rect 204904 41346 204956 41352
rect 182824 41336 182876 41342
rect 182824 41278 182876 41284
rect 194600 41336 194652 41342
rect 194600 41278 194652 41284
rect 166632 41268 166684 41274
rect 166632 41210 166684 41216
rect 177304 41268 177356 41274
rect 177304 41210 177356 41216
rect 205100 39438 205128 63174
rect 205192 41410 205220 63294
rect 205180 41404 205232 41410
rect 205180 41346 205232 41352
rect 206296 41342 206324 66234
rect 211264 55214 211292 66370
rect 222384 66360 222436 66366
rect 222384 66302 222436 66308
rect 211988 66292 212040 66298
rect 211988 66234 212040 66240
rect 212000 63866 212028 66234
rect 222396 63866 222424 66302
rect 212000 63838 212336 63866
rect 222396 63838 222640 63866
rect 232944 63294 233280 63322
rect 233252 59294 233280 63294
rect 233240 59288 233292 59294
rect 233240 59230 233292 59236
rect 211264 55186 211936 55214
rect 207018 53816 207074 53825
rect 207018 53751 207074 53760
rect 209686 53816 209742 53825
rect 209686 53751 209742 53760
rect 207032 45257 207060 53751
rect 209700 45257 209728 53751
rect 207018 45248 207074 45257
rect 207018 45183 207074 45192
rect 209686 45248 209742 45257
rect 209686 45183 209742 45192
rect 211908 43738 211936 55186
rect 211908 43710 212336 43738
rect 222640 43030 222976 43058
rect 222948 41342 222976 43030
rect 232608 43030 232944 43058
rect 232608 41410 232636 43030
rect 232596 41404 232648 41410
rect 232596 41346 232648 41352
rect 206284 41336 206336 41342
rect 206284 41278 206336 41284
rect 222936 41336 222988 41342
rect 222936 41278 222988 41284
rect 205088 39432 205140 39438
rect 205088 39374 205140 39380
rect 156328 38888 156380 38894
rect 156328 38830 156380 38836
rect 180064 38888 180116 38894
rect 180064 38830 180116 38836
rect 155224 38752 155276 38758
rect 155224 38694 155276 38700
rect 152464 38412 152516 38418
rect 152464 38354 152516 38360
rect 121092 36304 121144 36310
rect 121092 36246 121144 36252
rect 127084 36230 128018 36258
rect 148626 36230 148824 36258
rect 121000 36168 121052 36174
rect 121000 36110 121052 36116
rect 122838 34912 122894 34921
rect 122838 34847 122894 34856
rect 122852 26353 122880 34847
rect 122838 26344 122894 26353
rect 122838 26279 122894 26288
rect 120908 13252 120960 13258
rect 120908 13194 120960 13200
rect 100024 13184 100076 13190
rect 100024 13126 100076 13132
rect 110328 13184 110380 13190
rect 110328 13126 110380 13132
rect 127084 13122 127112 36230
rect 127716 18624 127768 18630
rect 127716 18566 127768 18572
rect 127728 16674 127756 18566
rect 127728 16646 128018 16674
rect 138308 13258 138336 16116
rect 148612 13802 148640 16116
rect 148600 13796 148652 13802
rect 148600 13738 148652 13744
rect 138296 13252 138348 13258
rect 138296 13194 138348 13200
rect 148796 13190 148824 36230
rect 150438 34776 150494 34785
rect 150438 34711 150494 34720
rect 154486 34776 154542 34785
rect 154486 34711 154542 34720
rect 150452 26353 150480 34711
rect 154500 26353 154528 34711
rect 150438 26344 150494 26353
rect 150438 26279 150494 26288
rect 154486 26344 154542 26353
rect 154486 26279 154542 26288
rect 155236 13802 155264 38694
rect 156340 36938 156368 38830
rect 176844 38820 176896 38826
rect 176844 38762 176896 38768
rect 165988 38752 166040 38758
rect 165988 38694 166040 38700
rect 156032 36910 156368 36938
rect 166000 36938 166028 38694
rect 166000 36910 166336 36938
rect 176640 36230 176792 36258
rect 176764 21418 176792 36230
rect 176752 21412 176804 21418
rect 176752 21354 176804 21360
rect 176856 16674 176884 38762
rect 178684 38684 178736 38690
rect 178684 38626 178736 38632
rect 178038 34912 178094 34921
rect 178038 34847 178094 34856
rect 178052 26353 178080 34847
rect 178038 26344 178094 26353
rect 178038 26279 178094 26288
rect 176936 21412 176988 21418
rect 176936 21354 176988 21360
rect 176640 16646 176884 16674
rect 156032 16102 156092 16130
rect 166336 16102 166672 16130
rect 155224 13796 155276 13802
rect 155224 13738 155276 13744
rect 148784 13184 148836 13190
rect 148784 13126 148836 13132
rect 156064 13122 156092 16102
rect 166644 13802 166672 16102
rect 166632 13796 166684 13802
rect 166632 13738 166684 13744
rect 176948 13258 176976 21354
rect 178696 13802 178724 38626
rect 180076 13802 180104 38830
rect 194324 38820 194376 38826
rect 194324 38762 194376 38768
rect 184020 38752 184072 38758
rect 184020 38694 184072 38700
rect 184032 36924 184060 38694
rect 194336 36924 194364 38762
rect 204904 38752 204956 38758
rect 204904 38694 204956 38700
rect 204628 38684 204680 38690
rect 204628 38626 204680 38632
rect 204812 38684 204864 38690
rect 204812 38626 204864 38632
rect 204640 36924 204668 38626
rect 182086 34912 182142 34921
rect 182086 34847 182142 34856
rect 182100 26353 182128 34847
rect 182086 26344 182142 26353
rect 182086 26279 182142 26288
rect 204824 16674 204852 38626
rect 204916 18018 204944 38694
rect 222200 38684 222252 38690
rect 222200 38626 222252 38632
rect 222212 36938 222240 38626
rect 222212 36910 222364 36938
rect 211264 36230 212060 36258
rect 232668 36230 232820 36258
rect 207018 34776 207074 34785
rect 207018 34711 207074 34720
rect 207032 26353 207060 34711
rect 207018 26344 207074 26353
rect 207018 26279 207074 26288
rect 204904 18012 204956 18018
rect 204904 17954 204956 17960
rect 204654 16646 204852 16674
rect 184032 13802 184060 16116
rect 178684 13796 178736 13802
rect 178684 13738 178736 13744
rect 180064 13796 180116 13802
rect 180064 13738 180116 13744
rect 184020 13796 184072 13802
rect 184020 13738 184072 13744
rect 194336 13258 194364 16116
rect 176936 13252 176988 13258
rect 176936 13194 176988 13200
rect 194324 13252 194376 13258
rect 194324 13194 194376 13200
rect 211264 13190 211292 36230
rect 211712 18012 211764 18018
rect 211712 17954 211764 17960
rect 211724 16674 211752 17954
rect 211724 16646 212060 16674
rect 222364 16102 222700 16130
rect 222672 13802 222700 16102
rect 232608 16102 232668 16130
rect 222660 13796 222712 13802
rect 222660 13738 222712 13744
rect 232608 13433 232636 16102
rect 232594 13424 232650 13433
rect 232594 13359 232650 13368
rect 232792 13258 232820 36230
rect 233896 15094 233924 700266
rect 233976 659728 234028 659734
rect 233976 659670 234028 659676
rect 233988 634710 234016 659670
rect 233976 634704 234028 634710
rect 233976 634646 234028 634652
rect 234068 605872 234120 605878
rect 234068 605814 234120 605820
rect 233976 599752 234028 599758
rect 233976 599694 234028 599700
rect 233988 580990 234016 599694
rect 233976 580984 234028 580990
rect 233976 580926 234028 580932
rect 234080 580922 234108 605814
rect 234068 580916 234120 580922
rect 234068 580858 234120 580864
rect 233976 550588 234028 550594
rect 233976 550530 234028 550536
rect 233988 527066 234016 550530
rect 234068 548548 234120 548554
rect 234068 548490 234120 548496
rect 234080 527134 234108 548490
rect 234068 527128 234120 527134
rect 234068 527070 234120 527076
rect 233976 527060 234028 527066
rect 233976 527002 234028 527008
rect 234068 498228 234120 498234
rect 234068 498170 234120 498176
rect 233976 492584 234028 492590
rect 233976 492526 234028 492532
rect 233988 473346 234016 492526
rect 233976 473340 234028 473346
rect 233976 473282 234028 473288
rect 234080 473278 234108 498170
rect 234068 473272 234120 473278
rect 234068 473214 234120 473220
rect 233976 436620 234028 436626
rect 233976 436562 234028 436568
rect 233988 419490 234016 436562
rect 233976 419484 234028 419490
rect 233976 419426 234028 419432
rect 233976 389224 234028 389230
rect 233976 389166 234028 389172
rect 233988 365634 234016 389166
rect 234068 385484 234120 385490
rect 234068 385426 234120 385432
rect 234080 365702 234108 385426
rect 234068 365696 234120 365702
rect 234068 365638 234120 365644
rect 233976 365628 234028 365634
rect 233976 365570 234028 365576
rect 233976 335368 234028 335374
rect 233976 335310 234028 335316
rect 233988 311778 234016 335310
rect 234068 329520 234120 329526
rect 234068 329462 234120 329468
rect 234080 311846 234108 329462
rect 234068 311840 234120 311846
rect 234068 311782 234120 311788
rect 233976 311772 234028 311778
rect 233976 311714 234028 311720
rect 233976 280152 234028 280158
rect 233976 280094 234028 280100
rect 233988 256630 234016 280094
rect 233976 256624 234028 256630
rect 233976 256566 234028 256572
rect 233976 227792 234028 227798
rect 233976 227734 234028 227740
rect 233988 202774 234016 227734
rect 234068 220720 234120 220726
rect 234068 220662 234120 220668
rect 234080 202842 234108 220662
rect 234068 202836 234120 202842
rect 234068 202778 234120 202784
rect 233976 202768 234028 202774
rect 233976 202710 234028 202716
rect 234068 173936 234120 173942
rect 234068 173878 234120 173884
rect 233976 166320 234028 166326
rect 233976 166262 234028 166268
rect 233988 149054 234016 166262
rect 233976 149048 234028 149054
rect 233976 148990 234028 148996
rect 234080 148986 234108 173878
rect 234068 148980 234120 148986
rect 234068 148922 234120 148928
rect 233976 146328 234028 146334
rect 233976 146270 234028 146276
rect 233988 122738 234016 146270
rect 233976 122732 234028 122738
rect 233976 122674 234028 122680
rect 233976 120148 234028 120154
rect 233976 120090 234028 120096
rect 233988 95130 234016 120090
rect 234068 114572 234120 114578
rect 234068 114514 234120 114520
rect 234080 95198 234108 114514
rect 234068 95192 234120 95198
rect 234068 95134 234120 95140
rect 233976 95124 234028 95130
rect 233976 95066 234028 95072
rect 233976 92540 234028 92546
rect 233976 92482 234028 92488
rect 233988 68950 234016 92482
rect 233976 68944 234028 68950
rect 233976 68886 234028 68892
rect 234068 66292 234120 66298
rect 234068 66234 234120 66240
rect 233976 59288 234028 59294
rect 233976 59230 234028 59236
rect 233988 41410 234016 59230
rect 233976 41404 234028 41410
rect 233976 41346 234028 41352
rect 234080 41342 234108 66234
rect 234068 41336 234120 41342
rect 234068 41278 234120 41284
rect 233976 38684 234028 38690
rect 233976 38626 234028 38632
rect 233884 15088 233936 15094
rect 233884 15030 233936 15036
rect 233988 13802 234016 38626
rect 234632 38350 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700738 267688 703520
rect 267648 700732 267700 700738
rect 267648 700674 267700 700680
rect 300136 700534 300164 703520
rect 332520 700670 332548 703520
rect 332508 700664 332560 700670
rect 332508 700606 332560 700612
rect 364996 700602 365024 703520
rect 364984 700596 365036 700602
rect 364984 700538 365036 700544
rect 397472 700534 397500 703520
rect 300124 700528 300176 700534
rect 300124 700470 300176 700476
rect 378784 700528 378836 700534
rect 378784 700470 378836 700476
rect 397460 700528 397512 700534
rect 397460 700470 397512 700476
rect 268016 687404 268068 687410
rect 268016 687346 268068 687352
rect 289084 687404 289136 687410
rect 289084 687346 289136 687352
rect 261484 687336 261536 687342
rect 261484 687278 261536 687284
rect 250352 687268 250404 687274
rect 250352 687210 250404 687216
rect 250364 684964 250392 687210
rect 260378 684584 260434 684593
rect 260434 684542 260682 684570
rect 260378 684519 260434 684528
rect 238864 684270 240074 684298
rect 234710 674248 234766 674257
rect 234710 674183 234766 674192
rect 238666 674248 238722 674257
rect 238666 674183 238722 674192
rect 234724 665961 234752 674183
rect 238680 665961 238708 674183
rect 234710 665952 234766 665961
rect 234710 665887 234766 665896
rect 238666 665952 238722 665961
rect 238666 665887 238722 665896
rect 238864 662386 238892 684270
rect 261496 673454 261524 687278
rect 268028 684964 268056 687346
rect 278320 687336 278372 687342
rect 278320 687278 278372 687284
rect 278332 684964 278360 687278
rect 288992 687268 289044 687274
rect 288992 687210 289044 687216
rect 288650 684270 288848 684298
rect 288820 683194 288848 684270
rect 288808 683188 288860 683194
rect 288808 683130 288860 683136
rect 288900 682984 288952 682990
rect 288900 682926 288952 682932
rect 288808 681080 288860 681086
rect 288808 681022 288860 681028
rect 262218 674248 262274 674257
rect 262218 674183 262274 674192
rect 266266 674248 266322 674257
rect 266266 674183 266322 674192
rect 261128 673426 261524 673454
rect 261128 664714 261156 673426
rect 262232 665174 262260 674183
rect 266280 665174 266308 674183
rect 262220 665168 262272 665174
rect 262220 665110 262272 665116
rect 266268 665168 266320 665174
rect 266268 665110 266320 665116
rect 288820 664714 288848 681022
rect 260682 664686 261156 664714
rect 288650 664686 288848 664714
rect 239784 664006 240074 664034
rect 250378 664006 250760 664034
rect 238852 662380 238904 662386
rect 238852 662322 238904 662328
rect 239784 662318 239812 664006
rect 239772 662312 239824 662318
rect 239772 662254 239824 662260
rect 250732 662250 250760 664006
rect 268028 662318 268056 664020
rect 278332 662318 278360 664020
rect 268016 662312 268068 662318
rect 268016 662254 268068 662260
rect 278320 662312 278372 662318
rect 278320 662254 278372 662260
rect 288912 662250 288940 682926
rect 289004 681086 289032 687210
rect 288992 681080 289044 681086
rect 288992 681022 289044 681028
rect 289096 667418 289124 687346
rect 317144 687336 317196 687342
rect 317144 687278 317196 687284
rect 334348 687336 334400 687342
rect 334348 687278 334400 687284
rect 372988 687336 373040 687342
rect 372988 687278 373040 687284
rect 306012 687268 306064 687274
rect 306012 687210 306064 687216
rect 317052 687268 317104 687274
rect 317052 687210 317104 687216
rect 306024 684978 306052 687210
rect 306024 684950 306360 684978
rect 316664 684542 317000 684570
rect 295444 684270 296056 684298
rect 316868 684276 316920 684282
rect 291198 674248 291254 674257
rect 291198 674183 291254 674192
rect 293866 674248 293922 674257
rect 293866 674183 293922 674192
rect 289084 667412 289136 667418
rect 289084 667354 289136 667360
rect 291212 665961 291240 674183
rect 293880 665961 293908 674183
rect 291198 665952 291254 665961
rect 291198 665887 291254 665896
rect 293866 665952 293922 665961
rect 293866 665887 293922 665896
rect 295444 662386 295472 684270
rect 316868 684218 316920 684224
rect 316776 684208 316828 684214
rect 316776 684150 316828 684156
rect 295708 667412 295760 667418
rect 295708 667354 295760 667360
rect 295720 664714 295748 667354
rect 316788 664714 316816 684150
rect 295720 664686 296056 664714
rect 316664 664686 316816 664714
rect 306300 664006 306360 664034
rect 295432 662380 295484 662386
rect 295432 662322 295484 662328
rect 306300 662250 306328 664006
rect 316880 662250 316908 684218
rect 316972 662318 317000 684542
rect 317064 684282 317092 687210
rect 317052 684276 317104 684282
rect 317052 684218 317104 684224
rect 317156 684214 317184 687278
rect 334360 684964 334388 687278
rect 344652 687268 344704 687274
rect 344652 687210 344704 687216
rect 352012 687268 352064 687274
rect 352012 687210 352064 687216
rect 344664 684964 344692 687210
rect 352024 684964 352052 687210
rect 361946 684584 362002 684593
rect 362002 684542 362342 684570
rect 372646 684542 372936 684570
rect 361946 684519 362002 684528
rect 323044 684270 324070 684298
rect 372804 684276 372856 684282
rect 317144 684208 317196 684214
rect 317144 684150 317196 684156
rect 318798 674248 318854 674257
rect 318798 674183 318854 674192
rect 322846 674248 322902 674257
rect 322846 674183 322902 674192
rect 318812 665174 318840 674183
rect 322860 665174 322888 674183
rect 318800 665168 318852 665174
rect 318800 665110 318852 665116
rect 322848 665168 322900 665174
rect 322848 665110 322900 665116
rect 323044 662318 323072 684270
rect 372804 684218 372856 684224
rect 346398 674248 346454 674257
rect 346398 674183 346454 674192
rect 350446 674248 350502 674257
rect 350446 674183 350502 674192
rect 346412 665961 346440 674183
rect 350460 665961 350488 674183
rect 346398 665952 346454 665961
rect 346398 665887 346454 665896
rect 350446 665952 350502 665961
rect 350446 665887 350502 665896
rect 372816 664714 372844 684218
rect 372646 664686 372844 664714
rect 323688 664006 324070 664034
rect 334374 664006 334664 664034
rect 344678 664006 344968 664034
rect 323688 662386 323716 664006
rect 334636 662386 334664 664006
rect 344940 662425 344968 664006
rect 344926 662416 344982 662425
rect 323676 662380 323728 662386
rect 323676 662322 323728 662328
rect 334624 662380 334676 662386
rect 344926 662351 344982 662360
rect 334624 662322 334676 662328
rect 352024 662318 352052 664020
rect 362328 662318 362356 664020
rect 372908 662386 372936 684542
rect 373000 684282 373028 687278
rect 373264 687268 373316 687274
rect 373264 687210 373316 687216
rect 372988 684276 373040 684282
rect 372988 684218 373040 684224
rect 373276 667214 373304 687210
rect 375378 674248 375434 674257
rect 375378 674183 375434 674192
rect 378046 674248 378102 674257
rect 378046 674183 378102 674192
rect 373264 667208 373316 667214
rect 373264 667150 373316 667156
rect 375392 665174 375420 674183
rect 378060 665174 378088 674183
rect 375380 665168 375432 665174
rect 375380 665110 375432 665116
rect 378048 665168 378100 665174
rect 378048 665110 378100 665116
rect 372896 662380 372948 662386
rect 372896 662322 372948 662328
rect 316960 662312 317012 662318
rect 316960 662254 317012 662260
rect 323032 662312 323084 662318
rect 323032 662254 323084 662260
rect 352012 662312 352064 662318
rect 352012 662254 352064 662260
rect 362316 662312 362368 662318
rect 362316 662254 362368 662260
rect 250720 662244 250772 662250
rect 250720 662186 250772 662192
rect 288900 662244 288952 662250
rect 288900 662186 288952 662192
rect 306288 662244 306340 662250
rect 306288 662186 306340 662192
rect 316868 662244 316920 662250
rect 316868 662186 316920 662192
rect 250628 659796 250680 659802
rect 250628 659738 250680 659744
rect 295432 659796 295484 659802
rect 295432 659738 295484 659744
rect 334624 659796 334676 659802
rect 334624 659738 334676 659744
rect 240324 659728 240376 659734
rect 240324 659670 240376 659676
rect 240336 657900 240364 659670
rect 250640 657900 250668 659738
rect 267832 659728 267884 659734
rect 267832 659670 267884 659676
rect 260958 657206 261064 657234
rect 234710 656024 234766 656033
rect 234710 655959 234766 655968
rect 238666 656024 238722 656033
rect 238666 655959 238722 655968
rect 234724 647737 234752 655959
rect 238680 647737 238708 655959
rect 234710 647728 234766 647737
rect 234710 647663 234766 647672
rect 238666 647728 238722 647737
rect 238666 647663 238722 647672
rect 240336 634817 240364 637092
rect 240322 634808 240378 634817
rect 240322 634743 240378 634752
rect 250640 634710 250668 637092
rect 260944 634778 260972 637092
rect 261036 634778 261064 657206
rect 262220 656940 262272 656946
rect 262220 656882 262272 656888
rect 266268 656940 266320 656946
rect 266268 656882 266320 656888
rect 262232 647737 262260 656882
rect 266280 647737 266308 656882
rect 267740 655716 267792 655722
rect 267740 655658 267792 655664
rect 262218 647728 262274 647737
rect 262218 647663 262274 647672
rect 266266 647728 266322 647737
rect 266266 647663 266322 647672
rect 260932 634772 260984 634778
rect 260932 634714 260984 634720
rect 261024 634772 261076 634778
rect 261024 634714 261076 634720
rect 267752 634710 267780 655658
rect 267844 637786 267872 659670
rect 278226 657384 278282 657393
rect 278282 657342 278622 657370
rect 278226 657319 278282 657328
rect 267936 657206 268318 657234
rect 288926 657206 289124 657234
rect 267936 655722 267964 657206
rect 267924 655716 267976 655722
rect 267924 655658 267976 655664
rect 267844 637758 268318 637786
rect 278608 634710 278636 637092
rect 288912 634778 288940 637092
rect 289096 634778 289124 657206
rect 291198 656024 291254 656033
rect 291198 655959 291254 655968
rect 293866 656024 293922 656033
rect 293866 655959 293922 655968
rect 291212 647737 291240 655959
rect 293880 647737 293908 655959
rect 295340 655716 295392 655722
rect 295340 655658 295392 655664
rect 291198 647728 291254 647737
rect 291198 647663 291254 647672
rect 293866 647728 293922 647737
rect 293866 647663 293922 647672
rect 288900 634772 288952 634778
rect 288900 634714 288952 634720
rect 289084 634772 289136 634778
rect 289084 634714 289136 634720
rect 295352 634710 295380 655658
rect 295444 654134 295472 659738
rect 306472 659728 306524 659734
rect 306472 659670 306524 659676
rect 318064 659728 318116 659734
rect 318064 659670 318116 659676
rect 324320 659728 324372 659734
rect 324320 659670 324372 659676
rect 306484 657914 306512 659670
rect 306484 657886 306636 657914
rect 295996 657206 296332 657234
rect 316940 657206 317092 657234
rect 295996 655722 296024 657206
rect 295984 655716 296036 655722
rect 295984 655658 296036 655664
rect 295444 654106 295932 654134
rect 295904 637786 295932 654106
rect 295904 637758 296332 637786
rect 306636 637078 306972 637106
rect 306944 634710 306972 637078
rect 316604 637078 316940 637106
rect 316604 634778 316632 637078
rect 317064 634778 317092 657206
rect 316592 634772 316644 634778
rect 316592 634714 316644 634720
rect 317052 634772 317104 634778
rect 317052 634714 317104 634720
rect 318076 634710 318104 659670
rect 324332 657900 324360 659670
rect 334636 657900 334664 659738
rect 345756 659728 345808 659734
rect 345756 659670 345808 659676
rect 362316 659728 362368 659734
rect 362316 659670 362368 659676
rect 344954 657206 345152 657234
rect 318800 656940 318852 656946
rect 318800 656882 318852 656888
rect 322848 656940 322900 656946
rect 322848 656882 322900 656888
rect 318812 647737 318840 656882
rect 322860 647737 322888 656882
rect 345124 654134 345152 657206
rect 345124 654106 345704 654134
rect 318798 647728 318854 647737
rect 318798 647663 318854 647672
rect 322846 647728 322902 647737
rect 322846 647663 322902 647672
rect 324332 634710 324360 637092
rect 250628 634704 250680 634710
rect 250628 634646 250680 634652
rect 267740 634704 267792 634710
rect 267740 634646 267792 634652
rect 278596 634704 278648 634710
rect 278596 634646 278648 634652
rect 295340 634704 295392 634710
rect 295340 634646 295392 634652
rect 306932 634704 306984 634710
rect 306932 634646 306984 634652
rect 318064 634704 318116 634710
rect 318064 634646 318116 634652
rect 324320 634704 324372 634710
rect 324320 634646 324372 634652
rect 334636 634642 334664 637092
rect 344940 634778 344968 637092
rect 345676 634778 345704 654106
rect 344928 634772 344980 634778
rect 344928 634714 344980 634720
rect 345664 634772 345716 634778
rect 345664 634714 345716 634720
rect 345768 634710 345796 659670
rect 362328 657914 362356 659670
rect 362328 657886 362664 657914
rect 351932 657206 352360 657234
rect 372968 657206 373120 657234
rect 346398 656024 346454 656033
rect 346398 655959 346454 655968
rect 350446 656024 350502 656033
rect 350446 655959 350502 655968
rect 346412 647737 346440 655959
rect 350460 647737 350488 655959
rect 346398 647728 346454 647737
rect 346398 647663 346454 647672
rect 350446 647728 350502 647737
rect 350446 647663 350502 647672
rect 345756 634704 345808 634710
rect 345756 634646 345808 634652
rect 351932 634642 351960 657206
rect 352360 637078 352696 637106
rect 362664 637078 362908 637106
rect 352668 634817 352696 637078
rect 352654 634808 352710 634817
rect 352654 634743 352710 634752
rect 362880 634710 362908 637078
rect 372632 637078 372968 637106
rect 372632 634778 372660 637078
rect 373092 634778 373120 657206
rect 375380 656940 375432 656946
rect 375380 656882 375432 656888
rect 378048 656940 378100 656946
rect 378048 656882 378100 656888
rect 375392 647737 375420 656882
rect 378060 647737 378088 656882
rect 375378 647728 375434 647737
rect 375378 647663 375434 647672
rect 378046 647728 378102 647737
rect 378046 647663 378102 647672
rect 372620 634772 372672 634778
rect 372620 634714 372672 634720
rect 373080 634772 373132 634778
rect 373080 634714 373132 634720
rect 362868 634704 362920 634710
rect 362868 634646 362920 634652
rect 334624 634636 334676 634642
rect 334624 634578 334676 634584
rect 351920 634636 351972 634642
rect 351920 634578 351972 634584
rect 268016 632256 268068 632262
rect 268016 632198 268068 632204
rect 289084 632256 289136 632262
rect 289084 632198 289136 632204
rect 261484 632188 261536 632194
rect 261484 632130 261536 632136
rect 250352 632120 250404 632126
rect 250352 632062 250404 632068
rect 250364 630972 250392 632062
rect 260378 630456 260434 630465
rect 260434 630414 260682 630442
rect 260378 630391 260434 630400
rect 238864 630278 240074 630306
rect 234710 620256 234766 620265
rect 234710 620191 234766 620200
rect 238666 620256 238722 620265
rect 238666 620191 238722 620200
rect 234724 611969 234752 620191
rect 238680 611969 238708 620191
rect 234710 611960 234766 611969
rect 234710 611895 234766 611904
rect 238666 611960 238722 611969
rect 238666 611895 238722 611904
rect 238864 608598 238892 630278
rect 261496 615494 261524 632130
rect 268028 630972 268056 632198
rect 278320 632188 278372 632194
rect 278320 632130 278372 632136
rect 278332 630972 278360 632130
rect 288900 632120 288952 632126
rect 288900 632062 288952 632068
rect 288650 630278 288848 630306
rect 262218 620256 262274 620265
rect 262218 620191 262274 620200
rect 266266 620256 266322 620265
rect 266266 620191 266322 620200
rect 261128 615466 261524 615494
rect 261128 610722 261156 615466
rect 262232 611318 262260 620191
rect 266280 611318 266308 620191
rect 262220 611312 262272 611318
rect 262220 611254 262272 611260
rect 266268 611312 266320 611318
rect 266268 611254 266320 611260
rect 288820 610842 288848 630278
rect 288808 610836 288860 610842
rect 288808 610778 288860 610784
rect 260682 610694 261156 610722
rect 288912 610450 288940 632062
rect 289096 612814 289124 632198
rect 317144 632188 317196 632194
rect 317144 632130 317196 632136
rect 334348 632188 334400 632194
rect 334348 632130 334400 632136
rect 372988 632188 373040 632194
rect 372988 632130 373040 632136
rect 306012 632120 306064 632126
rect 306012 632062 306064 632068
rect 317052 632120 317104 632126
rect 317052 632062 317104 632068
rect 306024 630986 306052 632062
rect 306024 630958 306360 630986
rect 316664 630550 317000 630578
rect 295444 630278 296056 630306
rect 291198 620256 291254 620265
rect 291198 620191 291254 620200
rect 293866 620256 293922 620265
rect 293866 620191 293922 620200
rect 289084 612808 289136 612814
rect 289084 612750 289136 612756
rect 291212 611969 291240 620191
rect 293880 611969 293908 620191
rect 291198 611960 291254 611969
rect 291198 611895 291254 611904
rect 293866 611960 293922 611969
rect 293866 611895 293922 611904
rect 288992 610836 289044 610842
rect 288992 610778 289044 610784
rect 288650 610422 288940 610450
rect 238852 608592 238904 608598
rect 238852 608534 238904 608540
rect 240060 608530 240088 610028
rect 240048 608524 240100 608530
rect 240048 608466 240100 608472
rect 250364 608462 250392 610028
rect 268028 608530 268056 610028
rect 278332 608530 278360 610028
rect 268016 608524 268068 608530
rect 268016 608466 268068 608472
rect 278320 608524 278372 608530
rect 278320 608466 278372 608472
rect 289004 608462 289032 610778
rect 295444 608598 295472 630278
rect 316776 628720 316828 628726
rect 316776 628662 316828 628668
rect 295708 612808 295760 612814
rect 295708 612750 295760 612756
rect 295720 610722 295748 612750
rect 316788 610722 316816 628662
rect 316868 628652 316920 628658
rect 316868 628594 316920 628600
rect 295720 610694 296056 610722
rect 316664 610694 316816 610722
rect 306300 610014 306360 610042
rect 295432 608592 295484 608598
rect 295432 608534 295484 608540
rect 306300 608462 306328 610014
rect 316880 608462 316908 628594
rect 316972 608530 317000 630550
rect 317064 628658 317092 632062
rect 317156 628726 317184 632130
rect 334360 630972 334388 632130
rect 344652 632120 344704 632126
rect 344652 632062 344704 632068
rect 352012 632120 352064 632126
rect 352012 632062 352064 632068
rect 344664 630972 344692 632062
rect 352024 630972 352052 632062
rect 372646 630550 372936 630578
rect 361946 630456 362002 630465
rect 362002 630414 362342 630442
rect 361946 630391 362002 630400
rect 323044 630278 324070 630306
rect 317144 628720 317196 628726
rect 317144 628662 317196 628668
rect 317052 628652 317104 628658
rect 317052 628594 317104 628600
rect 318798 620256 318854 620265
rect 318798 620191 318854 620200
rect 322846 620256 322902 620265
rect 322846 620191 322902 620200
rect 318812 611318 318840 620191
rect 322860 611318 322888 620191
rect 318800 611312 318852 611318
rect 318800 611254 318852 611260
rect 322848 611312 322900 611318
rect 322848 611254 322900 611260
rect 323044 608530 323072 630278
rect 372804 628652 372856 628658
rect 372804 628594 372856 628600
rect 346398 620256 346454 620265
rect 346398 620191 346454 620200
rect 350446 620256 350502 620265
rect 350446 620191 350502 620200
rect 346412 611969 346440 620191
rect 350460 611969 350488 620191
rect 346398 611960 346454 611969
rect 346398 611895 346454 611904
rect 350446 611960 350502 611969
rect 350446 611895 350502 611904
rect 372816 610722 372844 628594
rect 372646 610694 372844 610722
rect 324056 608598 324084 610028
rect 334360 608598 334388 610028
rect 324044 608592 324096 608598
rect 324044 608534 324096 608540
rect 334348 608592 334400 608598
rect 344664 608569 344692 610028
rect 334348 608534 334400 608540
rect 344650 608560 344706 608569
rect 316960 608524 317012 608530
rect 316960 608466 317012 608472
rect 323032 608524 323084 608530
rect 352024 608530 352052 610028
rect 362328 608530 362356 610028
rect 372908 608598 372936 630550
rect 373000 628658 373028 632130
rect 373264 632120 373316 632126
rect 373264 632062 373316 632068
rect 372988 628652 373040 628658
rect 372988 628594 373040 628600
rect 373276 613426 373304 632062
rect 375378 620256 375434 620265
rect 375378 620191 375434 620200
rect 378046 620256 378102 620265
rect 378046 620191 378102 620200
rect 373264 613420 373316 613426
rect 373264 613362 373316 613368
rect 375392 611318 375420 620191
rect 378060 611318 378088 620191
rect 375380 611312 375432 611318
rect 375380 611254 375432 611260
rect 378048 611312 378100 611318
rect 378048 611254 378100 611260
rect 372896 608592 372948 608598
rect 372896 608534 372948 608540
rect 344650 608495 344706 608504
rect 352012 608524 352064 608530
rect 323032 608466 323084 608472
rect 352012 608466 352064 608472
rect 362316 608524 362368 608530
rect 362316 608466 362368 608472
rect 250352 608456 250404 608462
rect 250352 608398 250404 608404
rect 288992 608456 289044 608462
rect 288992 608398 289044 608404
rect 306288 608456 306340 608462
rect 306288 608398 306340 608404
rect 316868 608456 316920 608462
rect 316868 608398 316920 608404
rect 250628 605940 250680 605946
rect 250628 605882 250680 605888
rect 267832 605940 267884 605946
rect 267832 605882 267884 605888
rect 306380 605940 306432 605946
rect 306380 605882 306432 605888
rect 318064 605940 318116 605946
rect 318064 605882 318116 605888
rect 324320 605940 324372 605946
rect 324320 605882 324372 605888
rect 345756 605940 345808 605946
rect 345756 605882 345808 605888
rect 362316 605940 362368 605946
rect 362316 605882 362368 605888
rect 240324 605872 240376 605878
rect 240324 605814 240376 605820
rect 240336 603908 240364 605814
rect 250640 603908 250668 605882
rect 261484 605872 261536 605878
rect 261484 605814 261536 605820
rect 260958 603214 261064 603242
rect 238666 602304 238722 602313
rect 238666 602239 238722 602248
rect 234710 602032 234766 602041
rect 234710 601967 234766 601976
rect 234724 593745 234752 601967
rect 238680 593745 238708 602239
rect 234710 593736 234766 593745
rect 234710 593671 234766 593680
rect 238666 593736 238722 593745
rect 238666 593671 238722 593680
rect 240336 580922 240364 583100
rect 240324 580916 240376 580922
rect 240324 580858 240376 580864
rect 250640 580854 250668 583100
rect 260944 580990 260972 583100
rect 261036 580990 261064 603214
rect 260932 580984 260984 580990
rect 260932 580926 260984 580932
rect 261024 580984 261076 580990
rect 261024 580926 261076 580932
rect 261496 580922 261524 605814
rect 266266 602032 266322 602041
rect 266266 601967 266322 601976
rect 266280 593745 266308 601967
rect 267740 599752 267792 599758
rect 267740 599694 267792 599700
rect 266266 593736 266322 593745
rect 266266 593671 266322 593680
rect 261484 580916 261536 580922
rect 261484 580858 261536 580864
rect 267752 580854 267780 599694
rect 267844 583794 267872 605882
rect 278596 605872 278648 605878
rect 278596 605814 278648 605820
rect 295340 605872 295392 605878
rect 295340 605814 295392 605820
rect 278608 603908 278636 605814
rect 267936 603214 268318 603242
rect 288926 603214 289124 603242
rect 267936 599758 267964 603214
rect 267924 599752 267976 599758
rect 267924 599694 267976 599700
rect 267844 583766 268318 583794
rect 278608 580922 278636 583100
rect 288912 580990 288940 583100
rect 289096 580990 289124 603214
rect 293866 602168 293922 602177
rect 293866 602103 293922 602112
rect 293880 593745 293908 602103
rect 293866 593736 293922 593745
rect 293866 593671 293922 593680
rect 289728 585200 289780 585206
rect 289728 585142 289780 585148
rect 288900 580984 288952 580990
rect 288900 580926 288952 580932
rect 289084 580984 289136 580990
rect 289084 580926 289136 580932
rect 289740 580922 289768 585142
rect 295352 583930 295380 605814
rect 306392 603922 306420 605882
rect 306392 603894 306636 603922
rect 295444 603214 296332 603242
rect 316940 603214 317092 603242
rect 295444 585206 295472 603214
rect 295432 585200 295484 585206
rect 295432 585142 295484 585148
rect 295352 583902 295932 583930
rect 295904 583794 295932 583902
rect 295904 583766 296332 583794
rect 306636 583086 306972 583114
rect 306944 580922 306972 583086
rect 316604 583086 316940 583114
rect 316604 580990 316632 583086
rect 317064 580990 317092 603214
rect 316592 580984 316644 580990
rect 316592 580926 316644 580932
rect 317052 580984 317104 580990
rect 317052 580926 317104 580932
rect 318076 580922 318104 605882
rect 324332 603908 324360 605882
rect 334624 605872 334676 605878
rect 334624 605814 334676 605820
rect 345664 605872 345716 605878
rect 345664 605814 345716 605820
rect 334636 603908 334664 605814
rect 345020 603288 345072 603294
rect 344954 603236 345020 603242
rect 344954 603230 345072 603236
rect 344954 603214 345060 603230
rect 318798 602032 318854 602041
rect 318798 601967 318854 601976
rect 322846 602032 322902 602041
rect 322846 601967 322902 601976
rect 318812 593745 318840 601967
rect 322860 593745 322888 601967
rect 318798 593736 318854 593745
rect 318798 593671 318854 593680
rect 322846 593736 322902 593745
rect 322846 593671 322902 593680
rect 324332 580922 324360 583100
rect 278596 580916 278648 580922
rect 278596 580858 278648 580864
rect 289728 580916 289780 580922
rect 289728 580858 289780 580864
rect 306932 580916 306984 580922
rect 306932 580858 306984 580864
rect 318064 580916 318116 580922
rect 318064 580858 318116 580864
rect 324320 580916 324372 580922
rect 324320 580858 324372 580864
rect 334636 580854 334664 583100
rect 344940 580990 344968 583100
rect 344928 580984 344980 580990
rect 344928 580926 344980 580932
rect 345676 580854 345704 605814
rect 345768 580922 345796 605882
rect 352012 605872 352064 605878
rect 352012 605814 352064 605820
rect 352024 603922 352052 605814
rect 362328 603922 362356 605882
rect 352024 603894 352360 603922
rect 362328 603894 362664 603922
rect 345848 603288 345900 603294
rect 345848 603230 345900 603236
rect 345860 580990 345888 603230
rect 372968 603214 373120 603242
rect 350446 602168 350502 602177
rect 350446 602103 350502 602112
rect 350460 593745 350488 602103
rect 350446 593736 350502 593745
rect 350446 593671 350502 593680
rect 352360 583086 352696 583114
rect 362664 583086 362908 583114
rect 345848 580984 345900 580990
rect 352668 580961 352696 583086
rect 345848 580926 345900 580932
rect 352654 580952 352710 580961
rect 345756 580916 345808 580922
rect 362880 580922 362908 583086
rect 372632 583086 372968 583114
rect 372632 580990 372660 583086
rect 373092 580990 373120 603214
rect 378046 602032 378102 602041
rect 378046 601967 378102 601976
rect 378060 593745 378088 601967
rect 378046 593736 378102 593745
rect 378046 593671 378102 593680
rect 373172 585812 373224 585818
rect 373172 585754 373224 585760
rect 372620 580984 372672 580990
rect 372620 580926 372672 580932
rect 373080 580984 373132 580990
rect 373080 580926 373132 580932
rect 373184 580922 373212 585754
rect 352654 580887 352710 580896
rect 362868 580916 362920 580922
rect 345756 580858 345808 580864
rect 362868 580858 362920 580864
rect 373172 580916 373224 580922
rect 373172 580858 373224 580864
rect 250628 580848 250680 580854
rect 250628 580790 250680 580796
rect 267740 580848 267792 580854
rect 267740 580790 267792 580796
rect 334624 580848 334676 580854
rect 334624 580790 334676 580796
rect 345664 580848 345716 580854
rect 345664 580790 345716 580796
rect 261484 578332 261536 578338
rect 261484 578274 261536 578280
rect 278320 578332 278372 578338
rect 278320 578274 278372 578280
rect 288900 578332 288952 578338
rect 288900 578274 288952 578280
rect 306012 578332 306064 578338
rect 306012 578274 306064 578280
rect 316776 578332 316828 578338
rect 316776 578274 316828 578280
rect 333980 578332 334032 578338
rect 333980 578274 334032 578280
rect 372896 578332 372948 578338
rect 372896 578274 372948 578280
rect 250076 578264 250128 578270
rect 250076 578206 250128 578212
rect 250088 576994 250116 578206
rect 250088 576966 250378 576994
rect 260378 576464 260434 576473
rect 260434 576422 260682 576450
rect 260378 576399 260434 576408
rect 238864 576286 240074 576314
rect 234710 574696 234766 574705
rect 234710 574631 234766 574640
rect 238666 574696 238722 574705
rect 238666 574631 238722 574640
rect 234724 566273 234752 574631
rect 238680 566273 238708 574631
rect 234710 566264 234766 566273
rect 234710 566199 234766 566208
rect 238666 566264 238722 566273
rect 238666 566199 238722 566208
rect 238864 554742 238892 576286
rect 261496 557534 261524 578274
rect 268016 578264 268068 578270
rect 268016 578206 268068 578212
rect 268028 576980 268056 578206
rect 278332 576980 278360 578274
rect 288650 576286 288848 576314
rect 262218 566264 262274 566273
rect 262218 566199 262274 566208
rect 266266 566264 266322 566273
rect 266266 566199 266322 566208
rect 261128 557506 261524 557534
rect 262232 557530 262260 566199
rect 266280 557530 266308 566199
rect 262220 557524 262272 557530
rect 261128 556730 261156 557506
rect 262220 557466 262272 557472
rect 266268 557524 266320 557530
rect 266268 557466 266320 557472
rect 288820 556850 288848 576286
rect 288808 556844 288860 556850
rect 288808 556786 288860 556792
rect 260682 556702 261156 556730
rect 288912 556458 288940 578274
rect 289084 578264 289136 578270
rect 289084 578206 289136 578212
rect 289096 560250 289124 578206
rect 306024 576994 306052 578274
rect 306024 576966 306360 576994
rect 316788 576434 316816 578274
rect 316868 578264 316920 578270
rect 316868 578206 316920 578212
rect 316880 576434 316908 578206
rect 333992 576994 334020 578274
rect 344284 578264 344336 578270
rect 344284 578206 344336 578212
rect 352012 578264 352064 578270
rect 352012 578206 352064 578212
rect 344296 576994 344324 578206
rect 333992 576966 334374 576994
rect 344296 576966 344678 576994
rect 352024 576980 352052 578206
rect 361946 576464 362002 576473
rect 316776 576428 316828 576434
rect 316776 576370 316828 576376
rect 316868 576428 316920 576434
rect 362002 576422 362342 576450
rect 361946 576399 362002 576408
rect 316868 576370 316920 576376
rect 295444 576286 296056 576314
rect 316664 576286 317000 576314
rect 291198 574696 291254 574705
rect 291198 574631 291254 574640
rect 293866 574696 293922 574705
rect 293866 574631 293922 574640
rect 291212 566273 291240 574631
rect 293880 566273 293908 574631
rect 291198 566264 291254 566273
rect 291198 566199 291254 566208
rect 293866 566264 293922 566273
rect 293866 566199 293922 566208
rect 289084 560244 289136 560250
rect 289084 560186 289136 560192
rect 288992 556844 289044 556850
rect 288992 556786 289044 556792
rect 288650 556430 288940 556458
rect 238852 554736 238904 554742
rect 238852 554678 238904 554684
rect 240060 554674 240088 556036
rect 240048 554668 240100 554674
rect 240048 554610 240100 554616
rect 250364 554606 250392 556036
rect 268028 554674 268056 556036
rect 278332 554674 278360 556036
rect 268016 554668 268068 554674
rect 268016 554610 268068 554616
rect 278320 554668 278372 554674
rect 278320 554610 278372 554616
rect 289004 554606 289032 556786
rect 295444 554742 295472 576286
rect 316776 576224 316828 576230
rect 316776 576166 316828 576172
rect 316868 576224 316920 576230
rect 316868 576166 316920 576172
rect 295708 560244 295760 560250
rect 295708 560186 295760 560192
rect 295720 556730 295748 560186
rect 316788 556730 316816 576166
rect 295720 556702 296056 556730
rect 316664 556702 316816 556730
rect 306300 556022 306360 556050
rect 295432 554736 295484 554742
rect 295432 554678 295484 554684
rect 306300 554606 306328 556022
rect 316880 554606 316908 576166
rect 316972 554674 317000 576286
rect 323044 576286 324070 576314
rect 372646 576286 372844 576314
rect 318798 566264 318854 566273
rect 318798 566199 318854 566208
rect 322846 566264 322902 566273
rect 322846 566199 322902 566208
rect 318812 557530 318840 566199
rect 322860 557530 322888 566199
rect 318800 557524 318852 557530
rect 318800 557466 318852 557472
rect 322848 557524 322900 557530
rect 322848 557466 322900 557472
rect 323044 554674 323072 576286
rect 346398 574696 346454 574705
rect 346398 574631 346454 574640
rect 350446 574696 350502 574705
rect 350446 574631 350502 574640
rect 346412 566273 346440 574631
rect 350460 566273 350488 574631
rect 346398 566264 346454 566273
rect 346398 566199 346454 566208
rect 350446 566264 350502 566273
rect 350446 566199 350502 566208
rect 372816 556850 372844 576286
rect 372804 556844 372856 556850
rect 372804 556786 372856 556792
rect 372908 556458 372936 578274
rect 373264 578264 373316 578270
rect 373264 578206 373316 578212
rect 373276 559570 373304 578206
rect 375378 566264 375434 566273
rect 375378 566199 375434 566208
rect 378046 566264 378102 566273
rect 378046 566199 378102 566208
rect 373264 559564 373316 559570
rect 373264 559506 373316 559512
rect 375392 557530 375420 566199
rect 378060 557530 378088 566199
rect 375380 557524 375432 557530
rect 375380 557466 375432 557472
rect 378048 557524 378100 557530
rect 378048 557466 378100 557472
rect 372988 556844 373040 556850
rect 372988 556786 373040 556792
rect 372646 556430 372936 556458
rect 324056 554742 324084 556036
rect 334360 554742 334388 556036
rect 324044 554736 324096 554742
rect 324044 554678 324096 554684
rect 334348 554736 334400 554742
rect 344664 554713 344692 556036
rect 334348 554678 334400 554684
rect 344650 554704 344706 554713
rect 316960 554668 317012 554674
rect 316960 554610 317012 554616
rect 323032 554668 323084 554674
rect 352024 554674 352052 556036
rect 362328 554674 362356 556036
rect 373000 554742 373028 556786
rect 372988 554736 373040 554742
rect 372988 554678 373040 554684
rect 344650 554639 344706 554648
rect 352012 554668 352064 554674
rect 323032 554610 323084 554616
rect 352012 554610 352064 554616
rect 362316 554668 362368 554674
rect 362316 554610 362368 554616
rect 250352 554600 250404 554606
rect 250352 554542 250404 554548
rect 288992 554600 289044 554606
rect 288992 554542 289044 554548
rect 306288 554600 306340 554606
rect 306288 554542 306340 554548
rect 316868 554600 316920 554606
rect 316868 554542 316920 554548
rect 250628 552152 250680 552158
rect 250628 552094 250680 552100
rect 261484 552152 261536 552158
rect 261484 552094 261536 552100
rect 278596 552152 278648 552158
rect 278596 552094 278648 552100
rect 295340 552152 295392 552158
rect 295340 552094 295392 552100
rect 334624 552152 334676 552158
rect 334624 552094 334676 552100
rect 345756 552152 345808 552158
rect 345756 552094 345808 552100
rect 362316 552152 362368 552158
rect 362316 552094 362368 552100
rect 240140 550588 240192 550594
rect 240140 550530 240192 550536
rect 240152 549930 240180 550530
rect 240152 549902 240350 549930
rect 250640 549916 250668 552094
rect 260958 549222 261064 549250
rect 238666 548312 238722 548321
rect 238666 548247 238722 548256
rect 234710 548040 234766 548049
rect 234710 547975 234766 547984
rect 234724 539753 234752 547975
rect 238680 539753 238708 548247
rect 234710 539744 234766 539753
rect 234710 539679 234766 539688
rect 238666 539744 238722 539753
rect 238666 539679 238722 539688
rect 240336 527066 240364 529108
rect 240324 527060 240376 527066
rect 240324 527002 240376 527008
rect 250640 526998 250668 529108
rect 260944 527134 260972 529108
rect 261036 527134 261064 549222
rect 260932 527128 260984 527134
rect 260932 527070 260984 527076
rect 261024 527128 261076 527134
rect 261024 527070 261076 527076
rect 261496 527066 261524 552094
rect 267740 552084 267792 552090
rect 267740 552026 267792 552032
rect 262218 548176 262274 548185
rect 262218 548111 262274 548120
rect 262232 539753 262260 548111
rect 266266 548040 266322 548049
rect 266266 547975 266322 547984
rect 266280 539753 266308 547975
rect 262218 539744 262274 539753
rect 262218 539679 262274 539688
rect 266266 539744 266322 539753
rect 266266 539679 266322 539688
rect 267752 533662 267780 552026
rect 278608 549916 278636 552094
rect 267844 549222 268318 549250
rect 288926 549222 289124 549250
rect 267740 533656 267792 533662
rect 267740 533598 267792 533604
rect 267844 530482 267872 549222
rect 268016 533656 268068 533662
rect 268016 533598 268068 533604
rect 267752 530454 267872 530482
rect 267752 528554 267780 530454
rect 268028 529666 268056 533598
rect 268028 529638 268318 529666
rect 267752 528526 267872 528554
rect 261484 527060 261536 527066
rect 261484 527002 261536 527008
rect 267844 526998 267872 528526
rect 278608 527066 278636 529108
rect 288912 527134 288940 529108
rect 289096 527134 289124 549222
rect 295352 533662 295380 552094
rect 306472 552084 306524 552090
rect 306472 552026 306524 552032
rect 318064 552084 318116 552090
rect 318064 552026 318116 552032
rect 324320 552084 324372 552090
rect 324320 552026 324372 552032
rect 306484 549930 306512 552026
rect 306484 549902 306636 549930
rect 295444 549222 296332 549250
rect 316940 549222 317092 549250
rect 295340 533656 295392 533662
rect 295340 533598 295392 533604
rect 288900 527128 288952 527134
rect 288900 527070 288952 527076
rect 289084 527128 289136 527134
rect 289084 527070 289136 527076
rect 295444 527066 295472 549222
rect 295984 533656 296036 533662
rect 295984 533598 296036 533604
rect 295996 529666 296024 533598
rect 295996 529638 296332 529666
rect 306636 529094 306972 529122
rect 306944 527066 306972 529094
rect 316604 529094 316940 529122
rect 316604 527134 316632 529094
rect 317064 527134 317092 549222
rect 316592 527128 316644 527134
rect 316592 527070 316644 527076
rect 317052 527128 317104 527134
rect 317052 527070 317104 527076
rect 318076 527066 318104 552026
rect 324332 549916 324360 552026
rect 334636 549916 334664 552094
rect 344954 549222 345152 549250
rect 322846 548312 322902 548321
rect 322846 548247 322902 548256
rect 318798 548040 318854 548049
rect 318798 547975 318854 547984
rect 318812 539753 318840 547975
rect 322860 539753 322888 548247
rect 345124 547874 345152 549222
rect 345124 547846 345704 547874
rect 318798 539744 318854 539753
rect 318798 539679 318854 539688
rect 322846 539744 322902 539753
rect 322846 539679 322902 539688
rect 324332 527066 324360 529108
rect 278596 527060 278648 527066
rect 278596 527002 278648 527008
rect 295432 527060 295484 527066
rect 295432 527002 295484 527008
rect 306932 527060 306984 527066
rect 306932 527002 306984 527008
rect 318064 527060 318116 527066
rect 318064 527002 318116 527008
rect 324320 527060 324372 527066
rect 324320 527002 324372 527008
rect 334636 526998 334664 529108
rect 344940 527134 344968 529108
rect 345676 527134 345704 547846
rect 344928 527128 344980 527134
rect 344928 527070 344980 527076
rect 345664 527128 345716 527134
rect 345664 527070 345716 527076
rect 345768 527066 345796 552094
rect 345848 552084 345900 552090
rect 345848 552026 345900 552032
rect 352012 552084 352064 552090
rect 352012 552026 352064 552032
rect 345756 527060 345808 527066
rect 345756 527002 345808 527008
rect 345860 526998 345888 552026
rect 352024 549930 352052 552026
rect 362328 549930 362356 552094
rect 352024 549902 352360 549930
rect 362328 549902 362664 549930
rect 372968 549222 373120 549250
rect 346398 548176 346454 548185
rect 346398 548111 346454 548120
rect 346412 539753 346440 548111
rect 350446 548040 350502 548049
rect 350446 547975 350502 547984
rect 350460 539753 350488 547975
rect 346398 539744 346454 539753
rect 346398 539679 346454 539688
rect 350446 539744 350502 539753
rect 350446 539679 350502 539688
rect 352360 529094 352696 529122
rect 362664 529094 362908 529122
rect 352668 527105 352696 529094
rect 352654 527096 352710 527105
rect 362880 527066 362908 529094
rect 372632 529094 372968 529122
rect 372632 527134 372660 529094
rect 373092 527134 373120 549222
rect 378046 548176 378102 548185
rect 378046 548111 378102 548120
rect 378060 539753 378088 548111
rect 378046 539744 378102 539753
rect 378046 539679 378102 539688
rect 372620 527128 372672 527134
rect 372620 527070 372672 527076
rect 373080 527128 373132 527134
rect 373080 527070 373132 527076
rect 352654 527031 352710 527040
rect 362868 527060 362920 527066
rect 362868 527002 362920 527008
rect 250628 526992 250680 526998
rect 250628 526934 250680 526940
rect 267832 526992 267884 526998
rect 267832 526934 267884 526940
rect 334624 526992 334676 526998
rect 334624 526934 334676 526940
rect 345848 526992 345900 526998
rect 345848 526934 345900 526940
rect 261484 524544 261536 524550
rect 261484 524486 261536 524492
rect 278320 524544 278372 524550
rect 278320 524486 278372 524492
rect 288992 524544 289044 524550
rect 288992 524486 289044 524492
rect 306012 524544 306064 524550
rect 306012 524486 306064 524492
rect 317144 524544 317196 524550
rect 317144 524486 317196 524492
rect 334348 524544 334400 524550
rect 334348 524486 334400 524492
rect 372988 524544 373040 524550
rect 372988 524486 373040 524492
rect 250352 524476 250404 524482
rect 250352 524418 250404 524424
rect 250364 522852 250392 524418
rect 260378 522472 260434 522481
rect 260434 522430 260682 522458
rect 260378 522407 260434 522416
rect 238864 522294 240074 522322
rect 238666 520976 238722 520985
rect 238666 520911 238722 520920
rect 234710 520704 234766 520713
rect 234710 520639 234766 520648
rect 234724 512281 234752 520639
rect 238680 512281 238708 520911
rect 234710 512272 234766 512281
rect 234710 512207 234766 512216
rect 238666 512272 238722 512281
rect 238666 512207 238722 512216
rect 238864 500954 238892 522294
rect 261496 509234 261524 524486
rect 268016 524476 268068 524482
rect 268016 524418 268068 524424
rect 268028 522852 268056 524418
rect 278332 522852 278360 524486
rect 288650 522430 288940 522458
rect 262218 520840 262274 520849
rect 262218 520775 262274 520784
rect 262232 512281 262260 520775
rect 266266 520704 266322 520713
rect 266266 520639 266322 520648
rect 266280 512281 266308 520639
rect 288912 519722 288940 522430
rect 288900 519716 288952 519722
rect 288900 519658 288952 519664
rect 289004 519602 289032 524486
rect 289084 524476 289136 524482
rect 289084 524418 289136 524424
rect 288820 519574 289032 519602
rect 262218 512272 262274 512281
rect 262218 512207 262274 512216
rect 266266 512272 266322 512281
rect 266266 512207 266322 512216
rect 261128 509206 261524 509234
rect 261128 502738 261156 509206
rect 288820 502738 288848 519574
rect 288900 519512 288952 519518
rect 288900 519454 288952 519460
rect 260682 502710 261156 502738
rect 288650 502710 288848 502738
rect 238852 500948 238904 500954
rect 238852 500890 238904 500896
rect 240060 500886 240088 502044
rect 240048 500880 240100 500886
rect 240048 500822 240100 500828
rect 250364 500818 250392 502044
rect 268028 500886 268056 502044
rect 278332 500886 278360 502044
rect 268016 500880 268068 500886
rect 268016 500822 268068 500828
rect 278320 500880 278372 500886
rect 278320 500822 278372 500828
rect 288912 500818 288940 519454
rect 289096 505646 289124 524418
rect 306024 522866 306052 524486
rect 317052 524476 317104 524482
rect 317052 524418 317104 524424
rect 306024 522838 306360 522866
rect 316664 522566 317000 522594
rect 295444 522294 296056 522322
rect 289084 505640 289136 505646
rect 289084 505582 289136 505588
rect 295444 500954 295472 522294
rect 316776 521756 316828 521762
rect 316776 521698 316828 521704
rect 295708 505640 295760 505646
rect 295708 505582 295760 505588
rect 295720 502738 295748 505582
rect 316788 502738 316816 521698
rect 316868 521688 316920 521694
rect 316868 521630 316920 521636
rect 295720 502710 296056 502738
rect 316664 502710 316816 502738
rect 306300 502030 306360 502058
rect 295432 500948 295484 500954
rect 295432 500890 295484 500896
rect 306300 500818 306328 502030
rect 316880 500818 316908 521630
rect 316972 500886 317000 522566
rect 317064 521694 317092 524418
rect 317156 521762 317184 524486
rect 334360 522852 334388 524486
rect 344652 524476 344704 524482
rect 344652 524418 344704 524424
rect 352012 524476 352064 524482
rect 352012 524418 352064 524424
rect 344664 522852 344692 524418
rect 352024 522852 352052 524418
rect 372646 522566 372936 522594
rect 361946 522472 362002 522481
rect 362002 522430 362342 522458
rect 361946 522407 362002 522416
rect 323044 522294 324070 522322
rect 317144 521756 317196 521762
rect 317144 521698 317196 521704
rect 317052 521688 317104 521694
rect 317052 521630 317104 521636
rect 317050 520704 317106 520713
rect 317050 520639 317106 520648
rect 322846 520704 322902 520713
rect 322846 520639 322902 520648
rect 317064 512825 317092 520639
rect 317050 512816 317106 512825
rect 317050 512751 317106 512760
rect 322860 512281 322888 520639
rect 322846 512272 322902 512281
rect 322846 512207 322902 512216
rect 323044 500886 323072 522294
rect 372804 521756 372856 521762
rect 372804 521698 372856 521704
rect 346398 520840 346454 520849
rect 346398 520775 346454 520784
rect 350446 520840 350502 520849
rect 350446 520775 350502 520784
rect 346412 512281 346440 520775
rect 350460 512281 350488 520775
rect 346398 512272 346454 512281
rect 346398 512207 346454 512216
rect 350446 512272 350502 512281
rect 350446 512207 350502 512216
rect 372816 502738 372844 521698
rect 372646 502710 372844 502738
rect 324056 500954 324084 502044
rect 334360 500954 334388 502044
rect 324044 500948 324096 500954
rect 324044 500890 324096 500896
rect 334348 500948 334400 500954
rect 334348 500890 334400 500896
rect 316960 500880 317012 500886
rect 316960 500822 317012 500828
rect 323032 500880 323084 500886
rect 344664 500857 344692 502044
rect 352024 500886 352052 502044
rect 362328 500886 362356 502044
rect 372908 500954 372936 522566
rect 373000 521762 373028 524486
rect 373264 524476 373316 524482
rect 373264 524418 373316 524424
rect 372988 521756 373040 521762
rect 372988 521698 373040 521704
rect 373276 505782 373304 524418
rect 378046 520704 378102 520713
rect 378046 520639 378102 520648
rect 378060 512281 378088 520639
rect 378046 512272 378102 512281
rect 378046 512207 378102 512216
rect 373264 505776 373316 505782
rect 373264 505718 373316 505724
rect 372896 500948 372948 500954
rect 372896 500890 372948 500896
rect 352012 500880 352064 500886
rect 323032 500822 323084 500828
rect 344650 500848 344706 500857
rect 250352 500812 250404 500818
rect 250352 500754 250404 500760
rect 288900 500812 288952 500818
rect 288900 500754 288952 500760
rect 306288 500812 306340 500818
rect 306288 500754 306340 500760
rect 316868 500812 316920 500818
rect 352012 500822 352064 500828
rect 362316 500880 362368 500886
rect 362316 500822 362368 500828
rect 344650 500783 344706 500792
rect 316868 500754 316920 500760
rect 250628 498296 250680 498302
rect 250628 498238 250680 498244
rect 267740 498296 267792 498302
rect 267740 498238 267792 498244
rect 306472 498296 306524 498302
rect 306472 498238 306524 498244
rect 318064 498296 318116 498302
rect 318064 498238 318116 498244
rect 324320 498296 324372 498302
rect 324320 498238 324372 498244
rect 345848 498296 345900 498302
rect 345848 498238 345900 498244
rect 362316 498296 362368 498302
rect 362316 498238 362368 498244
rect 240324 498228 240376 498234
rect 240324 498170 240376 498176
rect 240336 495924 240364 498170
rect 250640 495924 250668 498238
rect 261484 498228 261536 498234
rect 261484 498170 261536 498176
rect 260958 495230 261064 495258
rect 234710 485752 234766 485761
rect 234710 485687 234766 485696
rect 238666 485752 238722 485761
rect 238666 485687 238722 485696
rect 234724 477329 234752 485687
rect 234710 477320 234766 477329
rect 234710 477255 234766 477264
rect 238680 477057 238708 485687
rect 238666 477048 238722 477057
rect 238666 476983 238722 476992
rect 240336 473278 240364 475116
rect 240324 473272 240376 473278
rect 240324 473214 240376 473220
rect 250640 473210 250668 475116
rect 260944 473346 260972 475116
rect 261036 473346 261064 495230
rect 260932 473340 260984 473346
rect 260932 473282 260984 473288
rect 261024 473340 261076 473346
rect 261024 473282 261076 473288
rect 261496 473278 261524 498170
rect 262218 485752 262274 485761
rect 262218 485687 262274 485696
rect 266266 485752 266322 485761
rect 266266 485687 266322 485696
rect 262232 477193 262260 485687
rect 266280 477329 266308 485687
rect 267752 477698 267780 498238
rect 278596 498228 278648 498234
rect 278596 498170 278648 498176
rect 295340 498228 295392 498234
rect 295340 498170 295392 498176
rect 278608 495924 278636 498170
rect 267844 495230 268318 495258
rect 288926 495230 289124 495258
rect 267844 480254 267872 495230
rect 267844 480226 267964 480254
rect 267740 477692 267792 477698
rect 267740 477634 267792 477640
rect 266266 477320 266322 477329
rect 266266 477255 266322 477264
rect 262218 477184 262274 477193
rect 262218 477119 262274 477128
rect 261484 473272 261536 473278
rect 261484 473214 261536 473220
rect 267936 473210 267964 480226
rect 268016 477692 268068 477698
rect 268016 477634 268068 477640
rect 268028 475674 268056 477634
rect 268028 475646 268318 475674
rect 278608 473278 278636 475116
rect 288912 473346 288940 475116
rect 289096 473346 289124 495230
rect 295352 477698 295380 498170
rect 306484 495938 306512 498238
rect 306484 495910 306636 495938
rect 295444 495230 296332 495258
rect 316940 495230 317092 495258
rect 295340 477692 295392 477698
rect 295340 477634 295392 477640
rect 288900 473340 288952 473346
rect 288900 473282 288952 473288
rect 289084 473340 289136 473346
rect 289084 473282 289136 473288
rect 295444 473278 295472 495230
rect 295984 477692 296036 477698
rect 295984 477634 296036 477640
rect 295996 475674 296024 477634
rect 295996 475646 296332 475674
rect 306636 475102 306972 475130
rect 306944 473278 306972 475102
rect 316604 475102 316940 475130
rect 316604 473346 316632 475102
rect 317064 473346 317092 495230
rect 316592 473340 316644 473346
rect 316592 473282 316644 473288
rect 317052 473340 317104 473346
rect 317052 473282 317104 473288
rect 318076 473278 318104 498238
rect 324332 495924 324360 498238
rect 334624 498228 334676 498234
rect 334624 498170 334676 498176
rect 345756 498228 345808 498234
rect 345756 498170 345808 498176
rect 334636 495924 334664 498170
rect 344954 495230 345152 495258
rect 345124 489914 345152 495230
rect 345124 489886 345704 489914
rect 318798 485752 318854 485761
rect 318798 485687 318854 485696
rect 322846 485752 322902 485761
rect 322846 485687 322902 485696
rect 318812 477329 318840 485687
rect 318798 477320 318854 477329
rect 318798 477255 318854 477264
rect 322860 477057 322888 485687
rect 322846 477048 322902 477057
rect 322846 476983 322902 476992
rect 324332 473278 324360 475116
rect 278596 473272 278648 473278
rect 278596 473214 278648 473220
rect 295432 473272 295484 473278
rect 295432 473214 295484 473220
rect 306932 473272 306984 473278
rect 306932 473214 306984 473220
rect 318064 473272 318116 473278
rect 318064 473214 318116 473220
rect 324320 473272 324372 473278
rect 324320 473214 324372 473220
rect 334636 473210 334664 475116
rect 344940 473346 344968 475116
rect 345676 473346 345704 489886
rect 344928 473340 344980 473346
rect 344928 473282 344980 473288
rect 345664 473340 345716 473346
rect 345664 473282 345716 473288
rect 345768 473210 345796 498170
rect 345860 473278 345888 498238
rect 352012 498228 352064 498234
rect 352012 498170 352064 498176
rect 352024 495938 352052 498170
rect 362328 495938 362356 498238
rect 352024 495910 352360 495938
rect 362328 495910 362664 495938
rect 372968 495230 373120 495258
rect 346398 485752 346454 485761
rect 346398 485687 346454 485696
rect 350446 485752 350502 485761
rect 350446 485687 350502 485696
rect 346412 477193 346440 485687
rect 350460 477329 350488 485687
rect 350446 477320 350502 477329
rect 350446 477255 350502 477264
rect 346398 477184 346454 477193
rect 346398 477119 346454 477128
rect 352360 475102 352696 475130
rect 362664 475102 362908 475130
rect 345848 473272 345900 473278
rect 352668 473249 352696 475102
rect 362880 473278 362908 475102
rect 372632 475102 372968 475130
rect 372632 473346 372660 475102
rect 373092 473346 373120 495230
rect 378046 485752 378102 485761
rect 378046 485687 378102 485696
rect 378060 477193 378088 485687
rect 378046 477184 378102 477193
rect 378046 477119 378102 477128
rect 372620 473340 372672 473346
rect 372620 473282 372672 473288
rect 373080 473340 373132 473346
rect 373080 473282 373132 473288
rect 362868 473272 362920 473278
rect 345848 473214 345900 473220
rect 352654 473240 352710 473249
rect 250628 473204 250680 473210
rect 250628 473146 250680 473152
rect 267924 473204 267976 473210
rect 267924 473146 267976 473152
rect 334624 473204 334676 473210
rect 334624 473146 334676 473152
rect 345756 473204 345808 473210
rect 362868 473214 362920 473220
rect 352654 473175 352710 473184
rect 345756 473146 345808 473152
rect 268016 470824 268068 470830
rect 268016 470766 268068 470772
rect 289084 470824 289136 470830
rect 289084 470766 289136 470772
rect 261576 470756 261628 470762
rect 261576 470698 261628 470704
rect 250352 470688 250404 470694
rect 250352 470630 250404 470636
rect 250364 468860 250392 470630
rect 260378 468480 260434 468489
rect 260434 468438 260682 468466
rect 260378 468415 260434 468424
rect 238864 468302 240074 468330
rect 234710 466712 234766 466721
rect 234710 466647 234766 466656
rect 234724 458289 234752 466647
rect 234710 458280 234766 458289
rect 234710 458215 234766 458224
rect 238864 445738 238892 468302
rect 261588 451274 261616 470698
rect 268028 468860 268056 470766
rect 278320 470756 278372 470762
rect 278320 470698 278372 470704
rect 278332 468860 278360 470698
rect 288900 470688 288952 470694
rect 288900 470630 288952 470636
rect 288650 468302 288848 468330
rect 262218 466984 262274 466993
rect 262218 466919 262274 466928
rect 262232 458289 262260 466919
rect 266266 466712 266322 466721
rect 266266 466647 266322 466656
rect 266280 458289 266308 466647
rect 262218 458280 262274 458289
rect 262218 458215 262274 458224
rect 266266 458280 266322 458289
rect 266266 458215 266322 458224
rect 261128 451246 261616 451274
rect 261128 448746 261156 451246
rect 288820 448866 288848 468302
rect 288808 448860 288860 448866
rect 288808 448802 288860 448808
rect 260682 448718 261156 448746
rect 288912 448474 288940 470630
rect 289096 452606 289124 470766
rect 372896 470756 372948 470762
rect 372896 470698 372948 470704
rect 306012 470688 306064 470694
rect 306012 470630 306064 470636
rect 316776 470688 316828 470694
rect 316776 470630 316828 470636
rect 334348 470688 334400 470694
rect 334348 470630 334400 470636
rect 352012 470688 352064 470694
rect 352012 470630 352064 470636
rect 306024 468874 306052 470630
rect 306024 468846 306360 468874
rect 316788 468450 316816 470630
rect 334360 468860 334388 470630
rect 352024 468860 352052 470630
rect 361946 468480 362002 468489
rect 316776 468444 316828 468450
rect 362002 468438 362342 468466
rect 361946 468415 362002 468424
rect 316776 468386 316828 468392
rect 295444 468302 296056 468330
rect 316664 468302 316908 468330
rect 291198 466848 291254 466857
rect 291198 466783 291254 466792
rect 291212 458289 291240 466783
rect 291198 458280 291254 458289
rect 291198 458215 291254 458224
rect 289084 452600 289136 452606
rect 289084 452542 289136 452548
rect 288992 448860 289044 448866
rect 288992 448802 289044 448808
rect 288650 448446 288940 448474
rect 238852 445732 238904 445738
rect 238852 445674 238904 445680
rect 240060 445670 240088 448052
rect 240048 445664 240100 445670
rect 240048 445606 240100 445612
rect 250364 445534 250392 448052
rect 268028 445670 268056 448052
rect 268016 445664 268068 445670
rect 268016 445606 268068 445612
rect 278332 445602 278360 448052
rect 278320 445596 278372 445602
rect 278320 445538 278372 445544
rect 289004 445534 289032 448802
rect 295444 445738 295472 468302
rect 316776 468240 316828 468246
rect 316776 468182 316828 468188
rect 295708 452600 295760 452606
rect 295708 452542 295760 452548
rect 295720 448746 295748 452542
rect 316788 448746 316816 468182
rect 295720 448718 296056 448746
rect 316664 448718 316816 448746
rect 306300 448038 306360 448066
rect 295432 445732 295484 445738
rect 295432 445674 295484 445680
rect 306300 445670 306328 448038
rect 306288 445664 306340 445670
rect 306288 445606 306340 445612
rect 316880 445602 316908 468302
rect 323044 468302 324070 468330
rect 344678 468302 344784 468330
rect 372646 468302 372844 468330
rect 318798 466712 318854 466721
rect 318798 466647 318854 466656
rect 318812 458289 318840 466647
rect 318798 458280 318854 458289
rect 318798 458215 318854 458224
rect 323044 445602 323072 468302
rect 324056 445738 324084 448052
rect 334360 445738 334388 448052
rect 324044 445732 324096 445738
rect 324044 445674 324096 445680
rect 334348 445732 334400 445738
rect 334348 445674 334400 445680
rect 344664 445641 344692 448052
rect 344756 445670 344784 468302
rect 346398 466848 346454 466857
rect 346398 466783 346454 466792
rect 350446 466848 350502 466857
rect 350446 466783 350502 466792
rect 346412 458289 346440 466783
rect 350460 458289 350488 466783
rect 346398 458280 346454 458289
rect 346398 458215 346454 458224
rect 350446 458280 350502 458289
rect 350446 458215 350502 458224
rect 372816 448866 372844 468302
rect 372804 448860 372856 448866
rect 372804 448802 372856 448808
rect 372908 448474 372936 470698
rect 373264 470688 373316 470694
rect 373264 470630 373316 470636
rect 373276 451926 373304 470630
rect 375378 466712 375434 466721
rect 375378 466647 375434 466656
rect 378046 466712 378102 466721
rect 378046 466647 378102 466656
rect 375392 458289 375420 466647
rect 378060 458289 378088 466647
rect 375378 458280 375434 458289
rect 375378 458215 375434 458224
rect 378046 458280 378102 458289
rect 378046 458215 378102 458224
rect 373264 451920 373316 451926
rect 373264 451862 373316 451868
rect 372988 448860 373040 448866
rect 372988 448802 373040 448808
rect 372646 448446 372936 448474
rect 344744 445664 344796 445670
rect 344650 445632 344706 445641
rect 316868 445596 316920 445602
rect 316868 445538 316920 445544
rect 323032 445596 323084 445602
rect 344744 445606 344796 445612
rect 352024 445602 352052 448052
rect 362328 445670 362356 448052
rect 373000 445738 373028 448802
rect 372988 445732 373040 445738
rect 372988 445674 373040 445680
rect 362316 445664 362368 445670
rect 362316 445606 362368 445612
rect 344650 445567 344706 445576
rect 352012 445596 352064 445602
rect 323032 445538 323084 445544
rect 352012 445538 352064 445544
rect 250352 445528 250404 445534
rect 250352 445470 250404 445476
rect 288992 445528 289044 445534
rect 288992 445470 289044 445476
rect 250628 444508 250680 444514
rect 250628 444450 250680 444456
rect 261484 444508 261536 444514
rect 261484 444450 261536 444456
rect 278596 444508 278648 444514
rect 278596 444450 278648 444456
rect 295432 444508 295484 444514
rect 295432 444450 295484 444456
rect 334624 444508 334676 444514
rect 334624 444450 334676 444456
rect 345848 444508 345900 444514
rect 345848 444450 345900 444456
rect 362316 444508 362368 444514
rect 362316 444450 362368 444456
rect 250640 441932 250668 444450
rect 240152 441238 240350 441266
rect 260958 441238 261064 441266
rect 234710 431760 234766 431769
rect 234710 431695 234766 431704
rect 238666 431760 238722 431769
rect 238666 431695 238722 431704
rect 234724 423337 234752 431695
rect 234710 423328 234766 423337
rect 234710 423263 234766 423272
rect 238680 423065 238708 431695
rect 238666 423056 238722 423065
rect 238666 422991 238722 423000
rect 240152 419422 240180 441238
rect 240336 419422 240364 421124
rect 240140 419416 240192 419422
rect 240140 419358 240192 419364
rect 240324 419416 240376 419422
rect 240324 419358 240376 419364
rect 250640 419354 250668 421124
rect 260944 419490 260972 421124
rect 261036 419490 261064 441238
rect 260932 419484 260984 419490
rect 260932 419426 260984 419432
rect 261024 419484 261076 419490
rect 261024 419426 261076 419432
rect 261496 419422 261524 444450
rect 267832 444440 267884 444446
rect 267832 444382 267884 444388
rect 261576 438932 261628 438938
rect 261576 438874 261628 438880
rect 261484 419416 261536 419422
rect 261484 419358 261536 419364
rect 261588 419354 261616 438874
rect 266266 431760 266322 431769
rect 266266 431695 266322 431704
rect 266280 423337 266308 431695
rect 266266 423328 266322 423337
rect 266266 423263 266322 423272
rect 267844 421682 267872 444382
rect 278608 441932 278636 444450
rect 295444 441614 295472 444450
rect 306472 444440 306524 444446
rect 306472 444382 306524 444388
rect 318064 444440 318116 444446
rect 318064 444382 318116 444388
rect 324320 444440 324372 444446
rect 324320 444382 324372 444388
rect 306484 441946 306512 444382
rect 306484 441918 306636 441946
rect 295444 441586 295932 441614
rect 267936 441238 268318 441266
rect 288926 441238 289124 441266
rect 267936 438938 267964 441238
rect 267924 438932 267976 438938
rect 267924 438874 267976 438880
rect 267844 421654 268318 421682
rect 278608 419422 278636 421124
rect 288912 419490 288940 421124
rect 289096 419490 289124 441238
rect 289176 438932 289228 438938
rect 289176 438874 289228 438880
rect 288900 419484 288952 419490
rect 288900 419426 288952 419432
rect 289084 419484 289136 419490
rect 289084 419426 289136 419432
rect 289188 419422 289216 438874
rect 293866 431760 293922 431769
rect 293866 431695 293922 431704
rect 293880 423201 293908 431695
rect 293866 423192 293922 423201
rect 293866 423127 293922 423136
rect 295904 421682 295932 441586
rect 295996 441238 296332 441266
rect 316940 441238 317092 441266
rect 295996 438938 296024 441238
rect 295984 438932 296036 438938
rect 295984 438874 296036 438880
rect 295904 421654 296332 421682
rect 306636 421110 306972 421138
rect 306944 419422 306972 421110
rect 316604 421110 316940 421138
rect 316604 419490 316632 421110
rect 317064 419490 317092 441238
rect 316592 419484 316644 419490
rect 316592 419426 316644 419432
rect 317052 419484 317104 419490
rect 317052 419426 317104 419432
rect 318076 419422 318104 444382
rect 324332 441932 324360 444382
rect 334636 441932 334664 444450
rect 345664 444440 345716 444446
rect 345664 444382 345716 444388
rect 344954 441250 345060 441266
rect 344954 441244 345072 441250
rect 344954 441238 345020 441244
rect 345020 441186 345072 441192
rect 318798 431760 318854 431769
rect 318798 431695 318854 431704
rect 322846 431760 322902 431769
rect 322846 431695 322902 431704
rect 318812 423337 318840 431695
rect 322860 423337 322888 431695
rect 318798 423328 318854 423337
rect 318798 423263 318854 423272
rect 322846 423328 322902 423337
rect 322846 423263 322902 423272
rect 324332 419422 324360 421124
rect 278596 419416 278648 419422
rect 278596 419358 278648 419364
rect 289176 419416 289228 419422
rect 289176 419358 289228 419364
rect 306932 419416 306984 419422
rect 306932 419358 306984 419364
rect 318064 419416 318116 419422
rect 318064 419358 318116 419364
rect 324320 419416 324372 419422
rect 324320 419358 324372 419364
rect 334636 419354 334664 421124
rect 344940 419490 344968 421124
rect 344928 419484 344980 419490
rect 344928 419426 344980 419432
rect 345676 419354 345704 444382
rect 345756 441244 345808 441250
rect 345756 441186 345808 441192
rect 345768 419490 345796 441186
rect 345756 419484 345808 419490
rect 345756 419426 345808 419432
rect 345860 419422 345888 444450
rect 352012 444440 352064 444446
rect 352012 444382 352064 444388
rect 352024 441946 352052 444382
rect 362328 441946 362356 444450
rect 352024 441918 352360 441946
rect 362328 441918 362664 441946
rect 372968 441238 373120 441266
rect 350446 431760 350502 431769
rect 350446 431695 350502 431704
rect 350460 423201 350488 431695
rect 350446 423192 350502 423201
rect 350446 423127 350502 423136
rect 352360 421110 352696 421138
rect 362664 421110 362908 421138
rect 352668 419529 352696 421110
rect 352654 419520 352710 419529
rect 352654 419455 352710 419464
rect 362880 419422 362908 421110
rect 372632 421110 372968 421138
rect 372632 419490 372660 421110
rect 373092 419490 373120 441238
rect 373264 439544 373316 439550
rect 373264 439486 373316 439492
rect 372620 419484 372672 419490
rect 372620 419426 372672 419432
rect 373080 419484 373132 419490
rect 373080 419426 373132 419432
rect 373276 419422 373304 439486
rect 378046 431760 378102 431769
rect 378046 431695 378102 431704
rect 378060 423337 378088 431695
rect 378046 423328 378102 423337
rect 378046 423263 378102 423272
rect 345848 419416 345900 419422
rect 345848 419358 345900 419364
rect 362868 419416 362920 419422
rect 362868 419358 362920 419364
rect 373264 419416 373316 419422
rect 373264 419358 373316 419364
rect 250628 419348 250680 419354
rect 250628 419290 250680 419296
rect 261576 419348 261628 419354
rect 261576 419290 261628 419296
rect 334624 419348 334676 419354
rect 334624 419290 334676 419296
rect 345664 419348 345716 419354
rect 345664 419290 345716 419296
rect 268016 416968 268068 416974
rect 268016 416910 268068 416916
rect 289084 416968 289136 416974
rect 289084 416910 289136 416916
rect 261484 416900 261536 416906
rect 261484 416842 261536 416848
rect 250352 416832 250404 416838
rect 250352 416774 250404 416780
rect 250364 414868 250392 416774
rect 260378 414488 260434 414497
rect 260434 414446 260682 414474
rect 260378 414423 260434 414432
rect 238864 414310 240074 414338
rect 234710 404288 234766 404297
rect 234710 404223 234766 404232
rect 234724 396001 234752 404223
rect 234710 395992 234766 396001
rect 234710 395927 234766 395936
rect 238864 391950 238892 414310
rect 261496 402974 261524 416842
rect 268028 414868 268056 416910
rect 278320 416900 278372 416906
rect 278320 416842 278372 416848
rect 278332 414868 278360 416842
rect 288900 416832 288952 416838
rect 288900 416774 288952 416780
rect 288650 414310 288848 414338
rect 262218 404288 262274 404297
rect 262218 404223 262274 404232
rect 266266 404288 266322 404297
rect 266266 404223 266322 404232
rect 261128 402946 261524 402974
rect 261128 394618 261156 402946
rect 262232 395729 262260 404223
rect 266280 396001 266308 404223
rect 266266 395992 266322 396001
rect 266266 395927 266322 395936
rect 262218 395720 262274 395729
rect 262218 395655 262274 395664
rect 288820 394874 288848 414310
rect 288808 394868 288860 394874
rect 288808 394810 288860 394816
rect 288912 394754 288940 416774
rect 289096 396506 289124 416910
rect 372896 416900 372948 416906
rect 372896 416842 372948 416848
rect 306012 416832 306064 416838
rect 306012 416774 306064 416780
rect 316960 416832 317012 416838
rect 316960 416774 317012 416780
rect 334348 416832 334400 416838
rect 334348 416774 334400 416780
rect 352012 416832 352064 416838
rect 352012 416774 352064 416780
rect 306024 414882 306052 416774
rect 306024 414854 306360 414882
rect 295444 414310 296056 414338
rect 316664 414310 316908 414338
rect 291198 404288 291254 404297
rect 291198 404223 291254 404232
rect 289084 396500 289136 396506
rect 289084 396442 289136 396448
rect 291212 395865 291240 404223
rect 291198 395856 291254 395865
rect 291198 395791 291254 395800
rect 288650 394726 288940 394754
rect 260682 394590 261156 394618
rect 288808 394664 288860 394670
rect 288808 394606 288860 394612
rect 238852 391944 238904 391950
rect 238852 391886 238904 391892
rect 240060 391882 240088 394060
rect 240048 391876 240100 391882
rect 240048 391818 240100 391824
rect 250364 391746 250392 394060
rect 268028 391882 268056 394060
rect 268016 391876 268068 391882
rect 268016 391818 268068 391824
rect 278332 391814 278360 394060
rect 278320 391808 278372 391814
rect 278320 391750 278372 391756
rect 288820 391746 288848 394606
rect 295444 391950 295472 414310
rect 316880 412826 316908 414310
rect 316868 412820 316920 412826
rect 316868 412762 316920 412768
rect 316868 412616 316920 412622
rect 316868 412558 316920 412564
rect 316776 408740 316828 408746
rect 316776 408682 316828 408688
rect 295708 396500 295760 396506
rect 295708 396442 295760 396448
rect 295720 394754 295748 396442
rect 316788 394754 316816 408682
rect 295720 394726 296056 394754
rect 316664 394726 316816 394754
rect 306300 394046 306360 394074
rect 295432 391944 295484 391950
rect 295432 391886 295484 391892
rect 306300 391882 306328 394046
rect 306288 391876 306340 391882
rect 306288 391818 306340 391824
rect 316880 391814 316908 412558
rect 316972 408746 317000 416774
rect 334360 414868 334388 416774
rect 352024 414868 352052 416774
rect 361946 414488 362002 414497
rect 362002 414446 362342 414474
rect 361946 414423 362002 414432
rect 323044 414310 324070 414338
rect 344678 414310 344784 414338
rect 372646 414310 372844 414338
rect 316960 408740 317012 408746
rect 316960 408682 317012 408688
rect 318798 404288 318854 404297
rect 318798 404223 318854 404232
rect 318812 396001 318840 404223
rect 318798 395992 318854 396001
rect 318798 395927 318854 395936
rect 323044 391814 323072 414310
rect 324056 391950 324084 394060
rect 334360 391950 334388 394060
rect 324044 391944 324096 391950
rect 324044 391886 324096 391892
rect 334348 391944 334400 391950
rect 344664 391921 344692 394060
rect 334348 391886 334400 391892
rect 344650 391912 344706 391921
rect 344756 391882 344784 414310
rect 346398 404288 346454 404297
rect 346398 404223 346454 404232
rect 350446 404288 350502 404297
rect 350446 404223 350502 404232
rect 346412 395729 346440 404223
rect 350460 396001 350488 404223
rect 350446 395992 350502 396001
rect 350446 395927 350502 395936
rect 346398 395720 346454 395729
rect 346398 395655 346454 395664
rect 372816 394874 372844 414310
rect 372804 394868 372856 394874
rect 372804 394810 372856 394816
rect 372908 394754 372936 416842
rect 373264 416832 373316 416838
rect 373264 416774 373316 416780
rect 373276 396778 373304 416774
rect 375378 404288 375434 404297
rect 375378 404223 375434 404232
rect 378046 404288 378102 404297
rect 378046 404223 378102 404232
rect 373264 396772 373316 396778
rect 373264 396714 373316 396720
rect 375392 395865 375420 404223
rect 378060 395865 378088 404223
rect 375378 395856 375434 395865
rect 375378 395791 375434 395800
rect 378046 395856 378102 395865
rect 378046 395791 378102 395800
rect 372646 394726 372936 394754
rect 372804 394664 372856 394670
rect 372804 394606 372856 394612
rect 344650 391847 344706 391856
rect 344744 391876 344796 391882
rect 344744 391818 344796 391824
rect 352024 391814 352052 394060
rect 362328 391882 362356 394060
rect 372816 391950 372844 394606
rect 372804 391944 372856 391950
rect 372804 391886 372856 391892
rect 362316 391876 362368 391882
rect 362316 391818 362368 391824
rect 316868 391808 316920 391814
rect 316868 391750 316920 391756
rect 323032 391808 323084 391814
rect 323032 391750 323084 391756
rect 352012 391808 352064 391814
rect 352012 391750 352064 391756
rect 250352 391740 250404 391746
rect 250352 391682 250404 391688
rect 288808 391740 288860 391746
rect 288808 391682 288860 391688
rect 250628 389292 250680 389298
rect 250628 389234 250680 389240
rect 261484 389292 261536 389298
rect 261484 389234 261536 389240
rect 278596 389292 278648 389298
rect 278596 389234 278648 389240
rect 295432 389292 295484 389298
rect 295432 389234 295484 389240
rect 334624 389292 334676 389298
rect 334624 389234 334676 389240
rect 345756 389292 345808 389298
rect 345756 389234 345808 389240
rect 362316 389292 362368 389298
rect 362316 389234 362368 389240
rect 240324 389224 240376 389230
rect 240324 389166 240376 389172
rect 240336 387940 240364 389166
rect 250640 387940 250668 389234
rect 260958 387246 261064 387274
rect 234710 377768 234766 377777
rect 234710 377703 234766 377712
rect 238666 377768 238722 377777
rect 238666 377703 238722 377712
rect 234724 369345 234752 377703
rect 238680 369345 238708 377703
rect 234710 369336 234766 369345
rect 234710 369271 234766 369280
rect 238666 369336 238722 369345
rect 238666 369271 238722 369280
rect 240336 365634 240364 367132
rect 240324 365628 240376 365634
rect 240324 365570 240376 365576
rect 250640 365566 250668 367132
rect 260944 365702 260972 367132
rect 261036 365702 261064 387246
rect 260932 365696 260984 365702
rect 260932 365638 260984 365644
rect 261024 365696 261076 365702
rect 261024 365638 261076 365644
rect 261496 365634 261524 389234
rect 267832 389224 267884 389230
rect 267832 389166 267884 389172
rect 267740 384804 267792 384810
rect 267740 384746 267792 384752
rect 262218 377768 262274 377777
rect 262218 377703 262274 377712
rect 266266 377768 266322 377777
rect 266266 377703 266322 377712
rect 262232 368490 262260 377703
rect 266280 368490 266308 377703
rect 262220 368484 262272 368490
rect 262220 368426 262272 368432
rect 266268 368484 266320 368490
rect 266268 368426 266320 368432
rect 261484 365628 261536 365634
rect 261484 365570 261536 365576
rect 267752 365566 267780 384746
rect 267844 367690 267872 389166
rect 278608 387940 278636 389234
rect 267936 387246 268318 387274
rect 288926 387246 289124 387274
rect 267936 384810 267964 387246
rect 267924 384804 267976 384810
rect 267924 384746 267976 384752
rect 267844 367662 268318 367690
rect 278608 365634 278636 367132
rect 288912 365702 288940 367132
rect 289096 365702 289124 387246
rect 295340 385484 295392 385490
rect 295340 385426 295392 385432
rect 291198 377768 291254 377777
rect 291198 377703 291254 377712
rect 293866 377768 293922 377777
rect 293866 377703 293922 377712
rect 291212 369345 291240 377703
rect 293880 369345 293908 377703
rect 291198 369336 291254 369345
rect 291198 369271 291254 369280
rect 293866 369336 293922 369345
rect 293866 369271 293922 369280
rect 288900 365696 288952 365702
rect 288900 365638 288952 365644
rect 289084 365696 289136 365702
rect 289084 365638 289136 365644
rect 295352 365634 295380 385426
rect 295444 383654 295472 389234
rect 306472 389224 306524 389230
rect 306472 389166 306524 389172
rect 318064 389224 318116 389230
rect 318064 389166 318116 389172
rect 324320 389224 324372 389230
rect 324320 389166 324372 389172
rect 306484 387954 306512 389166
rect 306484 387926 306636 387954
rect 295996 387246 296332 387274
rect 316940 387246 317092 387274
rect 295996 385490 296024 387246
rect 295984 385484 296036 385490
rect 295984 385426 296036 385432
rect 295444 383626 295932 383654
rect 295904 367690 295932 383626
rect 295904 367662 296332 367690
rect 306636 367118 306972 367146
rect 306944 365634 306972 367118
rect 316604 367118 316940 367146
rect 316604 365702 316632 367118
rect 317064 365702 317092 387246
rect 316592 365696 316644 365702
rect 316592 365638 316644 365644
rect 317052 365696 317104 365702
rect 317052 365638 317104 365644
rect 318076 365634 318104 389166
rect 324332 387940 324360 389166
rect 334636 387940 334664 389234
rect 345664 389224 345716 389230
rect 345664 389166 345716 389172
rect 344954 387258 345060 387274
rect 344954 387252 345072 387258
rect 344954 387246 345020 387252
rect 345020 387194 345072 387200
rect 318798 377768 318854 377777
rect 318798 377703 318854 377712
rect 322846 377768 322902 377777
rect 322846 377703 322902 377712
rect 318812 368490 318840 377703
rect 322860 368490 322888 377703
rect 318800 368484 318852 368490
rect 318800 368426 318852 368432
rect 322848 368484 322900 368490
rect 322848 368426 322900 368432
rect 324332 365634 324360 367132
rect 278596 365628 278648 365634
rect 278596 365570 278648 365576
rect 295340 365628 295392 365634
rect 295340 365570 295392 365576
rect 306932 365628 306984 365634
rect 306932 365570 306984 365576
rect 318064 365628 318116 365634
rect 318064 365570 318116 365576
rect 324320 365628 324372 365634
rect 324320 365570 324372 365576
rect 334636 365566 334664 367132
rect 344940 365702 344968 367132
rect 344928 365696 344980 365702
rect 344928 365638 344980 365644
rect 345676 365566 345704 389166
rect 345768 365634 345796 389234
rect 352012 389224 352064 389230
rect 352012 389166 352064 389172
rect 352024 387954 352052 389166
rect 362328 387954 362356 389234
rect 352024 387926 352360 387954
rect 362328 387926 362664 387954
rect 345848 387252 345900 387258
rect 372968 387246 373120 387274
rect 345848 387194 345900 387200
rect 345860 365702 345888 387194
rect 346398 377768 346454 377777
rect 346398 377703 346454 377712
rect 350446 377768 350502 377777
rect 350446 377703 350502 377712
rect 346412 369345 346440 377703
rect 350460 369345 350488 377703
rect 346398 369336 346454 369345
rect 346398 369271 346454 369280
rect 350446 369336 350502 369345
rect 350446 369271 350502 369280
rect 352360 367118 352696 367146
rect 362664 367118 362908 367146
rect 345848 365696 345900 365702
rect 352668 365673 352696 367118
rect 345848 365638 345900 365644
rect 352654 365664 352710 365673
rect 345756 365628 345808 365634
rect 362880 365634 362908 367118
rect 372632 367118 372968 367146
rect 372632 365702 372660 367118
rect 373092 365702 373120 387246
rect 375378 377768 375434 377777
rect 375378 377703 375434 377712
rect 378046 377768 378102 377777
rect 378046 377703 378102 377712
rect 375392 368490 375420 377703
rect 378060 368490 378088 377703
rect 375380 368484 375432 368490
rect 375380 368426 375432 368432
rect 378048 368484 378100 368490
rect 378048 368426 378100 368432
rect 372620 365696 372672 365702
rect 372620 365638 372672 365644
rect 373080 365696 373132 365702
rect 373080 365638 373132 365644
rect 352654 365599 352710 365608
rect 362868 365628 362920 365634
rect 345756 365570 345808 365576
rect 362868 365570 362920 365576
rect 250628 365560 250680 365566
rect 250628 365502 250680 365508
rect 267740 365560 267792 365566
rect 267740 365502 267792 365508
rect 334624 365560 334676 365566
rect 334624 365502 334676 365508
rect 345664 365560 345716 365566
rect 345664 365502 345716 365508
rect 261484 363044 261536 363050
rect 261484 362986 261536 362992
rect 278320 363044 278372 363050
rect 278320 362986 278372 362992
rect 288900 363044 288952 363050
rect 288900 362986 288952 362992
rect 306012 363044 306064 363050
rect 306012 362986 306064 362992
rect 317144 363044 317196 363050
rect 317144 362986 317196 362992
rect 334348 363044 334400 363050
rect 334348 362986 334400 362992
rect 372896 363044 372948 363050
rect 372896 362986 372948 362992
rect 250352 362976 250404 362982
rect 250352 362918 250404 362924
rect 250364 360876 250392 362918
rect 260378 360496 260434 360505
rect 260434 360454 260682 360482
rect 260378 360431 260434 360440
rect 238864 360318 240074 360346
rect 234710 350296 234766 350305
rect 234710 350231 234766 350240
rect 234724 342009 234752 350231
rect 234710 342000 234766 342009
rect 234710 341935 234766 341944
rect 238864 338094 238892 360318
rect 261496 345014 261524 362986
rect 268016 362976 268068 362982
rect 268016 362918 268068 362924
rect 268028 360876 268056 362918
rect 278332 360876 278360 362986
rect 288650 360318 288848 360346
rect 262218 350296 262274 350305
rect 262218 350231 262274 350240
rect 266266 350296 266322 350305
rect 266266 350231 266322 350240
rect 261128 344986 261524 345014
rect 261128 340762 261156 344986
rect 262232 341737 262260 350231
rect 266280 342009 266308 350231
rect 266266 342000 266322 342009
rect 266266 341935 266322 341944
rect 262218 341728 262274 341737
rect 262218 341663 262274 341672
rect 288820 340950 288848 360318
rect 288808 340944 288860 340950
rect 288808 340886 288860 340892
rect 260682 340734 261156 340762
rect 288912 340490 288940 362986
rect 289084 362976 289136 362982
rect 289084 362918 289136 362924
rect 289096 342582 289124 362918
rect 306024 360890 306052 362986
rect 317052 362976 317104 362982
rect 317052 362918 317104 362924
rect 306024 360862 306360 360890
rect 316664 360590 317000 360618
rect 295444 360318 296056 360346
rect 291198 350296 291254 350305
rect 291198 350231 291254 350240
rect 289084 342576 289136 342582
rect 289084 342518 289136 342524
rect 291212 341873 291240 350231
rect 291198 341864 291254 341873
rect 291198 341799 291254 341808
rect 288992 340944 289044 340950
rect 288992 340886 289044 340892
rect 288650 340462 288940 340490
rect 238852 338088 238904 338094
rect 238852 338030 238904 338036
rect 240060 338026 240088 340068
rect 240048 338020 240100 338026
rect 240048 337962 240100 337968
rect 250364 337958 250392 340068
rect 268028 338026 268056 340068
rect 278332 338026 278360 340068
rect 268016 338020 268068 338026
rect 268016 337962 268068 337968
rect 278320 338020 278372 338026
rect 278320 337962 278372 337968
rect 289004 337958 289032 340886
rect 295444 338094 295472 360318
rect 316776 358896 316828 358902
rect 316776 358838 316828 358844
rect 295708 342576 295760 342582
rect 295708 342518 295760 342524
rect 295720 340762 295748 342518
rect 316788 340762 316816 358838
rect 316868 358828 316920 358834
rect 316868 358770 316920 358776
rect 295720 340734 296056 340762
rect 316664 340734 316816 340762
rect 306300 340054 306360 340082
rect 295432 338088 295484 338094
rect 295432 338030 295484 338036
rect 306300 337958 306328 340054
rect 316880 337958 316908 358770
rect 316972 338026 317000 360590
rect 317064 358834 317092 362918
rect 317156 358902 317184 362986
rect 334360 360876 334388 362986
rect 344652 362976 344704 362982
rect 344652 362918 344704 362924
rect 352012 362976 352064 362982
rect 352012 362918 352064 362924
rect 344664 360876 344692 362918
rect 352024 360876 352052 362918
rect 361946 360496 362002 360505
rect 362002 360454 362342 360482
rect 361946 360431 362002 360440
rect 323044 360318 324070 360346
rect 372646 360318 372844 360346
rect 317144 358896 317196 358902
rect 317144 358838 317196 358844
rect 317052 358828 317104 358834
rect 317052 358770 317104 358776
rect 318798 350296 318854 350305
rect 318798 350231 318854 350240
rect 318812 342009 318840 350231
rect 318798 342000 318854 342009
rect 318798 341935 318854 341944
rect 323044 338026 323072 360318
rect 346398 350296 346454 350305
rect 346398 350231 346454 350240
rect 350446 350296 350502 350305
rect 350446 350231 350502 350240
rect 346412 341737 346440 350231
rect 350460 342009 350488 350231
rect 372816 345710 372844 360318
rect 372804 345704 372856 345710
rect 372804 345646 372856 345652
rect 350446 342000 350502 342009
rect 350446 341935 350502 341944
rect 346398 341728 346454 341737
rect 346398 341663 346454 341672
rect 372908 340490 372936 362986
rect 373264 362976 373316 362982
rect 373264 362918 373316 362924
rect 372988 345704 373040 345710
rect 372988 345646 373040 345652
rect 372646 340462 372936 340490
rect 324056 338094 324084 340068
rect 334360 338094 334388 340068
rect 324044 338088 324096 338094
rect 324044 338030 324096 338036
rect 334348 338088 334400 338094
rect 344664 338065 344692 340068
rect 334348 338030 334400 338036
rect 344650 338056 344706 338065
rect 316960 338020 317012 338026
rect 316960 337962 317012 337968
rect 323032 338020 323084 338026
rect 352024 338026 352052 340068
rect 362328 338026 362356 340068
rect 373000 338094 373028 345646
rect 373276 342922 373304 362918
rect 375378 350296 375434 350305
rect 375378 350231 375434 350240
rect 378046 350296 378102 350305
rect 378046 350231 378102 350240
rect 373264 342916 373316 342922
rect 373264 342858 373316 342864
rect 375392 341873 375420 350231
rect 378060 341873 378088 350231
rect 375378 341864 375434 341873
rect 375378 341799 375434 341808
rect 378046 341864 378102 341873
rect 378046 341799 378102 341808
rect 372988 338088 373040 338094
rect 372988 338030 373040 338036
rect 344650 337991 344706 338000
rect 352012 338020 352064 338026
rect 323032 337962 323084 337968
rect 352012 337962 352064 337968
rect 362316 338020 362368 338026
rect 362316 337962 362368 337968
rect 250352 337952 250404 337958
rect 250352 337894 250404 337900
rect 288992 337952 289044 337958
rect 288992 337894 289044 337900
rect 306288 337952 306340 337958
rect 306288 337894 306340 337900
rect 316868 337952 316920 337958
rect 316868 337894 316920 337900
rect 250628 335436 250680 335442
rect 250628 335378 250680 335384
rect 267832 335436 267884 335442
rect 267832 335378 267884 335384
rect 306380 335436 306432 335442
rect 306380 335378 306432 335384
rect 318064 335436 318116 335442
rect 318064 335378 318116 335384
rect 324320 335436 324372 335442
rect 324320 335378 324372 335384
rect 345756 335436 345808 335442
rect 345756 335378 345808 335384
rect 362316 335436 362368 335442
rect 362316 335378 362368 335384
rect 240324 335368 240376 335374
rect 240324 335310 240376 335316
rect 240336 333948 240364 335310
rect 250640 333948 250668 335378
rect 261484 335368 261536 335374
rect 261484 335310 261536 335316
rect 260958 333254 261064 333282
rect 234710 323776 234766 323785
rect 234710 323711 234766 323720
rect 238666 323776 238722 323785
rect 238666 323711 238722 323720
rect 234724 315353 234752 323711
rect 238680 315353 238708 323711
rect 234710 315344 234766 315353
rect 234710 315279 234766 315288
rect 238666 315344 238722 315353
rect 238666 315279 238722 315288
rect 240336 311778 240364 313140
rect 240324 311772 240376 311778
rect 240324 311714 240376 311720
rect 250640 311710 250668 313140
rect 260944 311846 260972 313140
rect 261036 311846 261064 333254
rect 260932 311840 260984 311846
rect 260932 311782 260984 311788
rect 261024 311840 261076 311846
rect 261024 311782 261076 311788
rect 261496 311778 261524 335310
rect 262220 332648 262272 332654
rect 262220 332590 262272 332596
rect 266268 332648 266320 332654
rect 266268 332590 266320 332596
rect 262232 323785 262260 332590
rect 266280 323785 266308 332590
rect 267740 329520 267792 329526
rect 267740 329462 267792 329468
rect 262218 323776 262274 323785
rect 262218 323711 262274 323720
rect 266266 323776 266322 323785
rect 266266 323711 266322 323720
rect 261484 311772 261536 311778
rect 261484 311714 261536 311720
rect 267752 311710 267780 329462
rect 267844 313698 267872 335378
rect 278596 335368 278648 335374
rect 278596 335310 278648 335316
rect 295432 335368 295484 335374
rect 295432 335310 295484 335316
rect 278608 333948 278636 335310
rect 267936 333254 268318 333282
rect 288926 333254 289124 333282
rect 267936 329526 267964 333254
rect 267924 329520 267976 329526
rect 267924 329462 267976 329468
rect 267844 313670 268318 313698
rect 278608 311778 278636 313140
rect 288912 311846 288940 313140
rect 289096 311846 289124 333254
rect 295340 329520 295392 329526
rect 295340 329462 295392 329468
rect 291198 323776 291254 323785
rect 291198 323711 291254 323720
rect 293866 323776 293922 323785
rect 293866 323711 293922 323720
rect 291212 315353 291240 323711
rect 293880 315353 293908 323711
rect 291198 315344 291254 315353
rect 291198 315279 291254 315288
rect 293866 315344 293922 315353
rect 293866 315279 293922 315288
rect 288900 311840 288952 311846
rect 288900 311782 288952 311788
rect 289084 311840 289136 311846
rect 289084 311782 289136 311788
rect 295352 311778 295380 329462
rect 295444 325694 295472 335310
rect 306392 333962 306420 335378
rect 306392 333934 306636 333962
rect 295996 333254 296332 333282
rect 316940 333254 317092 333282
rect 295996 329526 296024 333254
rect 295984 329520 296036 329526
rect 295984 329462 296036 329468
rect 295444 325666 295932 325694
rect 295904 313698 295932 325666
rect 295904 313670 296332 313698
rect 306636 313126 306972 313154
rect 306944 311778 306972 313126
rect 316604 313126 316940 313154
rect 316604 311846 316632 313126
rect 317064 311846 317092 333254
rect 316592 311840 316644 311846
rect 316592 311782 316644 311788
rect 317052 311840 317104 311846
rect 317052 311782 317104 311788
rect 318076 311778 318104 335378
rect 324332 333948 324360 335378
rect 334624 335368 334676 335374
rect 334624 335310 334676 335316
rect 345664 335368 345716 335374
rect 345664 335310 345716 335316
rect 334636 333948 334664 335310
rect 344954 333266 345060 333282
rect 344954 333260 345072 333266
rect 344954 333254 345020 333260
rect 345020 333202 345072 333208
rect 318800 332648 318852 332654
rect 318800 332590 318852 332596
rect 322848 332648 322900 332654
rect 322848 332590 322900 332596
rect 318812 323785 318840 332590
rect 322860 323785 322888 332590
rect 318798 323776 318854 323785
rect 318798 323711 318854 323720
rect 322846 323776 322902 323785
rect 322846 323711 322902 323720
rect 324332 311778 324360 313140
rect 278596 311772 278648 311778
rect 278596 311714 278648 311720
rect 295340 311772 295392 311778
rect 295340 311714 295392 311720
rect 306932 311772 306984 311778
rect 306932 311714 306984 311720
rect 318064 311772 318116 311778
rect 318064 311714 318116 311720
rect 324320 311772 324372 311778
rect 324320 311714 324372 311720
rect 334636 311710 334664 313140
rect 344940 311846 344968 313140
rect 344928 311840 344980 311846
rect 344928 311782 344980 311788
rect 345676 311710 345704 335310
rect 345768 311778 345796 335378
rect 352012 335368 352064 335374
rect 352012 335310 352064 335316
rect 352024 333962 352052 335310
rect 362328 333962 362356 335378
rect 352024 333934 352360 333962
rect 362328 333934 362664 333962
rect 345848 333260 345900 333266
rect 372968 333254 373120 333282
rect 345848 333202 345900 333208
rect 345860 311846 345888 333202
rect 346398 323776 346454 323785
rect 346398 323711 346454 323720
rect 350446 323776 350502 323785
rect 350446 323711 350502 323720
rect 346412 315353 346440 323711
rect 350460 315353 350488 323711
rect 346398 315344 346454 315353
rect 346398 315279 346454 315288
rect 350446 315344 350502 315353
rect 350446 315279 350502 315288
rect 352360 313126 352696 313154
rect 362664 313126 362908 313154
rect 345848 311840 345900 311846
rect 352668 311817 352696 313126
rect 345848 311782 345900 311788
rect 352654 311808 352710 311817
rect 345756 311772 345808 311778
rect 362880 311778 362908 313126
rect 372632 313126 372968 313154
rect 372632 311846 372660 313126
rect 373092 311846 373120 333254
rect 375380 332648 375432 332654
rect 375380 332590 375432 332596
rect 378048 332648 378100 332654
rect 378048 332590 378100 332596
rect 375392 323785 375420 332590
rect 378060 323785 378088 332590
rect 375378 323776 375434 323785
rect 375378 323711 375434 323720
rect 378046 323776 378102 323785
rect 378046 323711 378102 323720
rect 372620 311840 372672 311846
rect 372620 311782 372672 311788
rect 373080 311840 373132 311846
rect 373080 311782 373132 311788
rect 352654 311743 352710 311752
rect 362868 311772 362920 311778
rect 345756 311714 345808 311720
rect 362868 311714 362920 311720
rect 250628 311704 250680 311710
rect 250628 311646 250680 311652
rect 267740 311704 267792 311710
rect 267740 311646 267792 311652
rect 334624 311704 334676 311710
rect 334624 311646 334676 311652
rect 345664 311704 345716 311710
rect 345664 311646 345716 311652
rect 268016 309324 268068 309330
rect 268016 309266 268068 309272
rect 289084 309324 289136 309330
rect 289084 309266 289136 309272
rect 261484 309256 261536 309262
rect 261484 309198 261536 309204
rect 250352 309188 250404 309194
rect 250352 309130 250404 309136
rect 250364 306884 250392 309130
rect 260378 306504 260434 306513
rect 260434 306462 260682 306490
rect 260378 306439 260434 306448
rect 238864 306326 240074 306354
rect 234710 296304 234766 296313
rect 234710 296239 234766 296248
rect 238666 296304 238722 296313
rect 238666 296239 238722 296248
rect 234724 288017 234752 296239
rect 234710 288008 234766 288017
rect 234710 287943 234766 287952
rect 238680 287745 238708 296239
rect 238666 287736 238722 287745
rect 238666 287671 238722 287680
rect 238864 284306 238892 306326
rect 261496 287054 261524 309198
rect 268028 306884 268056 309266
rect 278320 309256 278372 309262
rect 278320 309198 278372 309204
rect 278332 306884 278360 309198
rect 288808 309188 288860 309194
rect 288808 309130 288860 309136
rect 288650 306326 288756 306354
rect 288728 306270 288756 306326
rect 288716 306264 288768 306270
rect 288716 306206 288768 306212
rect 262218 296304 262274 296313
rect 262218 296239 262274 296248
rect 266266 296304 266322 296313
rect 266266 296239 266322 296248
rect 262232 287881 262260 296239
rect 266280 288017 266308 296239
rect 266266 288008 266322 288017
rect 266266 287943 266322 287952
rect 262218 287872 262274 287881
rect 262218 287807 262274 287816
rect 261128 287026 261524 287054
rect 261128 286770 261156 287026
rect 288820 286770 288848 309130
rect 288900 306264 288952 306270
rect 288900 306206 288952 306212
rect 260682 286742 261156 286770
rect 288650 286742 288848 286770
rect 238852 284300 238904 284306
rect 238852 284242 238904 284248
rect 240060 284238 240088 286076
rect 240048 284232 240100 284238
rect 240048 284174 240100 284180
rect 250364 284170 250392 286076
rect 268028 284238 268056 286076
rect 278332 284238 278360 286076
rect 268016 284232 268068 284238
rect 268016 284174 268068 284180
rect 278320 284232 278372 284238
rect 278320 284174 278372 284180
rect 288912 284170 288940 306206
rect 289096 289814 289124 309266
rect 317144 309256 317196 309262
rect 317144 309198 317196 309204
rect 334348 309256 334400 309262
rect 334348 309198 334400 309204
rect 372804 309256 372856 309262
rect 372804 309198 372856 309204
rect 306012 309188 306064 309194
rect 306012 309130 306064 309136
rect 317052 309188 317104 309194
rect 317052 309130 317104 309136
rect 306024 306898 306052 309130
rect 306024 306870 306360 306898
rect 316664 306598 317000 306626
rect 295628 306326 296056 306354
rect 295628 296714 295656 306326
rect 316776 305720 316828 305726
rect 316776 305662 316828 305668
rect 295444 296686 295656 296714
rect 289084 289808 289136 289814
rect 289084 289750 289136 289756
rect 295444 284306 295472 296686
rect 295708 289808 295760 289814
rect 295708 289750 295760 289756
rect 295720 286770 295748 289750
rect 316788 286770 316816 305662
rect 316868 301572 316920 301578
rect 316868 301514 316920 301520
rect 295720 286742 296056 286770
rect 316664 286742 316816 286770
rect 306300 286062 306360 286090
rect 295432 284300 295484 284306
rect 295432 284242 295484 284248
rect 306300 284170 306328 286062
rect 316880 284170 316908 301514
rect 316972 284238 317000 306598
rect 317064 301578 317092 309130
rect 317156 305726 317184 309198
rect 334360 306884 334388 309198
rect 344652 309188 344704 309194
rect 344652 309130 344704 309136
rect 352012 309188 352064 309194
rect 352012 309130 352064 309136
rect 344664 306884 344692 309130
rect 352024 306884 352052 309130
rect 361946 306504 362002 306513
rect 362002 306462 362342 306490
rect 361946 306439 362002 306448
rect 372816 306374 372844 309198
rect 373264 309188 373316 309194
rect 373264 309130 373316 309136
rect 323596 306326 324070 306354
rect 372646 306326 372752 306354
rect 372816 306346 373028 306374
rect 317144 305720 317196 305726
rect 317144 305662 317196 305668
rect 317052 301572 317104 301578
rect 317052 301514 317104 301520
rect 323596 296714 323624 306326
rect 372724 306218 372752 306326
rect 372724 306190 372936 306218
rect 372804 301572 372856 301578
rect 372804 301514 372856 301520
rect 323044 296686 323624 296714
rect 318798 296304 318854 296313
rect 318798 296239 318854 296248
rect 322846 296304 322902 296313
rect 322846 296239 322902 296248
rect 318812 288017 318840 296239
rect 322860 288017 322888 296239
rect 318798 288008 318854 288017
rect 318798 287943 318854 287952
rect 322846 288008 322902 288017
rect 322846 287943 322902 287952
rect 323044 284238 323072 296686
rect 346398 296304 346454 296313
rect 346398 296239 346454 296248
rect 350446 296304 350502 296313
rect 350446 296239 350502 296248
rect 346412 287881 346440 296239
rect 350460 287881 350488 296239
rect 346398 287872 346454 287881
rect 346398 287807 346454 287816
rect 350446 287872 350502 287881
rect 350446 287807 350502 287816
rect 372816 286770 372844 301514
rect 372646 286742 372844 286770
rect 324056 284306 324084 286076
rect 334360 284306 334388 286076
rect 324044 284300 324096 284306
rect 324044 284242 324096 284248
rect 334348 284300 334400 284306
rect 334348 284242 334400 284248
rect 316960 284232 317012 284238
rect 316960 284174 317012 284180
rect 323032 284232 323084 284238
rect 344664 284209 344692 286076
rect 352024 284238 352052 286076
rect 362328 284238 362356 286076
rect 372908 284306 372936 306190
rect 373000 301578 373028 306346
rect 372988 301572 373040 301578
rect 372988 301514 373040 301520
rect 373276 289134 373304 309130
rect 378046 296304 378102 296313
rect 378046 296239 378102 296248
rect 373264 289128 373316 289134
rect 373264 289070 373316 289076
rect 378060 288017 378088 296239
rect 378046 288008 378102 288017
rect 378046 287943 378102 287952
rect 372896 284300 372948 284306
rect 372896 284242 372948 284248
rect 352012 284232 352064 284238
rect 323032 284174 323084 284180
rect 344650 284200 344706 284209
rect 250352 284164 250404 284170
rect 250352 284106 250404 284112
rect 288900 284164 288952 284170
rect 288900 284106 288952 284112
rect 306288 284164 306340 284170
rect 306288 284106 306340 284112
rect 316868 284164 316920 284170
rect 352012 284174 352064 284180
rect 362316 284232 362368 284238
rect 362316 284174 362368 284180
rect 344650 284135 344706 284144
rect 316868 284106 316920 284112
rect 250628 281648 250680 281654
rect 250628 281590 250680 281596
rect 295432 281648 295484 281654
rect 295432 281590 295484 281596
rect 334624 281648 334676 281654
rect 334624 281590 334676 281596
rect 240140 280152 240192 280158
rect 240140 280094 240192 280100
rect 240152 279970 240180 280094
rect 240152 279942 240350 279970
rect 250640 279956 250668 281590
rect 267832 281580 267884 281586
rect 267832 281522 267884 281528
rect 260958 279262 261064 279290
rect 234710 278080 234766 278089
rect 234710 278015 234766 278024
rect 238666 278080 238722 278089
rect 238666 278015 238722 278024
rect 234724 269793 234752 278015
rect 238680 269793 238708 278015
rect 234710 269784 234766 269793
rect 234710 269719 234766 269728
rect 238666 269784 238722 269793
rect 238666 269719 238722 269728
rect 240336 256601 240364 259148
rect 250640 256630 250668 259148
rect 260944 256698 260972 259148
rect 261036 256698 261064 279262
rect 262220 278792 262272 278798
rect 262220 278734 262272 278740
rect 266268 278792 266320 278798
rect 266268 278734 266320 278740
rect 262232 269793 262260 278734
rect 266280 269793 266308 278734
rect 267740 272604 267792 272610
rect 267740 272546 267792 272552
rect 262218 269784 262274 269793
rect 262218 269719 262274 269728
rect 266266 269784 266322 269793
rect 266266 269719 266322 269728
rect 260932 256692 260984 256698
rect 260932 256634 260984 256640
rect 261024 256692 261076 256698
rect 261024 256634 261076 256640
rect 267752 256630 267780 272546
rect 267844 259706 267872 281522
rect 278226 279848 278282 279857
rect 278282 279806 278622 279834
rect 278226 279783 278282 279792
rect 267936 279262 268318 279290
rect 288926 279262 289124 279290
rect 267936 272610 267964 279262
rect 267924 272604 267976 272610
rect 267924 272546 267976 272552
rect 267844 259678 268318 259706
rect 278608 256630 278636 259148
rect 288912 256698 288940 259148
rect 289096 256698 289124 279262
rect 291198 278080 291254 278089
rect 291198 278015 291254 278024
rect 293866 278080 293922 278089
rect 293866 278015 293922 278024
rect 291212 269793 291240 278015
rect 293880 269793 293908 278015
rect 295340 272604 295392 272610
rect 295340 272546 295392 272552
rect 291198 269784 291254 269793
rect 291198 269719 291254 269728
rect 293866 269784 293922 269793
rect 293866 269719 293922 269728
rect 288900 256692 288952 256698
rect 288900 256634 288952 256640
rect 289084 256692 289136 256698
rect 289084 256634 289136 256640
rect 295352 256630 295380 272546
rect 295444 267734 295472 281590
rect 306472 281580 306524 281586
rect 306472 281522 306524 281528
rect 318064 281580 318116 281586
rect 318064 281522 318116 281528
rect 324320 281580 324372 281586
rect 324320 281522 324372 281528
rect 306484 279970 306512 281522
rect 306484 279942 306636 279970
rect 295996 279262 296332 279290
rect 316940 279262 317092 279290
rect 295996 272610 296024 279262
rect 295984 272604 296036 272610
rect 295984 272546 296036 272552
rect 295444 267706 295932 267734
rect 295904 259706 295932 267706
rect 295904 259678 296332 259706
rect 306636 259134 306972 259162
rect 306944 256630 306972 259134
rect 316604 259134 316940 259162
rect 316604 256698 316632 259134
rect 317064 256698 317092 279262
rect 316592 256692 316644 256698
rect 316592 256634 316644 256640
rect 317052 256692 317104 256698
rect 317052 256634 317104 256640
rect 318076 256630 318104 281522
rect 324332 279956 324360 281522
rect 334636 279956 334664 281590
rect 345756 281580 345808 281586
rect 345756 281522 345808 281528
rect 362316 281580 362368 281586
rect 362316 281522 362368 281528
rect 344954 279262 345152 279290
rect 318800 278792 318852 278798
rect 318800 278734 318852 278740
rect 322848 278792 322900 278798
rect 322848 278734 322900 278740
rect 318812 269793 318840 278734
rect 322860 269793 322888 278734
rect 345124 277394 345152 279262
rect 345124 277366 345704 277394
rect 318798 269784 318854 269793
rect 318798 269719 318854 269728
rect 322846 269784 322902 269793
rect 322846 269719 322902 269728
rect 324332 256630 324360 259148
rect 250628 256624 250680 256630
rect 240322 256592 240378 256601
rect 250628 256566 250680 256572
rect 267740 256624 267792 256630
rect 267740 256566 267792 256572
rect 278596 256624 278648 256630
rect 278596 256566 278648 256572
rect 295340 256624 295392 256630
rect 295340 256566 295392 256572
rect 306932 256624 306984 256630
rect 306932 256566 306984 256572
rect 318064 256624 318116 256630
rect 318064 256566 318116 256572
rect 324320 256624 324372 256630
rect 324320 256566 324372 256572
rect 334636 256562 334664 259148
rect 344940 256698 344968 259148
rect 345676 256698 345704 277366
rect 344928 256692 344980 256698
rect 344928 256634 344980 256640
rect 345664 256692 345716 256698
rect 345664 256634 345716 256640
rect 345768 256630 345796 281522
rect 362328 279970 362356 281522
rect 362328 279942 362664 279970
rect 351932 279262 352360 279290
rect 372968 279262 373120 279290
rect 346398 278080 346454 278089
rect 346398 278015 346454 278024
rect 350446 278080 350502 278089
rect 350446 278015 350502 278024
rect 346412 269793 346440 278015
rect 350460 269793 350488 278015
rect 346398 269784 346454 269793
rect 346398 269719 346454 269728
rect 350446 269784 350502 269793
rect 350446 269719 350502 269728
rect 345756 256624 345808 256630
rect 345756 256566 345808 256572
rect 351932 256562 351960 279262
rect 352360 259134 352696 259162
rect 362664 259134 362908 259162
rect 352668 256601 352696 259134
rect 362880 256630 362908 259134
rect 372632 259134 372968 259162
rect 372632 256698 372660 259134
rect 373092 256698 373120 279262
rect 375380 278792 375432 278798
rect 375380 278734 375432 278740
rect 378048 278792 378100 278798
rect 378048 278734 378100 278740
rect 375392 269793 375420 278734
rect 378060 269793 378088 278734
rect 375378 269784 375434 269793
rect 375378 269719 375434 269728
rect 378046 269784 378102 269793
rect 378046 269719 378102 269728
rect 372620 256692 372672 256698
rect 372620 256634 372672 256640
rect 373080 256692 373132 256698
rect 373080 256634 373132 256640
rect 362868 256624 362920 256630
rect 352654 256592 352710 256601
rect 240322 256527 240378 256536
rect 334624 256556 334676 256562
rect 334624 256498 334676 256504
rect 351920 256556 351972 256562
rect 362868 256566 362920 256572
rect 352654 256527 352710 256536
rect 351920 256498 351972 256504
rect 268016 255468 268068 255474
rect 268016 255410 268068 255416
rect 289176 255468 289228 255474
rect 289176 255410 289228 255416
rect 261484 255400 261536 255406
rect 261484 255342 261536 255348
rect 250352 255332 250404 255338
rect 250352 255274 250404 255280
rect 250364 252892 250392 255274
rect 260378 252648 260434 252657
rect 260434 252606 260682 252634
rect 260378 252583 260434 252592
rect 238864 252334 240074 252362
rect 234710 242312 234766 242321
rect 234710 242247 234766 242256
rect 238666 242312 238722 242321
rect 238666 242247 238722 242256
rect 234724 234025 234752 242247
rect 238680 234025 238708 242247
rect 234710 234016 234766 234025
rect 234710 233951 234766 233960
rect 238666 234016 238722 234025
rect 238666 233951 238722 233960
rect 238864 230450 238892 252334
rect 261496 238754 261524 255342
rect 268028 252892 268056 255410
rect 278320 255400 278372 255406
rect 278320 255342 278372 255348
rect 278332 252892 278360 255342
rect 289084 255332 289136 255338
rect 289084 255274 289136 255280
rect 289096 252362 289124 255274
rect 288650 252334 288848 252362
rect 288820 251326 288848 252334
rect 289004 252334 289124 252362
rect 288808 251320 288860 251326
rect 288808 251262 288860 251268
rect 289004 249098 289032 252334
rect 289084 251320 289136 251326
rect 289084 251262 289136 251268
rect 288820 249070 289032 249098
rect 262218 242312 262274 242321
rect 262218 242247 262274 242256
rect 266266 242312 266322 242321
rect 266266 242247 266322 242256
rect 261128 238726 261524 238754
rect 261128 232778 261156 238726
rect 262232 233238 262260 242247
rect 266280 233238 266308 242247
rect 262220 233232 262272 233238
rect 262220 233174 262272 233180
rect 266268 233232 266320 233238
rect 266268 233174 266320 233180
rect 288820 232778 288848 249070
rect 289096 244338 289124 251262
rect 260682 232750 261156 232778
rect 288650 232750 288848 232778
rect 288912 244310 289124 244338
rect 238852 230444 238904 230450
rect 238852 230386 238904 230392
rect 240060 230382 240088 232084
rect 240048 230376 240100 230382
rect 240048 230318 240100 230324
rect 250364 230314 250392 232084
rect 268028 230382 268056 232084
rect 278332 230382 278360 232084
rect 268016 230376 268068 230382
rect 268016 230318 268068 230324
rect 278320 230376 278372 230382
rect 278320 230318 278372 230324
rect 288912 230314 288940 244310
rect 289188 235074 289216 255410
rect 317144 255400 317196 255406
rect 317144 255342 317196 255348
rect 334348 255400 334400 255406
rect 334348 255342 334400 255348
rect 372988 255400 373040 255406
rect 372988 255342 373040 255348
rect 306012 255332 306064 255338
rect 306012 255274 306064 255280
rect 317052 255332 317104 255338
rect 317052 255274 317104 255280
rect 306024 252906 306052 255274
rect 306024 252878 306360 252906
rect 316664 252606 317000 252634
rect 295444 252334 296056 252362
rect 291198 242312 291254 242321
rect 291198 242247 291254 242256
rect 293866 242312 293922 242321
rect 293866 242247 293922 242256
rect 289176 235068 289228 235074
rect 289176 235010 289228 235016
rect 291212 234025 291240 242247
rect 293880 234025 293908 242247
rect 291198 234016 291254 234025
rect 291198 233951 291254 233960
rect 293866 234016 293922 234025
rect 293866 233951 293922 233960
rect 295444 230450 295472 252334
rect 316776 251932 316828 251938
rect 316776 251874 316828 251880
rect 295708 235068 295760 235074
rect 295708 235010 295760 235016
rect 295720 232778 295748 235010
rect 316788 232778 316816 251874
rect 316868 251864 316920 251870
rect 316868 251806 316920 251812
rect 295720 232750 296056 232778
rect 316664 232750 316816 232778
rect 306300 232070 306360 232098
rect 295432 230444 295484 230450
rect 295432 230386 295484 230392
rect 306300 230314 306328 232070
rect 316880 230314 316908 251806
rect 316972 230382 317000 252606
rect 317064 251870 317092 255274
rect 317156 251938 317184 255342
rect 334360 252892 334388 255342
rect 344652 255332 344704 255338
rect 344652 255274 344704 255280
rect 352012 255332 352064 255338
rect 352012 255274 352064 255280
rect 344664 252892 344692 255274
rect 352024 252892 352052 255274
rect 361946 252648 362002 252657
rect 362002 252606 362342 252634
rect 372646 252606 372936 252634
rect 361946 252583 362002 252592
rect 323044 252334 324070 252362
rect 317144 251932 317196 251938
rect 317144 251874 317196 251880
rect 317052 251864 317104 251870
rect 317052 251806 317104 251812
rect 318798 242312 318854 242321
rect 318798 242247 318854 242256
rect 322846 242312 322902 242321
rect 322846 242247 322902 242256
rect 318812 233238 318840 242247
rect 322860 233238 322888 242247
rect 318800 233232 318852 233238
rect 318800 233174 318852 233180
rect 322848 233232 322900 233238
rect 322848 233174 322900 233180
rect 323044 230382 323072 252334
rect 372804 250164 372856 250170
rect 372804 250106 372856 250112
rect 346398 242312 346454 242321
rect 346398 242247 346454 242256
rect 350446 242312 350502 242321
rect 350446 242247 350502 242256
rect 346412 234025 346440 242247
rect 350460 234025 350488 242247
rect 346398 234016 346454 234025
rect 346398 233951 346454 233960
rect 350446 234016 350502 234025
rect 350446 233951 350502 233960
rect 372816 232778 372844 250106
rect 372646 232750 372844 232778
rect 324056 230450 324084 232084
rect 334360 230450 334388 232084
rect 344664 230489 344692 232084
rect 344650 230480 344706 230489
rect 324044 230444 324096 230450
rect 324044 230386 324096 230392
rect 334348 230444 334400 230450
rect 344650 230415 344706 230424
rect 334348 230386 334400 230392
rect 352024 230382 352052 232084
rect 362328 230382 362356 232084
rect 372908 230450 372936 252606
rect 373000 250170 373028 255342
rect 373264 255332 373316 255338
rect 373264 255274 373316 255280
rect 372988 250164 373040 250170
rect 372988 250106 373040 250112
rect 373276 235278 373304 255274
rect 375378 242312 375434 242321
rect 375378 242247 375434 242256
rect 378046 242312 378102 242321
rect 378046 242247 378102 242256
rect 373264 235272 373316 235278
rect 373264 235214 373316 235220
rect 375392 233238 375420 242247
rect 378060 233238 378088 242247
rect 375380 233232 375432 233238
rect 375380 233174 375432 233180
rect 378048 233232 378100 233238
rect 378048 233174 378100 233180
rect 372896 230444 372948 230450
rect 372896 230386 372948 230392
rect 316960 230376 317012 230382
rect 316960 230318 317012 230324
rect 323032 230376 323084 230382
rect 323032 230318 323084 230324
rect 352012 230376 352064 230382
rect 352012 230318 352064 230324
rect 362316 230376 362368 230382
rect 362316 230318 362368 230324
rect 250352 230308 250404 230314
rect 250352 230250 250404 230256
rect 288900 230308 288952 230314
rect 288900 230250 288952 230256
rect 306288 230308 306340 230314
rect 306288 230250 306340 230256
rect 316868 230308 316920 230314
rect 316868 230250 316920 230256
rect 250628 227860 250680 227866
rect 250628 227802 250680 227808
rect 261484 227860 261536 227866
rect 261484 227802 261536 227808
rect 278596 227860 278648 227866
rect 278596 227802 278648 227808
rect 295892 227860 295944 227866
rect 295892 227802 295944 227808
rect 334624 227860 334676 227866
rect 334624 227802 334676 227808
rect 240324 227792 240376 227798
rect 240324 227734 240376 227740
rect 240336 225964 240364 227734
rect 250640 225964 250668 227802
rect 260958 225270 261064 225298
rect 238666 224360 238722 224369
rect 238666 224295 238722 224304
rect 234710 224088 234766 224097
rect 234710 224023 234766 224032
rect 234724 215801 234752 224023
rect 238680 215801 238708 224295
rect 234710 215792 234766 215801
rect 234710 215727 234766 215736
rect 238666 215792 238722 215801
rect 238666 215727 238722 215736
rect 240336 202774 240364 205020
rect 240324 202768 240376 202774
rect 240324 202710 240376 202716
rect 250640 202706 250668 205020
rect 260944 202842 260972 205020
rect 261036 202842 261064 225270
rect 260932 202836 260984 202842
rect 260932 202778 260984 202784
rect 261024 202836 261076 202842
rect 261024 202778 261076 202784
rect 261496 202774 261524 227802
rect 267832 227792 267884 227798
rect 267832 227734 267884 227740
rect 266266 224088 266322 224097
rect 266266 224023 266322 224032
rect 266280 215801 266308 224023
rect 267740 222352 267792 222358
rect 267740 222294 267792 222300
rect 266266 215792 266322 215801
rect 266266 215727 266322 215736
rect 261484 202768 261536 202774
rect 261484 202710 261536 202716
rect 267752 202706 267780 222294
rect 267844 205714 267872 227734
rect 278608 225964 278636 227802
rect 267936 225270 268318 225298
rect 288926 225270 289124 225298
rect 267936 222358 267964 225270
rect 267924 222352 267976 222358
rect 267924 222294 267976 222300
rect 267844 205686 268318 205714
rect 278516 205006 278622 205034
rect 288544 205006 288926 205034
rect 278516 202774 278544 205006
rect 288544 202842 288572 205006
rect 289096 202842 289124 225270
rect 293868 225004 293920 225010
rect 293868 224946 293920 224952
rect 293880 215801 293908 224946
rect 295340 222352 295392 222358
rect 295340 222294 295392 222300
rect 293866 215792 293922 215801
rect 293866 215727 293922 215736
rect 288532 202836 288584 202842
rect 288532 202778 288584 202784
rect 289084 202836 289136 202842
rect 289084 202778 289136 202784
rect 295352 202774 295380 222294
rect 295904 205714 295932 227802
rect 306472 227792 306524 227798
rect 306472 227734 306524 227740
rect 318064 227792 318116 227798
rect 318064 227734 318116 227740
rect 324320 227792 324372 227798
rect 324320 227734 324372 227740
rect 306484 225978 306512 227734
rect 306484 225950 306636 225978
rect 295996 225270 296332 225298
rect 316940 225270 317092 225298
rect 295996 222358 296024 225270
rect 295984 222352 296036 222358
rect 295984 222294 296036 222300
rect 295904 205686 296332 205714
rect 306636 205006 306972 205034
rect 306944 202774 306972 205006
rect 316604 205006 316940 205034
rect 316604 202842 316632 205006
rect 317064 202842 317092 225270
rect 316592 202836 316644 202842
rect 316592 202778 316644 202784
rect 317052 202836 317104 202842
rect 317052 202778 317104 202784
rect 318076 202774 318104 227734
rect 324332 225964 324360 227734
rect 334636 225964 334664 227802
rect 345664 227792 345716 227798
rect 345664 227734 345716 227740
rect 362316 227792 362368 227798
rect 362316 227734 362368 227740
rect 344954 225282 345060 225298
rect 344954 225276 345072 225282
rect 344954 225270 345020 225276
rect 345020 225218 345072 225224
rect 322848 225072 322900 225078
rect 322848 225014 322900 225020
rect 318798 224088 318854 224097
rect 318798 224023 318854 224032
rect 318812 215801 318840 224023
rect 322860 215801 322888 225014
rect 318798 215792 318854 215801
rect 318798 215727 318854 215736
rect 322846 215792 322902 215801
rect 322846 215727 322902 215736
rect 324332 202774 324360 205020
rect 278504 202768 278556 202774
rect 278504 202710 278556 202716
rect 295340 202768 295392 202774
rect 295340 202710 295392 202716
rect 306932 202768 306984 202774
rect 306932 202710 306984 202716
rect 318064 202768 318116 202774
rect 318064 202710 318116 202716
rect 324320 202768 324372 202774
rect 324320 202710 324372 202716
rect 334636 202706 334664 205020
rect 344940 202842 344968 205020
rect 344928 202836 344980 202842
rect 344928 202778 344980 202784
rect 345676 202774 345704 227734
rect 362328 225978 362356 227734
rect 362328 225950 362664 225978
rect 347044 225276 347096 225282
rect 347044 225218 347096 225224
rect 352024 225270 352360 225298
rect 372968 225270 373120 225298
rect 346400 225004 346452 225010
rect 346400 224946 346452 224952
rect 346412 215801 346440 224946
rect 346398 215792 346454 215801
rect 346398 215727 346454 215736
rect 347056 202842 347084 225218
rect 352024 225010 352052 225270
rect 348424 225004 348476 225010
rect 348424 224946 348476 224952
rect 352012 225004 352064 225010
rect 352012 224946 352064 224952
rect 347044 202836 347096 202842
rect 347044 202778 347096 202784
rect 345664 202768 345716 202774
rect 345664 202710 345716 202716
rect 348436 202706 348464 224946
rect 350446 224088 350502 224097
rect 350446 224023 350502 224032
rect 350460 215801 350488 224023
rect 350446 215792 350502 215801
rect 350446 215727 350502 215736
rect 352360 205006 352696 205034
rect 362664 205006 362908 205034
rect 352668 202774 352696 205006
rect 352656 202768 352708 202774
rect 352656 202710 352708 202716
rect 362880 202706 362908 205006
rect 372632 205006 372968 205034
rect 372632 202842 372660 205006
rect 373092 202842 373120 225270
rect 375380 225072 375432 225078
rect 375380 225014 375432 225020
rect 375392 215801 375420 225014
rect 378046 224224 378102 224233
rect 378046 224159 378102 224168
rect 378060 215801 378088 224159
rect 375378 215792 375434 215801
rect 375378 215727 375434 215736
rect 378046 215792 378102 215801
rect 378046 215727 378102 215736
rect 372620 202836 372672 202842
rect 372620 202778 372672 202784
rect 373080 202836 373132 202842
rect 373080 202778 373132 202784
rect 250628 202700 250680 202706
rect 250628 202642 250680 202648
rect 267740 202700 267792 202706
rect 267740 202642 267792 202648
rect 334624 202700 334676 202706
rect 334624 202642 334676 202648
rect 348424 202700 348476 202706
rect 348424 202642 348476 202648
rect 362868 202700 362920 202706
rect 362868 202642 362920 202648
rect 261484 200252 261536 200258
rect 261484 200194 261536 200200
rect 278320 200252 278372 200258
rect 278320 200194 278372 200200
rect 288900 200252 288952 200258
rect 288900 200194 288952 200200
rect 306012 200252 306064 200258
rect 306012 200194 306064 200200
rect 316776 200252 316828 200258
rect 316776 200194 316828 200200
rect 334348 200252 334400 200258
rect 334348 200194 334400 200200
rect 372896 200252 372948 200258
rect 372896 200194 372948 200200
rect 250352 200184 250404 200190
rect 250352 200126 250404 200132
rect 250364 198900 250392 200126
rect 260378 198520 260434 198529
rect 260434 198478 260682 198506
rect 260378 198455 260434 198464
rect 238864 198206 240074 198234
rect 234710 196752 234766 196761
rect 234710 196687 234766 196696
rect 238666 196752 238722 196761
rect 238666 196687 238722 196696
rect 234724 188329 234752 196687
rect 238680 188329 238708 196687
rect 234710 188320 234766 188329
rect 234710 188255 234766 188264
rect 238666 188320 238722 188329
rect 238666 188255 238722 188264
rect 238864 176594 238892 198206
rect 261496 180794 261524 200194
rect 268016 200184 268068 200190
rect 268016 200126 268068 200132
rect 268028 198900 268056 200126
rect 278332 198900 278360 200194
rect 288650 198206 288848 198234
rect 262218 188320 262274 188329
rect 262218 188255 262274 188264
rect 266266 188320 266322 188329
rect 266266 188255 266322 188264
rect 261128 180766 261524 180794
rect 261128 178786 261156 180766
rect 262232 179382 262260 188255
rect 266280 179382 266308 188255
rect 262220 179376 262272 179382
rect 262220 179318 262272 179324
rect 266268 179376 266320 179382
rect 266268 179318 266320 179324
rect 288820 178906 288848 198206
rect 288808 178900 288860 178906
rect 288808 178842 288860 178848
rect 260682 178758 261156 178786
rect 288912 178514 288940 200194
rect 289084 200184 289136 200190
rect 289084 200126 289136 200132
rect 290464 200184 290516 200190
rect 290464 200126 290516 200132
rect 289096 182170 289124 200126
rect 289084 182164 289136 182170
rect 289084 182106 289136 182112
rect 288992 178900 289044 178906
rect 288992 178842 289044 178848
rect 288650 178486 288940 178514
rect 240060 176662 240088 178092
rect 240048 176656 240100 176662
rect 240048 176598 240100 176604
rect 238852 176588 238904 176594
rect 238852 176530 238904 176536
rect 250364 176526 250392 178092
rect 268028 176594 268056 178092
rect 278332 176594 278360 178092
rect 268016 176588 268068 176594
rect 268016 176530 268068 176536
rect 278320 176588 278372 176594
rect 278320 176530 278372 176536
rect 289004 176526 289032 178842
rect 290476 176594 290504 200126
rect 306024 198914 306052 200194
rect 316316 200184 316368 200190
rect 316316 200126 316368 200132
rect 316328 198914 316356 200126
rect 306024 198886 306360 198914
rect 316328 198886 316664 198914
rect 295444 198206 296056 198234
rect 291198 196752 291254 196761
rect 291198 196687 291254 196696
rect 293866 196752 293922 196761
rect 293866 196687 293922 196696
rect 291212 188329 291240 196687
rect 293880 188329 293908 196687
rect 291198 188320 291254 188329
rect 291198 188255 291254 188264
rect 293866 188320 293922 188329
rect 293866 188255 293922 188264
rect 295444 176662 295472 198206
rect 295708 182164 295760 182170
rect 295708 182106 295760 182112
rect 295720 178786 295748 182106
rect 316788 178786 316816 200194
rect 318064 200184 318116 200190
rect 318064 200126 318116 200132
rect 295720 178758 296056 178786
rect 316664 178758 316816 178786
rect 306300 178078 306360 178106
rect 295432 176656 295484 176662
rect 295432 176598 295484 176604
rect 306300 176594 306328 178078
rect 318076 176594 318104 200126
rect 334360 198900 334388 200194
rect 344652 200184 344704 200190
rect 344652 200126 344704 200132
rect 352012 200184 352064 200190
rect 352012 200126 352064 200132
rect 344664 198900 344692 200126
rect 352024 198900 352052 200126
rect 361946 198520 362002 198529
rect 362002 198478 362342 198506
rect 361946 198455 362002 198464
rect 323044 198206 324070 198234
rect 372646 198206 372844 198234
rect 318798 188320 318854 188329
rect 318798 188255 318854 188264
rect 322846 188320 322902 188329
rect 322846 188255 322902 188264
rect 318812 179382 318840 188255
rect 322860 179382 322888 188255
rect 318800 179376 318852 179382
rect 318800 179318 318852 179324
rect 322848 179376 322900 179382
rect 322848 179318 322900 179324
rect 323044 176594 323072 198206
rect 346398 196752 346454 196761
rect 346398 196687 346454 196696
rect 350446 196752 350502 196761
rect 350446 196687 350502 196696
rect 346412 188329 346440 196687
rect 350460 188329 350488 196687
rect 346398 188320 346454 188329
rect 346398 188255 346454 188264
rect 350446 188320 350502 188329
rect 350446 188255 350502 188264
rect 372816 178906 372844 198206
rect 372804 178900 372856 178906
rect 372804 178842 372856 178848
rect 372908 178514 372936 200194
rect 373264 200184 373316 200190
rect 373264 200126 373316 200132
rect 373276 181490 373304 200126
rect 375378 188320 375434 188329
rect 375378 188255 375434 188264
rect 378046 188320 378102 188329
rect 378046 188255 378102 188264
rect 373264 181484 373316 181490
rect 373264 181426 373316 181432
rect 375392 179382 375420 188255
rect 378060 179382 378088 188255
rect 375380 179376 375432 179382
rect 375380 179318 375432 179324
rect 378048 179376 378100 179382
rect 378048 179318 378100 179324
rect 372988 178900 373040 178906
rect 372988 178842 373040 178848
rect 372646 178486 372936 178514
rect 324056 176662 324084 178092
rect 334360 176662 334388 178092
rect 324044 176656 324096 176662
rect 324044 176598 324096 176604
rect 334348 176656 334400 176662
rect 344664 176633 344692 178092
rect 334348 176598 334400 176604
rect 344650 176624 344706 176633
rect 290464 176588 290516 176594
rect 290464 176530 290516 176536
rect 306288 176588 306340 176594
rect 306288 176530 306340 176536
rect 318064 176588 318116 176594
rect 318064 176530 318116 176536
rect 323032 176588 323084 176594
rect 352024 176594 352052 178092
rect 362328 176594 362356 178092
rect 373000 176662 373028 178842
rect 372988 176656 373040 176662
rect 372988 176598 373040 176604
rect 344650 176559 344706 176568
rect 352012 176588 352064 176594
rect 323032 176530 323084 176536
rect 352012 176530 352064 176536
rect 362316 176588 362368 176594
rect 362316 176530 362368 176536
rect 250352 176520 250404 176526
rect 250352 176462 250404 176468
rect 288992 176520 289044 176526
rect 288992 176462 289044 176468
rect 374644 174072 374696 174078
rect 374644 174014 374696 174020
rect 250628 174004 250680 174010
rect 250628 173946 250680 173952
rect 262864 174004 262916 174010
rect 262864 173946 262916 173952
rect 267832 174004 267884 174010
rect 267832 173946 267884 173952
rect 306472 174004 306524 174010
rect 306472 173946 306524 173952
rect 318064 174004 318116 174010
rect 318064 173946 318116 173952
rect 324320 174004 324372 174010
rect 324320 173946 324372 173952
rect 345848 174004 345900 174010
rect 345848 173946 345900 173952
rect 362316 174004 362368 174010
rect 362316 173946 362368 173952
rect 373264 174004 373316 174010
rect 373264 173946 373316 173952
rect 240324 173936 240376 173942
rect 240324 173878 240376 173884
rect 240336 171972 240364 173878
rect 250640 171972 250668 173946
rect 238668 171488 238720 171494
rect 238668 171430 238720 171436
rect 234710 170096 234766 170105
rect 234710 170031 234766 170040
rect 234724 161809 234752 170031
rect 238680 161809 238708 171430
rect 262220 171420 262272 171426
rect 262220 171362 262272 171368
rect 260958 171278 261064 171306
rect 234710 161800 234766 161809
rect 234710 161735 234766 161744
rect 238666 161800 238722 161809
rect 238666 161735 238722 161744
rect 240336 148986 240364 151028
rect 240324 148980 240376 148986
rect 240324 148922 240376 148928
rect 250640 148918 250668 151028
rect 260944 149054 260972 151028
rect 261036 149054 261064 171278
rect 262232 161809 262260 171362
rect 262218 161800 262274 161809
rect 262218 161735 262274 161744
rect 260932 149048 260984 149054
rect 260932 148990 260984 148996
rect 261024 149048 261076 149054
rect 261024 148990 261076 148996
rect 262876 148986 262904 173946
rect 264244 173936 264296 173942
rect 264244 173878 264296 173884
rect 262864 148980 262916 148986
rect 262864 148922 262916 148928
rect 264256 148918 264284 173878
rect 266266 170096 266322 170105
rect 266266 170031 266322 170040
rect 266280 161809 266308 170031
rect 266266 161800 266322 161809
rect 266266 161735 266322 161744
rect 267844 151722 267872 173946
rect 278596 173936 278648 173942
rect 278596 173878 278648 173884
rect 295340 173936 295392 173942
rect 295340 173878 295392 173884
rect 267924 173868 267976 173874
rect 267924 173810 267976 173816
rect 267936 171986 267964 173810
rect 267936 171958 268318 171986
rect 278608 171972 278636 173878
rect 291200 171488 291252 171494
rect 291200 171430 291252 171436
rect 288926 171278 289124 171306
rect 267844 151694 268318 151722
rect 278608 148986 278636 151028
rect 288912 149054 288940 151028
rect 289096 149054 289124 171278
rect 291212 161809 291240 171430
rect 293866 170232 293922 170241
rect 293866 170167 293922 170176
rect 293880 161809 293908 170167
rect 291198 161800 291254 161809
rect 291198 161735 291254 161744
rect 293866 161800 293922 161809
rect 293866 161735 293922 161744
rect 289176 153740 289228 153746
rect 289176 153682 289228 153688
rect 288900 149048 288952 149054
rect 288900 148990 288952 148996
rect 289084 149048 289136 149054
rect 289084 148990 289136 148996
rect 289188 148986 289216 153682
rect 295352 151814 295380 173878
rect 306484 171986 306512 173946
rect 306484 171958 306636 171986
rect 295444 171278 296332 171306
rect 316940 171278 317092 171306
rect 295444 153746 295472 171278
rect 295432 153740 295484 153746
rect 295432 153682 295484 153688
rect 295352 151786 295932 151814
rect 295904 151722 295932 151786
rect 295904 151694 296332 151722
rect 306636 151014 306972 151042
rect 306944 148986 306972 151014
rect 316604 151014 316940 151042
rect 316604 149054 316632 151014
rect 317064 149054 317092 171278
rect 316592 149048 316644 149054
rect 316592 148990 316644 148996
rect 317052 149048 317104 149054
rect 317052 148990 317104 148996
rect 318076 148986 318104 173946
rect 324332 171972 324360 173946
rect 334624 173936 334676 173942
rect 334624 173878 334676 173884
rect 345756 173936 345808 173942
rect 345756 173878 345808 173884
rect 334636 171972 334664 173878
rect 344954 171278 345152 171306
rect 345124 171134 345152 171278
rect 345124 171106 345704 171134
rect 322846 170368 322902 170377
rect 322846 170303 322902 170312
rect 318798 170096 318854 170105
rect 318798 170031 318854 170040
rect 318812 161809 318840 170031
rect 322860 161809 322888 170303
rect 318798 161800 318854 161809
rect 318798 161735 318854 161744
rect 322846 161800 322902 161809
rect 322846 161735 322902 161744
rect 324332 148986 324360 151028
rect 278596 148980 278648 148986
rect 278596 148922 278648 148928
rect 289176 148980 289228 148986
rect 289176 148922 289228 148928
rect 306932 148980 306984 148986
rect 306932 148922 306984 148928
rect 318064 148980 318116 148986
rect 318064 148922 318116 148928
rect 324320 148980 324372 148986
rect 324320 148922 324372 148928
rect 334636 148918 334664 151028
rect 344940 149054 344968 151028
rect 345676 149054 345704 171106
rect 344928 149048 344980 149054
rect 344928 148990 344980 148996
rect 345664 149048 345716 149054
rect 345664 148990 345716 148996
rect 345768 148918 345796 173878
rect 345860 148986 345888 173946
rect 352012 173936 352064 173942
rect 352012 173878 352064 173884
rect 352024 171986 352052 173878
rect 362328 171986 362356 173946
rect 352024 171958 352360 171986
rect 362328 171958 362664 171986
rect 372968 171278 373120 171306
rect 350446 170096 350502 170105
rect 350446 170031 350502 170040
rect 350460 161809 350488 170031
rect 350446 161800 350502 161809
rect 350446 161735 350502 161744
rect 352360 151014 352696 151042
rect 362664 151014 362908 151042
rect 352668 148986 352696 151014
rect 345848 148980 345900 148986
rect 345848 148922 345900 148928
rect 352656 148980 352708 148986
rect 352656 148922 352708 148928
rect 362880 148918 362908 151014
rect 372632 151014 372968 151042
rect 372632 149054 372660 151014
rect 373092 149054 373120 171278
rect 372620 149048 372672 149054
rect 372620 148990 372672 148996
rect 373080 149048 373132 149054
rect 373080 148990 373132 148996
rect 373276 148986 373304 173946
rect 373264 148980 373316 148986
rect 373264 148922 373316 148928
rect 374656 148918 374684 174014
rect 378046 170232 378102 170241
rect 378046 170167 378102 170176
rect 378060 161809 378088 170167
rect 378046 161800 378102 161809
rect 378046 161735 378102 161744
rect 250628 148912 250680 148918
rect 250628 148854 250680 148860
rect 264244 148912 264296 148918
rect 264244 148854 264296 148860
rect 334624 148912 334676 148918
rect 334624 148854 334676 148860
rect 345756 148912 345808 148918
rect 345756 148854 345808 148860
rect 362868 148912 362920 148918
rect 362868 148854 362920 148860
rect 374644 148912 374696 148918
rect 374644 148854 374696 148860
rect 268016 146532 268068 146538
rect 268016 146474 268068 146480
rect 289084 146532 289136 146538
rect 289084 146474 289136 146480
rect 262864 146464 262916 146470
rect 262864 146406 262916 146412
rect 250352 146396 250404 146402
rect 250352 146338 250404 146344
rect 250364 144908 250392 146338
rect 260656 146328 260708 146334
rect 260656 146270 260708 146276
rect 261484 146328 261536 146334
rect 261484 146270 261536 146276
rect 260668 144908 260696 146270
rect 238864 144214 240074 144242
rect 234712 143608 234764 143614
rect 234712 143550 234764 143556
rect 234724 134337 234752 143550
rect 234710 134328 234766 134337
rect 234710 134263 234766 134272
rect 238666 134328 238722 134337
rect 238666 134263 238722 134272
rect 238680 125594 238708 134263
rect 238668 125588 238720 125594
rect 238668 125530 238720 125536
rect 238864 122670 238892 144214
rect 240060 122806 240088 124100
rect 240048 122800 240100 122806
rect 240048 122742 240100 122748
rect 250364 122738 250392 124100
rect 260668 122806 260696 124100
rect 260656 122800 260708 122806
rect 260656 122742 260708 122748
rect 261496 122738 261524 146270
rect 262218 142760 262274 142769
rect 262218 142695 262274 142704
rect 262232 134337 262260 142695
rect 262218 134328 262274 134337
rect 262218 134263 262274 134272
rect 262876 122806 262904 146406
rect 268028 144908 268056 146474
rect 278320 146464 278372 146470
rect 278320 146406 278372 146412
rect 278332 144908 278360 146406
rect 288808 146396 288860 146402
rect 288808 146338 288860 146344
rect 288624 146328 288676 146334
rect 288624 146270 288676 146276
rect 288636 144908 288664 146270
rect 266266 142760 266322 142769
rect 266266 142695 266322 142704
rect 266280 134337 266308 142695
rect 266266 134328 266322 134337
rect 266266 134263 266322 134272
rect 288820 124794 288848 146338
rect 289096 128042 289124 146474
rect 306012 146396 306064 146402
rect 306012 146338 306064 146344
rect 316776 146396 316828 146402
rect 316776 146338 316828 146344
rect 334348 146396 334400 146402
rect 334348 146338 334400 146344
rect 372896 146396 372948 146402
rect 372896 146338 372948 146344
rect 290464 146328 290516 146334
rect 290464 146270 290516 146276
rect 289084 128036 289136 128042
rect 289084 127978 289136 127984
rect 288650 124766 288848 124794
rect 262864 122800 262916 122806
rect 262864 122742 262916 122748
rect 250352 122732 250404 122738
rect 250352 122674 250404 122680
rect 261484 122732 261536 122738
rect 261484 122674 261536 122680
rect 268028 122670 268056 124100
rect 278332 122806 278360 124100
rect 290476 122806 290504 146270
rect 306024 144922 306052 146338
rect 316316 146328 316368 146334
rect 316316 146270 316368 146276
rect 316328 144922 316356 146270
rect 306024 144894 306360 144922
rect 316328 144894 316664 144922
rect 295444 144214 296056 144242
rect 291198 134328 291254 134337
rect 291198 134263 291254 134272
rect 293866 134328 293922 134337
rect 293866 134263 293922 134272
rect 291212 125594 291240 134263
rect 293880 125594 293908 134263
rect 291200 125588 291252 125594
rect 291200 125530 291252 125536
rect 293868 125588 293920 125594
rect 293868 125530 293920 125536
rect 295444 122806 295472 144214
rect 295708 128036 295760 128042
rect 295708 127978 295760 127984
rect 295720 124794 295748 127978
rect 316788 124794 316816 146338
rect 316868 146328 316920 146334
rect 316868 146270 316920 146276
rect 295720 124766 296056 124794
rect 316664 124766 316816 124794
rect 306300 124086 306360 124114
rect 278320 122800 278372 122806
rect 278320 122742 278372 122748
rect 290464 122800 290516 122806
rect 290464 122742 290516 122748
rect 295432 122800 295484 122806
rect 295432 122742 295484 122748
rect 306300 122738 306328 124086
rect 316880 122738 316908 146270
rect 334360 144908 334388 146338
rect 344652 146328 344704 146334
rect 344652 146270 344704 146276
rect 352012 146328 352064 146334
rect 352012 146270 352064 146276
rect 344664 144908 344692 146270
rect 352024 144908 352052 146270
rect 361946 144528 362002 144537
rect 362002 144486 362342 144514
rect 361946 144463 362002 144472
rect 323044 144214 324070 144242
rect 372646 144214 372844 144242
rect 318798 142760 318854 142769
rect 318798 142695 318854 142704
rect 322846 142760 322902 142769
rect 322846 142695 322902 142704
rect 318812 134337 318840 142695
rect 322860 134337 322888 142695
rect 318798 134328 318854 134337
rect 318798 134263 318854 134272
rect 322846 134328 322902 134337
rect 322846 134263 322902 134272
rect 323044 122738 323072 144214
rect 346398 134328 346454 134337
rect 346398 134263 346454 134272
rect 350446 134328 350502 134337
rect 350446 134263 350502 134272
rect 346412 125594 346440 134263
rect 350460 125594 350488 134263
rect 346400 125588 346452 125594
rect 346400 125530 346452 125536
rect 350448 125588 350500 125594
rect 350448 125530 350500 125536
rect 372816 124914 372844 144214
rect 372804 124908 372856 124914
rect 372804 124850 372856 124856
rect 372908 124794 372936 146338
rect 373264 146328 373316 146334
rect 373264 146270 373316 146276
rect 373276 127634 373304 146270
rect 375378 142760 375434 142769
rect 375378 142695 375434 142704
rect 378046 142760 378102 142769
rect 378046 142695 378102 142704
rect 375392 134337 375420 142695
rect 378060 134337 378088 142695
rect 375378 134328 375434 134337
rect 375378 134263 375434 134272
rect 378046 134328 378102 134337
rect 378046 134263 378102 134272
rect 373264 127628 373316 127634
rect 373264 127570 373316 127576
rect 372646 124766 372936 124794
rect 372804 124704 372856 124710
rect 372804 124646 372856 124652
rect 324056 122806 324084 124100
rect 334360 122806 334388 124100
rect 324044 122800 324096 122806
rect 324044 122742 324096 122748
rect 334348 122800 334400 122806
rect 344664 122777 344692 124100
rect 334348 122742 334400 122748
rect 344650 122768 344706 122777
rect 306288 122732 306340 122738
rect 306288 122674 306340 122680
rect 316868 122732 316920 122738
rect 316868 122674 316920 122680
rect 323032 122732 323084 122738
rect 352024 122738 352052 124100
rect 362328 122738 362356 124100
rect 372816 122806 372844 124646
rect 372804 122800 372856 122806
rect 372804 122742 372856 122748
rect 344650 122703 344706 122712
rect 352012 122732 352064 122738
rect 323032 122674 323084 122680
rect 352012 122674 352064 122680
rect 362316 122732 362368 122738
rect 362316 122674 362368 122680
rect 238852 122664 238904 122670
rect 238852 122606 238904 122612
rect 268016 122664 268068 122670
rect 268016 122606 268068 122612
rect 250628 120284 250680 120290
rect 250628 120226 250680 120232
rect 295432 120284 295484 120290
rect 295432 120226 295484 120232
rect 240324 120148 240376 120154
rect 240324 120090 240376 120096
rect 240336 117980 240364 120090
rect 250640 117980 250668 120226
rect 262864 120216 262916 120222
rect 262864 120158 262916 120164
rect 278228 120216 278280 120222
rect 278228 120158 278280 120164
rect 290464 120216 290516 120222
rect 290464 120158 290516 120164
rect 238668 117360 238720 117366
rect 238668 117302 238720 117308
rect 234710 116376 234766 116385
rect 234710 116311 234766 116320
rect 234724 107817 234752 116311
rect 238680 107817 238708 117302
rect 260958 117286 261064 117314
rect 234710 107808 234766 107817
rect 234710 107743 234766 107752
rect 238666 107808 238722 107817
rect 238666 107743 238722 107752
rect 240336 95130 240364 97036
rect 240324 95124 240376 95130
rect 240324 95066 240376 95072
rect 250640 95062 250668 97036
rect 260944 95198 260972 97036
rect 261036 95198 261064 117286
rect 260932 95192 260984 95198
rect 260932 95134 260984 95140
rect 261024 95192 261076 95198
rect 261024 95134 261076 95140
rect 262876 95130 262904 120158
rect 267832 120148 267884 120154
rect 267832 120090 267884 120096
rect 264244 117292 264296 117298
rect 264244 117234 264296 117240
rect 262864 95124 262916 95130
rect 262864 95066 262916 95072
rect 264256 95062 264284 117234
rect 266266 116104 266322 116113
rect 266266 116039 266322 116048
rect 266280 107817 266308 116039
rect 266266 107808 266322 107817
rect 266266 107743 266322 107752
rect 267844 97730 267872 120090
rect 278240 117994 278268 120158
rect 278240 117966 278622 117994
rect 267936 117298 268318 117314
rect 267924 117292 268318 117298
rect 267976 117286 268318 117292
rect 288926 117286 289124 117314
rect 267924 117234 267976 117240
rect 267844 97702 268318 97730
rect 278608 95130 278636 97036
rect 288912 95198 288940 97036
rect 289096 95198 289124 117286
rect 288900 95192 288952 95198
rect 288900 95134 288952 95140
rect 289084 95192 289136 95198
rect 289084 95134 289136 95140
rect 290476 95130 290504 120158
rect 293868 117428 293920 117434
rect 293868 117370 293920 117376
rect 291200 117360 291252 117366
rect 291200 117302 291252 117308
rect 291212 107817 291240 117302
rect 293880 107817 293908 117370
rect 295444 113174 295472 120226
rect 295984 120216 296036 120222
rect 295984 120158 296036 120164
rect 334624 120216 334676 120222
rect 334624 120158 334676 120164
rect 295996 117994 296024 120158
rect 306472 120148 306524 120154
rect 306472 120090 306524 120096
rect 306484 117994 306512 120090
rect 295996 117966 296332 117994
rect 306484 117966 306636 117994
rect 334636 117980 334664 120158
rect 345664 120148 345716 120154
rect 345664 120090 345716 120096
rect 362316 120148 362368 120154
rect 362316 120090 362368 120096
rect 322848 117360 322900 117366
rect 316940 117286 318104 117314
rect 322848 117302 322900 117308
rect 324226 117328 324282 117337
rect 295444 113146 295932 113174
rect 291198 107808 291254 107817
rect 291198 107743 291254 107752
rect 293866 107808 293922 107817
rect 293866 107743 293922 107752
rect 295904 97730 295932 113146
rect 295904 97702 296332 97730
rect 306636 97022 306972 97050
rect 306944 95169 306972 97022
rect 316604 97022 316940 97050
rect 316604 95198 316632 97022
rect 318076 95198 318104 117286
rect 318798 116104 318854 116113
rect 318798 116039 318854 116048
rect 318812 107817 318840 116039
rect 322860 107817 322888 117302
rect 324282 117286 324346 117314
rect 344954 117298 345060 117314
rect 344954 117292 345072 117298
rect 344954 117286 345020 117292
rect 324226 117263 324282 117272
rect 345020 117234 345072 117240
rect 318798 107808 318854 107817
rect 318798 107743 318854 107752
rect 322846 107808 322902 107817
rect 322846 107743 322902 107752
rect 316592 95192 316644 95198
rect 306930 95160 306986 95169
rect 278596 95124 278648 95130
rect 278596 95066 278648 95072
rect 290464 95124 290516 95130
rect 316592 95134 316644 95140
rect 318064 95192 318116 95198
rect 318064 95134 318116 95140
rect 324332 95130 324360 97036
rect 306930 95095 306986 95104
rect 324320 95124 324372 95130
rect 290464 95066 290516 95072
rect 324320 95066 324372 95072
rect 334636 95062 334664 97036
rect 344940 95198 344968 97036
rect 344928 95192 344980 95198
rect 344928 95134 344980 95140
rect 345676 95130 345704 120090
rect 362328 117994 362356 120090
rect 362328 117966 362664 117994
rect 346400 117428 346452 117434
rect 346400 117370 346452 117376
rect 346412 107817 346440 117370
rect 375380 117360 375432 117366
rect 352024 117298 352360 117314
rect 347044 117292 347096 117298
rect 347044 117234 347096 117240
rect 348424 117292 348476 117298
rect 348424 117234 348476 117240
rect 352012 117292 352360 117298
rect 352064 117286 352360 117292
rect 372968 117286 373120 117314
rect 375380 117302 375432 117308
rect 352012 117234 352064 117240
rect 346398 107808 346454 107817
rect 346398 107743 346454 107752
rect 347056 95198 347084 117234
rect 347044 95192 347096 95198
rect 347044 95134 347096 95140
rect 345664 95124 345716 95130
rect 345664 95066 345716 95072
rect 348436 95062 348464 117234
rect 350446 116104 350502 116113
rect 350446 116039 350502 116048
rect 350460 107817 350488 116039
rect 350446 107808 350502 107817
rect 350446 107743 350502 107752
rect 352360 97022 352696 97050
rect 362664 97022 362908 97050
rect 352668 95130 352696 97022
rect 352656 95124 352708 95130
rect 352656 95066 352708 95072
rect 362880 95062 362908 97022
rect 372632 97022 372968 97050
rect 372632 95198 372660 97022
rect 373092 95198 373120 117286
rect 375392 107817 375420 117302
rect 378046 116240 378102 116249
rect 378046 116175 378102 116184
rect 378060 107817 378088 116175
rect 375378 107808 375434 107817
rect 375378 107743 375434 107752
rect 378046 107808 378102 107817
rect 378046 107743 378102 107752
rect 372620 95192 372672 95198
rect 372620 95134 372672 95140
rect 373080 95192 373132 95198
rect 373080 95134 373132 95140
rect 250628 95056 250680 95062
rect 250628 94998 250680 95004
rect 264244 95056 264296 95062
rect 264244 94998 264296 95004
rect 334624 95056 334676 95062
rect 334624 94998 334676 95004
rect 348424 95056 348476 95062
rect 348424 94998 348476 95004
rect 362868 95056 362920 95062
rect 362868 94998 362920 95004
rect 268016 92744 268068 92750
rect 268016 92686 268068 92692
rect 289084 92744 289136 92750
rect 289084 92686 289136 92692
rect 261576 92676 261628 92682
rect 261576 92618 261628 92624
rect 250352 92608 250404 92614
rect 250352 92550 250404 92556
rect 250364 90916 250392 92550
rect 260656 92540 260708 92546
rect 260656 92482 260708 92488
rect 261484 92540 261536 92546
rect 261484 92482 261536 92488
rect 260668 90916 260696 92482
rect 238864 90222 240074 90250
rect 238666 88904 238722 88913
rect 238666 88839 238722 88848
rect 234710 88768 234766 88777
rect 234710 88703 234766 88712
rect 234724 80345 234752 88703
rect 238680 80345 238708 88839
rect 234710 80336 234766 80345
rect 234710 80271 234766 80280
rect 238666 80336 238722 80345
rect 238666 80271 238722 80280
rect 238864 68882 238892 90222
rect 261024 72344 261076 72350
rect 261024 72286 261076 72292
rect 261036 70666 261064 72286
rect 260682 70638 261064 70666
rect 240060 69018 240088 70108
rect 240048 69012 240100 69018
rect 240048 68954 240100 68960
rect 250364 68950 250392 70108
rect 261496 68950 261524 92482
rect 261588 72350 261616 92618
rect 268028 90916 268056 92686
rect 278320 92676 278372 92682
rect 278320 92618 278372 92624
rect 278332 90916 278360 92618
rect 288808 92608 288860 92614
rect 288808 92550 288860 92556
rect 288624 92540 288676 92546
rect 288624 92482 288676 92488
rect 288636 90916 288664 92482
rect 262220 89752 262272 89758
rect 262220 89694 262272 89700
rect 262232 80345 262260 89694
rect 266266 88768 266322 88777
rect 266266 88703 266322 88712
rect 266280 80345 266308 88703
rect 262218 80336 262274 80345
rect 262218 80271 262274 80280
rect 266266 80336 266322 80345
rect 266266 80271 266322 80280
rect 261576 72344 261628 72350
rect 261576 72286 261628 72292
rect 288820 70666 288848 92550
rect 289096 73234 289124 92686
rect 345756 92676 345808 92682
rect 345756 92618 345808 92624
rect 362316 92676 362368 92682
rect 362316 92618 362368 92624
rect 372804 92676 372856 92682
rect 372804 92618 372856 92624
rect 306012 92608 306064 92614
rect 306012 92550 306064 92556
rect 316776 92608 316828 92614
rect 316776 92550 316828 92556
rect 334348 92608 334400 92614
rect 334348 92550 334400 92556
rect 290464 92540 290516 92546
rect 290464 92482 290516 92488
rect 289084 73228 289136 73234
rect 289084 73170 289136 73176
rect 288650 70638 288848 70666
rect 250352 68944 250404 68950
rect 250352 68886 250404 68892
rect 261484 68944 261536 68950
rect 261484 68886 261536 68892
rect 268028 68882 268056 70108
rect 278332 69018 278360 70108
rect 290476 69018 290504 92482
rect 306024 90930 306052 92550
rect 316316 92540 316368 92546
rect 316316 92482 316368 92488
rect 316328 90930 316356 92482
rect 306024 90902 306360 90930
rect 316328 90902 316664 90930
rect 295444 90222 296056 90250
rect 295444 69018 295472 90222
rect 295708 73228 295760 73234
rect 295708 73170 295760 73176
rect 295720 70666 295748 73170
rect 316788 70666 316816 92550
rect 316868 92540 316920 92546
rect 316868 92482 316920 92488
rect 295720 70638 296056 70666
rect 316664 70638 316816 70666
rect 306300 70094 306360 70122
rect 278320 69012 278372 69018
rect 278320 68954 278372 68960
rect 290464 69012 290516 69018
rect 290464 68954 290516 68960
rect 295432 69012 295484 69018
rect 295432 68954 295484 68960
rect 306300 68950 306328 70094
rect 316880 68950 316908 92482
rect 334360 90916 334388 92550
rect 344652 92540 344704 92546
rect 344652 92482 344704 92488
rect 345664 92540 345716 92546
rect 345664 92482 345716 92488
rect 344664 90916 344692 92482
rect 323044 90222 324070 90250
rect 322846 89040 322902 89049
rect 322846 88975 322902 88984
rect 318798 88768 318854 88777
rect 318798 88703 318854 88712
rect 318812 80345 318840 88703
rect 322860 80345 322888 88975
rect 318798 80336 318854 80345
rect 318798 80271 318854 80280
rect 322846 80336 322902 80345
rect 322846 80271 322902 80280
rect 306288 68944 306340 68950
rect 306288 68886 306340 68892
rect 316868 68944 316920 68950
rect 316868 68886 316920 68892
rect 323044 68882 323072 90222
rect 344928 71732 344980 71738
rect 344928 71674 344980 71680
rect 344940 70666 344968 71674
rect 344678 70638 344968 70666
rect 324056 69018 324084 70108
rect 324044 69012 324096 69018
rect 324044 68954 324096 68960
rect 334360 68950 334388 70108
rect 345676 68950 345704 92482
rect 345768 71738 345796 92618
rect 352012 92608 352064 92614
rect 352012 92550 352064 92556
rect 352024 90916 352052 92550
rect 362328 90916 362356 92618
rect 372620 92540 372672 92546
rect 372620 92482 372672 92488
rect 372632 90916 372660 92482
rect 346398 88904 346454 88913
rect 346398 88839 346454 88848
rect 346412 80345 346440 88839
rect 350446 88768 350502 88777
rect 350446 88703 350502 88712
rect 350460 80345 350488 88703
rect 346398 80336 346454 80345
rect 346398 80271 346454 80280
rect 350446 80336 350502 80345
rect 350446 80271 350502 80280
rect 345756 71732 345808 71738
rect 345756 71674 345808 71680
rect 372816 70666 372844 92618
rect 376024 92608 376076 92614
rect 376024 92550 376076 92556
rect 374644 92540 374696 92546
rect 374644 92482 374696 92488
rect 372646 70638 372844 70666
rect 334348 68944 334400 68950
rect 334348 68886 334400 68892
rect 345664 68944 345716 68950
rect 345664 68886 345716 68892
rect 352024 68882 352052 70108
rect 362328 69018 362356 70108
rect 374656 69018 374684 92482
rect 376036 69018 376064 92550
rect 378046 88904 378102 88913
rect 378046 88839 378102 88848
rect 378060 80345 378088 88839
rect 378046 80336 378102 80345
rect 378046 80271 378102 80280
rect 362316 69012 362368 69018
rect 362316 68954 362368 68960
rect 374644 69012 374696 69018
rect 374644 68954 374696 68960
rect 376024 69012 376076 69018
rect 376024 68954 376076 68960
rect 238852 68876 238904 68882
rect 238852 68818 238904 68824
rect 268016 68876 268068 68882
rect 268016 68818 268068 68824
rect 323032 68876 323084 68882
rect 323032 68818 323084 68824
rect 352012 68876 352064 68882
rect 352012 68818 352064 68824
rect 250628 66428 250680 66434
rect 250628 66370 250680 66376
rect 345664 66428 345716 66434
rect 345664 66370 345716 66376
rect 362316 66428 362368 66434
rect 362316 66370 362368 66376
rect 374644 66428 374696 66434
rect 374644 66370 374696 66376
rect 240324 66292 240376 66298
rect 240324 66234 240376 66240
rect 240336 63852 240364 66234
rect 250640 63852 250668 66370
rect 267832 66360 267884 66366
rect 267832 66302 267884 66308
rect 306380 66360 306432 66366
rect 306380 66302 306432 66308
rect 318064 66360 318116 66366
rect 318064 66302 318116 66308
rect 324320 66360 324372 66366
rect 324320 66302 324372 66308
rect 261484 66292 261536 66298
rect 261484 66234 261536 66240
rect 260958 63294 261064 63322
rect 234710 53816 234766 53825
rect 234710 53751 234766 53760
rect 238666 53816 238722 53825
rect 238666 53751 238722 53760
rect 234724 45393 234752 53751
rect 234710 45384 234766 45393
rect 234710 45319 234766 45328
rect 238680 45121 238708 53751
rect 238666 45112 238722 45121
rect 238666 45047 238722 45056
rect 240336 41342 240364 43044
rect 240324 41336 240376 41342
rect 240324 41278 240376 41284
rect 250640 41274 250668 43044
rect 260944 41410 260972 43044
rect 261036 41410 261064 63294
rect 260932 41404 260984 41410
rect 260932 41346 260984 41352
rect 261024 41404 261076 41410
rect 261024 41346 261076 41352
rect 261496 41342 261524 66234
rect 261576 60784 261628 60790
rect 261576 60726 261628 60732
rect 261484 41336 261536 41342
rect 261484 41278 261536 41284
rect 261588 41274 261616 60726
rect 266266 53816 266322 53825
rect 266266 53751 266322 53760
rect 266280 45393 266308 53751
rect 266266 45384 266322 45393
rect 266266 45319 266322 45328
rect 267844 43738 267872 66302
rect 278596 66292 278648 66298
rect 278596 66234 278648 66240
rect 295432 66292 295484 66298
rect 295432 66234 295484 66240
rect 278608 63852 278636 66234
rect 267936 63294 268318 63322
rect 288926 63294 289124 63322
rect 267936 60790 267964 63294
rect 267924 60784 267976 60790
rect 267924 60726 267976 60732
rect 267844 43710 268318 43738
rect 278608 41342 278636 43044
rect 288912 41410 288940 43044
rect 289096 41410 289124 63294
rect 289176 60784 289228 60790
rect 289176 60726 289228 60732
rect 288900 41404 288952 41410
rect 288900 41346 288952 41352
rect 289084 41404 289136 41410
rect 289084 41346 289136 41352
rect 289188 41342 289216 60726
rect 295444 55214 295472 66234
rect 306392 63866 306420 66302
rect 306392 63838 306636 63866
rect 295996 63294 296332 63322
rect 316940 63294 317092 63322
rect 295996 60790 296024 63294
rect 295984 60784 296036 60790
rect 295984 60726 296036 60732
rect 295444 55186 295932 55214
rect 293866 53816 293922 53825
rect 293866 53751 293922 53760
rect 293880 45257 293908 53751
rect 293866 45248 293922 45257
rect 293866 45183 293922 45192
rect 295904 43738 295932 55186
rect 295904 43710 296332 43738
rect 306636 43030 306972 43058
rect 306944 41342 306972 43030
rect 316604 43030 316940 43058
rect 316604 41410 316632 43030
rect 317064 41410 317092 63294
rect 316592 41404 316644 41410
rect 316592 41346 316644 41352
rect 317052 41404 317104 41410
rect 317052 41346 317104 41352
rect 318076 41342 318104 66302
rect 324332 63852 324360 66302
rect 334624 66292 334676 66298
rect 334624 66234 334676 66240
rect 334636 63852 334664 66234
rect 344954 63306 345060 63322
rect 344954 63300 345072 63306
rect 344954 63294 345020 63300
rect 345020 63242 345072 63248
rect 318798 53816 318854 53825
rect 318798 53751 318854 53760
rect 322846 53816 322902 53825
rect 322846 53751 322902 53760
rect 318812 45393 318840 53751
rect 318798 45384 318854 45393
rect 318798 45319 318854 45328
rect 322860 45121 322888 53751
rect 322846 45112 322902 45121
rect 322846 45047 322902 45056
rect 324332 41342 324360 43044
rect 278596 41336 278648 41342
rect 278596 41278 278648 41284
rect 289176 41336 289228 41342
rect 289176 41278 289228 41284
rect 306932 41336 306984 41342
rect 306932 41278 306984 41284
rect 318064 41336 318116 41342
rect 318064 41278 318116 41284
rect 324320 41336 324372 41342
rect 324320 41278 324372 41284
rect 334636 41274 334664 43044
rect 344940 41410 344968 43044
rect 344928 41404 344980 41410
rect 344928 41346 344980 41352
rect 345676 41342 345704 66370
rect 362328 63866 362356 66370
rect 373264 66360 373316 66366
rect 373264 66302 373316 66308
rect 362328 63838 362664 63866
rect 352024 63578 352360 63594
rect 348424 63572 348476 63578
rect 348424 63514 348476 63520
rect 352012 63572 352360 63578
rect 352064 63566 352360 63572
rect 352012 63514 352064 63520
rect 347044 63300 347096 63306
rect 347044 63242 347096 63248
rect 347056 41410 347084 63242
rect 347044 41404 347096 41410
rect 347044 41346 347096 41352
rect 345664 41336 345716 41342
rect 345664 41278 345716 41284
rect 348436 41274 348464 63514
rect 372968 63294 373120 63322
rect 350446 53816 350502 53825
rect 350446 53751 350502 53760
rect 350460 45393 350488 53751
rect 350446 45384 350502 45393
rect 350446 45319 350502 45328
rect 352360 43030 352696 43058
rect 362664 43030 362908 43058
rect 352668 41342 352696 43030
rect 352656 41336 352708 41342
rect 352656 41278 352708 41284
rect 362880 41274 362908 43030
rect 372632 43030 372968 43058
rect 372632 41410 372660 43030
rect 373092 41410 373120 63294
rect 372620 41404 372672 41410
rect 372620 41346 372672 41352
rect 373080 41404 373132 41410
rect 373080 41346 373132 41352
rect 373276 41342 373304 66302
rect 373264 41336 373316 41342
rect 373264 41278 373316 41284
rect 374656 41274 374684 66370
rect 378046 53816 378102 53825
rect 378046 53751 378102 53760
rect 378060 45257 378088 53751
rect 378046 45248 378102 45257
rect 378046 45183 378102 45192
rect 250628 41268 250680 41274
rect 250628 41210 250680 41216
rect 261576 41268 261628 41274
rect 261576 41210 261628 41216
rect 334624 41268 334676 41274
rect 334624 41210 334676 41216
rect 348424 41268 348476 41274
rect 348424 41210 348476 41216
rect 362868 41268 362920 41274
rect 362868 41210 362920 41216
rect 374644 41268 374696 41274
rect 374644 41210 374696 41216
rect 352012 38888 352064 38894
rect 352012 38830 352064 38836
rect 373264 38888 373316 38894
rect 373264 38830 373316 38836
rect 268016 38820 268068 38826
rect 268016 38762 268068 38768
rect 289084 38820 289136 38826
rect 289084 38762 289136 38768
rect 345664 38820 345716 38826
rect 345664 38762 345716 38768
rect 261484 38752 261536 38758
rect 261484 38694 261536 38700
rect 260656 38684 260708 38690
rect 260656 38626 260708 38632
rect 234620 38344 234672 38350
rect 234620 38286 234672 38292
rect 260668 36924 260696 38626
rect 250074 36544 250130 36553
rect 250130 36502 250378 36530
rect 250074 36479 250130 36488
rect 238864 36230 240074 36258
rect 234618 34912 234674 34921
rect 234618 34847 234674 34856
rect 234632 26353 234660 34847
rect 234618 26344 234674 26353
rect 234618 26279 234674 26288
rect 233976 13796 234028 13802
rect 233976 13738 234028 13744
rect 238864 13258 238892 36230
rect 261496 16574 261524 38694
rect 268028 36924 268056 38762
rect 278320 38752 278372 38758
rect 278320 38694 278372 38700
rect 278332 36924 278360 38694
rect 288900 38684 288952 38690
rect 288900 38626 288952 38632
rect 288650 36230 288848 36258
rect 262218 34776 262274 34785
rect 262218 34711 262274 34720
rect 266266 34776 266322 34785
rect 266266 34711 266322 34720
rect 262232 26353 262260 34711
rect 266280 26353 266308 34711
rect 262218 26344 262274 26353
rect 262218 26279 262274 26288
rect 266266 26344 266322 26353
rect 266266 26279 266322 26288
rect 288532 16720 288584 16726
rect 288584 16668 288650 16674
rect 288532 16662 288650 16668
rect 288544 16646 288650 16662
rect 261128 16546 261524 16574
rect 261128 16538 261156 16546
rect 260682 16510 261156 16538
rect 232780 13252 232832 13258
rect 232780 13194 232832 13200
rect 238852 13252 238904 13258
rect 238852 13194 238904 13200
rect 240060 13190 240088 16116
rect 250364 13258 250392 16116
rect 250352 13252 250404 13258
rect 250352 13194 250404 13200
rect 268028 13190 268056 16116
rect 278332 13190 278360 16116
rect 288820 13258 288848 36230
rect 288912 16726 288940 38626
rect 289096 18698 289124 38762
rect 317144 38752 317196 38758
rect 317144 38694 317196 38700
rect 334348 38752 334400 38758
rect 334348 38694 334400 38700
rect 306012 38684 306064 38690
rect 306012 38626 306064 38632
rect 317052 38684 317104 38690
rect 317052 38626 317104 38632
rect 306024 36938 306052 38626
rect 306024 36910 306360 36938
rect 316664 36502 317000 36530
rect 295444 36230 296056 36258
rect 316868 36236 316920 36242
rect 291198 34912 291254 34921
rect 291198 34847 291254 34856
rect 291212 26353 291240 34847
rect 291198 26344 291254 26353
rect 291198 26279 291254 26288
rect 289084 18692 289136 18698
rect 289084 18634 289136 18640
rect 288900 16720 288952 16726
rect 288900 16662 288952 16668
rect 295444 13258 295472 36230
rect 316868 36178 316920 36184
rect 316776 36168 316828 36174
rect 316776 36110 316828 36116
rect 295708 18692 295760 18698
rect 295708 18634 295760 18640
rect 295720 16674 295748 18634
rect 316788 16674 316816 36110
rect 295720 16646 296056 16674
rect 316664 16646 316816 16674
rect 306300 16102 306360 16130
rect 306300 13802 306328 16102
rect 316880 13802 316908 36178
rect 306288 13796 306340 13802
rect 306288 13738 306340 13744
rect 316868 13796 316920 13802
rect 316868 13738 316920 13744
rect 288808 13252 288860 13258
rect 288808 13194 288860 13200
rect 295432 13252 295484 13258
rect 295432 13194 295484 13200
rect 316972 13190 317000 36502
rect 317064 36242 317092 38626
rect 317052 36236 317104 36242
rect 317052 36178 317104 36184
rect 317156 36174 317184 38694
rect 334360 36924 334388 38694
rect 344652 38684 344704 38690
rect 344652 38626 344704 38632
rect 344664 36924 344692 38626
rect 323044 36230 324070 36258
rect 317144 36168 317196 36174
rect 317144 36110 317196 36116
rect 318798 34776 318854 34785
rect 318798 34711 318854 34720
rect 318812 26353 318840 34711
rect 318798 26344 318854 26353
rect 318798 26279 318854 26288
rect 323044 13258 323072 36230
rect 345676 16574 345704 38762
rect 345756 38684 345808 38690
rect 345756 38626 345808 38632
rect 345032 16546 345704 16574
rect 345032 16538 345060 16546
rect 344678 16510 345060 16538
rect 323032 13252 323084 13258
rect 323032 13194 323084 13200
rect 324056 13190 324084 16116
rect 334360 13190 334388 16116
rect 345768 13190 345796 38626
rect 352024 36924 352052 38830
rect 362316 38820 362368 38826
rect 362316 38762 362368 38768
rect 362328 36924 362356 38762
rect 372804 38752 372856 38758
rect 372804 38694 372856 38700
rect 372620 38684 372672 38690
rect 372620 38626 372672 38632
rect 372632 36924 372660 38626
rect 346398 35048 346454 35057
rect 346398 34983 346454 34992
rect 346412 26353 346440 34983
rect 350446 34776 350502 34785
rect 350446 34711 350502 34720
rect 350460 26353 350488 34711
rect 346398 26344 346454 26353
rect 346398 26279 346454 26288
rect 350446 26344 350502 26353
rect 350446 26279 350502 26288
rect 372816 16674 372844 38694
rect 373276 18630 373304 38830
rect 375378 34912 375434 34921
rect 375378 34847 375434 34856
rect 378046 34912 378102 34921
rect 378046 34847 378102 34856
rect 375392 26353 375420 34847
rect 378060 26353 378088 34847
rect 375378 26344 375434 26353
rect 375378 26279 375434 26288
rect 378046 26344 378102 26353
rect 378046 26279 378102 26288
rect 373264 18624 373316 18630
rect 373264 18566 373316 18572
rect 372646 16646 372844 16674
rect 352024 13258 352052 16116
rect 362328 13258 362356 16116
rect 378796 13326 378824 700470
rect 380348 687404 380400 687410
rect 380348 687346 380400 687352
rect 401140 687404 401192 687410
rect 401140 687346 401192 687352
rect 380360 684978 380388 687346
rect 390008 687336 390060 687342
rect 390008 687278 390060 687284
rect 380052 684950 380388 684978
rect 390020 684978 390048 687278
rect 401048 687268 401100 687274
rect 401048 687210 401100 687216
rect 390020 684950 390356 684978
rect 400660 684542 400996 684570
rect 400772 684276 400824 684282
rect 400772 684218 400824 684224
rect 379704 667208 379756 667214
rect 379704 667150 379756 667156
rect 379716 664714 379744 667150
rect 400784 664714 400812 684218
rect 400864 684208 400916 684214
rect 400864 684150 400916 684156
rect 400876 667214 400904 684150
rect 400864 667208 400916 667214
rect 400864 667150 400916 667156
rect 379716 664686 380052 664714
rect 400660 664686 400812 664714
rect 390356 664006 390508 664034
rect 390480 662386 390508 664006
rect 390468 662380 390520 662386
rect 390468 662322 390520 662328
rect 400968 662318 400996 684542
rect 401060 684282 401088 687210
rect 401048 684276 401100 684282
rect 401048 684218 401100 684224
rect 401152 684214 401180 687346
rect 418344 687268 418396 687274
rect 418344 687210 418396 687216
rect 418356 684964 418384 687210
rect 407224 684270 408066 684298
rect 428674 684270 428780 684298
rect 401140 684208 401192 684214
rect 401140 684150 401192 684156
rect 402978 674248 403034 674257
rect 402978 674183 403034 674192
rect 405646 674248 405702 674257
rect 405646 674183 405702 674192
rect 402992 665961 403020 674183
rect 405660 665961 405688 674183
rect 402978 665952 403034 665961
rect 402978 665887 403034 665896
rect 405646 665952 405702 665961
rect 405646 665887 405702 665896
rect 407224 662318 407252 684270
rect 407764 667208 407816 667214
rect 407764 667150 407816 667156
rect 407776 664714 407804 667150
rect 407776 664686 408066 664714
rect 400956 662312 401008 662318
rect 400956 662254 401008 662260
rect 407212 662312 407264 662318
rect 407212 662254 407264 662260
rect 418356 662250 418384 664020
rect 428660 662425 428688 664020
rect 428646 662416 428702 662425
rect 428752 662386 428780 684270
rect 428646 662351 428702 662360
rect 428740 662380 428792 662386
rect 428740 662322 428792 662328
rect 418344 662244 418396 662250
rect 418344 662186 418396 662192
rect 407212 659796 407264 659802
rect 407212 659738 407264 659744
rect 379612 659728 379664 659734
rect 379612 659670 379664 659676
rect 379520 655716 379572 655722
rect 379520 655658 379572 655664
rect 379532 634710 379560 655658
rect 379624 654134 379652 659670
rect 390834 657384 390890 657393
rect 390678 657342 390834 657370
rect 390834 657319 390890 657328
rect 379992 657206 380374 657234
rect 400982 657206 401088 657234
rect 379992 655722 380020 657206
rect 379980 655716 380032 655722
rect 379980 655658 380032 655664
rect 379624 654106 379928 654134
rect 379900 637786 379928 654106
rect 379900 637758 380374 637786
rect 390664 634710 390692 637092
rect 400968 634778 400996 637092
rect 401060 634778 401088 657206
rect 402978 656024 403034 656033
rect 402978 655959 403034 655968
rect 402992 647737 403020 655959
rect 407120 655716 407172 655722
rect 407120 655658 407172 655664
rect 402978 647728 403034 647737
rect 402978 647663 403034 647672
rect 400956 634772 401008 634778
rect 400956 634714 401008 634720
rect 401048 634772 401100 634778
rect 401048 634714 401100 634720
rect 407132 634710 407160 655658
rect 407224 654134 407252 659738
rect 418620 659728 418672 659734
rect 418620 659670 418672 659676
rect 418632 657900 418660 659670
rect 407960 657206 408342 657234
rect 428950 657206 429148 657234
rect 407960 655722 407988 657206
rect 408130 656024 408186 656033
rect 408130 655959 408186 655968
rect 407948 655716 408000 655722
rect 407948 655658 408000 655664
rect 407224 654106 407896 654134
rect 407868 637786 407896 654106
rect 408144 648281 408172 655959
rect 408130 648272 408186 648281
rect 408130 648207 408186 648216
rect 407868 637758 408342 637786
rect 418632 634710 418660 637092
rect 428936 634778 428964 637092
rect 429120 634778 429148 657206
rect 428924 634772 428976 634778
rect 428924 634714 428976 634720
rect 429108 634772 429160 634778
rect 429108 634714 429160 634720
rect 379520 634704 379572 634710
rect 379520 634646 379572 634652
rect 390652 634704 390704 634710
rect 390652 634646 390704 634652
rect 407120 634704 407172 634710
rect 407120 634646 407172 634652
rect 418620 634704 418672 634710
rect 418620 634646 418672 634652
rect 380348 632256 380400 632262
rect 380348 632198 380400 632204
rect 401140 632256 401192 632262
rect 401140 632198 401192 632204
rect 380360 630986 380388 632198
rect 390008 632188 390060 632194
rect 390008 632130 390060 632136
rect 380052 630958 380388 630986
rect 390020 630986 390048 632130
rect 401048 632120 401100 632126
rect 401048 632062 401100 632068
rect 390020 630958 390356 630986
rect 400660 630550 400996 630578
rect 400864 630216 400916 630222
rect 400864 630158 400916 630164
rect 400772 628652 400824 628658
rect 400772 628594 400824 628600
rect 379704 613420 379756 613426
rect 379704 613362 379756 613368
rect 379716 610722 379744 613362
rect 400784 610722 400812 628594
rect 400876 613426 400904 630158
rect 400864 613420 400916 613426
rect 400864 613362 400916 613368
rect 379716 610694 380052 610722
rect 400660 610694 400812 610722
rect 390356 610014 390508 610042
rect 390480 608598 390508 610014
rect 390468 608592 390520 608598
rect 390468 608534 390520 608540
rect 400968 608530 400996 630550
rect 401060 628658 401088 632062
rect 401152 630222 401180 632198
rect 418344 632120 418396 632126
rect 418344 632062 418396 632068
rect 418356 630972 418384 632062
rect 407224 630278 408066 630306
rect 428674 630278 428780 630306
rect 401140 630216 401192 630222
rect 401140 630158 401192 630164
rect 401048 628652 401100 628658
rect 401048 628594 401100 628600
rect 402978 620256 403034 620265
rect 402978 620191 403034 620200
rect 405646 620256 405702 620265
rect 405646 620191 405702 620200
rect 402992 611969 403020 620191
rect 405660 611969 405688 620191
rect 402978 611960 403034 611969
rect 402978 611895 403034 611904
rect 405646 611960 405702 611969
rect 405646 611895 405702 611904
rect 407224 608530 407252 630278
rect 407764 613420 407816 613426
rect 407764 613362 407816 613368
rect 407776 610722 407804 613362
rect 407776 610694 408066 610722
rect 400956 608524 401008 608530
rect 400956 608466 401008 608472
rect 407212 608524 407264 608530
rect 407212 608466 407264 608472
rect 418356 608462 418384 610028
rect 428660 608569 428688 610028
rect 428752 608598 428780 630278
rect 428740 608592 428792 608598
rect 428646 608560 428702 608569
rect 428740 608534 428792 608540
rect 428646 608495 428702 608504
rect 418344 608456 418396 608462
rect 418344 608398 418396 608404
rect 407212 605940 407264 605946
rect 407212 605882 407264 605888
rect 379520 605872 379572 605878
rect 379520 605814 379572 605820
rect 379532 583930 379560 605814
rect 390834 603392 390890 603401
rect 390678 603350 390834 603378
rect 390834 603327 390890 603336
rect 379624 603214 380374 603242
rect 400982 603214 401088 603242
rect 379624 585818 379652 603214
rect 379612 585812 379664 585818
rect 379612 585754 379664 585760
rect 379532 583902 379928 583930
rect 379900 583794 379928 583902
rect 379900 583766 380374 583794
rect 390664 580922 390692 583100
rect 400968 580990 400996 583100
rect 401060 580990 401088 603214
rect 402978 602168 403034 602177
rect 402978 602103 403034 602112
rect 405646 602168 405702 602177
rect 405646 602103 405702 602112
rect 402992 593745 403020 602103
rect 405660 593745 405688 602103
rect 407120 599752 407172 599758
rect 407120 599694 407172 599700
rect 402978 593736 403034 593745
rect 402978 593671 403034 593680
rect 405646 593736 405702 593745
rect 405646 593671 405702 593680
rect 400956 580984 401008 580990
rect 400956 580926 401008 580932
rect 401048 580984 401100 580990
rect 401048 580926 401100 580932
rect 407132 580922 407160 599694
rect 407224 596174 407252 605882
rect 418620 605872 418672 605878
rect 418620 605814 418672 605820
rect 418632 603908 418660 605814
rect 407960 603214 408342 603242
rect 428950 603214 429148 603242
rect 407960 599758 407988 603214
rect 429120 603158 429148 603214
rect 429108 603152 429160 603158
rect 429108 603094 429160 603100
rect 407948 599752 408000 599758
rect 407948 599694 408000 599700
rect 407224 596146 407896 596174
rect 407868 583794 407896 596146
rect 407868 583766 408342 583794
rect 418632 580922 418660 583100
rect 428936 580990 428964 583100
rect 428924 580984 428976 580990
rect 428924 580926 428976 580932
rect 390652 580916 390704 580922
rect 390652 580858 390704 580864
rect 407120 580916 407172 580922
rect 407120 580858 407172 580864
rect 418620 580916 418672 580922
rect 418620 580858 418672 580864
rect 390008 578332 390060 578338
rect 390008 578274 390060 578280
rect 400772 578332 400824 578338
rect 400772 578274 400824 578280
rect 418344 578332 418396 578338
rect 418344 578274 418396 578280
rect 380348 578264 380400 578270
rect 380348 578206 380400 578212
rect 380360 576994 380388 578206
rect 380052 576966 380388 576994
rect 390020 576994 390048 578274
rect 390020 576966 390356 576994
rect 400784 576434 400812 578274
rect 400864 578264 400916 578270
rect 400864 578206 400916 578212
rect 400876 576434 400904 578206
rect 418356 576980 418384 578274
rect 400772 576428 400824 576434
rect 400772 576370 400824 576376
rect 400864 576428 400916 576434
rect 400864 576370 400916 576376
rect 400660 576286 400996 576314
rect 400772 576224 400824 576230
rect 400772 576166 400824 576172
rect 400864 576224 400916 576230
rect 400864 576166 400916 576172
rect 379704 559564 379756 559570
rect 379704 559506 379756 559512
rect 379716 556730 379744 559506
rect 400784 556730 400812 576166
rect 400876 559570 400904 576166
rect 400864 559564 400916 559570
rect 400864 559506 400916 559512
rect 379716 556702 380052 556730
rect 400660 556702 400812 556730
rect 390356 556022 390508 556050
rect 390480 554742 390508 556022
rect 390468 554736 390520 554742
rect 390468 554678 390520 554684
rect 400968 554674 400996 576286
rect 407224 576286 408066 576314
rect 428674 576286 428780 576314
rect 402978 574696 403034 574705
rect 402978 574631 403034 574640
rect 405646 574696 405702 574705
rect 405646 574631 405702 574640
rect 402992 566273 403020 574631
rect 405660 566273 405688 574631
rect 402978 566264 403034 566273
rect 402978 566199 403034 566208
rect 405646 566264 405702 566273
rect 405646 566199 405702 566208
rect 407224 554674 407252 576286
rect 407764 559564 407816 559570
rect 407764 559506 407816 559512
rect 407776 556730 407804 559506
rect 407776 556702 408066 556730
rect 400956 554668 401008 554674
rect 400956 554610 401008 554616
rect 407212 554668 407264 554674
rect 407212 554610 407264 554616
rect 418356 554606 418384 556036
rect 428660 554713 428688 556036
rect 428752 554742 428780 576286
rect 428740 554736 428792 554742
rect 428646 554704 428702 554713
rect 428740 554678 428792 554684
rect 428646 554639 428702 554648
rect 418344 554600 418396 554606
rect 418344 554542 418396 554548
rect 407120 552152 407172 552158
rect 407120 552094 407172 552100
rect 379520 552084 379572 552090
rect 379520 552026 379572 552032
rect 379532 533662 379560 552026
rect 390834 549400 390890 549409
rect 390678 549358 390834 549386
rect 390834 549335 390890 549344
rect 379624 549222 380374 549250
rect 400982 549222 401088 549250
rect 379520 533656 379572 533662
rect 379520 533598 379572 533604
rect 379624 527066 379652 549222
rect 379980 533656 380032 533662
rect 379980 533598 380032 533604
rect 379992 529666 380020 533598
rect 379992 529638 380374 529666
rect 390664 527066 390692 529108
rect 400968 527134 400996 529108
rect 401060 527134 401088 549222
rect 402978 548040 403034 548049
rect 402978 547975 403034 547984
rect 402992 539753 403020 547975
rect 402978 539744 403034 539753
rect 402978 539679 403034 539688
rect 407132 533662 407160 552094
rect 418620 552084 418672 552090
rect 418620 552026 418672 552032
rect 418632 549916 418660 552026
rect 428950 549358 429148 549386
rect 429120 549302 429148 549358
rect 429108 549296 429160 549302
rect 407224 549222 408342 549250
rect 429108 549238 429160 549244
rect 407120 533656 407172 533662
rect 407120 533598 407172 533604
rect 400956 527128 401008 527134
rect 400956 527070 401008 527076
rect 401048 527128 401100 527134
rect 401048 527070 401100 527076
rect 407224 527066 407252 549222
rect 407948 533656 408000 533662
rect 407948 533598 408000 533604
rect 407960 529666 407988 533598
rect 407960 529638 408342 529666
rect 418632 527066 418660 529108
rect 428936 527134 428964 529108
rect 428924 527128 428976 527134
rect 428924 527070 428976 527076
rect 379612 527060 379664 527066
rect 379612 527002 379664 527008
rect 390652 527060 390704 527066
rect 390652 527002 390704 527008
rect 407212 527060 407264 527066
rect 407212 527002 407264 527008
rect 418620 527060 418672 527066
rect 418620 527002 418672 527008
rect 390008 524544 390060 524550
rect 390008 524486 390060 524492
rect 401048 524544 401100 524550
rect 401048 524486 401100 524492
rect 418344 524544 418396 524550
rect 418344 524486 418396 524492
rect 380348 524476 380400 524482
rect 380348 524418 380400 524424
rect 380360 522866 380388 524418
rect 380052 522838 380388 522866
rect 390020 522866 390048 524486
rect 390020 522838 390356 522866
rect 400660 522566 400996 522594
rect 400864 522232 400916 522238
rect 400864 522174 400916 522180
rect 400772 521756 400824 521762
rect 400772 521698 400824 521704
rect 379704 505776 379756 505782
rect 379704 505718 379756 505724
rect 379716 502738 379744 505718
rect 400784 502738 400812 521698
rect 400876 505782 400904 522174
rect 400864 505776 400916 505782
rect 400864 505718 400916 505724
rect 379716 502710 380052 502738
rect 400660 502710 400812 502738
rect 390356 502030 390508 502058
rect 390480 500954 390508 502030
rect 390468 500948 390520 500954
rect 390468 500890 390520 500896
rect 400968 500886 400996 522566
rect 401060 521762 401088 524486
rect 401140 524476 401192 524482
rect 401140 524418 401192 524424
rect 401152 522238 401180 524418
rect 418356 522852 418384 524486
rect 407224 522294 408066 522322
rect 428674 522294 428780 522322
rect 401140 522232 401192 522238
rect 401140 522174 401192 522180
rect 401048 521756 401100 521762
rect 401048 521698 401100 521704
rect 402978 520840 403034 520849
rect 402978 520775 403034 520784
rect 402992 512281 403020 520775
rect 402978 512272 403034 512281
rect 402978 512207 403034 512216
rect 407224 500886 407252 522294
rect 407764 505776 407816 505782
rect 407764 505718 407816 505724
rect 407776 502738 407804 505718
rect 407776 502710 408066 502738
rect 400956 500880 401008 500886
rect 400956 500822 401008 500828
rect 407212 500880 407264 500886
rect 407212 500822 407264 500828
rect 418356 500818 418384 502044
rect 428660 500857 428688 502044
rect 428752 500954 428780 522294
rect 428740 500948 428792 500954
rect 428740 500890 428792 500896
rect 428646 500848 428702 500857
rect 418344 500812 418396 500818
rect 428646 500783 428702 500792
rect 418344 500754 418396 500760
rect 407120 498296 407172 498302
rect 407120 498238 407172 498244
rect 379520 498228 379572 498234
rect 379520 498170 379572 498176
rect 379532 477698 379560 498170
rect 390834 495544 390890 495553
rect 390678 495502 390834 495530
rect 390834 495479 390890 495488
rect 379624 495230 380374 495258
rect 400982 495230 401088 495258
rect 379520 477692 379572 477698
rect 379520 477634 379572 477640
rect 379624 473278 379652 495230
rect 379980 477692 380032 477698
rect 379980 477634 380032 477640
rect 379992 475674 380020 477634
rect 379992 475646 380374 475674
rect 390664 473278 390692 475116
rect 400968 473346 400996 475116
rect 401060 473346 401088 495230
rect 402978 485752 403034 485761
rect 402978 485687 403034 485696
rect 402992 477329 403020 485687
rect 407132 477698 407160 498238
rect 418620 498228 418672 498234
rect 418620 498170 418672 498176
rect 418632 495924 418660 498170
rect 407224 495230 408342 495258
rect 428950 495242 429148 495258
rect 428950 495236 429160 495242
rect 428950 495230 429108 495236
rect 407120 477692 407172 477698
rect 407120 477634 407172 477640
rect 402978 477320 403034 477329
rect 402978 477255 403034 477264
rect 400956 473340 401008 473346
rect 400956 473282 401008 473288
rect 401048 473340 401100 473346
rect 401048 473282 401100 473288
rect 407224 473278 407252 495230
rect 429108 495178 429160 495184
rect 407948 477692 408000 477698
rect 407948 477634 408000 477640
rect 407960 475674 407988 477634
rect 407960 475646 408342 475674
rect 418632 473278 418660 475116
rect 428936 473346 428964 475116
rect 428924 473340 428976 473346
rect 428924 473282 428976 473288
rect 379612 473272 379664 473278
rect 379612 473214 379664 473220
rect 390652 473272 390704 473278
rect 390652 473214 390704 473220
rect 407212 473272 407264 473278
rect 407212 473214 407264 473220
rect 418620 473272 418672 473278
rect 418620 473214 418672 473220
rect 380348 470824 380400 470830
rect 380348 470766 380400 470772
rect 400864 470824 400916 470830
rect 400864 470766 400916 470772
rect 380360 468874 380388 470766
rect 390008 470756 390060 470762
rect 390008 470698 390060 470704
rect 380052 468846 380388 468874
rect 390020 468874 390048 470698
rect 400772 470688 400824 470694
rect 400772 470630 400824 470636
rect 390020 468846 390356 468874
rect 400784 468450 400812 470630
rect 400876 468450 400904 470766
rect 418344 470688 418396 470694
rect 418344 470630 418396 470636
rect 418356 468860 418384 470630
rect 400772 468444 400824 468450
rect 400772 468386 400824 468392
rect 400864 468444 400916 468450
rect 400864 468386 400916 468392
rect 400660 468302 400996 468330
rect 400772 468240 400824 468246
rect 400772 468182 400824 468188
rect 400864 468240 400916 468246
rect 400864 468182 400916 468188
rect 379704 451920 379756 451926
rect 379704 451862 379756 451868
rect 379716 448746 379744 451862
rect 400784 448746 400812 468182
rect 400876 451926 400904 468182
rect 400864 451920 400916 451926
rect 400864 451862 400916 451868
rect 379716 448718 380052 448746
rect 400660 448718 400812 448746
rect 390356 448038 390508 448066
rect 390480 445738 390508 448038
rect 390468 445732 390520 445738
rect 390468 445674 390520 445680
rect 400968 445670 400996 468302
rect 407224 468302 408066 468330
rect 428674 468302 428780 468330
rect 402978 466848 403034 466857
rect 402978 466783 403034 466792
rect 402992 458289 403020 466783
rect 402978 458280 403034 458289
rect 402978 458215 403034 458224
rect 407224 445670 407252 468302
rect 407764 451920 407816 451926
rect 407764 451862 407816 451868
rect 407776 448746 407804 451862
rect 407776 448718 408066 448746
rect 400956 445664 401008 445670
rect 400956 445606 401008 445612
rect 407212 445664 407264 445670
rect 418356 445641 418384 448052
rect 407212 445606 407264 445612
rect 418342 445632 418398 445641
rect 418342 445567 418398 445576
rect 428660 445505 428688 448052
rect 428752 445738 428780 468302
rect 428740 445732 428792 445738
rect 428740 445674 428792 445680
rect 428646 445496 428702 445505
rect 428646 445431 428702 445440
rect 407120 444508 407172 444514
rect 407120 444450 407172 444456
rect 379612 444440 379664 444446
rect 379612 444382 379664 444388
rect 379624 441614 379652 444382
rect 390834 441688 390890 441697
rect 390678 441646 390834 441674
rect 390834 441623 390890 441632
rect 379624 441586 379928 441614
rect 379900 421682 379928 441586
rect 379992 441238 380374 441266
rect 400982 441238 401088 441266
rect 379992 439550 380020 441238
rect 379980 439544 380032 439550
rect 379980 439486 380032 439492
rect 379900 421654 380374 421682
rect 390664 419422 390692 421124
rect 400968 419490 400996 421124
rect 401060 419490 401088 441238
rect 402978 431760 403034 431769
rect 402978 431695 403034 431704
rect 405646 431760 405702 431769
rect 405646 431695 405702 431704
rect 402992 423201 403020 431695
rect 405660 423201 405688 431695
rect 407132 427174 407160 444450
rect 418620 444440 418672 444446
rect 418620 444382 418672 444388
rect 418632 441932 418660 444382
rect 428950 441658 429148 441674
rect 428950 441652 429160 441658
rect 428950 441646 429108 441652
rect 429108 441594 429160 441600
rect 407224 441238 408342 441266
rect 407120 427168 407172 427174
rect 407120 427110 407172 427116
rect 402978 423192 403034 423201
rect 402978 423127 403034 423136
rect 405646 423192 405702 423201
rect 405646 423127 405702 423136
rect 400956 419484 401008 419490
rect 400956 419426 401008 419432
rect 401048 419484 401100 419490
rect 401048 419426 401100 419432
rect 407224 419422 407252 441238
rect 407948 427168 408000 427174
rect 407948 427110 408000 427116
rect 407960 421682 407988 427110
rect 407960 421654 408342 421682
rect 418632 419422 418660 421124
rect 428936 419490 428964 421124
rect 428924 419484 428976 419490
rect 428924 419426 428976 419432
rect 390652 419416 390704 419422
rect 390652 419358 390704 419364
rect 407212 419416 407264 419422
rect 407212 419358 407264 419364
rect 418620 419416 418672 419422
rect 418620 419358 418672 419364
rect 380348 416968 380400 416974
rect 380348 416910 380400 416916
rect 401140 416968 401192 416974
rect 401140 416910 401192 416916
rect 380360 414882 380388 416910
rect 390008 416900 390060 416906
rect 390008 416842 390060 416848
rect 380052 414854 380388 414882
rect 390020 414882 390048 416842
rect 401048 416832 401100 416838
rect 401048 416774 401100 416780
rect 390020 414854 390356 414882
rect 400660 414582 400996 414610
rect 400772 414316 400824 414322
rect 400772 414258 400824 414264
rect 379704 396772 379756 396778
rect 379704 396714 379756 396720
rect 379716 394754 379744 396714
rect 400784 394754 400812 414258
rect 400864 414248 400916 414254
rect 400864 414190 400916 414196
rect 400876 396778 400904 414190
rect 400864 396772 400916 396778
rect 400864 396714 400916 396720
rect 379716 394726 380052 394754
rect 400660 394726 400812 394754
rect 390356 394046 390508 394074
rect 390480 391950 390508 394046
rect 390468 391944 390520 391950
rect 390468 391886 390520 391892
rect 400968 391882 400996 414582
rect 401060 414322 401088 416774
rect 401048 414316 401100 414322
rect 401048 414258 401100 414264
rect 401152 414254 401180 416910
rect 418344 416832 418396 416838
rect 418344 416774 418396 416780
rect 418356 414868 418384 416774
rect 407224 414310 408066 414338
rect 428674 414310 428780 414338
rect 401140 414248 401192 414254
rect 401140 414190 401192 414196
rect 402978 404288 403034 404297
rect 402978 404223 403034 404232
rect 402992 396001 403020 404223
rect 402978 395992 403034 396001
rect 402978 395927 403034 395936
rect 407224 391882 407252 414310
rect 407764 396772 407816 396778
rect 407764 396714 407816 396720
rect 407776 394754 407804 396714
rect 407776 394726 408066 394754
rect 418356 391921 418384 394060
rect 418342 391912 418398 391921
rect 400956 391876 401008 391882
rect 400956 391818 401008 391824
rect 407212 391876 407264 391882
rect 418342 391847 418398 391856
rect 407212 391818 407264 391824
rect 428660 391785 428688 394060
rect 428752 391950 428780 414310
rect 428740 391944 428792 391950
rect 428740 391886 428792 391892
rect 428646 391776 428702 391785
rect 428646 391711 428702 391720
rect 407212 389292 407264 389298
rect 407212 389234 407264 389240
rect 379612 389224 379664 389230
rect 379612 389166 379664 389172
rect 379520 385484 379572 385490
rect 379520 385426 379572 385432
rect 379532 365634 379560 385426
rect 379624 383654 379652 389166
rect 390834 387424 390890 387433
rect 390678 387382 390834 387410
rect 390834 387359 390890 387368
rect 379992 387246 380374 387274
rect 400982 387246 401088 387274
rect 379992 385490 380020 387246
rect 379980 385484 380032 385490
rect 379980 385426 380032 385432
rect 379624 383626 379928 383654
rect 379900 367690 379928 383626
rect 379900 367662 380374 367690
rect 390664 365634 390692 367132
rect 400968 365702 400996 367132
rect 401060 365702 401088 387246
rect 407120 385484 407172 385490
rect 407120 385426 407172 385432
rect 402978 377768 403034 377777
rect 402978 377703 403034 377712
rect 405646 377768 405702 377777
rect 405646 377703 405702 377712
rect 402992 369345 403020 377703
rect 405660 369345 405688 377703
rect 402978 369336 403034 369345
rect 402978 369271 403034 369280
rect 405646 369336 405702 369345
rect 405646 369271 405702 369280
rect 400956 365696 401008 365702
rect 400956 365638 401008 365644
rect 401048 365696 401100 365702
rect 401048 365638 401100 365644
rect 407132 365634 407160 385426
rect 407224 383654 407252 389234
rect 418620 389224 418672 389230
rect 418620 389166 418672 389172
rect 418632 387940 418660 389166
rect 407960 387246 408342 387274
rect 428950 387246 429148 387274
rect 407960 385490 407988 387246
rect 429120 386442 429148 387246
rect 429108 386436 429160 386442
rect 429108 386378 429160 386384
rect 407948 385484 408000 385490
rect 407948 385426 408000 385432
rect 407224 383626 407896 383654
rect 407868 367690 407896 383626
rect 407868 367662 408342 367690
rect 418632 365634 418660 367132
rect 428936 365702 428964 367132
rect 428924 365696 428976 365702
rect 428924 365638 428976 365644
rect 379520 365628 379572 365634
rect 379520 365570 379572 365576
rect 390652 365628 390704 365634
rect 390652 365570 390704 365576
rect 407120 365628 407172 365634
rect 407120 365570 407172 365576
rect 418620 365628 418672 365634
rect 418620 365570 418672 365576
rect 390008 363044 390060 363050
rect 390008 362986 390060 362992
rect 401048 363044 401100 363050
rect 401048 362986 401100 362992
rect 418344 363044 418396 363050
rect 418344 362986 418396 362992
rect 380348 362976 380400 362982
rect 380348 362918 380400 362924
rect 380360 360890 380388 362918
rect 380052 360862 380388 360890
rect 390020 360890 390048 362986
rect 390020 360862 390356 360890
rect 400660 360590 400996 360618
rect 400864 360256 400916 360262
rect 400864 360198 400916 360204
rect 400772 358896 400824 358902
rect 400772 358838 400824 358844
rect 379704 342916 379756 342922
rect 379704 342858 379756 342864
rect 379716 340762 379744 342858
rect 400784 340762 400812 358838
rect 400876 342922 400904 360198
rect 400864 342916 400916 342922
rect 400864 342858 400916 342864
rect 379716 340734 380052 340762
rect 400660 340734 400812 340762
rect 390356 340054 390508 340082
rect 390480 338094 390508 340054
rect 390468 338088 390520 338094
rect 390468 338030 390520 338036
rect 400968 338026 400996 360590
rect 401060 358902 401088 362986
rect 401140 362976 401192 362982
rect 401140 362918 401192 362924
rect 401152 360262 401180 362918
rect 418356 360876 418384 362986
rect 407224 360318 408066 360346
rect 428674 360318 428780 360346
rect 401140 360256 401192 360262
rect 401140 360198 401192 360204
rect 401048 358896 401100 358902
rect 401048 358838 401100 358844
rect 402978 350296 403034 350305
rect 402978 350231 403034 350240
rect 402992 342009 403020 350231
rect 402978 342000 403034 342009
rect 402978 341935 403034 341944
rect 407224 338026 407252 360318
rect 407764 342916 407816 342922
rect 407764 342858 407816 342864
rect 407776 340762 407804 342858
rect 407776 340734 408066 340762
rect 400956 338020 401008 338026
rect 400956 337962 401008 337968
rect 407212 338020 407264 338026
rect 407212 337962 407264 337968
rect 418356 337958 418384 340068
rect 428660 338065 428688 340068
rect 428752 338094 428780 360318
rect 428740 338088 428792 338094
rect 428646 338056 428702 338065
rect 428740 338030 428792 338036
rect 428646 337991 428702 338000
rect 418344 337952 418396 337958
rect 418344 337894 418396 337900
rect 407212 335436 407264 335442
rect 407212 335378 407264 335384
rect 379612 335368 379664 335374
rect 379612 335310 379664 335316
rect 379520 329520 379572 329526
rect 379520 329462 379572 329468
rect 379532 311778 379560 329462
rect 379624 325694 379652 335310
rect 390834 333296 390890 333305
rect 379992 333254 380374 333282
rect 390678 333254 390834 333282
rect 379992 329526 380020 333254
rect 400982 333254 401088 333282
rect 390834 333231 390890 333240
rect 379980 329520 380032 329526
rect 379980 329462 380032 329468
rect 379624 325666 379928 325694
rect 379900 313698 379928 325666
rect 379900 313670 380374 313698
rect 390664 311778 390692 313140
rect 400968 311846 400996 313140
rect 401060 311846 401088 333254
rect 407120 329520 407172 329526
rect 407120 329462 407172 329468
rect 402978 323776 403034 323785
rect 402978 323711 403034 323720
rect 405646 323776 405702 323785
rect 405646 323711 405702 323720
rect 402992 315353 403020 323711
rect 405660 315353 405688 323711
rect 402978 315344 403034 315353
rect 402978 315279 403034 315288
rect 405646 315344 405702 315353
rect 405646 315279 405702 315288
rect 400956 311840 401008 311846
rect 400956 311782 401008 311788
rect 401048 311840 401100 311846
rect 401048 311782 401100 311788
rect 407132 311778 407160 329462
rect 407224 325694 407252 335378
rect 418620 335368 418672 335374
rect 418620 335310 418672 335316
rect 418632 333948 418660 335310
rect 407960 333254 408342 333282
rect 428950 333254 429148 333282
rect 407960 329526 407988 333254
rect 429120 332654 429148 333254
rect 429108 332648 429160 332654
rect 429108 332590 429160 332596
rect 407948 329520 408000 329526
rect 407948 329462 408000 329468
rect 407224 325666 407896 325694
rect 407868 313698 407896 325666
rect 407868 313670 408342 313698
rect 418632 311778 418660 313140
rect 428936 311846 428964 313140
rect 428924 311840 428976 311846
rect 428924 311782 428976 311788
rect 379520 311772 379572 311778
rect 379520 311714 379572 311720
rect 390652 311772 390704 311778
rect 390652 311714 390704 311720
rect 407120 311772 407172 311778
rect 407120 311714 407172 311720
rect 418620 311772 418672 311778
rect 418620 311714 418672 311720
rect 380348 309324 380400 309330
rect 380348 309266 380400 309272
rect 401048 309324 401100 309330
rect 401048 309266 401100 309272
rect 380360 306898 380388 309266
rect 390008 309256 390060 309262
rect 390008 309198 390060 309204
rect 380052 306870 380388 306898
rect 390020 306898 390048 309198
rect 390020 306870 390356 306898
rect 400660 306598 400996 306626
rect 400772 305720 400824 305726
rect 400772 305662 400824 305668
rect 379704 289128 379756 289134
rect 379704 289070 379756 289076
rect 379716 286770 379744 289070
rect 400784 286770 400812 305662
rect 400968 297498 400996 306598
rect 400956 297492 401008 297498
rect 400956 297434 401008 297440
rect 400956 297288 401008 297294
rect 400956 297230 401008 297236
rect 400864 292528 400916 292534
rect 400864 292470 400916 292476
rect 400876 289134 400904 292470
rect 400864 289128 400916 289134
rect 400864 289070 400916 289076
rect 379716 286742 380052 286770
rect 400660 286742 400812 286770
rect 390356 286062 390508 286090
rect 390480 284306 390508 286062
rect 390468 284300 390520 284306
rect 390468 284242 390520 284248
rect 400968 284238 400996 297230
rect 401060 292534 401088 309266
rect 401140 309188 401192 309194
rect 401140 309130 401192 309136
rect 418344 309188 418396 309194
rect 418344 309130 418396 309136
rect 401152 305726 401180 309130
rect 418356 306884 418384 309130
rect 407224 306326 408066 306354
rect 428674 306326 428780 306354
rect 401140 305720 401192 305726
rect 401140 305662 401192 305668
rect 402978 296304 403034 296313
rect 402978 296239 403034 296248
rect 401048 292528 401100 292534
rect 401048 292470 401100 292476
rect 402992 287881 403020 296239
rect 402978 287872 403034 287881
rect 402978 287807 403034 287816
rect 407224 284238 407252 306326
rect 407764 289128 407816 289134
rect 407764 289070 407816 289076
rect 407776 286770 407804 289070
rect 407776 286742 408066 286770
rect 400956 284232 401008 284238
rect 400956 284174 401008 284180
rect 407212 284232 407264 284238
rect 407212 284174 407264 284180
rect 418356 284170 418384 286076
rect 428660 284209 428688 286076
rect 428752 284306 428780 306326
rect 428740 284300 428792 284306
rect 428740 284242 428792 284248
rect 428646 284200 428702 284209
rect 418344 284164 418396 284170
rect 428646 284135 428702 284144
rect 418344 284106 418396 284112
rect 407212 281648 407264 281654
rect 407212 281590 407264 281596
rect 379612 281580 379664 281586
rect 379612 281522 379664 281528
rect 379520 272604 379572 272610
rect 379520 272546 379572 272552
rect 379532 256630 379560 272546
rect 379624 267734 379652 281522
rect 390834 279304 390890 279313
rect 379992 279262 380374 279290
rect 390678 279262 390834 279290
rect 379992 272610 380020 279262
rect 400982 279262 401088 279290
rect 390834 279239 390890 279248
rect 379980 272604 380032 272610
rect 379980 272546 380032 272552
rect 379624 267706 379928 267734
rect 379900 259706 379928 267706
rect 379900 259678 380374 259706
rect 390664 256630 390692 259148
rect 400968 256698 400996 259148
rect 401060 256698 401088 279262
rect 402978 278080 403034 278089
rect 402978 278015 403034 278024
rect 405646 278080 405702 278089
rect 405646 278015 405702 278024
rect 402992 269793 403020 278015
rect 405660 269793 405688 278015
rect 407120 272604 407172 272610
rect 407120 272546 407172 272552
rect 402978 269784 403034 269793
rect 402978 269719 403034 269728
rect 405646 269784 405702 269793
rect 405646 269719 405702 269728
rect 400956 256692 401008 256698
rect 400956 256634 401008 256640
rect 401048 256692 401100 256698
rect 401048 256634 401100 256640
rect 407132 256630 407160 272546
rect 407224 267734 407252 281590
rect 418620 281580 418672 281586
rect 418620 281522 418672 281528
rect 418632 279956 418660 281522
rect 407960 279262 408342 279290
rect 428950 279262 429148 279290
rect 407960 272610 407988 279262
rect 407948 272604 408000 272610
rect 407948 272546 408000 272552
rect 407224 267706 407896 267734
rect 407868 259706 407896 267706
rect 407868 259678 408342 259706
rect 418632 256630 418660 259148
rect 428936 256698 428964 259148
rect 429120 256698 429148 279262
rect 428924 256692 428976 256698
rect 428924 256634 428976 256640
rect 429108 256692 429160 256698
rect 429108 256634 429160 256640
rect 379520 256624 379572 256630
rect 379520 256566 379572 256572
rect 390652 256624 390704 256630
rect 390652 256566 390704 256572
rect 407120 256624 407172 256630
rect 407120 256566 407172 256572
rect 418620 256624 418672 256630
rect 418620 256566 418672 256572
rect 380348 255468 380400 255474
rect 380348 255410 380400 255416
rect 401140 255468 401192 255474
rect 401140 255410 401192 255416
rect 380360 252906 380388 255410
rect 390008 255400 390060 255406
rect 390008 255342 390060 255348
rect 380052 252878 380388 252906
rect 390020 252906 390048 255342
rect 401048 255332 401100 255338
rect 401048 255274 401100 255280
rect 390020 252878 390356 252906
rect 400660 252606 400996 252634
rect 400864 252272 400916 252278
rect 400864 252214 400916 252220
rect 400772 249144 400824 249150
rect 400772 249086 400824 249092
rect 379704 235272 379756 235278
rect 379704 235214 379756 235220
rect 379716 232778 379744 235214
rect 400784 232778 400812 249086
rect 400876 235278 400904 252214
rect 400864 235272 400916 235278
rect 400864 235214 400916 235220
rect 379716 232750 380052 232778
rect 400660 232750 400812 232778
rect 390356 232070 390508 232098
rect 390480 230450 390508 232070
rect 390468 230444 390520 230450
rect 390468 230386 390520 230392
rect 400968 230382 400996 252606
rect 401060 249150 401088 255274
rect 401152 252278 401180 255410
rect 418344 255332 418396 255338
rect 418344 255274 418396 255280
rect 418356 252892 418384 255274
rect 407224 252334 408066 252362
rect 428674 252334 428780 252362
rect 401140 252272 401192 252278
rect 401140 252214 401192 252220
rect 401048 249144 401100 249150
rect 401048 249086 401100 249092
rect 402978 242312 403034 242321
rect 402978 242247 403034 242256
rect 405646 242312 405702 242321
rect 405646 242247 405702 242256
rect 402992 234025 403020 242247
rect 405660 234025 405688 242247
rect 402978 234016 403034 234025
rect 402978 233951 403034 233960
rect 405646 234016 405702 234025
rect 405646 233951 405702 233960
rect 407224 230382 407252 252334
rect 407764 235272 407816 235278
rect 407764 235214 407816 235220
rect 407776 232778 407804 235214
rect 407776 232750 408066 232778
rect 400956 230376 401008 230382
rect 400956 230318 401008 230324
rect 407212 230376 407264 230382
rect 407212 230318 407264 230324
rect 418356 230314 418384 232084
rect 428660 230489 428688 232084
rect 428646 230480 428702 230489
rect 428752 230450 428780 252334
rect 428646 230415 428702 230424
rect 428740 230444 428792 230450
rect 428740 230386 428792 230392
rect 418344 230308 418396 230314
rect 418344 230250 418396 230256
rect 407856 227928 407908 227934
rect 407856 227870 407908 227876
rect 379888 227860 379940 227866
rect 379888 227802 379940 227808
rect 378876 227792 378928 227798
rect 378876 227734 378928 227740
rect 378888 202774 378916 227734
rect 379520 222352 379572 222358
rect 379520 222294 379572 222300
rect 378876 202768 378928 202774
rect 378876 202710 378928 202716
rect 379532 202706 379560 222294
rect 379900 205714 379928 227802
rect 390652 227792 390704 227798
rect 390652 227734 390704 227740
rect 402244 227792 402296 227798
rect 402244 227734 402296 227740
rect 390664 225964 390692 227734
rect 379992 225270 380374 225298
rect 400982 225270 401088 225298
rect 379992 222358 380020 225270
rect 379980 222352 380032 222358
rect 379980 222294 380032 222300
rect 379900 205686 380374 205714
rect 390678 205006 390968 205034
rect 390940 202774 390968 205006
rect 400600 205006 400982 205034
rect 400600 202842 400628 205006
rect 401060 202842 401088 225270
rect 400588 202836 400640 202842
rect 400588 202778 400640 202784
rect 401048 202836 401100 202842
rect 401048 202778 401100 202784
rect 402256 202774 402284 227734
rect 405648 225072 405700 225078
rect 405648 225014 405700 225020
rect 402978 224088 403034 224097
rect 402978 224023 403034 224032
rect 402992 215801 403020 224023
rect 405660 215801 405688 225014
rect 402978 215792 403034 215801
rect 402978 215727 403034 215736
rect 405646 215792 405702 215801
rect 405646 215727 405702 215736
rect 407868 205714 407896 227870
rect 418620 227860 418672 227866
rect 418620 227802 418672 227808
rect 408316 227792 408368 227798
rect 408316 227734 408368 227740
rect 408328 225964 408356 227734
rect 418632 225964 418660 227802
rect 428950 225270 429148 225298
rect 429120 225010 429148 225270
rect 429108 225004 429160 225010
rect 429108 224946 429160 224952
rect 407868 205686 408342 205714
rect 418632 202774 418660 205020
rect 428936 202842 428964 205020
rect 428924 202836 428976 202842
rect 428924 202778 428976 202784
rect 390928 202768 390980 202774
rect 390928 202710 390980 202716
rect 402244 202768 402296 202774
rect 402244 202710 402296 202716
rect 418620 202768 418672 202774
rect 418620 202710 418672 202716
rect 379520 202700 379572 202706
rect 379520 202642 379572 202648
rect 390008 200252 390060 200258
rect 390008 200194 390060 200200
rect 400772 200252 400824 200258
rect 400772 200194 400824 200200
rect 418344 200252 418396 200258
rect 418344 200194 418396 200200
rect 380348 200184 380400 200190
rect 380348 200126 380400 200132
rect 380360 198914 380388 200126
rect 380052 198886 380388 198914
rect 390020 198914 390048 200194
rect 390020 198886 390356 198914
rect 400784 198354 400812 200194
rect 400864 200184 400916 200190
rect 400864 200126 400916 200132
rect 400876 198354 400904 200126
rect 418356 198900 418384 200194
rect 400772 198348 400824 198354
rect 400772 198290 400824 198296
rect 400864 198348 400916 198354
rect 400864 198290 400916 198296
rect 400660 198206 400996 198234
rect 400772 198144 400824 198150
rect 400772 198086 400824 198092
rect 400864 198144 400916 198150
rect 400864 198086 400916 198092
rect 379704 181484 379756 181490
rect 379704 181426 379756 181432
rect 379716 178786 379744 181426
rect 400784 178786 400812 198086
rect 400876 181490 400904 198086
rect 400864 181484 400916 181490
rect 400864 181426 400916 181432
rect 379716 178758 380052 178786
rect 400660 178758 400812 178786
rect 390356 178078 390508 178106
rect 390480 176662 390508 178078
rect 390468 176656 390520 176662
rect 390468 176598 390520 176604
rect 400968 176594 400996 198206
rect 407224 198206 408066 198234
rect 428674 198206 428780 198234
rect 402978 196752 403034 196761
rect 402978 196687 403034 196696
rect 405646 196752 405702 196761
rect 405646 196687 405702 196696
rect 402992 188329 403020 196687
rect 405660 188329 405688 196687
rect 402978 188320 403034 188329
rect 402978 188255 403034 188264
rect 405646 188320 405702 188329
rect 405646 188255 405702 188264
rect 407224 176594 407252 198206
rect 407764 181484 407816 181490
rect 407764 181426 407816 181432
rect 407776 178786 407804 181426
rect 407776 178758 408066 178786
rect 400956 176588 401008 176594
rect 400956 176530 401008 176536
rect 407212 176588 407264 176594
rect 407212 176530 407264 176536
rect 418356 176526 418384 178092
rect 428660 176633 428688 178092
rect 428752 176662 428780 198206
rect 428740 176656 428792 176662
rect 428646 176624 428702 176633
rect 428740 176598 428792 176604
rect 428646 176559 428702 176568
rect 418344 176520 418396 176526
rect 418344 176462 418396 176468
rect 380348 174072 380400 174078
rect 380348 174014 380400 174020
rect 407212 174072 407264 174078
rect 407212 174014 407264 174020
rect 379612 173936 379664 173942
rect 379612 173878 379664 173884
rect 379624 171134 379652 173878
rect 380360 171972 380388 174014
rect 390652 174004 390704 174010
rect 390652 173946 390704 173952
rect 402244 174004 402296 174010
rect 402244 173946 402296 173952
rect 390664 171972 390692 173946
rect 400982 171278 401088 171306
rect 379624 171106 379928 171134
rect 379900 151722 379928 171106
rect 379900 151694 380374 151722
rect 390664 148986 390692 151028
rect 400968 149054 400996 151028
rect 401060 149054 401088 171278
rect 400956 149048 401008 149054
rect 400956 148990 401008 148996
rect 401048 149048 401100 149054
rect 401048 148990 401100 148996
rect 402256 148986 402284 173946
rect 407224 171134 407252 174014
rect 408316 174004 408368 174010
rect 408316 173946 408368 173952
rect 408328 171972 408356 173946
rect 418620 173936 418672 173942
rect 418620 173878 418672 173884
rect 418632 171972 418660 173878
rect 428950 171278 429148 171306
rect 429120 171222 429148 171278
rect 429108 171216 429160 171222
rect 429108 171158 429160 171164
rect 407224 171106 407896 171134
rect 402978 170096 403034 170105
rect 402978 170031 403034 170040
rect 402992 161809 403020 170031
rect 402978 161800 403034 161809
rect 402978 161735 403034 161744
rect 407868 151722 407896 171106
rect 407868 151694 408342 151722
rect 418632 148986 418660 151028
rect 428936 149054 428964 151028
rect 428924 149048 428976 149054
rect 428924 148990 428976 148996
rect 390652 148980 390704 148986
rect 390652 148922 390704 148928
rect 402244 148980 402296 148986
rect 402244 148922 402296 148928
rect 418620 148980 418672 148986
rect 418620 148922 418672 148928
rect 380348 146464 380400 146470
rect 380348 146406 380400 146412
rect 401048 146464 401100 146470
rect 401048 146406 401100 146412
rect 380360 144922 380388 146406
rect 390008 146396 390060 146402
rect 390008 146338 390060 146344
rect 380052 144894 380388 144922
rect 390020 144922 390048 146338
rect 390020 144894 390356 144922
rect 400660 144486 400996 144514
rect 400772 144220 400824 144226
rect 400772 144162 400824 144168
rect 379704 127628 379756 127634
rect 379704 127570 379756 127576
rect 379716 124794 379744 127570
rect 400784 124794 400812 144162
rect 400864 144152 400916 144158
rect 400864 144094 400916 144100
rect 400876 127634 400904 144094
rect 400864 127628 400916 127634
rect 400864 127570 400916 127576
rect 379716 124766 380052 124794
rect 400660 124766 400812 124794
rect 390356 124086 390508 124114
rect 390480 122806 390508 124086
rect 390468 122800 390520 122806
rect 390468 122742 390520 122748
rect 400968 122738 400996 144486
rect 401060 144158 401088 146406
rect 401140 146328 401192 146334
rect 401140 146270 401192 146276
rect 418344 146328 418396 146334
rect 418344 146270 418396 146276
rect 401152 144226 401180 146270
rect 418356 144908 418384 146270
rect 401140 144220 401192 144226
rect 401140 144162 401192 144168
rect 407224 144214 408066 144242
rect 428674 144214 428780 144242
rect 401048 144152 401100 144158
rect 401048 144094 401100 144100
rect 402978 134328 403034 134337
rect 402978 134263 403034 134272
rect 405646 134328 405702 134337
rect 405646 134263 405702 134272
rect 402992 125594 403020 134263
rect 405660 125594 405688 134263
rect 402980 125588 403032 125594
rect 402980 125530 403032 125536
rect 405648 125588 405700 125594
rect 405648 125530 405700 125536
rect 407224 122738 407252 144214
rect 407764 127628 407816 127634
rect 407764 127570 407816 127576
rect 407776 124794 407804 127570
rect 407776 124766 408066 124794
rect 400956 122732 401008 122738
rect 400956 122674 401008 122680
rect 407212 122732 407264 122738
rect 407212 122674 407264 122680
rect 418356 122670 418384 124100
rect 428660 122777 428688 124100
rect 428752 122806 428780 144214
rect 428740 122800 428792 122806
rect 428646 122768 428702 122777
rect 428740 122742 428792 122748
rect 428646 122703 428702 122712
rect 418344 122664 418396 122670
rect 418344 122606 418396 122612
rect 407212 120284 407264 120290
rect 407212 120226 407264 120232
rect 378876 120216 378928 120222
rect 378876 120158 378928 120164
rect 390744 120216 390796 120222
rect 390744 120158 390796 120164
rect 402244 120216 402296 120222
rect 402244 120158 402296 120164
rect 378888 95130 378916 120158
rect 379520 120148 379572 120154
rect 379520 120090 379572 120096
rect 379532 100298 379560 120090
rect 390756 117858 390784 120158
rect 390678 117830 390784 117858
rect 379624 117286 380374 117314
rect 400982 117286 401088 117314
rect 379520 100292 379572 100298
rect 379520 100234 379572 100240
rect 378876 95124 378928 95130
rect 378876 95066 378928 95072
rect 379624 95062 379652 117286
rect 379980 100292 380032 100298
rect 379980 100234 380032 100240
rect 379992 97730 380020 100234
rect 379992 97702 380374 97730
rect 390664 95130 390692 97036
rect 400968 95198 400996 97036
rect 401060 95198 401088 117286
rect 400956 95192 401008 95198
rect 400956 95134 401008 95140
rect 401048 95192 401100 95198
rect 401048 95134 401100 95140
rect 402256 95130 402284 120158
rect 402978 116104 403034 116113
rect 402978 116039 403034 116048
rect 402992 107817 403020 116039
rect 407224 113174 407252 120226
rect 408316 120216 408368 120222
rect 408316 120158 408368 120164
rect 408328 117980 408356 120158
rect 418620 120148 418672 120154
rect 418620 120090 418672 120096
rect 418632 117980 418660 120090
rect 428950 117298 429148 117314
rect 428950 117292 429160 117298
rect 428950 117286 429108 117292
rect 429108 117234 429160 117240
rect 407224 113146 407896 113174
rect 402978 107808 403034 107817
rect 402978 107743 403034 107752
rect 407868 97730 407896 113146
rect 407868 97702 408342 97730
rect 418632 95130 418660 97036
rect 428936 95198 428964 97036
rect 428924 95192 428976 95198
rect 428924 95134 428976 95140
rect 390652 95124 390704 95130
rect 390652 95066 390704 95072
rect 402244 95124 402296 95130
rect 402244 95066 402296 95072
rect 418620 95124 418672 95130
rect 418620 95066 418672 95072
rect 379612 95056 379664 95062
rect 379612 94998 379664 95004
rect 390008 92676 390060 92682
rect 390008 92618 390060 92624
rect 380348 92608 380400 92614
rect 380348 92550 380400 92556
rect 380360 90930 380388 92550
rect 380052 90902 380388 90930
rect 390020 90930 390048 92618
rect 400864 92608 400916 92614
rect 400864 92550 400916 92556
rect 400312 92540 400364 92546
rect 400312 92482 400364 92488
rect 400772 92540 400824 92546
rect 400772 92482 400824 92488
rect 400324 90930 400352 92482
rect 390020 90902 390356 90930
rect 400324 90902 400660 90930
rect 400784 70666 400812 92482
rect 400876 73846 400904 92550
rect 418344 92540 418396 92546
rect 418344 92482 418396 92488
rect 418356 90916 418384 92482
rect 407224 90222 408066 90250
rect 428674 90222 428780 90250
rect 405648 89752 405700 89758
rect 405648 89694 405700 89700
rect 402978 88768 403034 88777
rect 402978 88703 403034 88712
rect 402992 80345 403020 88703
rect 405660 80345 405688 89694
rect 402978 80336 403034 80345
rect 402978 80271 403034 80280
rect 405646 80336 405702 80345
rect 405646 80271 405702 80280
rect 400864 73840 400916 73846
rect 400864 73782 400916 73788
rect 400660 70638 400812 70666
rect 379716 70094 380052 70122
rect 390356 70094 390508 70122
rect 379716 69018 379744 70094
rect 379704 69012 379756 69018
rect 379704 68954 379756 68960
rect 390480 68814 390508 70094
rect 407224 68950 407252 90222
rect 407764 73840 407816 73846
rect 407764 73782 407816 73788
rect 407776 70666 407804 73782
rect 407776 70638 408066 70666
rect 407212 68944 407264 68950
rect 407212 68886 407264 68892
rect 418356 68882 418384 70108
rect 428660 69018 428688 70108
rect 428648 69012 428700 69018
rect 428648 68954 428700 68960
rect 418344 68876 418396 68882
rect 418344 68818 418396 68824
rect 428752 68814 428780 90222
rect 390468 68808 390520 68814
rect 390468 68750 390520 68756
rect 428740 68808 428792 68814
rect 428740 68750 428792 68756
rect 380348 66428 380400 66434
rect 380348 66370 380400 66376
rect 379612 66292 379664 66298
rect 379612 66234 379664 66240
rect 379624 55214 379652 66234
rect 380360 63852 380388 66370
rect 390652 66360 390704 66366
rect 390652 66302 390704 66308
rect 407120 66360 407172 66366
rect 407120 66302 407172 66308
rect 390664 63852 390692 66302
rect 400982 63294 401088 63322
rect 379624 55186 379928 55214
rect 379900 43738 379928 55186
rect 379900 43710 380374 43738
rect 390664 41342 390692 43044
rect 400968 41410 400996 43044
rect 401060 41410 401088 63294
rect 402978 53816 403034 53825
rect 402978 53751 403034 53760
rect 405646 53816 405702 53825
rect 405646 53751 405702 53760
rect 402992 45393 403020 53751
rect 405660 45393 405688 53751
rect 407132 50386 407160 66302
rect 418620 66292 418672 66298
rect 418620 66234 418672 66240
rect 418632 63852 418660 66234
rect 407224 63294 408342 63322
rect 428950 63306 429148 63322
rect 428950 63300 429160 63306
rect 428950 63294 429108 63300
rect 407120 50380 407172 50386
rect 407120 50322 407172 50328
rect 402978 45384 403034 45393
rect 402978 45319 403034 45328
rect 405646 45384 405702 45393
rect 405646 45319 405702 45328
rect 400956 41404 401008 41410
rect 400956 41346 401008 41352
rect 401048 41404 401100 41410
rect 401048 41346 401100 41352
rect 407224 41342 407252 63294
rect 429108 63242 429160 63248
rect 407948 50380 408000 50386
rect 407948 50322 408000 50328
rect 407960 43738 407988 50322
rect 407960 43710 408342 43738
rect 418632 41342 418660 43044
rect 428936 41410 428964 43044
rect 428924 41404 428976 41410
rect 428924 41346 428976 41352
rect 390652 41336 390704 41342
rect 390652 41278 390704 41284
rect 407212 41336 407264 41342
rect 407212 41278 407264 41284
rect 418620 41336 418672 41342
rect 418620 41278 418672 41284
rect 390008 38752 390060 38758
rect 390008 38694 390060 38700
rect 401048 38752 401100 38758
rect 401048 38694 401100 38700
rect 418344 38752 418396 38758
rect 418344 38694 418396 38700
rect 380348 38684 380400 38690
rect 380348 38626 380400 38632
rect 380360 36938 380388 38626
rect 380052 36910 380388 36938
rect 390020 36938 390048 38694
rect 390020 36910 390356 36938
rect 400660 36502 400996 36530
rect 400772 36236 400824 36242
rect 400772 36178 400824 36184
rect 379704 18624 379756 18630
rect 379704 18566 379756 18572
rect 379716 16674 379744 18566
rect 400784 16674 400812 36178
rect 400864 36168 400916 36174
rect 400864 36110 400916 36116
rect 400876 18630 400904 36110
rect 400864 18624 400916 18630
rect 400864 18566 400916 18572
rect 379716 16646 380052 16674
rect 400660 16646 400812 16674
rect 390356 16102 390508 16130
rect 390480 13802 390508 16102
rect 390468 13796 390520 13802
rect 390468 13738 390520 13744
rect 378784 13320 378836 13326
rect 378784 13262 378836 13268
rect 400968 13258 400996 36502
rect 401060 36242 401088 38694
rect 401140 38684 401192 38690
rect 401140 38626 401192 38632
rect 402244 38684 402296 38690
rect 402244 38626 402296 38632
rect 401048 36236 401100 36242
rect 401048 36178 401100 36184
rect 401152 36174 401180 38626
rect 401140 36168 401192 36174
rect 401140 36110 401192 36116
rect 402256 13802 402284 38626
rect 418356 36924 418384 38694
rect 428648 38684 428700 38690
rect 428648 38626 428700 38632
rect 428740 38684 428792 38690
rect 428740 38626 428792 38632
rect 428660 36924 428688 38626
rect 407224 36230 408066 36258
rect 402978 34776 403034 34785
rect 402978 34711 403034 34720
rect 402992 26353 403020 34711
rect 402978 26344 403034 26353
rect 402978 26279 403034 26288
rect 402244 13796 402296 13802
rect 402244 13738 402296 13744
rect 407224 13326 407252 36230
rect 407764 18624 407816 18630
rect 407764 18566 407816 18572
rect 407776 16674 407804 18566
rect 428752 16674 428780 38626
rect 407776 16646 408066 16674
rect 428674 16646 428780 16674
rect 418356 13433 418384 16116
rect 429212 15162 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 700398 462360 703520
rect 494808 700466 494836 703520
rect 494796 700460 494848 700466
rect 494796 700402 494848 700408
rect 527192 700398 527220 703520
rect 462320 700392 462372 700398
rect 462320 700334 462372 700340
rect 518164 700392 518216 700398
rect 518164 700334 518216 700340
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 464344 687404 464396 687410
rect 464344 687346 464396 687352
rect 485044 687404 485096 687410
rect 485044 687346 485096 687352
rect 457444 687336 457496 687342
rect 457444 687278 457496 687284
rect 429844 687268 429896 687274
rect 429844 687210 429896 687216
rect 456616 687268 456668 687274
rect 456616 687210 456668 687216
rect 429856 662250 429884 687210
rect 456628 684964 456656 687210
rect 446034 684584 446090 684593
rect 446090 684542 446338 684570
rect 446034 684519 446090 684528
rect 434824 684270 436034 684298
rect 430578 674248 430634 674257
rect 430578 674183 430634 674192
rect 434626 674248 434682 674257
rect 434626 674183 434682 674192
rect 430592 665174 430620 674183
rect 434640 665174 434668 674183
rect 430580 665168 430632 665174
rect 430580 665110 430632 665116
rect 434628 665168 434680 665174
rect 434628 665110 434680 665116
rect 434824 662386 434852 684270
rect 457456 673454 457484 687278
rect 464356 684978 464384 687346
rect 474004 687336 474056 687342
rect 474004 687278 474056 687284
rect 464048 684950 464384 684978
rect 474016 684978 474044 687278
rect 484952 687268 485004 687274
rect 484952 687210 485004 687216
rect 474016 684950 474352 684978
rect 484656 684270 484900 684298
rect 484872 683194 484900 684270
rect 484860 683188 484912 683194
rect 484860 683130 484912 683136
rect 484860 682984 484912 682990
rect 484860 682926 484912 682932
rect 484768 677952 484820 677958
rect 484768 677894 484820 677900
rect 462226 674248 462282 674257
rect 462226 674183 462282 674192
rect 458178 673840 458234 673849
rect 458178 673775 458234 673784
rect 457088 673426 457484 673454
rect 457088 664714 457116 673426
rect 458192 665961 458220 673775
rect 462240 665961 462268 674183
rect 458178 665952 458234 665961
rect 458178 665887 458234 665896
rect 462226 665952 462282 665961
rect 462226 665887 462282 665896
rect 484780 664714 484808 677894
rect 456642 664686 457116 664714
rect 484656 664686 484808 664714
rect 434812 662380 434864 662386
rect 434812 662322 434864 662328
rect 436020 662318 436048 664020
rect 436008 662312 436060 662318
rect 436008 662254 436060 662260
rect 446324 662250 446352 664020
rect 463804 664006 464048 664034
rect 474352 664006 474688 664034
rect 463804 662318 463832 664006
rect 474660 662318 474688 664006
rect 463792 662312 463844 662318
rect 463792 662254 463844 662260
rect 474648 662312 474700 662318
rect 474648 662254 474700 662260
rect 484872 662250 484900 682926
rect 484964 677958 484992 687210
rect 484952 677952 485004 677958
rect 484952 677894 485004 677900
rect 485056 667894 485084 687346
rect 502340 687268 502392 687274
rect 502340 687210 502392 687216
rect 512920 687268 512972 687274
rect 512920 687210 512972 687216
rect 502352 684964 502380 687210
rect 491404 684270 492062 684298
rect 512670 684270 512868 684298
rect 487158 674248 487214 674257
rect 487158 674183 487214 674192
rect 489826 674248 489882 674257
rect 489826 674183 489882 674192
rect 485044 667888 485096 667894
rect 485044 667830 485096 667836
rect 487172 665174 487200 674183
rect 489840 665174 489868 674183
rect 487160 665168 487212 665174
rect 487160 665110 487212 665116
rect 489828 665168 489880 665174
rect 489828 665110 489880 665116
rect 491404 662386 491432 684270
rect 512840 683194 512868 684270
rect 512828 683188 512880 683194
rect 512828 683130 512880 683136
rect 512828 682984 512880 682990
rect 512828 682926 512880 682932
rect 512736 682644 512788 682650
rect 512736 682586 512788 682592
rect 491668 667888 491720 667894
rect 491668 667830 491720 667836
rect 491680 664714 491708 667830
rect 512748 664714 512776 682586
rect 491680 664686 492062 664714
rect 512670 664686 512776 664714
rect 491392 662380 491444 662386
rect 491392 662322 491444 662328
rect 502352 662250 502380 664020
rect 512840 662318 512868 682926
rect 512932 682650 512960 687210
rect 512920 682644 512972 682650
rect 512920 682586 512972 682592
rect 514758 674248 514814 674257
rect 514758 674183 514814 674192
rect 514772 665961 514800 674183
rect 514758 665952 514814 665961
rect 514758 665887 514814 665896
rect 512828 662312 512880 662318
rect 512828 662254 512880 662260
rect 429844 662244 429896 662250
rect 429844 662186 429896 662192
rect 446312 662244 446364 662250
rect 446312 662186 446364 662192
rect 484860 662244 484912 662250
rect 484860 662186 484912 662192
rect 502340 662244 502392 662250
rect 502340 662186 502392 662192
rect 446312 659796 446364 659802
rect 446312 659738 446364 659744
rect 491392 659796 491444 659802
rect 491392 659738 491444 659744
rect 429844 659728 429896 659734
rect 429844 659670 429896 659676
rect 436100 659728 436152 659734
rect 436100 659670 436152 659676
rect 429856 634710 429884 659670
rect 436112 657914 436140 659670
rect 446324 657914 446352 659738
rect 463792 659728 463844 659734
rect 463792 659670 463844 659676
rect 436112 657886 436356 657914
rect 446324 657886 446660 657914
rect 456964 657206 457116 657234
rect 430580 656940 430632 656946
rect 430580 656882 430632 656888
rect 434628 656940 434680 656946
rect 434628 656882 434680 656888
rect 430592 647737 430620 656882
rect 434640 647737 434668 656882
rect 430578 647728 430634 647737
rect 430578 647663 430634 647672
rect 434626 647728 434682 647737
rect 434626 647663 434682 647672
rect 436356 637078 436692 637106
rect 446660 637078 446996 637106
rect 436664 634817 436692 637078
rect 436650 634808 436706 634817
rect 436650 634743 436706 634752
rect 446968 634710 446996 637078
rect 456812 637078 456964 637106
rect 456812 634778 456840 637078
rect 457088 634778 457116 657206
rect 463700 655716 463752 655722
rect 463700 655658 463752 655664
rect 456800 634772 456852 634778
rect 456800 634714 456852 634720
rect 457076 634772 457128 634778
rect 457076 634714 457128 634720
rect 463712 634710 463740 655658
rect 463804 654134 463832 659670
rect 474278 657384 474334 657393
rect 474334 657342 474674 657370
rect 474278 657319 474334 657328
rect 464080 657206 464370 657234
rect 484978 657206 485084 657234
rect 464080 655722 464108 657206
rect 464158 656024 464214 656033
rect 464158 655959 464214 655968
rect 464068 655716 464120 655722
rect 464068 655658 464120 655664
rect 463804 654106 464016 654134
rect 463988 637786 464016 654106
rect 464172 648281 464200 655959
rect 464158 648272 464214 648281
rect 464158 648207 464214 648216
rect 463988 637758 464370 637786
rect 474660 634710 474688 637092
rect 484964 634778 484992 637092
rect 485056 634778 485084 657206
rect 487160 656940 487212 656946
rect 487160 656882 487212 656888
rect 489828 656940 489880 656946
rect 489828 656882 489880 656888
rect 487172 647737 487200 656882
rect 489840 647737 489868 656882
rect 491300 655716 491352 655722
rect 491300 655658 491352 655664
rect 487158 647728 487214 647737
rect 487158 647663 487214 647672
rect 489826 647728 489882 647737
rect 489826 647663 489882 647672
rect 484952 634772 485004 634778
rect 484952 634714 485004 634720
rect 485044 634772 485096 634778
rect 485044 634714 485096 634720
rect 491312 634710 491340 655658
rect 491404 654134 491432 659738
rect 502616 659728 502668 659734
rect 502616 659670 502668 659676
rect 502628 657900 502656 659670
rect 492048 657206 492338 657234
rect 512946 657206 513144 657234
rect 492048 655722 492076 657206
rect 492036 655716 492088 655722
rect 492036 655658 492088 655664
rect 491404 654106 491984 654134
rect 491956 637786 491984 654106
rect 491956 637758 492338 637786
rect 502628 634817 502656 637092
rect 502614 634808 502670 634817
rect 512932 634778 512960 637092
rect 513116 634778 513144 657206
rect 514758 656024 514814 656033
rect 514758 655959 514814 655968
rect 514772 647737 514800 655959
rect 514758 647728 514814 647737
rect 514758 647663 514814 647672
rect 502614 634743 502670 634752
rect 512920 634772 512972 634778
rect 512920 634714 512972 634720
rect 513104 634772 513156 634778
rect 513104 634714 513156 634720
rect 429844 634704 429896 634710
rect 429844 634646 429896 634652
rect 446956 634704 447008 634710
rect 446956 634646 447008 634652
rect 463700 634704 463752 634710
rect 463700 634646 463752 634652
rect 474648 634704 474700 634710
rect 474648 634646 474700 634652
rect 491300 634704 491352 634710
rect 491300 634646 491352 634652
rect 464344 632256 464396 632262
rect 464344 632198 464396 632204
rect 485044 632256 485096 632262
rect 485044 632198 485096 632204
rect 457444 632188 457496 632194
rect 457444 632130 457496 632136
rect 429844 632120 429896 632126
rect 429844 632062 429896 632068
rect 456616 632120 456668 632126
rect 456616 632062 456668 632068
rect 429856 608462 429884 632062
rect 456628 630972 456656 632062
rect 446034 630456 446090 630465
rect 446090 630414 446338 630442
rect 446034 630391 446090 630400
rect 434824 630278 436034 630306
rect 430578 620256 430634 620265
rect 430578 620191 430634 620200
rect 434626 620256 434682 620265
rect 434626 620191 434682 620200
rect 430592 611318 430620 620191
rect 434640 611318 434668 620191
rect 430580 611312 430632 611318
rect 430580 611254 430632 611260
rect 434628 611312 434680 611318
rect 434628 611254 434680 611260
rect 434824 608598 434852 630278
rect 457456 615494 457484 632130
rect 464356 630986 464384 632198
rect 474004 632188 474056 632194
rect 474004 632130 474056 632136
rect 464048 630958 464384 630986
rect 474016 630986 474044 632130
rect 484860 632120 484912 632126
rect 484860 632062 484912 632068
rect 474016 630958 474352 630986
rect 484656 630278 484808 630306
rect 458178 620256 458234 620265
rect 458178 620191 458234 620200
rect 462226 620256 462282 620265
rect 462226 620191 462282 620200
rect 457088 615466 457484 615494
rect 457088 610722 457116 615466
rect 458192 611969 458220 620191
rect 462240 611969 462268 620191
rect 458178 611960 458234 611969
rect 458178 611895 458234 611904
rect 462226 611960 462282 611969
rect 462226 611895 462282 611904
rect 484780 610842 484808 630278
rect 484768 610836 484820 610842
rect 484768 610778 484820 610784
rect 456642 610694 457116 610722
rect 484872 610450 484900 632062
rect 485056 613154 485084 632198
rect 502340 632120 502392 632126
rect 502340 632062 502392 632068
rect 514852 632120 514904 632126
rect 514852 632062 514904 632068
rect 502352 630972 502380 632062
rect 512670 630414 513052 630442
rect 491404 630278 492062 630306
rect 487158 620256 487214 620265
rect 487158 620191 487214 620200
rect 489826 620256 489882 620265
rect 489826 620191 489882 620200
rect 485044 613148 485096 613154
rect 485044 613090 485096 613096
rect 487172 611318 487200 620191
rect 489840 611318 489868 620191
rect 487160 611312 487212 611318
rect 487160 611254 487212 611260
rect 489828 611312 489880 611318
rect 489828 611254 489880 611260
rect 484952 610836 485004 610842
rect 484952 610778 485004 610784
rect 484656 610422 484900 610450
rect 434812 608592 434864 608598
rect 434812 608534 434864 608540
rect 436020 608530 436048 610028
rect 436008 608524 436060 608530
rect 436008 608466 436060 608472
rect 446324 608462 446352 610028
rect 463712 610014 464048 610042
rect 474352 610014 474688 610042
rect 463712 608530 463740 610014
rect 474660 608530 474688 610014
rect 463700 608524 463752 608530
rect 463700 608466 463752 608472
rect 474648 608524 474700 608530
rect 474648 608466 474700 608472
rect 484964 608462 484992 610778
rect 491404 608598 491432 630278
rect 512736 628652 512788 628658
rect 512736 628594 512788 628600
rect 491668 613148 491720 613154
rect 491668 613090 491720 613096
rect 491680 610722 491708 613090
rect 512748 610722 512776 628594
rect 513024 621058 513052 630414
rect 514864 628658 514892 632062
rect 514852 628652 514904 628658
rect 514852 628594 514904 628600
rect 491680 610694 492062 610722
rect 512670 610694 512776 610722
rect 512840 621030 513052 621058
rect 491392 608592 491444 608598
rect 491392 608534 491444 608540
rect 502352 608462 502380 610028
rect 512840 608530 512868 621030
rect 514758 620256 514814 620265
rect 514758 620191 514814 620200
rect 514772 611969 514800 620191
rect 514758 611960 514814 611969
rect 514758 611895 514814 611904
rect 512828 608524 512880 608530
rect 512828 608466 512880 608472
rect 429844 608456 429896 608462
rect 429844 608398 429896 608404
rect 446312 608456 446364 608462
rect 446312 608398 446364 608404
rect 484952 608456 485004 608462
rect 484952 608398 485004 608404
rect 502340 608456 502392 608462
rect 502340 608398 502392 608404
rect 446312 605940 446364 605946
rect 446312 605882 446364 605888
rect 463792 605940 463844 605946
rect 463792 605882 463844 605888
rect 502616 605940 502668 605946
rect 502616 605882 502668 605888
rect 514024 605940 514076 605946
rect 514024 605882 514076 605888
rect 429936 605872 429988 605878
rect 429936 605814 429988 605820
rect 436100 605872 436152 605878
rect 436100 605814 436152 605820
rect 429844 603152 429896 603158
rect 429844 603094 429896 603100
rect 429856 580990 429884 603094
rect 429844 580984 429896 580990
rect 429844 580926 429896 580932
rect 429948 580922 429976 605814
rect 436112 603922 436140 605814
rect 446324 603922 446352 605882
rect 457444 605872 457496 605878
rect 457444 605814 457496 605820
rect 436112 603894 436356 603922
rect 446324 603894 446660 603922
rect 456964 603214 457116 603242
rect 434626 602304 434682 602313
rect 434626 602239 434682 602248
rect 430578 602032 430634 602041
rect 430578 601967 430634 601976
rect 430592 593745 430620 601967
rect 434640 593745 434668 602239
rect 430578 593736 430634 593745
rect 430578 593671 430634 593680
rect 434626 593736 434682 593745
rect 434626 593671 434682 593680
rect 436356 583086 436692 583114
rect 446660 583086 446996 583114
rect 436664 580922 436692 583086
rect 429936 580916 429988 580922
rect 429936 580858 429988 580864
rect 436652 580916 436704 580922
rect 436652 580858 436704 580864
rect 446968 580854 446996 583086
rect 456812 583086 456964 583114
rect 456812 580990 456840 583086
rect 457088 580990 457116 603214
rect 456800 580984 456852 580990
rect 456800 580926 456852 580932
rect 457076 580984 457128 580990
rect 457076 580926 457128 580932
rect 457456 580922 457484 605814
rect 462226 602032 462282 602041
rect 462226 601967 462282 601976
rect 462240 593745 462268 601967
rect 463700 599752 463752 599758
rect 463700 599694 463752 599700
rect 462226 593736 462282 593745
rect 462226 593671 462282 593680
rect 457444 580916 457496 580922
rect 457444 580858 457496 580864
rect 463712 580854 463740 599694
rect 463804 596174 463832 605882
rect 474648 605872 474700 605878
rect 474648 605814 474700 605820
rect 491300 605872 491352 605878
rect 491300 605814 491352 605820
rect 474660 603908 474688 605814
rect 464080 603214 464370 603242
rect 484978 603214 485084 603242
rect 464080 599758 464108 603214
rect 464068 599752 464120 599758
rect 464068 599694 464120 599700
rect 463804 596146 464016 596174
rect 463988 583794 464016 596146
rect 463988 583766 464370 583794
rect 474660 580922 474688 583100
rect 484964 580990 484992 583100
rect 485056 580990 485084 603214
rect 485136 585200 485188 585206
rect 485136 585142 485188 585148
rect 484952 580984 485004 580990
rect 484952 580926 485004 580932
rect 485044 580984 485096 580990
rect 485044 580926 485096 580932
rect 485148 580922 485176 585142
rect 491312 584338 491340 605814
rect 502628 603908 502656 605882
rect 491404 603214 492338 603242
rect 512946 603214 513144 603242
rect 491404 585206 491432 603214
rect 491392 585200 491444 585206
rect 491392 585142 491444 585148
rect 491312 584310 491984 584338
rect 491956 583794 491984 584310
rect 491956 583766 492338 583794
rect 502628 580922 502656 583100
rect 512932 580990 512960 583100
rect 513116 580990 513144 603214
rect 512920 580984 512972 580990
rect 512920 580926 512972 580932
rect 513104 580984 513156 580990
rect 513104 580926 513156 580932
rect 514036 580922 514064 605882
rect 514758 602032 514814 602041
rect 514758 601967 514814 601976
rect 514772 593745 514800 601967
rect 514758 593736 514814 593745
rect 514758 593671 514814 593680
rect 474648 580916 474700 580922
rect 474648 580858 474700 580864
rect 485136 580916 485188 580922
rect 485136 580858 485188 580864
rect 502616 580916 502668 580922
rect 502616 580858 502668 580864
rect 514024 580916 514076 580922
rect 514024 580858 514076 580864
rect 446956 580848 447008 580854
rect 446956 580790 447008 580796
rect 463700 580848 463752 580854
rect 463700 580790 463752 580796
rect 457444 578332 457496 578338
rect 457444 578274 457496 578280
rect 474004 578332 474056 578338
rect 474004 578274 474056 578280
rect 484860 578332 484912 578338
rect 484860 578274 484912 578280
rect 502340 578332 502392 578338
rect 502340 578274 502392 578280
rect 429844 578264 429896 578270
rect 429844 578206 429896 578212
rect 456616 578264 456668 578270
rect 456616 578206 456668 578212
rect 429856 554606 429884 578206
rect 456628 576980 456656 578206
rect 446034 576464 446090 576473
rect 446090 576422 446338 576450
rect 446034 576399 446090 576408
rect 434824 576286 436034 576314
rect 430578 566264 430634 566273
rect 430578 566199 430634 566208
rect 434626 566264 434682 566273
rect 434626 566199 434682 566208
rect 430592 557530 430620 566199
rect 434640 557530 434668 566199
rect 430580 557524 430632 557530
rect 430580 557466 430632 557472
rect 434628 557524 434680 557530
rect 434628 557466 434680 557472
rect 434824 554742 434852 576286
rect 457456 557534 457484 578274
rect 464344 578264 464396 578270
rect 464344 578206 464396 578212
rect 464356 576994 464384 578206
rect 464048 576966 464384 576994
rect 474016 576994 474044 578274
rect 474016 576966 474352 576994
rect 484656 576286 484808 576314
rect 458178 574696 458234 574705
rect 458178 574631 458234 574640
rect 462226 574696 462282 574705
rect 462226 574631 462282 574640
rect 458192 566273 458220 574631
rect 462240 566273 462268 574631
rect 458178 566264 458234 566273
rect 458178 566199 458234 566208
rect 462226 566264 462282 566273
rect 462226 566199 462282 566208
rect 457088 557506 457484 557534
rect 457088 556730 457116 557506
rect 484780 556850 484808 576286
rect 484768 556844 484820 556850
rect 484768 556786 484820 556792
rect 456642 556702 457116 556730
rect 484872 556458 484900 578274
rect 485044 578264 485096 578270
rect 485044 578206 485096 578212
rect 485056 558958 485084 578206
rect 502352 576980 502380 578274
rect 512736 578264 512788 578270
rect 512736 578206 512788 578212
rect 512748 576434 512776 578206
rect 512736 576428 512788 576434
rect 512736 576370 512788 576376
rect 491404 576286 492062 576314
rect 512670 576286 512868 576314
rect 487158 566264 487214 566273
rect 487158 566199 487214 566208
rect 489826 566264 489882 566273
rect 489826 566199 489882 566208
rect 485044 558952 485096 558958
rect 485044 558894 485096 558900
rect 487172 557530 487200 566199
rect 489840 557530 489868 566199
rect 487160 557524 487212 557530
rect 487160 557466 487212 557472
rect 489828 557524 489880 557530
rect 489828 557466 489880 557472
rect 484952 556844 485004 556850
rect 484952 556786 485004 556792
rect 484656 556430 484900 556458
rect 434812 554736 434864 554742
rect 434812 554678 434864 554684
rect 436020 554674 436048 556036
rect 436008 554668 436060 554674
rect 436008 554610 436060 554616
rect 446324 554606 446352 556036
rect 463712 556022 464048 556050
rect 474352 556022 474688 556050
rect 463712 554674 463740 556022
rect 474660 554674 474688 556022
rect 463700 554668 463752 554674
rect 463700 554610 463752 554616
rect 474648 554668 474700 554674
rect 474648 554610 474700 554616
rect 484964 554606 484992 556786
rect 491404 554742 491432 576286
rect 512736 576224 512788 576230
rect 512736 576166 512788 576172
rect 491668 558952 491720 558958
rect 491668 558894 491720 558900
rect 491680 556730 491708 558894
rect 512748 556730 512776 576166
rect 491680 556702 492062 556730
rect 512670 556702 512776 556730
rect 491392 554736 491444 554742
rect 491392 554678 491444 554684
rect 502352 554606 502380 556036
rect 512840 554674 512868 576286
rect 514758 574696 514814 574705
rect 514758 574631 514814 574640
rect 514772 566273 514800 574631
rect 514758 566264 514814 566273
rect 514758 566199 514814 566208
rect 512828 554668 512880 554674
rect 512828 554610 512880 554616
rect 429844 554600 429896 554606
rect 429844 554542 429896 554548
rect 446312 554600 446364 554606
rect 446312 554542 446364 554548
rect 484952 554600 485004 554606
rect 484952 554542 485004 554548
rect 502340 554600 502392 554606
rect 502340 554542 502392 554548
rect 429844 552220 429896 552226
rect 429844 552162 429896 552168
rect 436100 552220 436152 552226
rect 436100 552162 436152 552168
rect 429856 527066 429884 552162
rect 436112 549930 436140 552162
rect 446312 552152 446364 552158
rect 446312 552094 446364 552100
rect 457444 552152 457496 552158
rect 457444 552094 457496 552100
rect 474648 552152 474700 552158
rect 474648 552094 474700 552100
rect 491300 552152 491352 552158
rect 491300 552094 491352 552100
rect 446324 549930 446352 552094
rect 436112 549902 436356 549930
rect 446324 549902 446660 549930
rect 429936 549296 429988 549302
rect 429936 549238 429988 549244
rect 429948 527134 429976 549238
rect 456964 549222 457116 549250
rect 430578 548176 430634 548185
rect 430578 548111 430634 548120
rect 434626 548176 434682 548185
rect 434626 548111 434682 548120
rect 430592 539753 430620 548111
rect 434640 539753 434668 548111
rect 430578 539744 430634 539753
rect 430578 539679 430634 539688
rect 434626 539744 434682 539753
rect 434626 539679 434682 539688
rect 436356 529094 436692 529122
rect 446660 529094 446996 529122
rect 429936 527128 429988 527134
rect 429936 527070 429988 527076
rect 436664 527066 436692 529094
rect 429844 527060 429896 527066
rect 429844 527002 429896 527008
rect 436652 527060 436704 527066
rect 436652 527002 436704 527008
rect 446968 526998 446996 529094
rect 456812 529094 456964 529122
rect 456812 527134 456840 529094
rect 457088 527134 457116 549222
rect 456800 527128 456852 527134
rect 456800 527070 456852 527076
rect 457076 527128 457128 527134
rect 457076 527070 457128 527076
rect 457456 527066 457484 552094
rect 463700 552084 463752 552090
rect 463700 552026 463752 552032
rect 458178 548040 458234 548049
rect 458178 547975 458234 547984
rect 462226 548040 462282 548049
rect 462226 547975 462282 547984
rect 458192 539753 458220 547975
rect 462240 539753 462268 547975
rect 458178 539744 458234 539753
rect 458178 539679 458234 539688
rect 462226 539744 462282 539753
rect 462226 539679 462282 539688
rect 463712 533662 463740 552026
rect 474660 549916 474688 552094
rect 463804 549222 464370 549250
rect 484978 549222 485084 549250
rect 463804 538214 463832 549222
rect 463804 538186 463924 538214
rect 463700 533656 463752 533662
rect 463700 533598 463752 533604
rect 463896 528554 463924 538186
rect 464068 533656 464120 533662
rect 464068 533598 464120 533604
rect 464080 529666 464108 533598
rect 464080 529638 464370 529666
rect 463804 528526 463924 528554
rect 457444 527060 457496 527066
rect 457444 527002 457496 527008
rect 463804 526998 463832 528526
rect 474660 527066 474688 529108
rect 484964 527134 484992 529108
rect 485056 527134 485084 549222
rect 489826 548176 489882 548185
rect 489826 548111 489882 548120
rect 489840 539753 489868 548111
rect 489826 539744 489882 539753
rect 489826 539679 489882 539688
rect 491312 531962 491340 552094
rect 502616 552084 502668 552090
rect 502616 552026 502668 552032
rect 502628 549916 502656 552026
rect 514024 550588 514076 550594
rect 514024 550530 514076 550536
rect 491404 549222 492338 549250
rect 512946 549222 513144 549250
rect 491300 531956 491352 531962
rect 491300 531898 491352 531904
rect 484952 527128 485004 527134
rect 484952 527070 485004 527076
rect 485044 527128 485096 527134
rect 485044 527070 485096 527076
rect 491404 527066 491432 549222
rect 492036 531956 492088 531962
rect 492036 531898 492088 531904
rect 492048 529666 492076 531898
rect 492048 529638 492338 529666
rect 502628 527066 502656 529108
rect 512932 527134 512960 529108
rect 513116 527134 513144 549222
rect 512920 527128 512972 527134
rect 512920 527070 512972 527076
rect 513104 527128 513156 527134
rect 513104 527070 513156 527076
rect 514036 527066 514064 550530
rect 514758 548040 514814 548049
rect 514758 547975 514814 547984
rect 514772 539753 514800 547975
rect 514758 539744 514814 539753
rect 514758 539679 514814 539688
rect 474648 527060 474700 527066
rect 474648 527002 474700 527008
rect 491392 527060 491444 527066
rect 491392 527002 491444 527008
rect 502616 527060 502668 527066
rect 502616 527002 502668 527008
rect 514024 527060 514076 527066
rect 514024 527002 514076 527008
rect 446956 526992 447008 526998
rect 446956 526934 447008 526940
rect 463792 526992 463844 526998
rect 463792 526934 463844 526940
rect 464344 524612 464396 524618
rect 464344 524554 464396 524560
rect 485044 524612 485096 524618
rect 485044 524554 485096 524560
rect 457444 524544 457496 524550
rect 457444 524486 457496 524492
rect 429844 524476 429896 524482
rect 429844 524418 429896 524424
rect 456616 524476 456668 524482
rect 456616 524418 456668 524424
rect 429856 500818 429884 524418
rect 456628 522852 456656 524418
rect 446034 522472 446090 522481
rect 446090 522430 446338 522458
rect 446034 522407 446090 522416
rect 434824 522294 436034 522322
rect 434626 520976 434682 520985
rect 434626 520911 434682 520920
rect 430578 520704 430634 520713
rect 430578 520639 430634 520648
rect 430592 512281 430620 520639
rect 434640 512281 434668 520911
rect 430578 512272 430634 512281
rect 430578 512207 430634 512216
rect 434626 512272 434682 512281
rect 434626 512207 434682 512216
rect 434824 500954 434852 522294
rect 457456 509234 457484 524486
rect 464356 522866 464384 524554
rect 474004 524544 474056 524550
rect 474004 524486 474056 524492
rect 464048 522838 464384 522866
rect 474016 522866 474044 524486
rect 484860 524476 484912 524482
rect 484860 524418 484912 524424
rect 474016 522838 474352 522866
rect 484656 522294 484808 522322
rect 458178 520840 458234 520849
rect 458178 520775 458234 520784
rect 458192 512281 458220 520775
rect 463882 520704 463938 520713
rect 463882 520639 463938 520648
rect 463896 518906 463924 520639
rect 462228 518900 462280 518906
rect 462228 518842 462280 518848
rect 463884 518900 463936 518906
rect 463884 518842 463936 518848
rect 462240 512281 462268 518842
rect 458178 512272 458234 512281
rect 458178 512207 458234 512216
rect 462226 512272 462282 512281
rect 462226 512207 462282 512216
rect 457088 509206 457484 509234
rect 457088 502738 457116 509206
rect 484780 502858 484808 522294
rect 484768 502852 484820 502858
rect 484768 502794 484820 502800
rect 456642 502710 457116 502738
rect 484872 502466 484900 524418
rect 485056 505578 485084 524554
rect 502340 524476 502392 524482
rect 502340 524418 502392 524424
rect 514484 524476 514536 524482
rect 514484 524418 514536 524424
rect 502352 522852 502380 524418
rect 512670 522430 513052 522458
rect 491404 522294 492062 522322
rect 512736 522300 512788 522306
rect 485044 505572 485096 505578
rect 485044 505514 485096 505520
rect 484952 502852 485004 502858
rect 484952 502794 485004 502800
rect 484656 502438 484900 502466
rect 434812 500948 434864 500954
rect 434812 500890 434864 500896
rect 436020 500886 436048 502044
rect 436008 500880 436060 500886
rect 436008 500822 436060 500828
rect 446324 500818 446352 502044
rect 463712 502030 464048 502058
rect 474352 502030 474688 502058
rect 463712 500886 463740 502030
rect 474660 500886 474688 502030
rect 463700 500880 463752 500886
rect 463700 500822 463752 500828
rect 474648 500880 474700 500886
rect 474648 500822 474700 500828
rect 484964 500818 484992 502794
rect 491404 500954 491432 522294
rect 512736 522242 512788 522248
rect 491668 505572 491720 505578
rect 491668 505514 491720 505520
rect 491680 502738 491708 505514
rect 512748 502738 512776 522242
rect 513024 514842 513052 522430
rect 514496 522306 514524 524418
rect 514484 522300 514536 522306
rect 514484 522242 514536 522248
rect 514758 520704 514814 520713
rect 514758 520639 514814 520648
rect 491680 502710 492062 502738
rect 512670 502710 512776 502738
rect 512840 514814 513052 514842
rect 491392 500948 491444 500954
rect 491392 500890 491444 500896
rect 502352 500818 502380 502044
rect 512840 500886 512868 514814
rect 514772 512281 514800 520639
rect 514758 512272 514814 512281
rect 514758 512207 514814 512216
rect 512828 500880 512880 500886
rect 512828 500822 512880 500828
rect 429844 500812 429896 500818
rect 429844 500754 429896 500760
rect 446312 500812 446364 500818
rect 446312 500754 446364 500760
rect 484952 500812 485004 500818
rect 484952 500754 485004 500760
rect 502340 500812 502392 500818
rect 502340 500754 502392 500760
rect 446312 498296 446364 498302
rect 446312 498238 446364 498244
rect 457444 498296 457496 498302
rect 457444 498238 457496 498244
rect 474648 498296 474700 498302
rect 474648 498238 474700 498244
rect 491300 498296 491352 498302
rect 491300 498238 491352 498244
rect 429936 498228 429988 498234
rect 429936 498170 429988 498176
rect 436100 498228 436152 498234
rect 436100 498170 436152 498176
rect 429844 495236 429896 495242
rect 429844 495178 429896 495184
rect 429856 473346 429884 495178
rect 429844 473340 429896 473346
rect 429844 473282 429896 473288
rect 429948 473278 429976 498170
rect 436112 495938 436140 498170
rect 446324 495938 446352 498238
rect 436112 495910 436356 495938
rect 446324 495910 446660 495938
rect 456964 495230 457116 495258
rect 430578 485752 430634 485761
rect 430578 485687 430634 485696
rect 434626 485752 434682 485761
rect 434626 485687 434682 485696
rect 430592 477193 430620 485687
rect 434640 477193 434668 485687
rect 430578 477184 430634 477193
rect 430578 477119 430634 477128
rect 434626 477184 434682 477193
rect 434626 477119 434682 477128
rect 436356 475102 436692 475130
rect 446660 475102 446996 475130
rect 436664 473278 436692 475102
rect 429936 473272 429988 473278
rect 429936 473214 429988 473220
rect 436652 473272 436704 473278
rect 436652 473214 436704 473220
rect 446968 473210 446996 475102
rect 456812 475102 456964 475130
rect 456812 473346 456840 475102
rect 457088 473346 457116 495230
rect 456800 473340 456852 473346
rect 456800 473282 456852 473288
rect 457076 473340 457128 473346
rect 457076 473282 457128 473288
rect 457456 473278 457484 498238
rect 463700 498228 463752 498234
rect 463700 498170 463752 498176
rect 458178 485752 458234 485761
rect 458178 485687 458234 485696
rect 462226 485752 462282 485761
rect 462226 485687 462282 485696
rect 458192 477329 458220 485687
rect 462240 477329 462268 485687
rect 463712 485110 463740 498170
rect 474660 495924 474688 498238
rect 463804 495230 464370 495258
rect 484978 495230 485084 495258
rect 463700 485104 463752 485110
rect 463700 485046 463752 485052
rect 458178 477320 458234 477329
rect 458178 477255 458234 477264
rect 462226 477320 462282 477329
rect 462226 477255 462282 477264
rect 457444 473272 457496 473278
rect 457444 473214 457496 473220
rect 463804 473210 463832 495230
rect 463976 485104 464028 485110
rect 463976 485046 464028 485052
rect 463988 475674 464016 485046
rect 463988 475646 464370 475674
rect 474660 473278 474688 475116
rect 484964 473346 484992 475116
rect 485056 473346 485084 495230
rect 489826 485752 489882 485761
rect 489826 485687 489882 485696
rect 489840 477193 489868 485687
rect 491312 477698 491340 498238
rect 502616 498228 502668 498234
rect 502616 498170 502668 498176
rect 514024 498228 514076 498234
rect 514024 498170 514076 498176
rect 502628 495924 502656 498170
rect 491404 495230 492338 495258
rect 512946 495230 513144 495258
rect 491300 477692 491352 477698
rect 491300 477634 491352 477640
rect 489826 477184 489882 477193
rect 489826 477119 489882 477128
rect 484952 473340 485004 473346
rect 484952 473282 485004 473288
rect 485044 473340 485096 473346
rect 485044 473282 485096 473288
rect 491404 473278 491432 495230
rect 492036 477692 492088 477698
rect 492036 477634 492088 477640
rect 492048 475674 492076 477634
rect 492048 475646 492338 475674
rect 502628 473278 502656 475116
rect 512932 473346 512960 475116
rect 513116 473346 513144 495230
rect 512920 473340 512972 473346
rect 512920 473282 512972 473288
rect 513104 473340 513156 473346
rect 513104 473282 513156 473288
rect 514036 473278 514064 498170
rect 514758 485752 514814 485761
rect 514758 485687 514814 485696
rect 514772 477329 514800 485687
rect 514758 477320 514814 477329
rect 514758 477255 514814 477264
rect 474648 473272 474700 473278
rect 474648 473214 474700 473220
rect 491392 473272 491444 473278
rect 491392 473214 491444 473220
rect 502616 473272 502668 473278
rect 502616 473214 502668 473220
rect 514024 473272 514076 473278
rect 514024 473214 514076 473220
rect 446956 473204 447008 473210
rect 446956 473146 447008 473152
rect 463792 473204 463844 473210
rect 463792 473146 463844 473152
rect 464344 470824 464396 470830
rect 464344 470766 464396 470772
rect 485044 470824 485096 470830
rect 485044 470766 485096 470772
rect 457536 470756 457588 470762
rect 457536 470698 457588 470704
rect 446034 468480 446090 468489
rect 456338 468480 456394 468489
rect 446090 468438 446338 468466
rect 446034 468415 446090 468424
rect 456394 468438 456642 468466
rect 456338 468415 456394 468424
rect 434824 468302 436034 468330
rect 430578 466712 430634 466721
rect 430578 466647 430634 466656
rect 430592 458289 430620 466647
rect 430578 458280 430634 458289
rect 430578 458215 430634 458224
rect 434824 445738 434852 468302
rect 457548 451274 457576 470698
rect 464356 468874 464384 470766
rect 474004 470756 474056 470762
rect 474004 470698 474056 470704
rect 464048 468846 464384 468874
rect 474016 468874 474044 470698
rect 484860 470688 484912 470694
rect 484860 470630 484912 470636
rect 474016 468846 474352 468874
rect 484656 468302 484808 468330
rect 458178 466984 458234 466993
rect 458178 466919 458234 466928
rect 458192 458289 458220 466919
rect 462226 466712 462282 466721
rect 462226 466647 462282 466656
rect 462240 458289 462268 466647
rect 458178 458280 458234 458289
rect 458178 458215 458234 458224
rect 462226 458280 462282 458289
rect 462226 458215 462282 458224
rect 457088 451246 457576 451274
rect 457088 448746 457116 451246
rect 484780 448866 484808 468302
rect 484768 448860 484820 448866
rect 484768 448802 484820 448808
rect 456642 448718 457116 448746
rect 484872 448474 484900 470630
rect 485056 451314 485084 470766
rect 502340 470688 502392 470694
rect 502340 470630 502392 470636
rect 512736 470688 512788 470694
rect 512736 470630 512788 470636
rect 502352 468860 502380 470630
rect 512748 468450 512776 470630
rect 512736 468444 512788 468450
rect 512736 468386 512788 468392
rect 491404 468302 492062 468330
rect 512670 468302 512868 468330
rect 487158 466848 487214 466857
rect 487158 466783 487214 466792
rect 487172 458289 487200 466783
rect 487158 458280 487214 458289
rect 487158 458215 487214 458224
rect 485044 451308 485096 451314
rect 485044 451250 485096 451256
rect 484952 448860 485004 448866
rect 484952 448802 485004 448808
rect 484656 448446 484900 448474
rect 434812 445732 434864 445738
rect 434812 445674 434864 445680
rect 436020 445670 436048 448052
rect 436008 445664 436060 445670
rect 436008 445606 436060 445612
rect 446324 445602 446352 448052
rect 463712 448038 464048 448066
rect 474352 448038 474688 448066
rect 463712 445670 463740 448038
rect 474660 445670 474688 448038
rect 463700 445664 463752 445670
rect 463700 445606 463752 445612
rect 474648 445664 474700 445670
rect 474648 445606 474700 445612
rect 484964 445602 484992 448802
rect 491404 445738 491432 468302
rect 512736 468240 512788 468246
rect 512736 468182 512788 468188
rect 491668 451308 491720 451314
rect 491668 451250 491720 451256
rect 491680 448746 491708 451250
rect 512748 448746 512776 468182
rect 491680 448718 492062 448746
rect 512670 448718 512776 448746
rect 491392 445732 491444 445738
rect 491392 445674 491444 445680
rect 502352 445602 502380 448052
rect 512840 445670 512868 468302
rect 514758 466712 514814 466721
rect 514758 466647 514814 466656
rect 514772 458289 514800 466647
rect 514758 458280 514814 458289
rect 514758 458215 514814 458224
rect 512828 445664 512880 445670
rect 512828 445606 512880 445612
rect 446312 445596 446364 445602
rect 446312 445538 446364 445544
rect 484952 445596 485004 445602
rect 484952 445538 485004 445544
rect 502340 445596 502392 445602
rect 502340 445538 502392 445544
rect 446312 444508 446364 444514
rect 446312 444450 446364 444456
rect 457444 444508 457496 444514
rect 457444 444450 457496 444456
rect 474648 444508 474700 444514
rect 474648 444450 474700 444456
rect 491392 444508 491444 444514
rect 491392 444450 491444 444456
rect 446324 441946 446352 444450
rect 446324 441918 446660 441946
rect 429844 441652 429896 441658
rect 429844 441594 429896 441600
rect 429856 419490 429884 441594
rect 436112 441238 436356 441266
rect 456964 441238 457116 441266
rect 430578 431760 430634 431769
rect 430578 431695 430634 431704
rect 434626 431760 434682 431769
rect 434626 431695 434682 431704
rect 430592 423337 430620 431695
rect 430578 423328 430634 423337
rect 430578 423263 430634 423272
rect 434640 423065 434668 431695
rect 434626 423056 434682 423065
rect 434626 422991 434682 423000
rect 429844 419484 429896 419490
rect 429844 419426 429896 419432
rect 436112 419422 436140 441238
rect 436356 421110 436692 421138
rect 446660 421110 446996 421138
rect 436664 419422 436692 421110
rect 436100 419416 436152 419422
rect 436100 419358 436152 419364
rect 436652 419416 436704 419422
rect 436652 419358 436704 419364
rect 446968 419354 446996 421110
rect 456812 421110 456964 421138
rect 456812 419490 456840 421110
rect 457088 419490 457116 441238
rect 456800 419484 456852 419490
rect 456800 419426 456852 419432
rect 457076 419484 457128 419490
rect 457076 419426 457128 419432
rect 457456 419422 457484 444450
rect 463792 444440 463844 444446
rect 463792 444382 463844 444388
rect 463804 441614 463832 444382
rect 474660 441932 474688 444450
rect 491404 441614 491432 444450
rect 502616 444440 502668 444446
rect 502616 444382 502668 444388
rect 514024 444440 514076 444446
rect 514024 444382 514076 444388
rect 502628 441932 502656 444382
rect 463804 441586 464016 441614
rect 491404 441586 491984 441614
rect 457536 439544 457588 439550
rect 457536 439486 457588 439492
rect 457444 419416 457496 419422
rect 457444 419358 457496 419364
rect 457548 419354 457576 439486
rect 462226 431760 462282 431769
rect 462226 431695 462282 431704
rect 462240 423337 462268 431695
rect 462226 423328 462282 423337
rect 462226 423263 462282 423272
rect 463988 421682 464016 441586
rect 464080 441238 464370 441266
rect 484978 441238 485084 441266
rect 464080 439550 464108 441238
rect 464068 439544 464120 439550
rect 464068 439486 464120 439492
rect 463988 421654 464370 421682
rect 474660 419422 474688 421124
rect 484964 419490 484992 421124
rect 485056 419490 485084 441238
rect 485136 438932 485188 438938
rect 485136 438874 485188 438880
rect 484952 419484 485004 419490
rect 484952 419426 485004 419432
rect 485044 419484 485096 419490
rect 485044 419426 485096 419432
rect 485148 419422 485176 438874
rect 491956 421682 491984 441586
rect 492048 441238 492338 441266
rect 512946 441238 513144 441266
rect 492048 438938 492076 441238
rect 492036 438932 492088 438938
rect 492036 438874 492088 438880
rect 491956 421654 492338 421682
rect 502628 419422 502656 421124
rect 512932 419490 512960 421124
rect 513116 419490 513144 441238
rect 512920 419484 512972 419490
rect 512920 419426 512972 419432
rect 513104 419484 513156 419490
rect 513104 419426 513156 419432
rect 514036 419422 514064 444382
rect 514758 431760 514814 431769
rect 514758 431695 514814 431704
rect 514772 423337 514800 431695
rect 514758 423328 514814 423337
rect 514758 423263 514814 423272
rect 474648 419416 474700 419422
rect 474648 419358 474700 419364
rect 485136 419416 485188 419422
rect 485136 419358 485188 419364
rect 502616 419416 502668 419422
rect 502616 419358 502668 419364
rect 514024 419416 514076 419422
rect 514024 419358 514076 419364
rect 446956 419348 447008 419354
rect 446956 419290 447008 419296
rect 457536 419348 457588 419354
rect 457536 419290 457588 419296
rect 464344 416968 464396 416974
rect 464344 416910 464396 416916
rect 485044 416968 485096 416974
rect 485044 416910 485096 416916
rect 457444 416900 457496 416906
rect 457444 416842 457496 416848
rect 446034 414488 446090 414497
rect 456338 414488 456394 414497
rect 446090 414446 446338 414474
rect 446034 414423 446090 414432
rect 456394 414446 456642 414474
rect 456338 414423 456394 414432
rect 434824 414310 436034 414338
rect 430578 404288 430634 404297
rect 430578 404223 430634 404232
rect 430592 395865 430620 404223
rect 430578 395856 430634 395865
rect 430578 395791 430634 395800
rect 434824 391950 434852 414310
rect 457456 402974 457484 416842
rect 464356 414882 464384 416910
rect 474004 416900 474056 416906
rect 474004 416842 474056 416848
rect 464048 414854 464384 414882
rect 474016 414882 474044 416842
rect 484860 416832 484912 416838
rect 484860 416774 484912 416780
rect 474016 414854 474352 414882
rect 484656 414310 484808 414338
rect 458178 404288 458234 404297
rect 458178 404223 458234 404232
rect 462226 404288 462282 404297
rect 462226 404223 462282 404232
rect 457088 402946 457484 402974
rect 457088 394618 457116 402946
rect 458192 396001 458220 404223
rect 462240 396001 462268 404223
rect 458178 395992 458234 396001
rect 458178 395927 458234 395936
rect 462226 395992 462282 396001
rect 462226 395927 462282 395936
rect 484780 394874 484808 414310
rect 484768 394868 484820 394874
rect 484768 394810 484820 394816
rect 484872 394754 484900 416774
rect 485056 397458 485084 416910
rect 502340 416832 502392 416838
rect 502340 416774 502392 416780
rect 512920 416832 512972 416838
rect 512920 416774 512972 416780
rect 502352 414868 502380 416774
rect 491404 414310 492062 414338
rect 512670 414310 512868 414338
rect 487158 404288 487214 404297
rect 487158 404223 487214 404232
rect 485044 397452 485096 397458
rect 485044 397394 485096 397400
rect 487172 395865 487200 404223
rect 487158 395856 487214 395865
rect 487158 395791 487214 395800
rect 484656 394726 484900 394754
rect 456642 394590 457116 394618
rect 484768 394664 484820 394670
rect 484768 394606 484820 394612
rect 434812 391944 434864 391950
rect 434812 391886 434864 391892
rect 436020 391882 436048 394060
rect 436008 391876 436060 391882
rect 436008 391818 436060 391824
rect 446324 391814 446352 394060
rect 463804 394046 464048 394074
rect 474352 394046 474688 394074
rect 463804 391882 463832 394046
rect 474660 391882 474688 394046
rect 463792 391876 463844 391882
rect 463792 391818 463844 391824
rect 474648 391876 474700 391882
rect 474648 391818 474700 391824
rect 484780 391814 484808 394606
rect 491404 391950 491432 414310
rect 512736 412888 512788 412894
rect 512736 412830 512788 412836
rect 491668 397452 491720 397458
rect 491668 397394 491720 397400
rect 491680 394754 491708 397394
rect 512748 394754 512776 412830
rect 512840 412826 512868 414310
rect 512932 412894 512960 416774
rect 512920 412888 512972 412894
rect 512920 412830 512972 412836
rect 512828 412820 512880 412826
rect 512828 412762 512880 412768
rect 512828 412616 512880 412622
rect 512828 412558 512880 412564
rect 491680 394726 492062 394754
rect 512670 394726 512776 394754
rect 491392 391944 491444 391950
rect 491392 391886 491444 391892
rect 502352 391814 502380 394060
rect 512840 391882 512868 412558
rect 514758 404288 514814 404297
rect 514758 404223 514814 404232
rect 514772 396001 514800 404223
rect 514758 395992 514814 396001
rect 514758 395927 514814 395936
rect 512828 391876 512880 391882
rect 512828 391818 512880 391824
rect 446312 391808 446364 391814
rect 446312 391750 446364 391756
rect 484768 391808 484820 391814
rect 484768 391750 484820 391756
rect 502340 391808 502392 391814
rect 502340 391750 502392 391756
rect 446312 389292 446364 389298
rect 446312 389234 446364 389240
rect 457444 389292 457496 389298
rect 457444 389234 457496 389240
rect 474648 389292 474700 389298
rect 474648 389234 474700 389240
rect 491392 389292 491444 389298
rect 491392 389234 491444 389240
rect 429844 389224 429896 389230
rect 429844 389166 429896 389172
rect 436100 389224 436152 389230
rect 436100 389166 436152 389172
rect 429856 365634 429884 389166
rect 436112 387954 436140 389166
rect 446324 387954 446352 389234
rect 436112 387926 436356 387954
rect 446324 387926 446660 387954
rect 456964 387246 457116 387274
rect 429936 386436 429988 386442
rect 429936 386378 429988 386384
rect 429948 365702 429976 386378
rect 430578 377768 430634 377777
rect 430578 377703 430634 377712
rect 434626 377768 434682 377777
rect 434626 377703 434682 377712
rect 430592 368490 430620 377703
rect 434640 368490 434668 377703
rect 430580 368484 430632 368490
rect 430580 368426 430632 368432
rect 434628 368484 434680 368490
rect 434628 368426 434680 368432
rect 436356 367118 436692 367146
rect 446660 367118 446996 367146
rect 429936 365696 429988 365702
rect 429936 365638 429988 365644
rect 436664 365634 436692 367118
rect 429844 365628 429896 365634
rect 429844 365570 429896 365576
rect 436652 365628 436704 365634
rect 436652 365570 436704 365576
rect 446968 365566 446996 367118
rect 456812 367118 456964 367146
rect 456812 365702 456840 367118
rect 457088 365702 457116 387246
rect 456800 365696 456852 365702
rect 456800 365638 456852 365644
rect 457076 365696 457128 365702
rect 457076 365638 457128 365644
rect 457456 365634 457484 389234
rect 463700 389224 463752 389230
rect 463700 389166 463752 389172
rect 463712 378826 463740 389166
rect 474660 387940 474688 389234
rect 463804 387246 464370 387274
rect 484978 387246 485084 387274
rect 463700 378820 463752 378826
rect 463700 378762 463752 378768
rect 462226 377768 462282 377777
rect 462226 377703 462282 377712
rect 462240 369345 462268 377703
rect 462226 369336 462282 369345
rect 462226 369271 462282 369280
rect 457444 365628 457496 365634
rect 457444 365570 457496 365576
rect 463804 365566 463832 387246
rect 463976 378820 464028 378826
rect 463976 378762 464028 378768
rect 463988 367690 464016 378762
rect 463988 367662 464370 367690
rect 474660 365634 474688 367132
rect 484964 365702 484992 367132
rect 485056 365702 485084 387246
rect 491300 385484 491352 385490
rect 491300 385426 491352 385432
rect 487158 377768 487214 377777
rect 487158 377703 487214 377712
rect 489826 377768 489882 377777
rect 489826 377703 489882 377712
rect 487172 368490 487200 377703
rect 489840 368490 489868 377703
rect 487160 368484 487212 368490
rect 487160 368426 487212 368432
rect 489828 368484 489880 368490
rect 489828 368426 489880 368432
rect 484952 365696 485004 365702
rect 484952 365638 485004 365644
rect 485044 365696 485096 365702
rect 485044 365638 485096 365644
rect 491312 365634 491340 385426
rect 491404 383654 491432 389234
rect 502616 389224 502668 389230
rect 502616 389166 502668 389172
rect 514024 389224 514076 389230
rect 514024 389166 514076 389172
rect 502628 387940 502656 389166
rect 492048 387246 492338 387274
rect 512946 387246 513144 387274
rect 492048 385490 492076 387246
rect 492036 385484 492088 385490
rect 492036 385426 492088 385432
rect 491404 383626 491984 383654
rect 491956 367690 491984 383626
rect 491956 367662 492338 367690
rect 502628 365634 502656 367132
rect 512932 365702 512960 367132
rect 513116 365702 513144 387246
rect 512920 365696 512972 365702
rect 512920 365638 512972 365644
rect 513104 365696 513156 365702
rect 513104 365638 513156 365644
rect 514036 365634 514064 389166
rect 514758 377768 514814 377777
rect 514758 377703 514814 377712
rect 514772 369345 514800 377703
rect 514758 369336 514814 369345
rect 514758 369271 514814 369280
rect 474648 365628 474700 365634
rect 474648 365570 474700 365576
rect 491300 365628 491352 365634
rect 491300 365570 491352 365576
rect 502616 365628 502668 365634
rect 502616 365570 502668 365576
rect 514024 365628 514076 365634
rect 514024 365570 514076 365576
rect 446956 365560 447008 365566
rect 446956 365502 447008 365508
rect 463792 365560 463844 365566
rect 463792 365502 463844 365508
rect 464344 363112 464396 363118
rect 464344 363054 464396 363060
rect 485044 363112 485096 363118
rect 485044 363054 485096 363060
rect 457444 363044 457496 363050
rect 457444 362986 457496 362992
rect 429844 362976 429896 362982
rect 429844 362918 429896 362924
rect 456616 362976 456668 362982
rect 456616 362918 456668 362924
rect 429856 337958 429884 362918
rect 456628 360876 456656 362918
rect 446034 360496 446090 360505
rect 446090 360454 446338 360482
rect 446034 360431 446090 360440
rect 434824 360318 436034 360346
rect 430578 350296 430634 350305
rect 430578 350231 430634 350240
rect 430592 341873 430620 350231
rect 430578 341864 430634 341873
rect 430578 341799 430634 341808
rect 434824 338094 434852 360318
rect 457456 345014 457484 362986
rect 464356 360890 464384 363054
rect 474004 363044 474056 363050
rect 474004 362986 474056 362992
rect 464048 360862 464384 360890
rect 474016 360890 474044 362986
rect 484952 362976 485004 362982
rect 484952 362918 485004 362924
rect 474016 360862 474352 360890
rect 484656 360590 484900 360618
rect 484872 355434 484900 360590
rect 484860 355428 484912 355434
rect 484860 355370 484912 355376
rect 484860 355224 484912 355230
rect 484860 355166 484912 355172
rect 484768 352300 484820 352306
rect 484768 352242 484820 352248
rect 458178 350296 458234 350305
rect 458178 350231 458234 350240
rect 462226 350296 462282 350305
rect 462226 350231 462282 350240
rect 457088 344986 457484 345014
rect 457088 340762 457116 344986
rect 458192 342009 458220 350231
rect 462240 342009 462268 350231
rect 458178 342000 458234 342009
rect 458178 341935 458234 341944
rect 462226 342000 462282 342009
rect 462226 341935 462282 341944
rect 484780 340762 484808 352242
rect 456642 340734 457116 340762
rect 484656 340734 484808 340762
rect 434812 338088 434864 338094
rect 434812 338030 434864 338036
rect 436020 338026 436048 340068
rect 436008 338020 436060 338026
rect 436008 337962 436060 337968
rect 446324 337958 446352 340068
rect 463712 340054 464048 340082
rect 474352 340054 474688 340082
rect 463712 338026 463740 340054
rect 474660 338026 474688 340054
rect 463700 338020 463752 338026
rect 463700 337962 463752 337968
rect 474648 338020 474700 338026
rect 474648 337962 474700 337968
rect 484872 337958 484900 355166
rect 484964 352306 484992 362918
rect 484952 352300 485004 352306
rect 484952 352242 485004 352248
rect 485056 342650 485084 363054
rect 502340 362976 502392 362982
rect 502340 362918 502392 362924
rect 512920 362976 512972 362982
rect 512920 362918 512972 362924
rect 502352 360876 502380 362918
rect 512670 360590 512868 360618
rect 491404 360318 492062 360346
rect 487158 350296 487214 350305
rect 487158 350231 487214 350240
rect 485044 342644 485096 342650
rect 485044 342586 485096 342592
rect 487172 341873 487200 350231
rect 487158 341864 487214 341873
rect 487158 341799 487214 341808
rect 491404 338094 491432 360318
rect 512840 355434 512868 360590
rect 512828 355428 512880 355434
rect 512828 355370 512880 355376
rect 512932 352594 512960 362918
rect 513012 355428 513064 355434
rect 513012 355370 513064 355376
rect 512748 352566 512960 352594
rect 491668 342644 491720 342650
rect 491668 342586 491720 342592
rect 491680 340762 491708 342586
rect 512748 340762 512776 352566
rect 513024 347818 513052 355370
rect 514758 350296 514814 350305
rect 514758 350231 514814 350240
rect 512828 347812 512880 347818
rect 512828 347754 512880 347760
rect 513012 347812 513064 347818
rect 513012 347754 513064 347760
rect 491680 340734 492062 340762
rect 512670 340734 512776 340762
rect 491392 338088 491444 338094
rect 491392 338030 491444 338036
rect 502352 337958 502380 340068
rect 512840 338026 512868 347754
rect 514772 342009 514800 350231
rect 514758 342000 514814 342009
rect 514758 341935 514814 341944
rect 512828 338020 512880 338026
rect 512828 337962 512880 337968
rect 429844 337952 429896 337958
rect 429844 337894 429896 337900
rect 446312 337952 446364 337958
rect 446312 337894 446364 337900
rect 484860 337952 484912 337958
rect 484860 337894 484912 337900
rect 502340 337952 502392 337958
rect 502340 337894 502392 337900
rect 429844 335504 429896 335510
rect 429844 335446 429896 335452
rect 436100 335504 436152 335510
rect 436100 335446 436152 335452
rect 429856 311778 429884 335446
rect 436112 333962 436140 335446
rect 446312 335436 446364 335442
rect 446312 335378 446364 335384
rect 457444 335436 457496 335442
rect 457444 335378 457496 335384
rect 474648 335436 474700 335442
rect 474648 335378 474700 335384
rect 491392 335436 491444 335442
rect 491392 335378 491444 335384
rect 446324 333962 446352 335378
rect 436112 333934 436356 333962
rect 446324 333934 446660 333962
rect 456964 333254 457116 333282
rect 430580 332716 430632 332722
rect 430580 332658 430632 332664
rect 429936 332648 429988 332654
rect 429936 332590 429988 332596
rect 429948 311846 429976 332590
rect 430592 323785 430620 332658
rect 434628 332648 434680 332654
rect 434628 332590 434680 332596
rect 434640 323785 434668 332590
rect 430578 323776 430634 323785
rect 430578 323711 430634 323720
rect 434626 323776 434682 323785
rect 434626 323711 434682 323720
rect 436356 313126 436692 313154
rect 446660 313126 446996 313154
rect 429936 311840 429988 311846
rect 429936 311782 429988 311788
rect 436664 311778 436692 313126
rect 429844 311772 429896 311778
rect 429844 311714 429896 311720
rect 436652 311772 436704 311778
rect 436652 311714 436704 311720
rect 446968 311710 446996 313126
rect 456812 313126 456964 313154
rect 456812 311846 456840 313126
rect 457088 311846 457116 333254
rect 456800 311840 456852 311846
rect 456800 311782 456852 311788
rect 457076 311840 457128 311846
rect 457076 311782 457128 311788
rect 457456 311778 457484 335378
rect 463792 335368 463844 335374
rect 463792 335310 463844 335316
rect 463700 325780 463752 325786
rect 463700 325722 463752 325728
rect 462226 323776 462282 323785
rect 462226 323711 462282 323720
rect 462240 315353 462268 323711
rect 462226 315344 462282 315353
rect 462226 315279 462282 315288
rect 457444 311772 457496 311778
rect 457444 311714 457496 311720
rect 463712 311710 463740 325722
rect 463804 325694 463832 335310
rect 474660 333948 474688 335378
rect 464080 333254 464370 333282
rect 484978 333254 485084 333282
rect 464080 325786 464108 333254
rect 464068 325780 464120 325786
rect 464068 325722 464120 325728
rect 463804 325666 464016 325694
rect 463988 313698 464016 325666
rect 463988 313670 464370 313698
rect 474660 311778 474688 313140
rect 484964 311846 484992 313140
rect 485056 311846 485084 333254
rect 487160 332648 487212 332654
rect 487160 332590 487212 332596
rect 489828 332648 489880 332654
rect 489828 332590 489880 332596
rect 487172 323785 487200 332590
rect 489840 323785 489868 332590
rect 491300 329520 491352 329526
rect 491300 329462 491352 329468
rect 487158 323776 487214 323785
rect 487158 323711 487214 323720
rect 489826 323776 489882 323785
rect 489826 323711 489882 323720
rect 484952 311840 485004 311846
rect 484952 311782 485004 311788
rect 485044 311840 485096 311846
rect 485044 311782 485096 311788
rect 491312 311778 491340 329462
rect 491404 325694 491432 335378
rect 502616 335368 502668 335374
rect 502616 335310 502668 335316
rect 514024 335368 514076 335374
rect 514024 335310 514076 335316
rect 502628 333948 502656 335310
rect 492048 333254 492338 333282
rect 512946 333254 513144 333282
rect 492048 329526 492076 333254
rect 492036 329520 492088 329526
rect 492036 329462 492088 329468
rect 491404 325666 491984 325694
rect 491956 313698 491984 325666
rect 491956 313670 492338 313698
rect 502628 311778 502656 313140
rect 512932 311846 512960 313140
rect 513116 311846 513144 333254
rect 512920 311840 512972 311846
rect 512920 311782 512972 311788
rect 513104 311840 513156 311846
rect 513104 311782 513156 311788
rect 514036 311778 514064 335310
rect 514758 323776 514814 323785
rect 514758 323711 514814 323720
rect 514772 315353 514800 323711
rect 514758 315344 514814 315353
rect 514758 315279 514814 315288
rect 474648 311772 474700 311778
rect 474648 311714 474700 311720
rect 491300 311772 491352 311778
rect 491300 311714 491352 311720
rect 502616 311772 502668 311778
rect 502616 311714 502668 311720
rect 514024 311772 514076 311778
rect 514024 311714 514076 311720
rect 446956 311704 447008 311710
rect 446956 311646 447008 311652
rect 463700 311704 463752 311710
rect 463700 311646 463752 311652
rect 464344 309324 464396 309330
rect 464344 309266 464396 309272
rect 485044 309324 485096 309330
rect 485044 309266 485096 309272
rect 457444 309256 457496 309262
rect 457444 309198 457496 309204
rect 429844 309188 429896 309194
rect 429844 309130 429896 309136
rect 456616 309188 456668 309194
rect 456616 309130 456668 309136
rect 429856 284170 429884 309130
rect 456628 306884 456656 309130
rect 446034 306504 446090 306513
rect 446090 306462 446338 306490
rect 446034 306439 446090 306448
rect 434824 306326 436034 306354
rect 430578 296304 430634 296313
rect 430578 296239 430634 296248
rect 434626 296304 434682 296313
rect 434626 296239 434682 296248
rect 430592 288017 430620 296239
rect 430578 288008 430634 288017
rect 430578 287943 430634 287952
rect 434640 287745 434668 296239
rect 434626 287736 434682 287745
rect 434626 287671 434682 287680
rect 434824 284306 434852 306326
rect 457456 287054 457484 309198
rect 464356 306898 464384 309266
rect 474004 309256 474056 309262
rect 474004 309198 474056 309204
rect 464048 306870 464384 306898
rect 474016 306898 474044 309198
rect 484952 309188 485004 309194
rect 484952 309130 485004 309136
rect 474016 306870 474352 306898
rect 484656 306326 484808 306354
rect 484780 305794 484808 306326
rect 484768 305788 484820 305794
rect 484768 305730 484820 305736
rect 484860 305584 484912 305590
rect 484860 305526 484912 305532
rect 484768 302728 484820 302734
rect 484768 302670 484820 302676
rect 458178 296304 458234 296313
rect 458178 296239 458234 296248
rect 462226 296304 462282 296313
rect 462226 296239 462282 296248
rect 458192 287881 458220 296239
rect 462240 288017 462268 296239
rect 462226 288008 462282 288017
rect 462226 287943 462282 287952
rect 458178 287872 458234 287881
rect 458178 287807 458234 287816
rect 457088 287026 457484 287054
rect 457088 286770 457116 287026
rect 484780 286770 484808 302670
rect 456642 286742 457116 286770
rect 484656 286742 484808 286770
rect 434812 284300 434864 284306
rect 434812 284242 434864 284248
rect 436020 284238 436048 286076
rect 436008 284232 436060 284238
rect 436008 284174 436060 284180
rect 446324 284170 446352 286076
rect 463712 286062 464048 286090
rect 474352 286062 474688 286090
rect 463712 284238 463740 286062
rect 474660 284238 474688 286062
rect 463700 284232 463752 284238
rect 463700 284174 463752 284180
rect 474648 284232 474700 284238
rect 474648 284174 474700 284180
rect 484872 284170 484900 305526
rect 484964 302734 484992 309130
rect 484952 302728 485004 302734
rect 484952 302670 485004 302676
rect 485056 288454 485084 309266
rect 502340 309188 502392 309194
rect 502340 309130 502392 309136
rect 512920 309188 512972 309194
rect 512920 309130 512972 309136
rect 502352 306884 502380 309130
rect 491404 306326 492062 306354
rect 512670 306326 512776 306354
rect 485044 288448 485096 288454
rect 485044 288390 485096 288396
rect 491404 284306 491432 306326
rect 512748 305794 512776 306326
rect 512736 305788 512788 305794
rect 512736 305730 512788 305736
rect 512828 305584 512880 305590
rect 512828 305526 512880 305532
rect 512736 304632 512788 304638
rect 512736 304574 512788 304580
rect 491668 288448 491720 288454
rect 491668 288390 491720 288396
rect 491680 286770 491708 288390
rect 512748 286770 512776 304574
rect 491680 286742 492062 286770
rect 512670 286742 512776 286770
rect 491392 284300 491444 284306
rect 491392 284242 491444 284248
rect 502352 284170 502380 286076
rect 512840 284238 512868 305526
rect 512932 304638 512960 309130
rect 512920 304632 512972 304638
rect 512920 304574 512972 304580
rect 514758 296304 514814 296313
rect 514758 296239 514814 296248
rect 514772 288017 514800 296239
rect 514758 288008 514814 288017
rect 514758 287943 514814 287952
rect 512828 284232 512880 284238
rect 512828 284174 512880 284180
rect 429844 284164 429896 284170
rect 429844 284106 429896 284112
rect 446312 284164 446364 284170
rect 446312 284106 446364 284112
rect 484860 284164 484912 284170
rect 484860 284106 484912 284112
rect 502340 284164 502392 284170
rect 502340 284106 502392 284112
rect 446312 281648 446364 281654
rect 446312 281590 446364 281596
rect 491392 281648 491444 281654
rect 491392 281590 491444 281596
rect 429936 281580 429988 281586
rect 429936 281522 429988 281528
rect 436100 281580 436152 281586
rect 436100 281522 436152 281528
rect 429948 256630 429976 281522
rect 436112 279970 436140 281522
rect 446324 279970 446352 281590
rect 463792 281580 463844 281586
rect 463792 281522 463844 281528
rect 436112 279942 436356 279970
rect 446324 279942 446660 279970
rect 456964 279262 457116 279290
rect 430580 278792 430632 278798
rect 430580 278734 430632 278740
rect 434628 278792 434680 278798
rect 434628 278734 434680 278740
rect 430592 269793 430620 278734
rect 434640 269793 434668 278734
rect 430578 269784 430634 269793
rect 430578 269719 430634 269728
rect 434626 269784 434682 269793
rect 434626 269719 434682 269728
rect 436356 259134 436692 259162
rect 446660 259134 446996 259162
rect 429936 256624 429988 256630
rect 436664 256601 436692 259134
rect 446968 256630 446996 259134
rect 456812 259134 456964 259162
rect 456812 256698 456840 259134
rect 457088 256698 457116 279262
rect 462226 278080 462282 278089
rect 462226 278015 462282 278024
rect 462240 269793 462268 278015
rect 463700 272604 463752 272610
rect 463700 272546 463752 272552
rect 462226 269784 462282 269793
rect 462226 269719 462282 269728
rect 456800 256692 456852 256698
rect 456800 256634 456852 256640
rect 457076 256692 457128 256698
rect 457076 256634 457128 256640
rect 463712 256630 463740 272546
rect 463804 267734 463832 281522
rect 474278 279304 474334 279313
rect 464080 279262 464370 279290
rect 464080 272610 464108 279262
rect 474334 279262 474674 279290
rect 484978 279262 485084 279290
rect 474278 279239 474334 279248
rect 464068 272604 464120 272610
rect 464068 272546 464120 272552
rect 463804 267706 464016 267734
rect 463988 259706 464016 267706
rect 463988 259678 464370 259706
rect 474660 256630 474688 259148
rect 484964 256698 484992 259148
rect 485056 256698 485084 279262
rect 487160 278792 487212 278798
rect 487160 278734 487212 278740
rect 489828 278792 489880 278798
rect 489828 278734 489880 278740
rect 487172 269793 487200 278734
rect 489840 269793 489868 278734
rect 491300 272604 491352 272610
rect 491300 272546 491352 272552
rect 487158 269784 487214 269793
rect 487158 269719 487214 269728
rect 489826 269784 489882 269793
rect 489826 269719 489882 269728
rect 484952 256692 485004 256698
rect 484952 256634 485004 256640
rect 485044 256692 485096 256698
rect 485044 256634 485096 256640
rect 491312 256630 491340 272546
rect 491404 267734 491432 281590
rect 502616 281580 502668 281586
rect 502616 281522 502668 281528
rect 502628 279956 502656 281522
rect 492048 279262 492338 279290
rect 512946 279262 513144 279290
rect 492048 272610 492076 279262
rect 492036 272604 492088 272610
rect 492036 272546 492088 272552
rect 491404 267706 491984 267734
rect 491956 259706 491984 267706
rect 491956 259678 492338 259706
rect 446956 256624 447008 256630
rect 429936 256566 429988 256572
rect 436650 256592 436706 256601
rect 446956 256566 447008 256572
rect 463700 256624 463752 256630
rect 463700 256566 463752 256572
rect 474648 256624 474700 256630
rect 474648 256566 474700 256572
rect 491300 256624 491352 256630
rect 502628 256601 502656 259148
rect 512932 256698 512960 259148
rect 513116 256698 513144 279262
rect 514758 278080 514814 278089
rect 514758 278015 514814 278024
rect 514772 269793 514800 278015
rect 514758 269784 514814 269793
rect 514758 269719 514814 269728
rect 512920 256692 512972 256698
rect 512920 256634 512972 256640
rect 513104 256692 513156 256698
rect 513104 256634 513156 256640
rect 491300 256566 491352 256572
rect 502614 256592 502670 256601
rect 436650 256527 436706 256536
rect 502614 256527 502670 256536
rect 464344 255468 464396 255474
rect 464344 255410 464396 255416
rect 485136 255468 485188 255474
rect 485136 255410 485188 255416
rect 457444 255400 457496 255406
rect 457444 255342 457496 255348
rect 429844 255332 429896 255338
rect 429844 255274 429896 255280
rect 456616 255332 456668 255338
rect 456616 255274 456668 255280
rect 429856 230314 429884 255274
rect 456628 252892 456656 255274
rect 446034 252648 446090 252657
rect 446090 252606 446338 252634
rect 446034 252583 446090 252592
rect 434824 252334 436034 252362
rect 430578 242312 430634 242321
rect 430578 242247 430634 242256
rect 434626 242312 434682 242321
rect 434626 242247 434682 242256
rect 430592 233238 430620 242247
rect 434640 233238 434668 242247
rect 430580 233232 430632 233238
rect 430580 233174 430632 233180
rect 434628 233232 434680 233238
rect 434628 233174 434680 233180
rect 434824 230450 434852 252334
rect 457456 238754 457484 255342
rect 464356 252906 464384 255410
rect 474004 255400 474056 255406
rect 474004 255342 474056 255348
rect 464048 252878 464384 252906
rect 474016 252906 474044 255342
rect 485044 255332 485096 255338
rect 485044 255274 485096 255280
rect 474016 252878 474352 252906
rect 485056 252362 485084 255274
rect 484656 252334 484808 252362
rect 484780 251394 484808 252334
rect 484964 252334 485084 252362
rect 484768 251388 484820 251394
rect 484768 251330 484820 251336
rect 484964 249098 484992 252334
rect 485044 251388 485096 251394
rect 485044 251330 485096 251336
rect 484780 249070 484992 249098
rect 458178 242312 458234 242321
rect 458178 242247 458234 242256
rect 462226 242312 462282 242321
rect 462226 242247 462282 242256
rect 457088 238726 457484 238754
rect 457088 232778 457116 238726
rect 458192 234025 458220 242247
rect 462240 234025 462268 242247
rect 458178 234016 458234 234025
rect 458178 233951 458234 233960
rect 462226 234016 462282 234025
rect 462226 233951 462282 233960
rect 484780 232778 484808 249070
rect 485056 244338 485084 251330
rect 456642 232750 457116 232778
rect 484656 232750 484808 232778
rect 484872 244310 485084 244338
rect 434812 230444 434864 230450
rect 434812 230386 434864 230392
rect 436020 230382 436048 232084
rect 436008 230376 436060 230382
rect 436008 230318 436060 230324
rect 446324 230314 446352 232084
rect 463712 232070 464048 232098
rect 474352 232070 474688 232098
rect 463712 230382 463740 232070
rect 474660 230382 474688 232070
rect 463700 230376 463752 230382
rect 463700 230318 463752 230324
rect 474648 230376 474700 230382
rect 474648 230318 474700 230324
rect 484872 230314 484900 244310
rect 485148 235346 485176 255410
rect 502340 255332 502392 255338
rect 502340 255274 502392 255280
rect 513104 255332 513156 255338
rect 513104 255274 513156 255280
rect 502352 252892 502380 255274
rect 512670 252470 513052 252498
rect 491404 252334 492062 252362
rect 487158 242312 487214 242321
rect 487158 242247 487214 242256
rect 489826 242312 489882 242321
rect 489826 242247 489882 242256
rect 485136 235340 485188 235346
rect 485136 235282 485188 235288
rect 487172 233238 487200 242247
rect 489840 233238 489868 242247
rect 487160 233232 487212 233238
rect 487160 233174 487212 233180
rect 489828 233232 489880 233238
rect 489828 233174 489880 233180
rect 491404 230450 491432 252334
rect 512736 252068 512788 252074
rect 512736 252010 512788 252016
rect 491668 235340 491720 235346
rect 491668 235282 491720 235288
rect 491680 232778 491708 235282
rect 512748 232778 512776 252010
rect 513024 248282 513052 252470
rect 513116 252074 513144 255274
rect 513104 252068 513156 252074
rect 513104 252010 513156 252016
rect 491680 232750 492062 232778
rect 512670 232750 512776 232778
rect 512840 248254 513052 248282
rect 491392 230444 491444 230450
rect 491392 230386 491444 230392
rect 502352 230314 502380 232084
rect 512840 230382 512868 248254
rect 514758 242312 514814 242321
rect 514758 242247 514814 242256
rect 514772 234025 514800 242247
rect 514758 234016 514814 234025
rect 514758 233951 514814 233960
rect 512828 230376 512880 230382
rect 512828 230318 512880 230324
rect 429844 230308 429896 230314
rect 429844 230250 429896 230256
rect 446312 230308 446364 230314
rect 446312 230250 446364 230256
rect 484860 230308 484912 230314
rect 484860 230250 484912 230256
rect 502340 230308 502392 230314
rect 502340 230250 502392 230256
rect 446312 227928 446364 227934
rect 446312 227870 446364 227876
rect 491944 227928 491996 227934
rect 491944 227870 491996 227876
rect 429844 227860 429896 227866
rect 429844 227802 429896 227808
rect 436100 227860 436152 227866
rect 436100 227802 436152 227808
rect 429856 202774 429884 227802
rect 436112 225978 436140 227802
rect 446324 225978 446352 227870
rect 458824 227860 458876 227866
rect 458824 227802 458876 227808
rect 474648 227860 474700 227866
rect 474648 227802 474700 227808
rect 486424 227860 486476 227866
rect 486424 227802 486476 227808
rect 436112 225950 436356 225978
rect 446324 225950 446660 225978
rect 456964 225270 457116 225298
rect 434628 225140 434680 225146
rect 434628 225082 434680 225088
rect 429936 225004 429988 225010
rect 429936 224946 429988 224952
rect 429948 202842 429976 224946
rect 430578 224224 430634 224233
rect 430578 224159 430634 224168
rect 430592 215801 430620 224159
rect 434640 215801 434668 225082
rect 430578 215792 430634 215801
rect 430578 215727 430634 215736
rect 434626 215792 434682 215801
rect 434626 215727 434682 215736
rect 436356 205006 436692 205034
rect 446660 205006 446996 205034
rect 429936 202836 429988 202842
rect 429936 202778 429988 202784
rect 436664 202774 436692 205006
rect 429844 202768 429896 202774
rect 429844 202710 429896 202716
rect 436652 202768 436704 202774
rect 436652 202710 436704 202716
rect 446968 202706 446996 205006
rect 456812 205006 456964 205034
rect 456812 202842 456840 205006
rect 457088 202842 457116 225270
rect 458180 225072 458232 225078
rect 458180 225014 458232 225020
rect 458192 215801 458220 225014
rect 458178 215792 458234 215801
rect 458178 215727 458234 215736
rect 456800 202836 456852 202842
rect 456800 202778 456852 202784
rect 457076 202836 457128 202842
rect 457076 202778 457128 202784
rect 458836 202774 458864 227802
rect 460204 227792 460256 227798
rect 460204 227734 460256 227740
rect 464344 227792 464396 227798
rect 464344 227734 464396 227740
rect 458824 202768 458876 202774
rect 458824 202710 458876 202716
rect 460216 202706 460244 227734
rect 463976 227724 464028 227730
rect 463976 227666 464028 227672
rect 462226 224088 462282 224097
rect 462226 224023 462282 224032
rect 462240 215801 462268 224023
rect 462226 215792 462282 215801
rect 462226 215727 462282 215736
rect 463988 205714 464016 227666
rect 464356 225964 464384 227734
rect 474660 225964 474688 227802
rect 484978 225270 485084 225298
rect 463988 205686 464370 205714
rect 474476 205142 474674 205170
rect 474476 202774 474504 205142
rect 484688 205006 484978 205034
rect 484688 202842 484716 205006
rect 485056 202842 485084 225270
rect 484676 202836 484728 202842
rect 484676 202778 484728 202784
rect 485044 202836 485096 202842
rect 485044 202778 485096 202784
rect 486436 202774 486464 227802
rect 487160 225140 487212 225146
rect 487160 225082 487212 225088
rect 487172 215801 487200 225082
rect 487158 215792 487214 215801
rect 487158 215727 487214 215736
rect 491956 205714 491984 227870
rect 492312 227860 492364 227866
rect 492312 227802 492364 227808
rect 492324 225964 492352 227802
rect 502616 227792 502668 227798
rect 502616 227734 502668 227740
rect 514024 227792 514076 227798
rect 514024 227734 514076 227740
rect 502628 225964 502656 227734
rect 512946 225270 513144 225298
rect 491956 205686 492338 205714
rect 502628 202774 502656 205020
rect 512932 202842 512960 205020
rect 513116 202842 513144 225270
rect 512920 202836 512972 202842
rect 512920 202778 512972 202784
rect 513104 202836 513156 202842
rect 513104 202778 513156 202784
rect 514036 202774 514064 227734
rect 514758 224088 514814 224097
rect 514758 224023 514814 224032
rect 514772 215801 514800 224023
rect 514758 215792 514814 215801
rect 514758 215727 514814 215736
rect 474464 202768 474516 202774
rect 474464 202710 474516 202716
rect 486424 202768 486476 202774
rect 486424 202710 486476 202716
rect 502616 202768 502668 202774
rect 502616 202710 502668 202716
rect 514024 202768 514076 202774
rect 514024 202710 514076 202716
rect 446956 202700 447008 202706
rect 446956 202642 447008 202648
rect 460204 202700 460256 202706
rect 460204 202642 460256 202648
rect 464344 200320 464396 200326
rect 464344 200262 464396 200268
rect 485044 200320 485096 200326
rect 485044 200262 485096 200268
rect 457444 200252 457496 200258
rect 457444 200194 457496 200200
rect 429844 200184 429896 200190
rect 429844 200126 429896 200132
rect 456616 200184 456668 200190
rect 456616 200126 456668 200132
rect 429856 176526 429884 200126
rect 456628 198900 456656 200126
rect 446034 198520 446090 198529
rect 446090 198478 446338 198506
rect 446034 198455 446090 198464
rect 434824 198206 436034 198234
rect 430578 188320 430634 188329
rect 430578 188255 430634 188264
rect 434626 188320 434682 188329
rect 434626 188255 434682 188264
rect 430592 179382 430620 188255
rect 434640 179382 434668 188255
rect 430580 179376 430632 179382
rect 430580 179318 430632 179324
rect 434628 179376 434680 179382
rect 434628 179318 434680 179324
rect 434824 176662 434852 198206
rect 457456 180794 457484 200194
rect 464356 198914 464384 200262
rect 474004 200252 474056 200258
rect 474004 200194 474056 200200
rect 464048 198886 464384 198914
rect 474016 198914 474044 200194
rect 484860 200184 484912 200190
rect 484860 200126 484912 200132
rect 474016 198886 474352 198914
rect 484656 198206 484808 198234
rect 458178 196752 458234 196761
rect 458178 196687 458234 196696
rect 462226 196752 462282 196761
rect 462226 196687 462282 196696
rect 458192 188329 458220 196687
rect 462240 188329 462268 196687
rect 458178 188320 458234 188329
rect 458178 188255 458234 188264
rect 462226 188320 462282 188329
rect 462226 188255 462282 188264
rect 457088 180766 457484 180794
rect 457088 178786 457116 180766
rect 484780 178906 484808 198206
rect 484768 178900 484820 178906
rect 484768 178842 484820 178848
rect 456642 178758 457116 178786
rect 484872 178514 484900 200126
rect 485056 180878 485084 200262
rect 502340 200184 502392 200190
rect 502340 200126 502392 200132
rect 512736 200184 512788 200190
rect 512736 200126 512788 200132
rect 502352 198900 502380 200126
rect 512748 198354 512776 200126
rect 512736 198348 512788 198354
rect 512736 198290 512788 198296
rect 491404 198206 492062 198234
rect 512670 198206 512868 198234
rect 487158 188320 487214 188329
rect 487158 188255 487214 188264
rect 489826 188320 489882 188329
rect 489826 188255 489882 188264
rect 485044 180872 485096 180878
rect 485044 180814 485096 180820
rect 487172 179382 487200 188255
rect 489840 179382 489868 188255
rect 487160 179376 487212 179382
rect 487160 179318 487212 179324
rect 489828 179376 489880 179382
rect 489828 179318 489880 179324
rect 484952 178900 485004 178906
rect 484952 178842 485004 178848
rect 484656 178486 484900 178514
rect 434812 176656 434864 176662
rect 434812 176598 434864 176604
rect 436020 176594 436048 178092
rect 436008 176588 436060 176594
rect 436008 176530 436060 176536
rect 446324 176526 446352 178092
rect 463712 178078 464048 178106
rect 474352 178078 474688 178106
rect 463712 176594 463740 178078
rect 474660 176594 474688 178078
rect 463700 176588 463752 176594
rect 463700 176530 463752 176536
rect 474648 176588 474700 176594
rect 474648 176530 474700 176536
rect 484964 176526 484992 178842
rect 491404 176662 491432 198206
rect 512736 198144 512788 198150
rect 512736 198086 512788 198092
rect 491668 180872 491720 180878
rect 491668 180814 491720 180820
rect 491680 178786 491708 180814
rect 512748 178786 512776 198086
rect 491680 178758 492062 178786
rect 512670 178758 512776 178786
rect 491392 176656 491444 176662
rect 491392 176598 491444 176604
rect 502352 176526 502380 178092
rect 512840 176594 512868 198206
rect 514758 196752 514814 196761
rect 514758 196687 514814 196696
rect 514772 188329 514800 196687
rect 514758 188320 514814 188329
rect 514758 188255 514814 188264
rect 512828 176588 512880 176594
rect 512828 176530 512880 176536
rect 429844 176520 429896 176526
rect 429844 176462 429896 176468
rect 446312 176520 446364 176526
rect 446312 176462 446364 176468
rect 484952 176520 485004 176526
rect 484952 176462 485004 176468
rect 502340 176520 502392 176526
rect 502340 176462 502392 176468
rect 491392 174072 491444 174078
rect 491392 174014 491444 174020
rect 492404 174072 492456 174078
rect 492404 174014 492456 174020
rect 446312 174004 446364 174010
rect 446312 173946 446364 173952
rect 463792 174004 463844 174010
rect 463792 173946 463844 173952
rect 429936 173936 429988 173942
rect 429936 173878 429988 173884
rect 436100 173936 436152 173942
rect 436100 173878 436152 173884
rect 429844 171216 429896 171222
rect 429844 171158 429896 171164
rect 429856 149054 429884 171158
rect 429844 149048 429896 149054
rect 429844 148990 429896 148996
rect 429948 148986 429976 173878
rect 436112 171986 436140 173878
rect 446324 171986 446352 173946
rect 457444 173936 457496 173942
rect 457444 173878 457496 173884
rect 436112 171958 436356 171986
rect 446324 171958 446660 171986
rect 434628 171420 434680 171426
rect 434628 171362 434680 171368
rect 430578 170232 430634 170241
rect 430578 170167 430634 170176
rect 430592 161809 430620 170167
rect 434640 161809 434668 171362
rect 456964 171278 457116 171306
rect 430578 161800 430634 161809
rect 430578 161735 430634 161744
rect 434626 161800 434682 161809
rect 434626 161735 434682 161744
rect 436356 151014 436692 151042
rect 446660 151014 446996 151042
rect 436664 148986 436692 151014
rect 429936 148980 429988 148986
rect 429936 148922 429988 148928
rect 436652 148980 436704 148986
rect 436652 148922 436704 148928
rect 446968 148918 446996 151014
rect 456812 151014 456964 151042
rect 456812 149054 456840 151014
rect 457088 149054 457116 171278
rect 456800 149048 456852 149054
rect 456800 148990 456852 148996
rect 457076 149048 457128 149054
rect 457076 148990 457128 148996
rect 457456 148986 457484 173878
rect 462228 171488 462280 171494
rect 462228 171430 462280 171436
rect 458178 170096 458234 170105
rect 458178 170031 458234 170040
rect 458192 161809 458220 170031
rect 462240 161809 462268 171430
rect 463804 171134 463832 173946
rect 474648 173936 474700 173942
rect 474648 173878 474700 173884
rect 486424 173936 486476 173942
rect 486424 173878 486476 173884
rect 474660 171972 474688 173878
rect 464080 171278 464370 171306
rect 484978 171278 485084 171306
rect 463804 171106 464016 171134
rect 463700 166320 463752 166326
rect 463700 166262 463752 166268
rect 458178 161800 458234 161809
rect 458178 161735 458234 161744
rect 462226 161800 462282 161809
rect 462226 161735 462282 161744
rect 457444 148980 457496 148986
rect 457444 148922 457496 148928
rect 463712 148918 463740 166262
rect 463988 151722 464016 171106
rect 464080 166326 464108 171278
rect 464068 166320 464120 166326
rect 464068 166262 464120 166268
rect 463988 151694 464370 151722
rect 474660 148986 474688 151028
rect 484964 149054 484992 151028
rect 485056 149054 485084 171278
rect 484952 149048 485004 149054
rect 484952 148990 485004 148996
rect 485044 149048 485096 149054
rect 485044 148990 485096 148996
rect 486436 148986 486464 173878
rect 487160 171420 487212 171426
rect 487160 171362 487212 171368
rect 487172 161809 487200 171362
rect 491404 171134 491432 174014
rect 492416 173942 492444 174014
rect 502616 174004 502668 174010
rect 502616 173946 502668 173952
rect 492312 173936 492364 173942
rect 492312 173878 492364 173884
rect 492404 173936 492456 173942
rect 492404 173878 492456 173884
rect 492324 171972 492352 173878
rect 502628 171972 502656 173946
rect 514024 173936 514076 173942
rect 514024 173878 514076 173884
rect 512946 171278 513144 171306
rect 491404 171106 491984 171134
rect 489826 170232 489882 170241
rect 489826 170167 489882 170176
rect 489840 161809 489868 170167
rect 487158 161800 487214 161809
rect 487158 161735 487214 161744
rect 489826 161800 489882 161809
rect 489826 161735 489882 161744
rect 491956 151722 491984 171106
rect 491956 151694 492338 151722
rect 502628 148986 502656 151028
rect 512932 149054 512960 151028
rect 513116 149054 513144 171278
rect 512920 149048 512972 149054
rect 512920 148990 512972 148996
rect 513104 149048 513156 149054
rect 513104 148990 513156 148996
rect 514036 148986 514064 173878
rect 514760 171488 514812 171494
rect 514760 171430 514812 171436
rect 514772 161809 514800 171430
rect 514758 161800 514814 161809
rect 514758 161735 514814 161744
rect 474648 148980 474700 148986
rect 474648 148922 474700 148928
rect 486424 148980 486476 148986
rect 486424 148922 486476 148928
rect 502616 148980 502668 148986
rect 502616 148922 502668 148928
rect 514024 148980 514076 148986
rect 514024 148922 514076 148928
rect 446956 148912 447008 148918
rect 446956 148854 447008 148860
rect 463700 148912 463752 148918
rect 463700 148854 463752 148860
rect 457444 146396 457496 146402
rect 457444 146338 457496 146344
rect 474004 146396 474056 146402
rect 474004 146338 474056 146344
rect 484860 146396 484912 146402
rect 484860 146338 484912 146344
rect 502340 146396 502392 146402
rect 502340 146338 502392 146344
rect 512736 146396 512788 146402
rect 512736 146338 512788 146344
rect 429844 146328 429896 146334
rect 429844 146270 429896 146276
rect 456616 146328 456668 146334
rect 456616 146270 456668 146276
rect 429856 122670 429884 146270
rect 456628 144908 456656 146270
rect 446034 144528 446090 144537
rect 446090 144486 446338 144514
rect 446034 144463 446090 144472
rect 434824 144214 436034 144242
rect 430578 142760 430634 142769
rect 430578 142695 430634 142704
rect 434626 142760 434682 142769
rect 434626 142695 434682 142704
rect 430592 134337 430620 142695
rect 434640 134337 434668 142695
rect 430578 134328 430634 134337
rect 430578 134263 430634 134272
rect 434626 134328 434682 134337
rect 434626 134263 434682 134272
rect 434824 122806 434852 144214
rect 457456 132494 457484 146338
rect 464344 146328 464396 146334
rect 464344 146270 464396 146276
rect 464356 144922 464384 146270
rect 464048 144894 464384 144922
rect 474016 144922 474044 146338
rect 474016 144894 474352 144922
rect 484656 144214 484808 144242
rect 458178 134328 458234 134337
rect 458178 134263 458234 134272
rect 462226 134328 462282 134337
rect 462226 134263 462282 134272
rect 457088 132466 457484 132494
rect 457088 124794 457116 132466
rect 458192 125594 458220 134263
rect 462240 125594 462268 134263
rect 458180 125588 458232 125594
rect 458180 125530 458232 125536
rect 462228 125588 462280 125594
rect 462228 125530 462280 125536
rect 484780 124914 484808 144214
rect 484768 124908 484820 124914
rect 484768 124850 484820 124856
rect 484872 124794 484900 146338
rect 485044 146328 485096 146334
rect 485044 146270 485096 146276
rect 486424 146328 486476 146334
rect 486424 146270 486476 146276
rect 485056 128314 485084 146270
rect 485044 128308 485096 128314
rect 485044 128250 485096 128256
rect 456642 124766 457116 124794
rect 484656 124766 484900 124794
rect 484768 124704 484820 124710
rect 484768 124646 484820 124652
rect 434812 122800 434864 122806
rect 434812 122742 434864 122748
rect 436020 122738 436048 124100
rect 436008 122732 436060 122738
rect 436008 122674 436060 122680
rect 446324 122670 446352 124100
rect 463804 124086 464048 124114
rect 474352 124086 474688 124114
rect 463804 122738 463832 124086
rect 474660 122738 474688 124086
rect 463792 122732 463844 122738
rect 463792 122674 463844 122680
rect 474648 122732 474700 122738
rect 474648 122674 474700 122680
rect 484780 122670 484808 124646
rect 486436 122738 486464 146270
rect 502352 144908 502380 146338
rect 512644 146328 512696 146334
rect 512644 146270 512696 146276
rect 512656 144908 512684 146270
rect 491404 144214 492062 144242
rect 487158 142760 487214 142769
rect 487158 142695 487214 142704
rect 489826 142760 489882 142769
rect 489826 142695 489882 142704
rect 487172 134337 487200 142695
rect 489840 134337 489868 142695
rect 487158 134328 487214 134337
rect 487158 134263 487214 134272
rect 489826 134328 489882 134337
rect 489826 134263 489882 134272
rect 491404 122806 491432 144214
rect 491668 128308 491720 128314
rect 491668 128250 491720 128256
rect 491680 124794 491708 128250
rect 512748 124794 512776 146338
rect 514024 146328 514076 146334
rect 514024 146270 514076 146276
rect 491680 124766 492062 124794
rect 512670 124766 512776 124794
rect 491392 122800 491444 122806
rect 491392 122742 491444 122748
rect 502352 122738 502380 124100
rect 514036 122738 514064 146270
rect 514758 134328 514814 134337
rect 514758 134263 514814 134272
rect 514772 125594 514800 134263
rect 514760 125588 514812 125594
rect 514760 125530 514812 125536
rect 486424 122732 486476 122738
rect 486424 122674 486476 122680
rect 502340 122732 502392 122738
rect 502340 122674 502392 122680
rect 514024 122732 514076 122738
rect 514024 122674 514076 122680
rect 429844 122664 429896 122670
rect 429844 122606 429896 122612
rect 446312 122664 446364 122670
rect 446312 122606 446364 122612
rect 484768 122664 484820 122670
rect 484768 122606 484820 122612
rect 429844 120284 429896 120290
rect 429844 120226 429896 120232
rect 436100 120284 436152 120290
rect 436100 120226 436152 120232
rect 491392 120284 491444 120290
rect 491392 120226 491444 120232
rect 429856 95130 429884 120226
rect 436112 117994 436140 120226
rect 446312 120216 446364 120222
rect 446312 120158 446364 120164
rect 457444 120216 457496 120222
rect 457444 120158 457496 120164
rect 474372 120216 474424 120222
rect 474372 120158 474424 120164
rect 486424 120216 486476 120222
rect 486424 120158 486476 120164
rect 446324 117994 446352 120158
rect 436112 117966 436356 117994
rect 446324 117966 446660 117994
rect 434628 117360 434680 117366
rect 434628 117302 434680 117308
rect 429936 117292 429988 117298
rect 429936 117234 429988 117240
rect 429948 95198 429976 117234
rect 430578 116240 430634 116249
rect 430578 116175 430634 116184
rect 430592 107817 430620 116175
rect 434640 107817 434668 117302
rect 456964 117286 457116 117314
rect 430578 107808 430634 107817
rect 430578 107743 430634 107752
rect 434626 107808 434682 107817
rect 434626 107743 434682 107752
rect 436356 97022 436692 97050
rect 446660 97022 446996 97050
rect 429936 95192 429988 95198
rect 429936 95134 429988 95140
rect 436664 95130 436692 97022
rect 429844 95124 429896 95130
rect 429844 95066 429896 95072
rect 436652 95124 436704 95130
rect 436652 95066 436704 95072
rect 446968 95062 446996 97022
rect 456812 97022 456964 97050
rect 456812 95198 456840 97022
rect 457088 95198 457116 117286
rect 456800 95192 456852 95198
rect 456800 95134 456852 95140
rect 457076 95192 457128 95198
rect 457076 95134 457128 95140
rect 457456 95130 457484 120158
rect 458824 120148 458876 120154
rect 458824 120090 458876 120096
rect 464068 120148 464120 120154
rect 464068 120090 464120 120096
rect 458178 116104 458234 116113
rect 458178 116039 458234 116048
rect 458192 108361 458220 116039
rect 458178 108352 458234 108361
rect 458178 108287 458234 108296
rect 457444 95124 457496 95130
rect 457444 95066 457496 95072
rect 458836 95062 458864 120090
rect 463792 120080 463844 120086
rect 463792 120022 463844 120028
rect 462226 116104 462282 116113
rect 462226 116039 462282 116048
rect 462240 107817 462268 116039
rect 463804 113174 463832 120022
rect 464080 117994 464108 120090
rect 474384 117994 474412 120158
rect 464080 117966 464370 117994
rect 474384 117966 474674 117994
rect 484978 117286 485084 117314
rect 463804 113146 464016 113174
rect 462226 107808 462282 107817
rect 462226 107743 462282 107752
rect 463988 97730 464016 113146
rect 463988 97702 464370 97730
rect 474660 95130 474688 97036
rect 484964 95198 484992 97036
rect 485056 95198 485084 117286
rect 484952 95192 485004 95198
rect 484952 95134 485004 95140
rect 485044 95192 485096 95198
rect 485044 95134 485096 95140
rect 486436 95130 486464 120158
rect 487160 117360 487212 117366
rect 487160 117302 487212 117308
rect 487172 107817 487200 117302
rect 489826 116240 489882 116249
rect 489826 116175 489882 116184
rect 489840 107817 489868 116175
rect 491404 113174 491432 120226
rect 492312 120216 492364 120222
rect 492312 120158 492364 120164
rect 492324 117980 492352 120158
rect 502616 120148 502668 120154
rect 502616 120090 502668 120096
rect 514024 120148 514076 120154
rect 514024 120090 514076 120096
rect 502628 117980 502656 120090
rect 512946 117286 513144 117314
rect 491404 113146 491984 113174
rect 487158 107808 487214 107817
rect 487158 107743 487214 107752
rect 489826 107808 489882 107817
rect 489826 107743 489882 107752
rect 491956 97730 491984 113146
rect 491956 97702 492338 97730
rect 502628 95130 502656 97036
rect 512932 95198 512960 97036
rect 513116 95198 513144 117286
rect 512920 95192 512972 95198
rect 512920 95134 512972 95140
rect 513104 95192 513156 95198
rect 513104 95134 513156 95140
rect 514036 95130 514064 120090
rect 514758 116104 514814 116113
rect 514758 116039 514814 116048
rect 514772 107817 514800 116039
rect 514758 107808 514814 107817
rect 514758 107743 514814 107752
rect 474648 95124 474700 95130
rect 474648 95066 474700 95072
rect 486424 95124 486476 95130
rect 486424 95066 486476 95072
rect 502616 95124 502668 95130
rect 502616 95066 502668 95072
rect 514024 95124 514076 95130
rect 514024 95066 514076 95072
rect 446956 95056 447008 95062
rect 446956 94998 447008 95004
rect 458824 95056 458876 95062
rect 458824 94998 458876 95004
rect 458824 92676 458876 92682
rect 458824 92618 458876 92624
rect 474004 92676 474056 92682
rect 474004 92618 474056 92624
rect 435364 92608 435416 92614
rect 435364 92550 435416 92556
rect 446312 92608 446364 92614
rect 446312 92550 446364 92556
rect 429844 92540 429896 92546
rect 429844 92482 429896 92488
rect 429856 68882 429884 92482
rect 430578 88904 430634 88913
rect 430578 88839 430634 88848
rect 434626 88904 434682 88913
rect 434626 88839 434682 88848
rect 430592 80345 430620 88839
rect 434640 80345 434668 88839
rect 434720 87236 434772 87242
rect 434720 87178 434772 87184
rect 430578 80336 430634 80345
rect 430578 80271 430634 80280
rect 434626 80336 434682 80345
rect 434626 80271 434682 80280
rect 434732 68882 434760 87178
rect 435376 69018 435404 92550
rect 446324 90916 446352 92550
rect 456616 92540 456668 92546
rect 456616 92482 456668 92488
rect 457444 92540 457496 92546
rect 457444 92482 457496 92488
rect 456628 90916 456656 92482
rect 435744 90222 436034 90250
rect 435744 87242 435772 90222
rect 435732 87236 435784 87242
rect 435732 87178 435784 87184
rect 435364 69012 435416 69018
rect 435364 68954 435416 68960
rect 436020 68950 436048 70108
rect 446324 68950 446352 70108
rect 456628 69018 456656 70108
rect 456616 69012 456668 69018
rect 456616 68954 456668 68960
rect 457456 68950 457484 92482
rect 458180 89752 458232 89758
rect 458180 89694 458232 89700
rect 458192 80345 458220 89694
rect 458178 80336 458234 80345
rect 458178 80271 458234 80280
rect 458836 69018 458864 92618
rect 464344 92608 464396 92614
rect 464344 92550 464396 92556
rect 464356 90930 464384 92550
rect 464048 90902 464384 90930
rect 474016 90930 474044 92618
rect 485044 92608 485096 92614
rect 485044 92550 485096 92556
rect 512920 92608 512972 92614
rect 512920 92550 512972 92556
rect 484400 92540 484452 92546
rect 484400 92482 484452 92488
rect 484768 92540 484820 92546
rect 484768 92482 484820 92488
rect 484412 90930 484440 92482
rect 474016 90902 474352 90930
rect 484412 90902 484656 90930
rect 462226 88768 462282 88777
rect 462226 88703 462282 88712
rect 462240 80345 462268 88703
rect 462226 80336 462282 80345
rect 462226 80271 462282 80280
rect 484780 70666 484808 92482
rect 485056 73710 485084 92550
rect 502340 92540 502392 92546
rect 502340 92482 502392 92488
rect 502352 90916 502380 92482
rect 512670 90494 512868 90522
rect 491404 90222 492062 90250
rect 489828 89752 489880 89758
rect 489828 89694 489880 89700
rect 489840 80345 489868 89694
rect 489826 80336 489882 80345
rect 489826 80271 489882 80280
rect 485044 73704 485096 73710
rect 485044 73646 485096 73652
rect 484656 70638 484808 70666
rect 463712 70094 464048 70122
rect 474352 70094 474688 70122
rect 458824 69012 458876 69018
rect 458824 68954 458876 68960
rect 436008 68944 436060 68950
rect 436008 68886 436060 68892
rect 446312 68944 446364 68950
rect 446312 68886 446364 68892
rect 457444 68944 457496 68950
rect 457444 68886 457496 68892
rect 463712 68882 463740 70094
rect 474660 69018 474688 70094
rect 474648 69012 474700 69018
rect 474648 68954 474700 68960
rect 491404 68950 491432 90222
rect 512840 85066 512868 90494
rect 512828 85060 512880 85066
rect 512828 85002 512880 85008
rect 512932 82090 512960 92550
rect 514024 92540 514076 92546
rect 514024 92482 514076 92488
rect 513012 85060 513064 85066
rect 513012 85002 513064 85008
rect 512748 82062 512960 82090
rect 491668 73704 491720 73710
rect 491668 73646 491720 73652
rect 491680 70666 491708 73646
rect 512748 70666 512776 82062
rect 513024 77314 513052 85002
rect 512828 77308 512880 77314
rect 512828 77250 512880 77256
rect 513012 77308 513064 77314
rect 513012 77250 513064 77256
rect 491680 70638 492062 70666
rect 512670 70638 512776 70666
rect 491392 68944 491444 68950
rect 491392 68886 491444 68892
rect 502352 68882 502380 70108
rect 512840 69018 512868 77250
rect 512828 69012 512880 69018
rect 512828 68954 512880 68960
rect 514036 68882 514064 92482
rect 514758 88768 514814 88777
rect 514758 88703 514814 88712
rect 514772 80345 514800 88703
rect 514758 80336 514814 80345
rect 514758 80271 514814 80280
rect 429844 68876 429896 68882
rect 429844 68818 429896 68824
rect 434720 68876 434772 68882
rect 434720 68818 434772 68824
rect 463700 68876 463752 68882
rect 463700 68818 463752 68824
rect 502340 68876 502392 68882
rect 502340 68818 502392 68824
rect 514024 68876 514076 68882
rect 514024 68818 514076 68824
rect 491392 66428 491444 66434
rect 491392 66370 491444 66376
rect 446312 66360 446364 66366
rect 446312 66302 446364 66308
rect 457444 66360 457496 66366
rect 457444 66302 457496 66308
rect 474648 66360 474700 66366
rect 474648 66302 474700 66308
rect 486424 66360 486476 66366
rect 486424 66302 486476 66308
rect 446324 63866 446352 66302
rect 446324 63838 446660 63866
rect 429844 63300 429896 63306
rect 429844 63242 429896 63248
rect 436112 63294 436356 63322
rect 456964 63294 457116 63322
rect 429856 41410 429884 63242
rect 430578 53816 430634 53825
rect 430578 53751 430634 53760
rect 434626 53816 434682 53825
rect 434626 53751 434682 53760
rect 430592 45257 430620 53751
rect 434640 45257 434668 53751
rect 430578 45248 430634 45257
rect 430578 45183 430634 45192
rect 434626 45248 434682 45257
rect 434626 45183 434682 45192
rect 429844 41404 429896 41410
rect 429844 41346 429896 41352
rect 436112 41342 436140 63294
rect 436356 43030 436692 43058
rect 446660 43030 446996 43058
rect 436664 41342 436692 43030
rect 436100 41336 436152 41342
rect 436100 41278 436152 41284
rect 436652 41336 436704 41342
rect 436652 41278 436704 41284
rect 446968 41274 446996 43030
rect 456812 43030 456964 43058
rect 456812 41410 456840 43030
rect 457088 41410 457116 63294
rect 456800 41404 456852 41410
rect 456800 41346 456852 41352
rect 457076 41404 457128 41410
rect 457076 41346 457128 41352
rect 457456 41342 457484 66302
rect 458824 66292 458876 66298
rect 458824 66234 458876 66240
rect 464344 66292 464396 66298
rect 464344 66234 464396 66240
rect 457444 41336 457496 41342
rect 457444 41278 457496 41284
rect 458836 41274 458864 66234
rect 463792 66224 463844 66230
rect 463792 66166 463844 66172
rect 463804 55214 463832 66166
rect 464356 63852 464384 66234
rect 474660 63852 474688 66302
rect 484978 63294 485084 63322
rect 463804 55186 464016 55214
rect 462226 53816 462282 53825
rect 462226 53751 462282 53760
rect 462240 45393 462268 53751
rect 462226 45384 462282 45393
rect 462226 45319 462282 45328
rect 463988 43738 464016 55186
rect 463988 43710 464370 43738
rect 474660 41342 474688 43044
rect 484964 41410 484992 43044
rect 485056 41410 485084 63294
rect 484952 41404 485004 41410
rect 484952 41346 485004 41352
rect 485044 41404 485096 41410
rect 485044 41346 485096 41352
rect 486436 41342 486464 66302
rect 491404 55214 491432 66370
rect 492312 66360 492364 66366
rect 492312 66302 492364 66308
rect 492324 63852 492352 66302
rect 502616 66292 502668 66298
rect 502616 66234 502668 66240
rect 514024 66292 514076 66298
rect 514024 66234 514076 66240
rect 502628 63852 502656 66234
rect 512946 63294 513144 63322
rect 491404 55186 491984 55214
rect 489826 53816 489882 53825
rect 489826 53751 489882 53760
rect 489840 44130 489868 53751
rect 489828 44124 489880 44130
rect 489828 44066 489880 44072
rect 491956 43738 491984 55186
rect 491956 43710 492338 43738
rect 502628 41342 502656 43044
rect 512932 41410 512960 43044
rect 513116 41410 513144 63294
rect 512920 41404 512972 41410
rect 512920 41346 512972 41352
rect 513104 41404 513156 41410
rect 513104 41346 513156 41352
rect 514036 41342 514064 66234
rect 514758 53816 514814 53825
rect 514758 53751 514814 53760
rect 514772 45393 514800 53751
rect 514758 45384 514814 45393
rect 514758 45319 514814 45328
rect 474648 41336 474700 41342
rect 474648 41278 474700 41284
rect 486424 41336 486476 41342
rect 486424 41278 486476 41284
rect 502616 41336 502668 41342
rect 502616 41278 502668 41284
rect 514024 41336 514076 41342
rect 514024 41278 514076 41284
rect 446956 41268 447008 41274
rect 446956 41210 447008 41216
rect 458824 41268 458876 41274
rect 458824 41210 458876 41216
rect 457444 38752 457496 38758
rect 457444 38694 457496 38700
rect 474004 38752 474056 38758
rect 474004 38694 474056 38700
rect 484860 38752 484912 38758
rect 484860 38694 484912 38700
rect 502340 38752 502392 38758
rect 502340 38694 502392 38700
rect 512736 38752 512788 38758
rect 512736 38694 512788 38700
rect 446312 38684 446364 38690
rect 446312 38626 446364 38632
rect 446324 36924 446352 38626
rect 456338 36544 456394 36553
rect 456394 36502 456642 36530
rect 456338 36479 456394 36488
rect 434824 36230 436034 36258
rect 430578 34912 430634 34921
rect 430578 34847 430634 34856
rect 430592 26353 430620 34847
rect 430578 26344 430634 26353
rect 430578 26279 430634 26288
rect 429200 15156 429252 15162
rect 429200 15098 429252 15104
rect 418342 13424 418398 13433
rect 418342 13359 418398 13368
rect 407212 13320 407264 13326
rect 407212 13262 407264 13268
rect 434824 13258 434852 36230
rect 457456 16574 457484 38694
rect 464344 38684 464396 38690
rect 464344 38626 464396 38632
rect 464356 36938 464384 38626
rect 464048 36910 464384 36938
rect 474016 36938 474044 38694
rect 474016 36910 474352 36938
rect 484656 36230 484808 36258
rect 458178 34776 458234 34785
rect 458178 34711 458234 34720
rect 462226 34776 462282 34785
rect 462226 34711 462282 34720
rect 458192 26897 458220 34711
rect 458178 26888 458234 26897
rect 458178 26823 458234 26832
rect 462240 26353 462268 34711
rect 462226 26344 462282 26353
rect 462226 26279 462282 26288
rect 484780 21418 484808 36230
rect 484768 21412 484820 21418
rect 484768 21354 484820 21360
rect 484872 16674 484900 38694
rect 485044 38684 485096 38690
rect 485044 38626 485096 38632
rect 486424 38684 486476 38690
rect 486424 38626 486476 38632
rect 484952 21412 485004 21418
rect 484952 21354 485004 21360
rect 484656 16646 484900 16674
rect 457088 16546 457484 16574
rect 457088 16538 457116 16546
rect 456642 16510 457116 16538
rect 436020 13326 436048 16116
rect 446324 13326 446352 16116
rect 463712 16102 464048 16130
rect 474352 16102 474688 16130
rect 436008 13320 436060 13326
rect 436008 13262 436060 13268
rect 446312 13320 446364 13326
rect 446312 13262 446364 13268
rect 463712 13258 463740 16102
rect 474660 13802 474688 16102
rect 474648 13796 474700 13802
rect 474648 13738 474700 13744
rect 484964 13326 484992 21354
rect 485056 18018 485084 38626
rect 485044 18012 485096 18018
rect 485044 17954 485096 17960
rect 486436 13802 486464 38626
rect 502352 36924 502380 38694
rect 512644 38684 512696 38690
rect 512644 38626 512696 38632
rect 512656 36924 512684 38626
rect 491404 36230 492062 36258
rect 487158 34912 487214 34921
rect 487158 34847 487214 34856
rect 487172 26353 487200 34847
rect 487158 26344 487214 26353
rect 487158 26279 487214 26288
rect 486424 13796 486476 13802
rect 486424 13738 486476 13744
rect 491404 13326 491432 36230
rect 491668 18012 491720 18018
rect 491668 17954 491720 17960
rect 491680 16674 491708 17954
rect 512748 16674 512776 38694
rect 512828 38684 512880 38690
rect 512828 38626 512880 38632
rect 491680 16646 492062 16674
rect 512670 16646 512776 16674
rect 502352 13802 502380 16116
rect 512840 13802 512868 38626
rect 514758 34776 514814 34785
rect 514758 34711 514814 34720
rect 514772 26353 514800 34711
rect 514758 26344 514814 26353
rect 514758 26279 514814 26288
rect 502340 13796 502392 13802
rect 502340 13738 502392 13744
rect 512828 13796 512880 13802
rect 512828 13738 512880 13744
rect 518176 13394 518204 700334
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 530308 687268 530360 687274
rect 530308 687210 530360 687216
rect 530320 684964 530348 687210
rect 557998 684584 558054 684593
rect 558054 684542 558348 684570
rect 557998 684519 558054 684528
rect 519004 684270 520030 684298
rect 540638 684270 540836 684298
rect 568652 684270 568804 684298
rect 518806 674248 518862 674257
rect 518806 674183 518862 674192
rect 518820 665961 518848 674183
rect 518806 665952 518862 665961
rect 518806 665887 518862 665896
rect 519004 662318 519032 684270
rect 520016 662386 520044 664020
rect 530320 662386 530348 664020
rect 540624 662425 540652 664020
rect 540610 662416 540666 662425
rect 520004 662380 520056 662386
rect 520004 662322 520056 662328
rect 530308 662380 530360 662386
rect 540610 662351 540666 662360
rect 530308 662322 530360 662328
rect 518992 662312 519044 662318
rect 518992 662254 519044 662260
rect 540808 662250 540836 684270
rect 542358 674248 542414 674257
rect 542358 674183 542414 674192
rect 545762 674248 545818 674257
rect 545762 674183 545818 674192
rect 542372 665174 542400 674183
rect 542360 665168 542412 665174
rect 542360 665110 542412 665116
rect 540796 662244 540848 662250
rect 540796 662186 540848 662192
rect 530308 659796 530360 659802
rect 530308 659738 530360 659744
rect 530320 657914 530348 659738
rect 541624 659728 541676 659734
rect 541624 659670 541676 659676
rect 530320 657886 530656 657914
rect 520186 657248 520242 657257
rect 520242 657206 520352 657234
rect 540960 657206 541112 657234
rect 520186 657183 520242 657192
rect 518806 656024 518862 656033
rect 518806 655959 518862 655968
rect 518820 647737 518848 655959
rect 518806 647728 518862 647737
rect 518806 647663 518862 647672
rect 520352 637078 520688 637106
rect 530656 637078 530992 637106
rect 520660 634710 520688 637078
rect 520648 634704 520700 634710
rect 520648 634646 520700 634652
rect 530964 634642 530992 637078
rect 540624 637078 540960 637106
rect 540624 634778 540652 637078
rect 541084 634778 541112 657206
rect 540612 634772 540664 634778
rect 540612 634714 540664 634720
rect 541072 634772 541124 634778
rect 541072 634714 541124 634720
rect 541636 634710 541664 659670
rect 542360 656940 542412 656946
rect 542360 656882 542412 656888
rect 542372 647737 542400 656882
rect 542358 647728 542414 647737
rect 542358 647663 542414 647672
rect 541624 634704 541676 634710
rect 541624 634646 541676 634652
rect 530952 634636 531004 634642
rect 530952 634578 531004 634584
rect 530308 632120 530360 632126
rect 530308 632062 530360 632068
rect 530320 630972 530348 632062
rect 519004 630278 520030 630306
rect 540638 630278 540836 630306
rect 518806 620256 518862 620265
rect 518806 620191 518862 620200
rect 518820 611969 518848 620191
rect 518806 611960 518862 611969
rect 518806 611895 518862 611904
rect 519004 608394 519032 630278
rect 520016 608598 520044 610028
rect 530320 608598 530348 610028
rect 520004 608592 520056 608598
rect 520004 608534 520056 608540
rect 530308 608592 530360 608598
rect 540624 608569 540652 610028
rect 530308 608534 530360 608540
rect 540610 608560 540666 608569
rect 540610 608495 540666 608504
rect 540808 608462 540836 630278
rect 542358 620256 542414 620265
rect 542358 620191 542414 620200
rect 542372 611318 542400 620191
rect 542360 611312 542412 611318
rect 542360 611254 542412 611260
rect 540796 608456 540848 608462
rect 540796 608398 540848 608404
rect 518992 608388 519044 608394
rect 518992 608330 519044 608336
rect 520280 605940 520332 605946
rect 520280 605882 520332 605888
rect 520292 603922 520320 605882
rect 530308 605872 530360 605878
rect 530308 605814 530360 605820
rect 541624 605872 541676 605878
rect 541624 605814 541676 605820
rect 530320 603922 530348 605814
rect 520292 603894 520352 603922
rect 530320 603894 530656 603922
rect 540960 603214 541112 603242
rect 520352 583086 520688 583114
rect 530656 583086 530992 583114
rect 520660 580922 520688 583086
rect 520648 580916 520700 580922
rect 520648 580858 520700 580864
rect 530964 580854 530992 583086
rect 540624 583086 540960 583114
rect 540624 580990 540652 583086
rect 541084 580990 541112 603214
rect 540612 580984 540664 580990
rect 540612 580926 540664 580932
rect 541072 580984 541124 580990
rect 541072 580926 541124 580932
rect 541636 580922 541664 605814
rect 542358 602168 542414 602177
rect 542358 602103 542414 602112
rect 542372 593745 542400 602103
rect 542358 593736 542414 593745
rect 542358 593671 542414 593680
rect 541624 580916 541676 580922
rect 541624 580858 541676 580864
rect 530952 580848 531004 580854
rect 530952 580790 531004 580796
rect 530308 578264 530360 578270
rect 530308 578206 530360 578212
rect 530320 576980 530348 578206
rect 519004 576286 520030 576314
rect 540638 576286 540836 576314
rect 518806 574696 518862 574705
rect 518806 574631 518862 574640
rect 518820 566273 518848 574631
rect 518806 566264 518862 566273
rect 518806 566199 518862 566208
rect 519004 554538 519032 576286
rect 520016 554742 520044 556036
rect 530320 554742 530348 556036
rect 520004 554736 520056 554742
rect 520004 554678 520056 554684
rect 530308 554736 530360 554742
rect 540624 554713 540652 556036
rect 530308 554678 530360 554684
rect 540610 554704 540666 554713
rect 540610 554639 540666 554648
rect 540808 554606 540836 576286
rect 542358 566264 542414 566273
rect 542358 566199 542414 566208
rect 542372 557530 542400 566199
rect 542360 557524 542412 557530
rect 542360 557466 542412 557472
rect 540796 554600 540848 554606
rect 540796 554542 540848 554548
rect 518992 554532 519044 554538
rect 518992 554474 519044 554480
rect 530308 552152 530360 552158
rect 530308 552094 530360 552100
rect 520280 550588 520332 550594
rect 520280 550530 520332 550536
rect 520292 549930 520320 550530
rect 530320 549930 530348 552094
rect 541624 552084 541676 552090
rect 541624 552026 541676 552032
rect 520292 549902 520352 549930
rect 530320 549902 530656 549930
rect 540960 549222 541112 549250
rect 520352 529094 520688 529122
rect 530656 529094 530992 529122
rect 520660 527066 520688 529094
rect 520648 527060 520700 527066
rect 520648 527002 520700 527008
rect 530964 526998 530992 529094
rect 540624 529094 540960 529122
rect 540624 527134 540652 529094
rect 541084 527134 541112 549222
rect 540612 527128 540664 527134
rect 540612 527070 540664 527076
rect 541072 527128 541124 527134
rect 541072 527070 541124 527076
rect 541636 527066 541664 552026
rect 541624 527060 541676 527066
rect 541624 527002 541676 527008
rect 530952 526992 531004 526998
rect 530952 526934 531004 526940
rect 530308 524476 530360 524482
rect 530308 524418 530360 524424
rect 530320 522852 530348 524418
rect 519004 522294 520030 522322
rect 540638 522294 540836 522322
rect 519004 500750 519032 522294
rect 520016 500954 520044 502044
rect 530320 500954 530348 502044
rect 520004 500948 520056 500954
rect 520004 500890 520056 500896
rect 530308 500948 530360 500954
rect 530308 500890 530360 500896
rect 540624 500857 540652 502044
rect 540610 500848 540666 500857
rect 540808 500818 540836 522294
rect 542358 520840 542414 520849
rect 542358 520775 542414 520784
rect 542372 512281 542400 520775
rect 542358 512272 542414 512281
rect 542358 512207 542414 512216
rect 540610 500783 540666 500792
rect 540796 500812 540848 500818
rect 540796 500754 540848 500760
rect 518992 500744 519044 500750
rect 518992 500686 519044 500692
rect 530308 498296 530360 498302
rect 530308 498238 530360 498244
rect 520280 498228 520332 498234
rect 520280 498170 520332 498176
rect 520292 495938 520320 498170
rect 530320 495938 530348 498238
rect 541624 498228 541676 498234
rect 541624 498170 541676 498176
rect 520292 495910 520352 495938
rect 530320 495910 530656 495938
rect 540960 495230 541112 495258
rect 520352 475102 520688 475130
rect 530656 475102 530992 475130
rect 520660 473278 520688 475102
rect 520648 473272 520700 473278
rect 520648 473214 520700 473220
rect 530964 473210 530992 475102
rect 540624 475102 540960 475130
rect 540624 473346 540652 475102
rect 541084 473346 541112 495230
rect 540612 473340 540664 473346
rect 540612 473282 540664 473288
rect 541072 473340 541124 473346
rect 541072 473282 541124 473288
rect 541636 473278 541664 498170
rect 541624 473272 541676 473278
rect 541624 473214 541676 473220
rect 530952 473204 531004 473210
rect 530952 473146 531004 473152
rect 530308 470688 530360 470694
rect 530308 470630 530360 470636
rect 530320 468860 530348 470630
rect 519004 468302 520030 468330
rect 540638 468302 540836 468330
rect 519004 445670 519032 468302
rect 520016 445738 520044 448052
rect 530320 445738 530348 448052
rect 520004 445732 520056 445738
rect 520004 445674 520056 445680
rect 530308 445732 530360 445738
rect 530308 445674 530360 445680
rect 518992 445664 519044 445670
rect 540624 445641 540652 448052
rect 518992 445606 519044 445612
rect 540610 445632 540666 445641
rect 540808 445602 540836 468302
rect 542358 466848 542414 466857
rect 542358 466783 542414 466792
rect 542372 458289 542400 466783
rect 542358 458280 542414 458289
rect 542358 458215 542414 458224
rect 540610 445567 540666 445576
rect 540796 445596 540848 445602
rect 540796 445538 540848 445544
rect 530308 444508 530360 444514
rect 530308 444450 530360 444456
rect 520280 444440 520332 444446
rect 520280 444382 520332 444388
rect 520292 441946 520320 444382
rect 530320 441946 530348 444450
rect 541624 444440 541676 444446
rect 541624 444382 541676 444388
rect 520292 441918 520352 441946
rect 530320 441918 530656 441946
rect 540960 441238 541112 441266
rect 520352 421110 520688 421138
rect 530656 421110 530992 421138
rect 520660 419422 520688 421110
rect 520648 419416 520700 419422
rect 520648 419358 520700 419364
rect 530964 419354 530992 421110
rect 540624 421110 540960 421138
rect 540624 419490 540652 421110
rect 541084 419490 541112 441238
rect 540612 419484 540664 419490
rect 540612 419426 540664 419432
rect 541072 419484 541124 419490
rect 541072 419426 541124 419432
rect 541636 419422 541664 444382
rect 542358 431760 542414 431769
rect 542358 431695 542414 431704
rect 542372 423201 542400 431695
rect 542358 423192 542414 423201
rect 542358 423127 542414 423136
rect 541624 419416 541676 419422
rect 541624 419358 541676 419364
rect 530952 419348 531004 419354
rect 530952 419290 531004 419296
rect 530308 416832 530360 416838
rect 530308 416774 530360 416780
rect 530320 414868 530348 416774
rect 519004 414310 520030 414338
rect 540638 414310 540836 414338
rect 519004 391746 519032 414310
rect 520016 391950 520044 394060
rect 530320 391950 530348 394060
rect 520004 391944 520056 391950
rect 520004 391886 520056 391892
rect 530308 391944 530360 391950
rect 540624 391921 540652 394060
rect 530308 391886 530360 391892
rect 540610 391912 540666 391921
rect 540610 391847 540666 391856
rect 540808 391814 540836 414310
rect 542358 404288 542414 404297
rect 542358 404223 542414 404232
rect 542372 395865 542400 404223
rect 542358 395856 542414 395865
rect 542358 395791 542414 395800
rect 540796 391808 540848 391814
rect 540796 391750 540848 391756
rect 518992 391740 519044 391746
rect 518992 391682 519044 391688
rect 530308 389292 530360 389298
rect 530308 389234 530360 389240
rect 520280 389224 520332 389230
rect 520280 389166 520332 389172
rect 520292 387954 520320 389166
rect 530320 387954 530348 389234
rect 541624 389224 541676 389230
rect 541624 389166 541676 389172
rect 520292 387926 520352 387954
rect 530320 387926 530656 387954
rect 540960 387246 541112 387274
rect 518806 377768 518862 377777
rect 518806 377703 518862 377712
rect 518820 369345 518848 377703
rect 518806 369336 518862 369345
rect 518806 369271 518862 369280
rect 520352 367118 520688 367146
rect 530656 367118 530992 367146
rect 520660 365634 520688 367118
rect 520648 365628 520700 365634
rect 520648 365570 520700 365576
rect 530964 365566 530992 367118
rect 540624 367118 540960 367146
rect 540624 365702 540652 367118
rect 541084 365702 541112 387246
rect 540612 365696 540664 365702
rect 540612 365638 540664 365644
rect 541072 365696 541124 365702
rect 541072 365638 541124 365644
rect 541636 365634 541664 389166
rect 542358 377768 542414 377777
rect 542358 377703 542414 377712
rect 542372 368490 542400 377703
rect 542360 368484 542412 368490
rect 542360 368426 542412 368432
rect 541624 365628 541676 365634
rect 541624 365570 541676 365576
rect 530952 365560 531004 365566
rect 530952 365502 531004 365508
rect 530308 362976 530360 362982
rect 530308 362918 530360 362924
rect 530320 360876 530348 362918
rect 519004 360318 520030 360346
rect 540638 360318 540836 360346
rect 519004 337890 519032 360318
rect 520016 338094 520044 340068
rect 530320 338094 530348 340068
rect 520004 338088 520056 338094
rect 520004 338030 520056 338036
rect 530308 338088 530360 338094
rect 540624 338065 540652 340068
rect 530308 338030 530360 338036
rect 540610 338056 540666 338065
rect 540610 337991 540666 338000
rect 540808 337958 540836 360318
rect 542358 350296 542414 350305
rect 542358 350231 542414 350240
rect 542372 341873 542400 350231
rect 542358 341864 542414 341873
rect 542358 341799 542414 341808
rect 540796 337952 540848 337958
rect 540796 337894 540848 337900
rect 518992 337884 519044 337890
rect 518992 337826 519044 337832
rect 530308 335436 530360 335442
rect 530308 335378 530360 335384
rect 520280 335368 520332 335374
rect 520280 335310 520332 335316
rect 520292 333962 520320 335310
rect 530320 333962 530348 335378
rect 541624 335368 541676 335374
rect 541624 335310 541676 335316
rect 520292 333934 520352 333962
rect 530320 333934 530656 333962
rect 540960 333254 541112 333282
rect 518806 323776 518862 323785
rect 518806 323711 518862 323720
rect 518820 315353 518848 323711
rect 518806 315344 518862 315353
rect 518806 315279 518862 315288
rect 520352 313126 520688 313154
rect 530656 313126 530992 313154
rect 520660 311778 520688 313126
rect 520648 311772 520700 311778
rect 520648 311714 520700 311720
rect 530964 311710 530992 313126
rect 540624 313126 540960 313154
rect 540624 311846 540652 313126
rect 541084 311846 541112 333254
rect 540612 311840 540664 311846
rect 540612 311782 540664 311788
rect 541072 311840 541124 311846
rect 541072 311782 541124 311788
rect 541636 311778 541664 335310
rect 542360 332648 542412 332654
rect 542360 332590 542412 332596
rect 542372 323785 542400 332590
rect 542358 323776 542414 323785
rect 542358 323711 542414 323720
rect 541624 311772 541676 311778
rect 541624 311714 541676 311720
rect 530952 311704 531004 311710
rect 530952 311646 531004 311652
rect 530308 309188 530360 309194
rect 530308 309130 530360 309136
rect 530320 306884 530348 309130
rect 519004 306326 520030 306354
rect 540638 306326 540836 306354
rect 519004 284238 519032 306326
rect 520016 284306 520044 286076
rect 530320 284306 530348 286076
rect 520004 284300 520056 284306
rect 520004 284242 520056 284248
rect 530308 284300 530360 284306
rect 530308 284242 530360 284248
rect 518992 284232 519044 284238
rect 540624 284209 540652 286076
rect 518992 284174 519044 284180
rect 540610 284200 540666 284209
rect 540808 284170 540836 306326
rect 542358 296304 542414 296313
rect 542358 296239 542414 296248
rect 542372 287881 542400 296239
rect 542358 287872 542414 287881
rect 542358 287807 542414 287816
rect 540610 284135 540666 284144
rect 540796 284164 540848 284170
rect 540796 284106 540848 284112
rect 530308 281648 530360 281654
rect 530308 281590 530360 281596
rect 530320 279970 530348 281590
rect 541624 281580 541676 281586
rect 541624 281522 541676 281528
rect 530320 279942 530656 279970
rect 520186 279304 520242 279313
rect 520242 279262 520352 279290
rect 540960 279262 541112 279290
rect 520186 279239 520242 279248
rect 518806 278080 518862 278089
rect 518806 278015 518862 278024
rect 518820 269793 518848 278015
rect 518806 269784 518862 269793
rect 518806 269719 518862 269728
rect 520352 259134 520688 259162
rect 530656 259134 530992 259162
rect 520660 256630 520688 259134
rect 520648 256624 520700 256630
rect 520648 256566 520700 256572
rect 530964 256562 530992 259134
rect 540624 259134 540960 259162
rect 540624 256698 540652 259134
rect 541084 256698 541112 279262
rect 540612 256692 540664 256698
rect 540612 256634 540664 256640
rect 541072 256692 541124 256698
rect 541072 256634 541124 256640
rect 541636 256630 541664 281522
rect 542360 278792 542412 278798
rect 542360 278734 542412 278740
rect 542372 269793 542400 278734
rect 542358 269784 542414 269793
rect 542358 269719 542414 269728
rect 541624 256624 541676 256630
rect 541624 256566 541676 256572
rect 530952 256556 531004 256562
rect 530952 256498 531004 256504
rect 530308 255332 530360 255338
rect 530308 255274 530360 255280
rect 530320 252892 530348 255274
rect 519004 252334 520030 252362
rect 540638 252334 540836 252362
rect 518806 242312 518862 242321
rect 518806 242247 518862 242256
rect 518820 234025 518848 242247
rect 518806 234016 518862 234025
rect 518806 233951 518862 233960
rect 519004 230246 519032 252334
rect 520016 230450 520044 232084
rect 530320 230450 530348 232084
rect 540624 230489 540652 232084
rect 540610 230480 540666 230489
rect 520004 230444 520056 230450
rect 520004 230386 520056 230392
rect 530308 230444 530360 230450
rect 540610 230415 540666 230424
rect 530308 230386 530360 230392
rect 540808 230314 540836 252334
rect 542358 242312 542414 242321
rect 542358 242247 542414 242256
rect 542372 233238 542400 242247
rect 542360 233232 542412 233238
rect 542360 233174 542412 233180
rect 540796 230308 540848 230314
rect 540796 230250 540848 230256
rect 518992 230240 519044 230246
rect 518992 230182 519044 230188
rect 530308 227860 530360 227866
rect 530308 227802 530360 227808
rect 520280 227792 520332 227798
rect 520280 227734 520332 227740
rect 520292 225978 520320 227734
rect 530320 225978 530348 227802
rect 541624 227792 541676 227798
rect 541624 227734 541676 227740
rect 520292 225950 520352 225978
rect 530320 225950 530656 225978
rect 540960 225270 541112 225298
rect 520352 205006 520688 205034
rect 530656 205006 530992 205034
rect 520660 202774 520688 205006
rect 520648 202768 520700 202774
rect 520648 202710 520700 202716
rect 530964 202706 530992 205006
rect 540624 205006 540960 205034
rect 540624 202842 540652 205006
rect 541084 202842 541112 225270
rect 540612 202836 540664 202842
rect 540612 202778 540664 202784
rect 541072 202836 541124 202842
rect 541072 202778 541124 202784
rect 541636 202774 541664 227734
rect 542358 224224 542414 224233
rect 542358 224159 542414 224168
rect 542372 215801 542400 224159
rect 542358 215792 542414 215801
rect 542358 215727 542414 215736
rect 541624 202768 541676 202774
rect 541624 202710 541676 202716
rect 530952 202700 531004 202706
rect 530952 202642 531004 202648
rect 530308 200184 530360 200190
rect 530308 200126 530360 200132
rect 530320 198900 530348 200126
rect 519004 198206 520030 198234
rect 540638 198206 540836 198234
rect 518806 196752 518862 196761
rect 518806 196687 518862 196696
rect 518820 188329 518848 196687
rect 518806 188320 518862 188329
rect 518806 188255 518862 188264
rect 519004 176594 519032 198206
rect 520016 176662 520044 178092
rect 530320 176662 530348 178092
rect 520004 176656 520056 176662
rect 520004 176598 520056 176604
rect 530308 176656 530360 176662
rect 530308 176598 530360 176604
rect 518992 176588 519044 176594
rect 518992 176530 519044 176536
rect 540624 176526 540652 178092
rect 540612 176520 540664 176526
rect 540612 176462 540664 176468
rect 540808 176458 540836 198206
rect 542358 188320 542414 188329
rect 542358 188255 542414 188264
rect 542372 179382 542400 188255
rect 542360 179376 542412 179382
rect 542360 179318 542412 179324
rect 540796 176452 540848 176458
rect 540796 176394 540848 176400
rect 530308 174072 530360 174078
rect 530308 174014 530360 174020
rect 541624 174072 541676 174078
rect 541624 174014 541676 174020
rect 520280 173936 520332 173942
rect 520280 173878 520332 173884
rect 520292 171986 520320 173878
rect 530320 171986 530348 174014
rect 520292 171958 520352 171986
rect 530320 171958 530656 171986
rect 540960 171290 541204 171306
rect 540960 171284 541216 171290
rect 540960 171278 541164 171284
rect 541164 171226 541216 171232
rect 520352 151014 520688 151042
rect 530656 151014 530992 151042
rect 520660 148986 520688 151014
rect 520648 148980 520700 148986
rect 520648 148922 520700 148928
rect 530964 148918 530992 151014
rect 540624 151014 540960 151042
rect 540624 149054 540652 151014
rect 540612 149048 540664 149054
rect 540612 148990 540664 148996
rect 541636 148986 541664 174014
rect 544384 171284 544436 171290
rect 544384 171226 544436 171232
rect 544396 149054 544424 171226
rect 544384 149048 544436 149054
rect 544384 148990 544436 148996
rect 541624 148980 541676 148986
rect 541624 148922 541676 148928
rect 530952 148912 531004 148918
rect 530952 148854 531004 148860
rect 530308 146396 530360 146402
rect 530308 146338 530360 146344
rect 530320 144908 530348 146338
rect 540612 146328 540664 146334
rect 540612 146270 540664 146276
rect 540624 144908 540652 146270
rect 519004 144214 520030 144242
rect 518806 134328 518862 134337
rect 518806 134263 518862 134272
rect 518820 125594 518848 134263
rect 518808 125588 518860 125594
rect 518808 125530 518860 125536
rect 519004 122602 519032 144214
rect 542358 142760 542414 142769
rect 542358 142695 542414 142704
rect 542372 134337 542400 142695
rect 542358 134328 542414 134337
rect 542358 134263 542414 134272
rect 520016 122806 520044 124100
rect 530320 122806 530348 124100
rect 520004 122800 520056 122806
rect 520004 122742 520056 122748
rect 530308 122800 530360 122806
rect 530308 122742 530360 122748
rect 540624 122738 540652 124100
rect 540612 122732 540664 122738
rect 540612 122674 540664 122680
rect 518992 122596 519044 122602
rect 518992 122538 519044 122544
rect 541624 120284 541676 120290
rect 541624 120226 541676 120232
rect 530308 120216 530360 120222
rect 530308 120158 530360 120164
rect 520280 120148 520332 120154
rect 520280 120090 520332 120096
rect 520292 117994 520320 120090
rect 530320 117994 530348 120158
rect 520292 117966 520352 117994
rect 530320 117966 530656 117994
rect 540960 117298 541204 117314
rect 540960 117292 541216 117298
rect 540960 117286 541164 117292
rect 541164 117234 541216 117240
rect 520352 97022 520688 97050
rect 530656 97022 530992 97050
rect 520660 95130 520688 97022
rect 520648 95124 520700 95130
rect 520648 95066 520700 95072
rect 530964 95062 530992 97022
rect 540624 97022 540960 97050
rect 540624 95198 540652 97022
rect 540612 95192 540664 95198
rect 540612 95134 540664 95140
rect 541636 95130 541664 120226
rect 544384 117292 544436 117298
rect 544384 117234 544436 117240
rect 544396 95198 544424 117234
rect 544384 95192 544436 95198
rect 544384 95134 544436 95140
rect 541624 95124 541676 95130
rect 541624 95066 541676 95072
rect 530952 95056 531004 95062
rect 530952 94998 531004 95004
rect 530308 92608 530360 92614
rect 530308 92550 530360 92556
rect 541716 92608 541768 92614
rect 541716 92550 541768 92556
rect 530320 90916 530348 92550
rect 540612 92540 540664 92546
rect 540612 92482 540664 92488
rect 541624 92540 541676 92546
rect 541624 92482 541676 92488
rect 540624 90916 540652 92482
rect 518912 90222 520030 90250
rect 518912 68882 518940 90222
rect 540888 71732 540940 71738
rect 540888 71674 540940 71680
rect 540900 70666 540928 71674
rect 540638 70638 540928 70666
rect 520016 68950 520044 70108
rect 530320 68950 530348 70108
rect 541636 68950 541664 92482
rect 541728 71738 541756 92550
rect 542360 89752 542412 89758
rect 542360 89694 542412 89700
rect 542372 80345 542400 89694
rect 542358 80336 542414 80345
rect 542358 80271 542414 80280
rect 541716 71732 541768 71738
rect 541716 71674 541768 71680
rect 520004 68944 520056 68950
rect 520004 68886 520056 68892
rect 530308 68944 530360 68950
rect 530308 68886 530360 68892
rect 541624 68944 541676 68950
rect 541624 68886 541676 68892
rect 518900 68876 518952 68882
rect 518900 68818 518952 68824
rect 530308 66360 530360 66366
rect 530308 66302 530360 66308
rect 520280 66292 520332 66298
rect 520280 66234 520332 66240
rect 520292 63866 520320 66234
rect 530320 63866 530348 66302
rect 541624 66292 541676 66298
rect 541624 66234 541676 66240
rect 520292 63838 520352 63866
rect 530320 63838 530656 63866
rect 540960 63294 541112 63322
rect 520352 43030 520688 43058
rect 530656 43030 530992 43058
rect 520660 41342 520688 43030
rect 520648 41336 520700 41342
rect 520648 41278 520700 41284
rect 530964 41274 530992 43030
rect 540624 43030 540960 43058
rect 540624 41410 540652 43030
rect 541084 41410 541112 63294
rect 540612 41404 540664 41410
rect 540612 41346 540664 41352
rect 541072 41404 541124 41410
rect 541072 41346 541124 41352
rect 541636 41342 541664 66234
rect 541716 60784 541768 60790
rect 541716 60726 541768 60732
rect 541624 41336 541676 41342
rect 541624 41278 541676 41284
rect 541728 41274 541756 60726
rect 542358 53816 542414 53825
rect 542358 53751 542414 53760
rect 542372 44130 542400 53751
rect 542360 44124 542412 44130
rect 542360 44066 542412 44072
rect 530952 41268 531004 41274
rect 530952 41210 531004 41216
rect 541716 41268 541768 41274
rect 541716 41210 541768 41216
rect 530308 38752 530360 38758
rect 530308 38694 530360 38700
rect 530320 36924 530348 38694
rect 540612 38684 540664 38690
rect 540612 38626 540664 38632
rect 540624 36924 540652 38626
rect 545776 38214 545804 674183
rect 547892 664006 548044 664034
rect 558012 664006 558348 664034
rect 547892 662318 547920 664006
rect 547880 662312 547932 662318
rect 547880 662254 547932 662260
rect 558012 661706 558040 664006
rect 568776 662386 568804 684270
rect 571338 674248 571394 674257
rect 571338 674183 571394 674192
rect 571352 665961 571380 674183
rect 571338 665952 571394 665961
rect 571338 665887 571394 665896
rect 568764 662380 568816 662386
rect 568764 662322 568816 662328
rect 558000 661700 558052 661706
rect 558000 661642 558052 661648
rect 558644 659728 558696 659734
rect 558644 659670 558696 659676
rect 558656 657900 558684 659670
rect 547984 657206 548366 657234
rect 568974 657206 569080 657234
rect 546406 647728 546462 647737
rect 546406 647663 546462 647672
rect 546420 620265 546448 647663
rect 547984 634642 548012 657206
rect 548076 637078 548366 637106
rect 547972 634636 548024 634642
rect 547972 634578 548024 634584
rect 548076 631122 548104 637078
rect 558656 634098 558684 637092
rect 568960 634778 568988 637092
rect 568948 634772 569000 634778
rect 568948 634714 569000 634720
rect 558644 634092 558696 634098
rect 558644 634034 558696 634040
rect 568948 634092 569000 634098
rect 568948 634034 569000 634040
rect 548340 632732 548392 632738
rect 548340 632674 548392 632680
rect 547892 631094 548104 631122
rect 546406 620256 546462 620265
rect 546406 620191 546462 620200
rect 547892 610706 547920 631094
rect 548352 630986 548380 632674
rect 548044 630958 548380 630986
rect 557998 630456 558054 630465
rect 558054 630414 558348 630442
rect 557998 630391 558054 630400
rect 568652 630278 568896 630306
rect 568764 625864 568816 625870
rect 568764 625806 568816 625812
rect 568776 610722 568804 625806
rect 547880 610700 547932 610706
rect 547880 610642 547932 610648
rect 548156 610700 548208 610706
rect 568652 610694 568804 610722
rect 548156 610642 548208 610648
rect 547892 610014 548044 610042
rect 547892 608394 547920 610014
rect 548168 608530 548196 610642
rect 558012 610014 558348 610042
rect 558012 608530 558040 610014
rect 568868 608598 568896 630278
rect 568960 625870 568988 634034
rect 569052 632738 569080 657206
rect 569040 632732 569092 632738
rect 569040 632674 569092 632680
rect 568948 625864 569000 625870
rect 568948 625806 569000 625812
rect 571338 620256 571394 620265
rect 571338 620191 571394 620200
rect 571352 611969 571380 620191
rect 580262 617536 580318 617545
rect 580262 617471 580318 617480
rect 571338 611960 571394 611969
rect 571338 611895 571394 611904
rect 568856 608592 568908 608598
rect 568856 608534 568908 608540
rect 548156 608524 548208 608530
rect 548156 608466 548208 608472
rect 558000 608524 558052 608530
rect 558000 608466 558052 608472
rect 547880 608388 547932 608394
rect 547880 608330 547932 608336
rect 558644 605872 558696 605878
rect 558644 605814 558696 605820
rect 558656 603908 558684 605814
rect 547984 603214 548366 603242
rect 568974 603214 569080 603242
rect 546406 593736 546462 593745
rect 546406 593671 546462 593680
rect 546420 566273 546448 593671
rect 547984 580854 548012 603214
rect 548076 583086 548366 583114
rect 547972 580848 548024 580854
rect 547972 580790 548024 580796
rect 548076 579986 548104 583086
rect 558656 580310 558684 583100
rect 568960 580990 568988 583100
rect 568948 580984 569000 580990
rect 568948 580926 569000 580932
rect 558644 580304 558696 580310
rect 558644 580246 558696 580252
rect 568764 580304 568816 580310
rect 568764 580246 568816 580252
rect 547892 579958 548104 579986
rect 546406 566264 546462 566273
rect 546406 566199 546462 566208
rect 547892 556170 547920 579958
rect 548340 578944 548392 578950
rect 548340 578886 548392 578892
rect 548352 576994 548380 578886
rect 548044 576966 548380 576994
rect 557998 576464 558054 576473
rect 558054 576422 558348 576450
rect 568776 576434 568804 580246
rect 569052 578950 569080 603214
rect 571338 602032 571394 602041
rect 571338 601967 571394 601976
rect 571352 593745 571380 601967
rect 571338 593736 571394 593745
rect 571338 593671 571394 593680
rect 569040 578944 569092 578950
rect 569040 578886 569092 578892
rect 568764 576428 568816 576434
rect 557998 576399 558054 576408
rect 568764 576370 568816 576376
rect 568652 576286 568896 576314
rect 568764 576224 568816 576230
rect 568764 576166 568816 576172
rect 568776 556730 568804 576166
rect 568652 556702 568804 556730
rect 547880 556164 547932 556170
rect 547880 556106 547932 556112
rect 548156 556164 548208 556170
rect 548156 556106 548208 556112
rect 547892 556022 548044 556050
rect 547892 554538 547920 556022
rect 548168 554674 548196 556106
rect 558012 556022 558348 556050
rect 558012 554674 558040 556022
rect 568868 554742 568896 576286
rect 571338 574696 571394 574705
rect 571338 574631 571394 574640
rect 571352 566273 571380 574631
rect 571338 566264 571394 566273
rect 571338 566199 571394 566208
rect 568856 554736 568908 554742
rect 568856 554678 568908 554684
rect 548156 554668 548208 554674
rect 548156 554610 548208 554616
rect 558000 554668 558052 554674
rect 558000 554610 558052 554616
rect 547880 554532 547932 554538
rect 547880 554474 547932 554480
rect 558644 552084 558696 552090
rect 558644 552026 558696 552032
rect 558656 549916 558684 552026
rect 547984 549222 548366 549250
rect 568974 549222 569080 549250
rect 546406 539744 546462 539753
rect 546406 539679 546462 539688
rect 546420 512281 546448 539679
rect 547984 526998 548012 549222
rect 548076 529094 548366 529122
rect 547972 526992 548024 526998
rect 547972 526934 548024 526940
rect 548076 523682 548104 529094
rect 558656 526454 558684 529108
rect 568960 527134 568988 529108
rect 568948 527128 569000 527134
rect 568948 527070 569000 527076
rect 558644 526448 558696 526454
rect 558644 526390 558696 526396
rect 568948 526448 569000 526454
rect 568948 526390 569000 526396
rect 548340 525088 548392 525094
rect 548340 525030 548392 525036
rect 547892 523654 548104 523682
rect 546406 512272 546462 512281
rect 546406 512207 546462 512216
rect 547892 502722 547920 523654
rect 548352 522866 548380 525030
rect 548044 522838 548380 522866
rect 568652 522566 568896 522594
rect 557998 522472 558054 522481
rect 558054 522430 558348 522458
rect 557998 522407 558054 522416
rect 568868 522306 568896 522566
rect 568856 522300 568908 522306
rect 568856 522242 568908 522248
rect 568960 522186 568988 526390
rect 569052 525094 569080 549222
rect 571338 548040 571394 548049
rect 571338 547975 571394 547984
rect 571352 539753 571380 547975
rect 571338 539744 571394 539753
rect 571338 539679 571394 539688
rect 569040 525088 569092 525094
rect 569040 525030 569092 525036
rect 568776 522158 568988 522186
rect 568776 502738 568804 522158
rect 568856 522096 568908 522102
rect 568856 522038 568908 522044
rect 547880 502716 547932 502722
rect 547880 502658 547932 502664
rect 548156 502716 548208 502722
rect 568652 502710 568804 502738
rect 548156 502658 548208 502664
rect 547892 502030 548044 502058
rect 547892 500750 547920 502030
rect 548168 500886 548196 502658
rect 558012 502030 558348 502058
rect 558012 500886 558040 502030
rect 568868 500954 568896 522038
rect 568946 520704 569002 520713
rect 568946 520639 569002 520648
rect 568960 512825 568988 520639
rect 568946 512816 569002 512825
rect 568946 512751 569002 512760
rect 568856 500948 568908 500954
rect 568856 500890 568908 500896
rect 548156 500880 548208 500886
rect 548156 500822 548208 500828
rect 558000 500880 558052 500886
rect 558000 500822 558052 500828
rect 547880 500744 547932 500750
rect 547880 500686 547932 500692
rect 558644 498228 558696 498234
rect 558644 498170 558696 498176
rect 558656 495924 558684 498170
rect 547984 495230 548366 495258
rect 568974 495230 569080 495258
rect 546406 485752 546462 485761
rect 546406 485687 546462 485696
rect 546420 458289 546448 485687
rect 547984 473210 548012 495230
rect 548076 475102 548366 475130
rect 547972 473204 548024 473210
rect 547972 473146 548024 473152
rect 548076 470594 548104 475102
rect 558656 472666 558684 475116
rect 568960 473346 568988 475116
rect 568948 473340 569000 473346
rect 568948 473282 569000 473288
rect 558644 472660 558696 472666
rect 558644 472602 558696 472608
rect 568764 472660 568816 472666
rect 568764 472602 568816 472608
rect 548340 471300 548392 471306
rect 548340 471242 548392 471248
rect 547892 470566 548104 470594
rect 546406 458280 546462 458289
rect 546406 458215 546462 458224
rect 547892 448458 547920 470566
rect 548352 468874 548380 471242
rect 548044 468846 548380 468874
rect 557998 468480 558054 468489
rect 558054 468438 558348 468466
rect 568776 468450 568804 472602
rect 569052 471306 569080 495230
rect 571338 485752 571394 485761
rect 571338 485687 571394 485696
rect 571352 477329 571380 485687
rect 571338 477320 571394 477329
rect 571338 477255 571394 477264
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 569040 471300 569092 471306
rect 569040 471242 569092 471248
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 568764 468444 568816 468450
rect 557998 468415 558054 468424
rect 568764 468386 568816 468392
rect 568652 468302 568896 468330
rect 568764 468240 568816 468246
rect 568764 468182 568816 468188
rect 568776 448746 568804 468182
rect 568652 448718 568804 448746
rect 547880 448452 547932 448458
rect 547880 448394 547932 448400
rect 548156 448452 548208 448458
rect 548156 448394 548208 448400
rect 547892 448038 548044 448066
rect 547892 445670 547920 448038
rect 547880 445664 547932 445670
rect 547880 445606 547932 445612
rect 548168 445602 548196 448394
rect 558012 448038 558348 448066
rect 558012 445602 558040 448038
rect 568868 445738 568896 468302
rect 571338 466712 571394 466721
rect 571338 466647 571394 466656
rect 571352 458289 571380 466647
rect 571338 458280 571394 458289
rect 571338 458215 571394 458224
rect 568856 445732 568908 445738
rect 568856 445674 568908 445680
rect 548156 445596 548208 445602
rect 548156 445538 548208 445544
rect 558000 445596 558052 445602
rect 558000 445538 558052 445544
rect 558644 444440 558696 444446
rect 558644 444382 558696 444388
rect 558656 441932 558684 444382
rect 547984 441238 548366 441266
rect 568974 441238 569080 441266
rect 546406 431760 546462 431769
rect 546406 431695 546462 431704
rect 546420 404297 546448 431695
rect 547984 419354 548012 441238
rect 548076 421110 548366 421138
rect 547972 419348 548024 419354
rect 547972 419290 548024 419296
rect 548076 416922 548104 421110
rect 558656 418810 558684 421124
rect 568960 419490 568988 421124
rect 568948 419484 569000 419490
rect 568948 419426 569000 419432
rect 558644 418804 558696 418810
rect 558644 418746 558696 418752
rect 568948 418804 569000 418810
rect 568948 418746 569000 418752
rect 548340 417444 548392 417450
rect 548340 417386 548392 417392
rect 547892 416894 548104 416922
rect 546406 404288 546462 404297
rect 546406 404223 546462 404232
rect 547892 394738 547920 416894
rect 548352 414882 548380 417386
rect 548044 414854 548380 414882
rect 557998 414488 558054 414497
rect 558054 414446 558348 414474
rect 557998 414423 558054 414432
rect 568652 414310 568896 414338
rect 568764 410916 568816 410922
rect 568764 410858 568816 410864
rect 568776 394754 568804 410858
rect 547880 394732 547932 394738
rect 547880 394674 547932 394680
rect 548156 394732 548208 394738
rect 568652 394726 568804 394754
rect 548156 394674 548208 394680
rect 547892 394046 548044 394074
rect 547892 391746 547920 394046
rect 548168 391882 548196 394674
rect 558012 394046 558348 394074
rect 558012 391882 558040 394046
rect 568868 391950 568896 414310
rect 568960 410922 568988 418746
rect 569052 417450 569080 441238
rect 571338 431760 571394 431769
rect 571338 431695 571394 431704
rect 571352 423337 571380 431695
rect 571338 423328 571394 423337
rect 571338 423263 571394 423272
rect 569040 417444 569092 417450
rect 569040 417386 569092 417392
rect 568948 410916 569000 410922
rect 568948 410858 569000 410864
rect 571338 404288 571394 404297
rect 571338 404223 571394 404232
rect 571352 396001 571380 404223
rect 571338 395992 571394 396001
rect 571338 395927 571394 395936
rect 568856 391944 568908 391950
rect 568856 391886 568908 391892
rect 548156 391876 548208 391882
rect 548156 391818 548208 391824
rect 558000 391876 558052 391882
rect 558000 391818 558052 391824
rect 547880 391740 547932 391746
rect 547880 391682 547932 391688
rect 558644 389224 558696 389230
rect 558644 389166 558696 389172
rect 558656 387940 558684 389166
rect 547984 387246 548366 387274
rect 568974 387246 569080 387274
rect 546406 377768 546462 377777
rect 546406 377703 546462 377712
rect 546420 350305 546448 377703
rect 547984 365566 548012 387246
rect 548076 367118 548366 367146
rect 547972 365560 548024 365566
rect 547972 365502 548024 365508
rect 548076 364334 548104 367118
rect 558656 365022 558684 367132
rect 568960 365702 568988 367132
rect 568948 365696 569000 365702
rect 568948 365638 569000 365644
rect 558644 365016 558696 365022
rect 558644 364958 558696 364964
rect 568764 365016 568816 365022
rect 568764 364958 568816 364964
rect 547892 364306 548104 364334
rect 546406 350296 546462 350305
rect 546406 350231 546462 350240
rect 547892 340746 547920 364306
rect 548340 363656 548392 363662
rect 548340 363598 548392 363604
rect 548352 360890 548380 363598
rect 548044 360862 548380 360890
rect 557998 360496 558054 360505
rect 558054 360454 558348 360482
rect 568776 360466 568804 364958
rect 569052 363662 569080 387246
rect 579802 378448 579858 378457
rect 579802 378383 579858 378392
rect 579816 378214 579844 378383
rect 569224 378208 569276 378214
rect 569224 378150 569276 378156
rect 579804 378208 579856 378214
rect 579804 378150 579856 378156
rect 569040 363656 569092 363662
rect 569040 363598 569092 363604
rect 568764 360460 568816 360466
rect 557998 360431 558054 360440
rect 568764 360402 568816 360408
rect 568652 360318 568896 360346
rect 568764 360256 568816 360262
rect 568764 360198 568816 360204
rect 568776 340762 568804 360198
rect 547880 340740 547932 340746
rect 547880 340682 547932 340688
rect 548156 340740 548208 340746
rect 568652 340734 568804 340762
rect 548156 340682 548208 340688
rect 547892 340054 548044 340082
rect 547892 337890 547920 340054
rect 548168 338026 548196 340682
rect 558012 340054 558348 340082
rect 558012 338026 558040 340054
rect 568868 338094 568896 360318
rect 568856 338088 568908 338094
rect 568856 338030 568908 338036
rect 548156 338020 548208 338026
rect 548156 337962 548208 337968
rect 558000 338020 558052 338026
rect 558000 337962 558052 337968
rect 547880 337884 547932 337890
rect 547880 337826 547932 337832
rect 558644 335368 558696 335374
rect 558644 335310 558696 335316
rect 558656 333948 558684 335310
rect 547984 333254 548366 333282
rect 568974 333254 569080 333282
rect 546406 323776 546462 323785
rect 546406 323711 546462 323720
rect 546420 296313 546448 323711
rect 547984 311710 548012 333254
rect 548076 313126 548366 313154
rect 547972 311704 548024 311710
rect 547972 311646 548024 311652
rect 548076 309754 548104 313126
rect 558656 311166 558684 313140
rect 568960 311846 568988 313140
rect 568948 311840 569000 311846
rect 568948 311782 569000 311788
rect 558644 311160 558696 311166
rect 558644 311102 558696 311108
rect 568948 311160 569000 311166
rect 568948 311102 569000 311108
rect 547892 309726 548104 309754
rect 548340 309800 548392 309806
rect 548340 309742 548392 309748
rect 546406 296304 546462 296313
rect 546406 296239 546462 296248
rect 547892 286210 547920 309726
rect 548352 306898 548380 309742
rect 548044 306870 548380 306898
rect 557998 306504 558054 306513
rect 558054 306462 558348 306490
rect 557998 306439 558054 306448
rect 568652 306338 568896 306354
rect 568652 306332 568908 306338
rect 568652 306326 568856 306332
rect 568856 306274 568908 306280
rect 568856 306128 568908 306134
rect 568856 306070 568908 306076
rect 568764 304292 568816 304298
rect 568764 304234 568816 304240
rect 568776 286770 568804 304234
rect 568652 286742 568804 286770
rect 547880 286204 547932 286210
rect 547880 286146 547932 286152
rect 548156 286204 548208 286210
rect 548156 286146 548208 286152
rect 547892 286062 548044 286090
rect 547892 284238 547920 286062
rect 547880 284232 547932 284238
rect 547880 284174 547932 284180
rect 548168 284170 548196 286146
rect 558012 286062 558348 286090
rect 558012 284170 558040 286062
rect 568868 284306 568896 306070
rect 568960 304298 568988 311102
rect 569052 309806 569080 333254
rect 569040 309800 569092 309806
rect 569040 309742 569092 309748
rect 568948 304292 569000 304298
rect 568948 304234 569000 304240
rect 568856 284300 568908 284306
rect 568856 284242 568908 284248
rect 548156 284164 548208 284170
rect 548156 284106 548208 284112
rect 558000 284164 558052 284170
rect 558000 284106 558052 284112
rect 558644 281580 558696 281586
rect 558644 281522 558696 281528
rect 558656 279956 558684 281522
rect 547984 279262 548366 279290
rect 568974 279262 569080 279290
rect 546406 269784 546462 269793
rect 546406 269719 546462 269728
rect 546420 242321 546448 269719
rect 547984 256562 548012 279262
rect 548076 259134 548366 259162
rect 547972 256556 548024 256562
rect 547972 256498 548024 256504
rect 548076 253178 548104 259134
rect 558656 256086 558684 259148
rect 568960 256698 568988 259148
rect 568948 256692 569000 256698
rect 568948 256634 569000 256640
rect 558644 256080 558696 256086
rect 558644 256022 558696 256028
rect 568948 256080 569000 256086
rect 568948 256022 569000 256028
rect 548340 256012 548392 256018
rect 548340 255954 548392 255960
rect 547892 253150 548104 253178
rect 546406 242312 546462 242321
rect 546406 242247 546462 242256
rect 547892 232762 547920 253150
rect 548352 252906 548380 255954
rect 548044 252878 548380 252906
rect 557998 252648 558054 252657
rect 558054 252606 558348 252634
rect 557998 252583 558054 252592
rect 568652 252334 568896 252362
rect 568764 249144 568816 249150
rect 568764 249086 568816 249092
rect 568776 232778 568804 249086
rect 547880 232756 547932 232762
rect 547880 232698 547932 232704
rect 548156 232756 548208 232762
rect 568652 232750 568804 232778
rect 548156 232698 548208 232704
rect 547892 232070 548044 232098
rect 547892 230246 547920 232070
rect 548168 230382 548196 232698
rect 558012 232070 558348 232098
rect 558012 230382 558040 232070
rect 568868 230450 568896 252334
rect 568960 249150 568988 256022
rect 569052 256018 569080 279262
rect 569040 256012 569092 256018
rect 569040 255954 569092 255960
rect 568948 249144 569000 249150
rect 568948 249086 569000 249092
rect 568856 230444 568908 230450
rect 568856 230386 568908 230392
rect 548156 230376 548208 230382
rect 548156 230318 548208 230324
rect 558000 230376 558052 230382
rect 558000 230318 558052 230324
rect 547880 230240 547932 230246
rect 547880 230182 547932 230188
rect 558644 227792 558696 227798
rect 558644 227734 558696 227740
rect 558656 225964 558684 227734
rect 547984 225270 548366 225298
rect 568974 225270 569080 225298
rect 546406 215792 546462 215801
rect 546406 215727 546462 215736
rect 546420 188329 546448 215727
rect 547984 202706 548012 225270
rect 548076 205006 548366 205034
rect 547972 202700 548024 202706
rect 547972 202642 548024 202648
rect 547144 200184 547196 200190
rect 547144 200126 547196 200132
rect 546406 188320 546462 188329
rect 546406 188255 546462 188264
rect 547156 176526 547184 200126
rect 548076 200114 548104 205006
rect 558656 202162 558684 205020
rect 568960 202842 568988 205020
rect 568948 202836 569000 202842
rect 568948 202778 569000 202784
rect 558644 202156 558696 202162
rect 558644 202098 558696 202104
rect 568764 202156 568816 202162
rect 568764 202098 568816 202104
rect 548340 200796 548392 200802
rect 548340 200738 548392 200744
rect 547892 200086 548104 200114
rect 547892 178702 547920 200086
rect 548352 198914 548380 200738
rect 558000 200184 558052 200190
rect 558000 200126 558052 200132
rect 548044 198886 548380 198914
rect 558012 198914 558040 200126
rect 558012 198886 558348 198914
rect 568776 198354 568804 202098
rect 569052 200802 569080 225270
rect 569040 200796 569092 200802
rect 569040 200738 569092 200744
rect 568764 198348 568816 198354
rect 568764 198290 568816 198296
rect 568652 198206 568896 198234
rect 568764 198144 568816 198150
rect 568764 198086 568816 198092
rect 568776 178786 568804 198086
rect 568652 178758 568804 178786
rect 547880 178696 547932 178702
rect 547880 178638 547932 178644
rect 548156 178696 548208 178702
rect 548156 178638 548208 178644
rect 547892 178078 548044 178106
rect 547892 176594 547920 178078
rect 547880 176588 547932 176594
rect 547880 176530 547932 176536
rect 548168 176526 548196 178638
rect 558012 178078 558348 178106
rect 558012 176526 558040 178078
rect 568868 176662 568896 198206
rect 568856 176656 568908 176662
rect 568856 176598 568908 176604
rect 547144 176520 547196 176526
rect 547144 176462 547196 176468
rect 548156 176520 548208 176526
rect 548156 176462 548208 176468
rect 558000 176520 558052 176526
rect 558000 176462 558052 176468
rect 558644 174072 558696 174078
rect 558644 174014 558696 174020
rect 558656 171972 558684 174014
rect 547892 171278 548366 171306
rect 568974 171278 569080 171306
rect 547892 171170 547920 171278
rect 547800 171142 547920 171170
rect 546406 161800 546462 161809
rect 546406 161735 546462 161744
rect 546420 134337 546448 161735
rect 547800 161474 547828 171142
rect 547156 161446 547828 161474
rect 547156 148918 547184 161446
rect 547892 151014 548366 151042
rect 547144 148912 547196 148918
rect 547144 148854 547196 148860
rect 547144 146328 547196 146334
rect 547144 146270 547196 146276
rect 546406 134328 546462 134337
rect 546406 134263 546462 134272
rect 547156 122738 547184 146270
rect 547892 124710 547920 151014
rect 558656 148374 558684 151028
rect 568960 149054 568988 151028
rect 568948 149048 569000 149054
rect 568948 148990 569000 148996
rect 558644 148368 558696 148374
rect 558644 148310 558696 148316
rect 568948 148368 569000 148374
rect 568948 148310 569000 148316
rect 548340 146940 548392 146946
rect 548340 146882 548392 146888
rect 548352 144922 548380 146882
rect 558000 146328 558052 146334
rect 558000 146270 558052 146276
rect 548044 144894 548380 144922
rect 558012 144922 558040 146270
rect 558012 144894 558348 144922
rect 568652 144214 568896 144242
rect 568764 142860 568816 142866
rect 568764 142802 568816 142808
rect 568776 124794 568804 142802
rect 568652 124766 568804 124794
rect 547880 124704 547932 124710
rect 547880 124646 547932 124652
rect 548156 124704 548208 124710
rect 548156 124646 548208 124652
rect 547892 124086 548044 124114
rect 547144 122732 547196 122738
rect 547144 122674 547196 122680
rect 547892 122602 547920 124086
rect 548168 122738 548196 124646
rect 558012 124086 558348 124114
rect 558012 122738 558040 124086
rect 568868 122806 568896 144214
rect 568960 142866 568988 148310
rect 569052 146946 569080 171278
rect 569040 146940 569092 146946
rect 569040 146882 569092 146888
rect 568948 142860 569000 142866
rect 568948 142802 569000 142808
rect 568856 122800 568908 122806
rect 568856 122742 568908 122748
rect 548156 122732 548208 122738
rect 548156 122674 548208 122680
rect 558000 122732 558052 122738
rect 558000 122674 558052 122680
rect 547880 122596 547932 122602
rect 547880 122538 547932 122544
rect 558644 120284 558696 120290
rect 558644 120226 558696 120232
rect 558656 117980 558684 120226
rect 547156 117286 548366 117314
rect 568974 117286 569080 117314
rect 546406 107808 546462 107817
rect 546406 107743 546462 107752
rect 546420 80345 546448 107743
rect 547156 95062 547184 117286
rect 547892 97022 548366 97050
rect 547144 95056 547196 95062
rect 547144 94998 547196 95004
rect 546406 80336 546462 80345
rect 546406 80271 546462 80280
rect 547892 70718 547920 97022
rect 558656 94518 558684 97036
rect 568960 95198 568988 97036
rect 568948 95192 569000 95198
rect 568948 95134 569000 95140
rect 558644 94512 558696 94518
rect 558644 94454 558696 94460
rect 568764 94512 568816 94518
rect 568764 94454 568816 94460
rect 548340 93152 548392 93158
rect 548340 93094 548392 93100
rect 548352 90930 548380 93094
rect 558000 92608 558052 92614
rect 558000 92550 558052 92556
rect 548044 90902 548380 90930
rect 558012 90930 558040 92550
rect 568580 92540 568632 92546
rect 568580 92482 568632 92488
rect 568592 91066 568620 92482
rect 568592 91038 568666 91066
rect 558012 90902 558348 90930
rect 568638 90916 568666 91038
rect 547880 70712 547932 70718
rect 547880 70654 547932 70660
rect 548156 70712 548208 70718
rect 568776 70666 568804 94454
rect 569052 93158 569080 117286
rect 569040 93152 569092 93158
rect 569040 93094 569092 93100
rect 548156 70654 548208 70660
rect 547892 70094 548044 70122
rect 547892 68882 547920 70094
rect 548168 69018 548196 70654
rect 568652 70638 568804 70666
rect 558012 70094 558348 70122
rect 558012 69018 558040 70094
rect 548156 69012 548208 69018
rect 548156 68954 548208 68960
rect 558000 69012 558052 69018
rect 558000 68954 558052 68960
rect 547880 68876 547932 68882
rect 547880 68818 547932 68824
rect 558644 66292 558696 66298
rect 558644 66234 558696 66240
rect 558656 63852 558684 66234
rect 548076 63294 548366 63322
rect 568974 63294 569080 63322
rect 548076 60790 548104 63294
rect 548064 60784 548116 60790
rect 548064 60726 548116 60732
rect 546406 53272 546462 53281
rect 546406 53207 546462 53216
rect 545764 38208 545816 38214
rect 545764 38150 545816 38156
rect 519004 36230 520030 36258
rect 518164 13388 518216 13394
rect 518164 13330 518216 13336
rect 519004 13326 519032 36230
rect 542358 34912 542414 34921
rect 542358 34847 542414 34856
rect 542372 26353 542400 34847
rect 546420 26353 546448 53207
rect 547892 43030 548366 43058
rect 542358 26344 542414 26353
rect 542358 26279 542414 26288
rect 546406 26344 546462 26353
rect 546406 26279 546462 26288
rect 520016 13394 520044 16116
rect 530320 13394 530348 16116
rect 540624 13433 540652 16116
rect 547892 13802 547920 43030
rect 558656 40730 558684 43044
rect 568960 41410 568988 43044
rect 568948 41404 569000 41410
rect 568948 41346 569000 41352
rect 558644 40724 558696 40730
rect 558644 40666 558696 40672
rect 568856 40724 568908 40730
rect 568856 40666 568908 40672
rect 548340 39432 548392 39438
rect 548340 39374 548392 39380
rect 548352 36938 548380 39374
rect 548044 36910 548380 36938
rect 557998 36544 558054 36553
rect 558054 36502 558348 36530
rect 557998 36479 558054 36488
rect 568652 36230 568804 36258
rect 568776 16946 568804 36230
rect 568868 35894 568896 40666
rect 569052 39438 569080 63294
rect 569040 39432 569092 39438
rect 569040 39374 569092 39380
rect 569236 36786 569264 378150
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 571338 350296 571394 350305
rect 571338 350231 571394 350240
rect 571352 342009 571380 350231
rect 571338 342000 571394 342009
rect 571338 341935 571394 341944
rect 580078 325272 580134 325281
rect 580078 325207 580134 325216
rect 580092 324358 580120 325207
rect 574744 324352 574796 324358
rect 574744 324294 574796 324300
rect 580080 324352 580132 324358
rect 580080 324294 580132 324300
rect 571338 296304 571394 296313
rect 571338 296239 571394 296248
rect 571352 288017 571380 296239
rect 571338 288008 571394 288017
rect 571338 287943 571394 287952
rect 571338 242312 571394 242321
rect 571338 242247 571394 242256
rect 571352 234025 571380 242247
rect 571338 234016 571394 234025
rect 571338 233951 571394 233960
rect 571338 224088 571394 224097
rect 571338 224023 571394 224032
rect 571352 215801 571380 224023
rect 571338 215792 571394 215801
rect 571338 215727 571394 215736
rect 571338 196752 571394 196761
rect 571338 196687 571394 196696
rect 569316 191888 569368 191894
rect 569316 191830 569368 191836
rect 569328 39370 569356 191830
rect 571352 188329 571380 196687
rect 571338 188320 571394 188329
rect 571338 188255 571394 188264
rect 571338 170096 571394 170105
rect 571338 170031 571394 170040
rect 571352 161809 571380 170031
rect 571338 161800 571394 161809
rect 571338 161735 571394 161744
rect 569408 151836 569460 151842
rect 569408 151778 569460 151784
rect 569316 39364 569368 39370
rect 569316 39306 569368 39312
rect 569420 38146 569448 151778
rect 571338 134328 571394 134337
rect 571338 134263 571394 134272
rect 571352 125594 571380 134263
rect 571340 125588 571392 125594
rect 571340 125530 571392 125536
rect 571338 116104 571394 116113
rect 571338 116039 571394 116048
rect 569500 111852 569552 111858
rect 569500 111794 569552 111800
rect 569512 38282 569540 111794
rect 571352 107817 571380 116039
rect 571338 107808 571394 107817
rect 571338 107743 571394 107752
rect 571338 88768 571394 88777
rect 571338 88703 571394 88712
rect 571352 80345 571380 88703
rect 571338 80336 571394 80345
rect 571338 80271 571394 80280
rect 571338 53816 571394 53825
rect 571338 53751 571394 53760
rect 571352 45393 571380 53751
rect 571338 45384 571394 45393
rect 571338 45319 571394 45328
rect 569500 38276 569552 38282
rect 569500 38218 569552 38224
rect 569408 38140 569460 38146
rect 569408 38082 569460 38088
rect 569224 36780 569276 36786
rect 569224 36722 569276 36728
rect 568868 35866 569080 35894
rect 568776 16918 568988 16946
rect 568488 16720 568540 16726
rect 568540 16668 568652 16674
rect 568488 16662 568652 16668
rect 568500 16646 568652 16662
rect 548030 15858 548058 16116
rect 547984 15830 548058 15858
rect 558012 16102 558348 16130
rect 547880 13796 547932 13802
rect 547880 13738 547932 13744
rect 540610 13424 540666 13433
rect 520004 13388 520056 13394
rect 520004 13330 520056 13336
rect 530308 13388 530360 13394
rect 540610 13359 540666 13368
rect 530308 13330 530360 13336
rect 547984 13326 548012 15830
rect 558012 13802 558040 16102
rect 558000 13796 558052 13802
rect 558000 13738 558052 13744
rect 568960 13394 568988 16918
rect 569052 16726 569080 35866
rect 571338 34776 571394 34785
rect 571338 34711 571394 34720
rect 571352 26353 571380 34711
rect 571338 26344 571394 26353
rect 571338 26279 571394 26288
rect 569040 16720 569092 16726
rect 569040 16662 569092 16668
rect 574756 13734 574784 324294
rect 578882 272232 578938 272241
rect 578882 272167 578938 272176
rect 574744 13728 574796 13734
rect 574744 13670 574796 13676
rect 568948 13388 569000 13394
rect 568948 13330 569000 13336
rect 484952 13320 485004 13326
rect 484952 13262 485004 13268
rect 491392 13320 491444 13326
rect 491392 13262 491444 13268
rect 518992 13320 519044 13326
rect 518992 13262 519044 13268
rect 547972 13320 548024 13326
rect 547972 13262 548024 13268
rect 352012 13252 352064 13258
rect 352012 13194 352064 13200
rect 362316 13252 362368 13258
rect 362316 13194 362368 13200
rect 400956 13252 401008 13258
rect 400956 13194 401008 13200
rect 434812 13252 434864 13258
rect 434812 13194 434864 13200
rect 463700 13252 463752 13258
rect 463700 13194 463752 13200
rect 211252 13184 211304 13190
rect 211252 13126 211304 13132
rect 240048 13184 240100 13190
rect 240048 13126 240100 13132
rect 268016 13184 268068 13190
rect 268016 13126 268068 13132
rect 278320 13184 278372 13190
rect 278320 13126 278372 13132
rect 316960 13184 317012 13190
rect 316960 13126 317012 13132
rect 324044 13184 324096 13190
rect 324044 13126 324096 13132
rect 334348 13184 334400 13190
rect 334348 13126 334400 13132
rect 345756 13184 345808 13190
rect 345756 13126 345808 13132
rect 72056 13116 72108 13122
rect 72056 13058 72108 13064
rect 127072 13116 127124 13122
rect 127072 13058 127124 13064
rect 156052 13116 156104 13122
rect 156052 13058 156104 13064
rect 68284 13048 68336 13054
rect 68284 12990 68336 12996
rect 578896 12986 578924 272167
rect 580078 232384 580134 232393
rect 580078 232319 580134 232328
rect 580092 231878 580120 232319
rect 580080 231872 580132 231878
rect 580080 231814 580132 231820
rect 580078 192536 580134 192545
rect 580078 192471 580134 192480
rect 580092 191894 580120 192471
rect 580080 191888 580132 191894
rect 580080 191830 580132 191836
rect 580078 152688 580134 152697
rect 580078 152623 580134 152632
rect 580092 151842 580120 152623
rect 580080 151836 580132 151842
rect 580080 151778 580132 151784
rect 580078 112840 580134 112849
rect 580078 112775 580134 112784
rect 580092 111858 580120 112775
rect 580080 111852 580132 111858
rect 580080 111794 580132 111800
rect 580078 72992 580134 73001
rect 580078 72927 580134 72936
rect 580092 13666 580120 72927
rect 580080 13660 580132 13666
rect 580080 13602 580132 13608
rect 580184 13530 580212 351863
rect 580172 13524 580224 13530
rect 580172 13466 580224 13472
rect 580276 13462 580304 617471
rect 580354 591016 580410 591025
rect 580354 590951 580410 590960
rect 580368 36718 580396 590951
rect 580446 564360 580502 564369
rect 580446 564295 580502 564304
rect 580460 38010 580488 564295
rect 580538 537840 580594 537849
rect 580538 537775 580594 537784
rect 580448 38004 580500 38010
rect 580448 37946 580500 37952
rect 580356 36712 580408 36718
rect 580356 36654 580408 36660
rect 580552 36650 580580 537775
rect 580630 511320 580686 511329
rect 580630 511255 580686 511264
rect 580644 38078 580672 511255
rect 580722 484664 580778 484673
rect 580722 484599 580778 484608
rect 580632 38072 580684 38078
rect 580632 38014 580684 38020
rect 580540 36644 580592 36650
rect 580540 36586 580592 36592
rect 580736 13598 580764 484599
rect 580814 431624 580870 431633
rect 580814 431559 580870 431568
rect 580828 36582 580856 431559
rect 580906 404968 580962 404977
rect 580906 404903 580962 404912
rect 580920 37942 580948 404903
rect 580908 37936 580960 37942
rect 580908 37878 580960 37884
rect 580816 36576 580868 36582
rect 580816 36518 580868 36524
rect 580908 35964 580960 35970
rect 580908 35906 580960 35912
rect 580920 33153 580948 35906
rect 580906 33144 580962 33153
rect 580906 33079 580962 33088
rect 580724 13592 580776 13598
rect 580724 13534 580776 13540
rect 580264 13456 580316 13462
rect 580264 13398 580316 13404
rect 578884 12980 578936 12986
rect 578884 12922 578936 12928
rect 64236 3732 64288 3738
rect 64236 3674 64288 3680
rect 125876 3732 125928 3738
rect 125876 3674 125928 3680
rect 64144 3664 64196 3670
rect 64144 3606 64196 3612
rect 61476 3596 61528 3602
rect 61476 3538 61528 3544
rect 48320 3460 48372 3466
rect 48320 3402 48372 3408
rect 61384 3460 61436 3466
rect 61384 3402 61436 3408
rect 125888 480 125916 3674
rect 126980 3664 127032 3670
rect 126980 3606 127032 3612
rect 126992 480 127020 3606
rect 132960 3596 133012 3602
rect 132960 3538 133012 3544
rect 129372 3528 129424 3534
rect 129372 3470 129424 3476
rect 129384 480 129412 3470
rect 132972 480 133000 3538
rect 136456 3460 136508 3466
rect 136456 3402 136508 3408
rect 136468 480 136496 3402
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 2778 606056 2834 606112
rect 2962 527856 3018 527912
rect 2778 449520 2834 449576
rect 3146 410488 3202 410544
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 2778 345344 2834 345400
rect 3146 293120 3202 293176
rect 3238 241032 3294 241088
rect 2778 188808 2834 188864
rect 2778 149776 2834 149832
rect 3330 136740 3386 136776
rect 3330 136720 3332 136740
rect 3332 136720 3384 136740
rect 3384 136720 3386 136740
rect 3330 84652 3386 84688
rect 3330 84632 3332 84652
rect 3332 84632 3384 84652
rect 3384 84632 3386 84652
rect 3330 58520 3386 58576
rect 2962 45464 3018 45520
rect 3514 658144 3570 658200
rect 3514 579944 3570 580000
rect 3606 553832 3662 553888
rect 3606 501744 3662 501800
rect 3698 475632 3754 475688
rect 3790 358400 3846 358456
rect 3882 306176 3938 306232
rect 3790 19352 3846 19408
rect 3974 254088 4030 254144
rect 4066 97552 4122 97608
rect 11886 34448 11942 34504
rect 13634 674192 13690 674248
rect 13634 665896 13690 665952
rect 13542 620200 13598 620256
rect 13542 611904 13598 611960
rect 13542 601976 13598 602032
rect 13542 593680 13598 593736
rect 13542 574640 13598 574696
rect 13542 566208 13598 566264
rect 13542 547984 13598 548040
rect 13542 539688 13598 539744
rect 13542 485696 13598 485752
rect 13542 477264 13598 477320
rect 13542 466656 13598 466712
rect 13542 458224 13598 458280
rect 13542 404232 13598 404288
rect 13542 395936 13598 395992
rect 13542 377712 13598 377768
rect 13542 369280 13598 369336
rect 13542 350240 13598 350296
rect 13542 341944 13598 342000
rect 13542 323720 13598 323776
rect 13542 315288 13598 315344
rect 13542 278024 13598 278080
rect 13542 269728 13598 269784
rect 13542 242256 13598 242312
rect 13542 233960 13598 234016
rect 13542 224032 13598 224088
rect 13542 215736 13598 215792
rect 13542 196696 13598 196752
rect 13542 188264 13598 188320
rect 13542 161744 13598 161800
rect 13542 142704 13598 142760
rect 13542 134272 13598 134328
rect 13542 116048 13598 116104
rect 13542 107752 13598 107808
rect 13542 88712 13598 88768
rect 13542 80280 13598 80336
rect 13542 53760 13598 53816
rect 13542 45328 13598 45384
rect 13450 33088 13506 33144
rect 12438 31048 12494 31104
rect 13542 29688 13598 29744
rect 13726 655968 13782 656024
rect 13726 647672 13782 647728
rect 13726 520648 13782 520704
rect 13726 512216 13782 512272
rect 13726 431704 13782 431760
rect 13726 423272 13782 423328
rect 13726 296248 13782 296304
rect 13726 287952 13782 288008
rect 13634 27648 13690 27704
rect 38658 674192 38714 674248
rect 38658 647672 38714 647728
rect 38658 620200 38714 620256
rect 38658 593680 38714 593736
rect 38658 566208 38714 566264
rect 38658 539688 38714 539744
rect 38658 512216 38714 512272
rect 38658 485696 38714 485752
rect 38658 458224 38714 458280
rect 38658 431704 38714 431760
rect 38658 404232 38714 404288
rect 38658 377712 38714 377768
rect 38658 350240 38714 350296
rect 38658 323720 38714 323776
rect 38658 296248 38714 296304
rect 38658 269728 38714 269784
rect 38658 242256 38714 242312
rect 38658 215736 38714 215792
rect 38658 188264 38714 188320
rect 38658 161744 38714 161800
rect 38658 134272 38714 134328
rect 38658 107752 38714 107808
rect 38658 80280 38714 80336
rect 38658 53760 38714 53816
rect 42706 674192 42762 674248
rect 42706 647672 42762 647728
rect 44638 634752 44694 634808
rect 42706 620200 42762 620256
rect 42706 602112 42762 602168
rect 42706 593680 42762 593736
rect 42706 566208 42762 566264
rect 42706 548120 42762 548176
rect 42706 539688 42762 539744
rect 42706 485696 42762 485752
rect 42706 477128 42762 477184
rect 64602 445576 64658 445632
rect 42706 431704 42762 431760
rect 42706 423136 42762 423192
rect 64602 391856 64658 391912
rect 42706 377712 42762 377768
rect 42706 323720 42762 323776
rect 42706 269728 42762 269784
rect 44638 256536 44694 256592
rect 42706 242256 42762 242312
rect 42706 224168 42762 224224
rect 42706 215736 42762 215792
rect 42706 188264 42762 188320
rect 42706 170040 42762 170096
rect 42706 161744 42762 161800
rect 42706 134272 42762 134328
rect 42706 116184 42762 116240
rect 42706 107752 42762 107808
rect 42706 53760 42762 53816
rect 42706 45192 42762 45248
rect 53378 37848 53434 37904
rect 61290 34312 61346 34368
rect 13726 26288 13782 26344
rect 13726 24112 13782 24168
rect 12438 22888 12494 22944
rect 12438 20848 12494 20904
rect 12438 19488 12494 19544
rect 12438 17448 12494 17504
rect 3422 6432 3478 6488
rect 45006 13640 45062 13696
rect 61106 13504 61162 13560
rect 64234 35128 64290 35184
rect 64418 31592 64474 31648
rect 64142 30232 64198 30288
rect 63498 26968 63554 27024
rect 63590 21392 63646 21448
rect 63498 18128 63554 18184
rect 64234 28328 64290 28384
rect 64234 24928 64290 24984
rect 64418 23568 64474 23624
rect 64326 16768 64382 16824
rect 66258 674192 66314 674248
rect 66258 665896 66314 665952
rect 66258 655968 66314 656024
rect 66258 647672 66314 647728
rect 66258 620200 66314 620256
rect 66258 611904 66314 611960
rect 66258 574640 66314 574696
rect 66258 566208 66314 566264
rect 66258 520648 66314 520704
rect 66258 512216 66314 512272
rect 66258 466656 66314 466712
rect 66258 458224 66314 458280
rect 66258 404232 66314 404288
rect 66258 395936 66314 395992
rect 66258 377712 66314 377768
rect 66258 369280 66314 369336
rect 66258 350240 66314 350296
rect 66258 341944 66314 342000
rect 66258 323720 66314 323776
rect 66258 315288 66314 315344
rect 66258 296248 66314 296304
rect 66258 287952 66314 288008
rect 66258 278024 66314 278080
rect 66258 269728 66314 269784
rect 66258 242256 66314 242312
rect 66258 233960 66314 234016
rect 66258 196696 66314 196752
rect 66258 188264 66314 188320
rect 66258 161744 66314 161800
rect 66258 142704 66314 142760
rect 66258 134272 66314 134328
rect 66258 88712 66314 88768
rect 66258 80280 66314 80336
rect 70306 673784 70362 673840
rect 70306 665896 70362 665952
rect 70306 655968 70362 656024
rect 70306 647672 70362 647728
rect 70306 620200 70362 620256
rect 70306 611904 70362 611960
rect 70306 601976 70362 602032
rect 70306 593680 70362 593736
rect 70306 574640 70362 574696
rect 70306 566208 70362 566264
rect 70306 547984 70362 548040
rect 70306 539688 70362 539744
rect 70306 520784 70362 520840
rect 70306 512216 70362 512272
rect 70306 485696 70362 485752
rect 70306 477264 70362 477320
rect 70306 466656 70362 466712
rect 70306 458224 70362 458280
rect 70306 431704 70362 431760
rect 70306 423272 70362 423328
rect 70306 404232 70362 404288
rect 70306 395936 70362 395992
rect 70306 377712 70362 377768
rect 70306 369280 70362 369336
rect 70306 350240 70362 350296
rect 70306 341808 70362 341864
rect 70306 323720 70362 323776
rect 70306 315288 70362 315344
rect 70306 296248 70362 296304
rect 70306 287952 70362 288008
rect 70306 278024 70362 278080
rect 70306 269728 70362 269784
rect 70306 242256 70362 242312
rect 70306 233960 70362 234016
rect 70306 224032 70362 224088
rect 70306 215736 70362 215792
rect 70306 196696 70362 196752
rect 70306 188264 70362 188320
rect 70306 161744 70362 161800
rect 70306 142704 70362 142760
rect 70306 134272 70362 134328
rect 70306 116048 70362 116104
rect 70306 108296 70362 108352
rect 70306 88712 70362 88768
rect 70306 80280 70362 80336
rect 70306 53216 70362 53272
rect 70306 45328 70362 45384
rect 70306 34856 70362 34912
rect 70306 26832 70362 26888
rect 95238 674192 95294 674248
rect 82266 657328 82322 657384
rect 95238 647672 95294 647728
rect 95238 620200 95294 620256
rect 95238 566208 95294 566264
rect 95238 520920 95294 520976
rect 95238 512216 95294 512272
rect 81990 468424 82046 468480
rect 95238 466792 95294 466848
rect 95238 458224 95294 458280
rect 81990 414432 82046 414488
rect 95238 404232 95294 404288
rect 95238 395800 95294 395856
rect 95238 377712 95294 377768
rect 95238 350240 95294 350296
rect 95238 341672 95294 341728
rect 95238 323720 95294 323776
rect 95238 296248 95294 296304
rect 95238 287816 95294 287872
rect 82266 279248 82322 279304
rect 95238 269728 95294 269784
rect 95238 242256 95294 242312
rect 95238 188264 95294 188320
rect 95238 170040 95294 170096
rect 95238 161744 95294 161800
rect 95238 134272 95294 134328
rect 95238 88848 95294 88904
rect 95238 80280 95294 80336
rect 97906 674192 97962 674248
rect 122838 674192 122894 674248
rect 126886 674192 126942 674248
rect 122838 665896 122894 665952
rect 126886 665896 126942 665952
rect 148690 662360 148746 662416
rect 150438 674192 150494 674248
rect 97906 647672 97962 647728
rect 128450 657328 128506 657384
rect 110602 634752 110658 634808
rect 122838 655968 122894 656024
rect 126886 655968 126942 656024
rect 122838 647672 122894 647728
rect 126886 647672 126942 647728
rect 150438 647672 150494 647728
rect 97906 620200 97962 620256
rect 122838 620200 122894 620256
rect 126886 620200 126942 620256
rect 122838 611904 122894 611960
rect 126886 611904 126942 611960
rect 148598 608504 148654 608560
rect 150438 620200 150494 620256
rect 97906 602112 97962 602168
rect 97906 593680 97962 593736
rect 128450 603336 128506 603392
rect 122838 601976 122894 602032
rect 126886 601976 126942 602032
rect 122838 593680 122894 593736
rect 126886 593680 126942 593736
rect 110602 580896 110658 580952
rect 97906 566208 97962 566264
rect 122838 574640 122894 574696
rect 126886 574640 126942 574696
rect 122838 566208 122894 566264
rect 126886 566208 126942 566264
rect 148598 554648 148654 554704
rect 150438 566208 150494 566264
rect 97906 548120 97962 548176
rect 97906 539688 97962 539744
rect 128450 549344 128506 549400
rect 122838 547984 122894 548040
rect 126886 547984 126942 548040
rect 122838 539688 122894 539744
rect 126886 539688 126942 539744
rect 110602 527040 110658 527096
rect 97906 520648 97962 520704
rect 97906 512216 97962 512272
rect 126886 520920 126942 520976
rect 122838 520784 122894 520840
rect 122838 512216 122894 512272
rect 126886 512216 126942 512272
rect 150438 520648 150494 520704
rect 150438 512216 150494 512272
rect 148598 500792 148654 500848
rect 97906 485696 97962 485752
rect 97906 477128 97962 477184
rect 128174 495216 128230 495272
rect 122838 485696 122894 485752
rect 126886 485696 126942 485752
rect 122838 477264 122894 477320
rect 126886 477264 126942 477320
rect 110602 473184 110658 473240
rect 97906 466792 97962 466848
rect 97906 458224 97962 458280
rect 122838 466656 122894 466712
rect 122838 458224 122894 458280
rect 150438 466792 150494 466848
rect 150438 458224 150494 458280
rect 148598 445576 148654 445632
rect 128450 441632 128506 441688
rect 97906 431704 97962 431760
rect 97906 423136 97962 423192
rect 110602 419464 110658 419520
rect 122838 431704 122894 431760
rect 126886 431704 126942 431760
rect 122838 423272 122894 423328
rect 126886 423272 126942 423328
rect 97906 404232 97962 404288
rect 97906 395800 97962 395856
rect 122838 404232 122894 404288
rect 122838 395936 122894 395992
rect 148598 391856 148654 391912
rect 150438 404232 150494 404288
rect 150438 395800 150494 395856
rect 97906 377712 97962 377768
rect 128450 387368 128506 387424
rect 122838 377712 122894 377768
rect 126886 377712 126942 377768
rect 122838 369280 122894 369336
rect 126886 369280 126942 369336
rect 110602 365608 110658 365664
rect 150438 377712 150494 377768
rect 97906 350240 97962 350296
rect 97906 341944 97962 342000
rect 122838 350240 122894 350296
rect 122838 341808 122894 341864
rect 148598 338000 148654 338056
rect 150438 350240 150494 350296
rect 150438 341944 150494 342000
rect 97906 323720 97962 323776
rect 128450 333240 128506 333296
rect 122838 323720 122894 323776
rect 126886 323720 126942 323776
rect 122838 315288 122894 315344
rect 126886 315288 126942 315344
rect 110602 311752 110658 311808
rect 150438 323720 150494 323776
rect 97906 296248 97962 296304
rect 97906 287816 97962 287872
rect 122838 296248 122894 296304
rect 126886 296248 126942 296304
rect 122838 287952 122894 288008
rect 126886 287952 126942 288008
rect 150438 296248 150494 296304
rect 150438 287816 150494 287872
rect 148598 284144 148654 284200
rect 97906 269728 97962 269784
rect 128450 279248 128506 279304
rect 122838 278024 122894 278080
rect 126886 278024 126942 278080
rect 122838 269728 122894 269784
rect 126886 269728 126942 269784
rect 110602 256536 110658 256592
rect 150438 269728 150494 269784
rect 97906 242256 97962 242312
rect 122838 242256 122894 242312
rect 126886 242256 126942 242312
rect 122838 233960 122894 234016
rect 126886 233960 126942 234016
rect 148598 230424 148654 230480
rect 150438 242256 150494 242312
rect 97906 224168 97962 224224
rect 97906 215736 97962 215792
rect 110602 202816 110658 202872
rect 128450 225256 128506 225312
rect 122838 224032 122894 224088
rect 126886 224032 126942 224088
rect 122838 215736 122894 215792
rect 126886 215736 126942 215792
rect 97906 188264 97962 188320
rect 122838 196696 122894 196752
rect 126886 196696 126942 196752
rect 122838 188264 122894 188320
rect 126886 188264 126942 188320
rect 150438 188264 150494 188320
rect 97906 170584 97962 170640
rect 97906 161744 97962 161800
rect 122838 161744 122894 161800
rect 97906 134272 97962 134328
rect 122838 142704 122894 142760
rect 126886 142704 126942 142760
rect 122838 134272 122894 134328
rect 126886 134272 126942 134328
rect 150438 134272 150494 134328
rect 97906 116184 97962 116240
rect 97906 107752 97962 107808
rect 126886 116320 126942 116376
rect 122838 116048 122894 116104
rect 122838 107752 122894 107808
rect 126886 107752 126942 107808
rect 97906 88848 97962 88904
rect 97906 80280 97962 80336
rect 122838 88712 122894 88768
rect 126886 88712 126942 88768
rect 122838 80280 122894 80336
rect 126886 80280 126942 80336
rect 150438 88848 150494 88904
rect 150438 80280 150494 80336
rect 97906 53760 97962 53816
rect 97906 45192 97962 45248
rect 122838 53760 122894 53816
rect 126886 53760 126942 53816
rect 122838 45328 122894 45384
rect 126886 45328 126942 45384
rect 97906 34720 97962 34776
rect 95238 26288 95294 26344
rect 97906 26288 97962 26344
rect 165986 684528 166042 684584
rect 154486 674192 154542 674248
rect 178038 674192 178094 674248
rect 182086 674192 182142 674248
rect 178038 665896 178094 665952
rect 182086 665896 182142 665952
rect 154486 647672 154542 647728
rect 156326 634752 156382 634808
rect 194782 657328 194838 657384
rect 207018 674192 207074 674248
rect 209686 674192 209742 674248
rect 222658 662360 222714 662416
rect 184202 655968 184258 656024
rect 184202 648216 184258 648272
rect 165986 630400 166042 630456
rect 154486 620200 154542 620256
rect 178038 620200 178094 620256
rect 182086 620200 182142 620256
rect 178038 611904 178094 611960
rect 182086 611904 182142 611960
rect 154486 602112 154542 602168
rect 154486 593680 154542 593736
rect 156326 580896 156382 580952
rect 182086 601976 182142 602032
rect 182086 593680 182142 593736
rect 194782 603336 194838 603392
rect 207018 647672 207074 647728
rect 209686 647672 209742 647728
rect 207018 620200 207074 620256
rect 209686 620200 209742 620256
rect 222658 608504 222714 608560
rect 165986 576408 166042 576464
rect 154486 566208 154542 566264
rect 178038 574640 178094 574696
rect 182086 574640 182142 574696
rect 178038 566208 178094 566264
rect 182086 566208 182142 566264
rect 154486 548120 154542 548176
rect 154486 539688 154542 539744
rect 156326 527040 156382 527096
rect 182086 547984 182142 548040
rect 182086 539688 182142 539744
rect 194782 549344 194838 549400
rect 207018 602112 207074 602168
rect 209686 602112 209742 602168
rect 207018 593680 207074 593736
rect 209686 593680 209742 593736
rect 207018 566208 207074 566264
rect 209686 566208 209742 566264
rect 222658 554648 222714 554704
rect 165986 522416 166042 522472
rect 155866 520784 155922 520840
rect 154486 512216 154542 512272
rect 182086 520648 182142 520704
rect 182086 512216 182142 512272
rect 154486 485696 154542 485752
rect 154486 477128 154542 477184
rect 182086 485696 182142 485752
rect 194782 495488 194838 495544
rect 207018 548120 207074 548176
rect 207018 539688 207074 539744
rect 207018 520784 207074 520840
rect 207018 512216 207074 512272
rect 222658 500792 222714 500848
rect 182086 477264 182142 477320
rect 156326 473184 156382 473240
rect 165986 468424 166042 468480
rect 154486 466792 154542 466848
rect 154486 458224 154542 458280
rect 178038 466656 178094 466712
rect 182086 466656 182142 466712
rect 178038 458224 178094 458280
rect 182086 458224 182142 458280
rect 194782 441632 194838 441688
rect 154486 431704 154542 431760
rect 154486 423136 154542 423192
rect 156326 419464 156382 419520
rect 182086 431704 182142 431760
rect 182086 423272 182142 423328
rect 207018 485696 207074 485752
rect 207018 477128 207074 477184
rect 207018 466792 207074 466848
rect 207018 458224 207074 458280
rect 222658 445576 222714 445632
rect 165986 414432 166042 414488
rect 154486 404232 154542 404288
rect 154486 395800 154542 395856
rect 178038 404232 178094 404288
rect 182086 404232 182142 404288
rect 178038 395936 178094 395992
rect 182086 395936 182142 395992
rect 154486 377712 154542 377768
rect 156326 365608 156382 365664
rect 182086 377712 182142 377768
rect 194782 387368 194838 387424
rect 207018 431704 207074 431760
rect 209686 431704 209742 431760
rect 207018 423136 207074 423192
rect 209686 423136 209742 423192
rect 207018 404232 207074 404288
rect 207018 395800 207074 395856
rect 222658 391856 222714 391912
rect 182086 369280 182142 369336
rect 165986 360440 166042 360496
rect 154486 350240 154542 350296
rect 154486 341808 154542 341864
rect 178038 350240 178094 350296
rect 182086 350240 182142 350296
rect 182086 341944 182142 342000
rect 178038 341672 178094 341728
rect 154486 323720 154542 323776
rect 156326 311752 156382 311808
rect 182086 323720 182142 323776
rect 182086 315288 182142 315344
rect 207018 377712 207074 377768
rect 209686 377712 209742 377768
rect 207018 350240 207074 350296
rect 207018 341808 207074 341864
rect 222658 338000 222714 338056
rect 194782 333240 194838 333296
rect 165986 306448 166042 306504
rect 154486 296248 154542 296304
rect 154486 287816 154542 287872
rect 182086 296248 182142 296304
rect 182086 287952 182142 288008
rect 154486 269728 154542 269784
rect 182086 278024 182142 278080
rect 182086 269728 182142 269784
rect 207018 323720 207074 323776
rect 209686 323720 209742 323776
rect 207018 296248 207074 296304
rect 207018 287816 207074 287872
rect 222658 284144 222714 284200
rect 194782 279248 194838 279304
rect 156326 256536 156382 256592
rect 165986 252592 166042 252648
rect 154486 242256 154542 242312
rect 178038 242256 178094 242312
rect 182086 242256 182142 242312
rect 178038 233960 178094 234016
rect 182086 233960 182142 234016
rect 154486 224168 154542 224224
rect 154486 215736 154542 215792
rect 156326 202816 156382 202872
rect 182086 224032 182142 224088
rect 182086 215736 182142 215792
rect 207018 269728 207074 269784
rect 209686 269728 209742 269784
rect 207018 242256 207074 242312
rect 209686 242256 209742 242312
rect 222658 230424 222714 230480
rect 194782 225256 194838 225312
rect 154486 188264 154542 188320
rect 178038 196696 178094 196752
rect 182086 196696 182142 196752
rect 178038 188264 178094 188320
rect 182086 188264 182142 188320
rect 154486 170176 154542 170232
rect 154486 161744 154542 161800
rect 178038 170312 178094 170368
rect 178038 161744 178094 161800
rect 207018 224168 207074 224224
rect 209686 224168 209742 224224
rect 207018 215736 207074 215792
rect 209686 215736 209742 215792
rect 207018 188264 207074 188320
rect 209686 188264 209742 188320
rect 222658 176568 222714 176624
rect 182086 170040 182142 170096
rect 182086 161744 182142 161800
rect 154486 134272 154542 134328
rect 178038 142704 178094 142760
rect 178038 134272 178094 134328
rect 182086 134272 182142 134328
rect 154486 116048 154542 116104
rect 154486 107752 154542 107808
rect 156326 95104 156382 95160
rect 182086 116320 182142 116376
rect 182086 107752 182142 107808
rect 207018 170176 207074 170232
rect 207018 161744 207074 161800
rect 209686 161744 209742 161800
rect 209686 142704 209742 142760
rect 207018 134272 207074 134328
rect 209686 134272 209742 134328
rect 194782 117272 194838 117328
rect 154486 88848 154542 88904
rect 154486 80280 154542 80336
rect 182086 88712 182142 88768
rect 182086 80280 182142 80336
rect 154486 53760 154542 53816
rect 154486 45192 154542 45248
rect 182086 53760 182142 53816
rect 182086 45328 182142 45384
rect 209686 116456 209742 116512
rect 207018 116048 207074 116104
rect 207018 107752 207074 107808
rect 209686 107752 209742 107808
rect 207018 88848 207074 88904
rect 207018 80280 207074 80336
rect 209686 80280 209742 80336
rect 207018 53760 207074 53816
rect 209686 53760 209742 53816
rect 207018 45192 207074 45248
rect 209686 45192 209742 45248
rect 122838 34856 122894 34912
rect 122838 26288 122894 26344
rect 150438 34720 150494 34776
rect 154486 34720 154542 34776
rect 150438 26288 150494 26344
rect 154486 26288 154542 26344
rect 178038 34856 178094 34912
rect 178038 26288 178094 26344
rect 182086 34856 182142 34912
rect 182086 26288 182142 26344
rect 207018 34720 207074 34776
rect 207018 26288 207074 26344
rect 232594 13368 232650 13424
rect 260378 684528 260434 684584
rect 234710 674192 234766 674248
rect 238666 674192 238722 674248
rect 234710 665896 234766 665952
rect 238666 665896 238722 665952
rect 262218 674192 262274 674248
rect 266266 674192 266322 674248
rect 291198 674192 291254 674248
rect 293866 674192 293922 674248
rect 291198 665896 291254 665952
rect 293866 665896 293922 665952
rect 361946 684528 362002 684584
rect 318798 674192 318854 674248
rect 322846 674192 322902 674248
rect 346398 674192 346454 674248
rect 350446 674192 350502 674248
rect 346398 665896 346454 665952
rect 350446 665896 350502 665952
rect 344926 662360 344982 662416
rect 375378 674192 375434 674248
rect 378046 674192 378102 674248
rect 234710 655968 234766 656024
rect 238666 655968 238722 656024
rect 234710 647672 234766 647728
rect 238666 647672 238722 647728
rect 240322 634752 240378 634808
rect 262218 647672 262274 647728
rect 266266 647672 266322 647728
rect 278226 657328 278282 657384
rect 291198 655968 291254 656024
rect 293866 655968 293922 656024
rect 291198 647672 291254 647728
rect 293866 647672 293922 647728
rect 318798 647672 318854 647728
rect 322846 647672 322902 647728
rect 346398 655968 346454 656024
rect 350446 655968 350502 656024
rect 346398 647672 346454 647728
rect 350446 647672 350502 647728
rect 352654 634752 352710 634808
rect 375378 647672 375434 647728
rect 378046 647672 378102 647728
rect 260378 630400 260434 630456
rect 234710 620200 234766 620256
rect 238666 620200 238722 620256
rect 234710 611904 234766 611960
rect 238666 611904 238722 611960
rect 262218 620200 262274 620256
rect 266266 620200 266322 620256
rect 291198 620200 291254 620256
rect 293866 620200 293922 620256
rect 291198 611904 291254 611960
rect 293866 611904 293922 611960
rect 361946 630400 362002 630456
rect 318798 620200 318854 620256
rect 322846 620200 322902 620256
rect 346398 620200 346454 620256
rect 350446 620200 350502 620256
rect 346398 611904 346454 611960
rect 350446 611904 350502 611960
rect 344650 608504 344706 608560
rect 375378 620200 375434 620256
rect 378046 620200 378102 620256
rect 238666 602248 238722 602304
rect 234710 601976 234766 602032
rect 234710 593680 234766 593736
rect 238666 593680 238722 593736
rect 266266 601976 266322 602032
rect 266266 593680 266322 593736
rect 293866 602112 293922 602168
rect 293866 593680 293922 593736
rect 318798 601976 318854 602032
rect 322846 601976 322902 602032
rect 318798 593680 318854 593736
rect 322846 593680 322902 593736
rect 350446 602112 350502 602168
rect 350446 593680 350502 593736
rect 352654 580896 352710 580952
rect 378046 601976 378102 602032
rect 378046 593680 378102 593736
rect 260378 576408 260434 576464
rect 234710 574640 234766 574696
rect 238666 574640 238722 574696
rect 234710 566208 234766 566264
rect 238666 566208 238722 566264
rect 262218 566208 262274 566264
rect 266266 566208 266322 566264
rect 361946 576408 362002 576464
rect 291198 574640 291254 574696
rect 293866 574640 293922 574696
rect 291198 566208 291254 566264
rect 293866 566208 293922 566264
rect 318798 566208 318854 566264
rect 322846 566208 322902 566264
rect 346398 574640 346454 574696
rect 350446 574640 350502 574696
rect 346398 566208 346454 566264
rect 350446 566208 350502 566264
rect 375378 566208 375434 566264
rect 378046 566208 378102 566264
rect 344650 554648 344706 554704
rect 238666 548256 238722 548312
rect 234710 547984 234766 548040
rect 234710 539688 234766 539744
rect 238666 539688 238722 539744
rect 262218 548120 262274 548176
rect 266266 547984 266322 548040
rect 262218 539688 262274 539744
rect 266266 539688 266322 539744
rect 322846 548256 322902 548312
rect 318798 547984 318854 548040
rect 318798 539688 318854 539744
rect 322846 539688 322902 539744
rect 346398 548120 346454 548176
rect 350446 547984 350502 548040
rect 346398 539688 346454 539744
rect 350446 539688 350502 539744
rect 352654 527040 352710 527096
rect 378046 548120 378102 548176
rect 378046 539688 378102 539744
rect 260378 522416 260434 522472
rect 238666 520920 238722 520976
rect 234710 520648 234766 520704
rect 234710 512216 234766 512272
rect 238666 512216 238722 512272
rect 262218 520784 262274 520840
rect 266266 520648 266322 520704
rect 262218 512216 262274 512272
rect 266266 512216 266322 512272
rect 361946 522416 362002 522472
rect 317050 520648 317106 520704
rect 322846 520648 322902 520704
rect 317050 512760 317106 512816
rect 322846 512216 322902 512272
rect 346398 520784 346454 520840
rect 350446 520784 350502 520840
rect 346398 512216 346454 512272
rect 350446 512216 350502 512272
rect 378046 520648 378102 520704
rect 378046 512216 378102 512272
rect 344650 500792 344706 500848
rect 234710 485696 234766 485752
rect 238666 485696 238722 485752
rect 234710 477264 234766 477320
rect 238666 476992 238722 477048
rect 262218 485696 262274 485752
rect 266266 485696 266322 485752
rect 266266 477264 266322 477320
rect 262218 477128 262274 477184
rect 318798 485696 318854 485752
rect 322846 485696 322902 485752
rect 318798 477264 318854 477320
rect 322846 476992 322902 477048
rect 346398 485696 346454 485752
rect 350446 485696 350502 485752
rect 350446 477264 350502 477320
rect 346398 477128 346454 477184
rect 378046 485696 378102 485752
rect 378046 477128 378102 477184
rect 352654 473184 352710 473240
rect 260378 468424 260434 468480
rect 234710 466656 234766 466712
rect 234710 458224 234766 458280
rect 262218 466928 262274 466984
rect 266266 466656 266322 466712
rect 262218 458224 262274 458280
rect 266266 458224 266322 458280
rect 361946 468424 362002 468480
rect 291198 466792 291254 466848
rect 291198 458224 291254 458280
rect 318798 466656 318854 466712
rect 318798 458224 318854 458280
rect 346398 466792 346454 466848
rect 350446 466792 350502 466848
rect 346398 458224 346454 458280
rect 350446 458224 350502 458280
rect 375378 466656 375434 466712
rect 378046 466656 378102 466712
rect 375378 458224 375434 458280
rect 378046 458224 378102 458280
rect 344650 445576 344706 445632
rect 234710 431704 234766 431760
rect 238666 431704 238722 431760
rect 234710 423272 234766 423328
rect 238666 423000 238722 423056
rect 266266 431704 266322 431760
rect 266266 423272 266322 423328
rect 293866 431704 293922 431760
rect 293866 423136 293922 423192
rect 318798 431704 318854 431760
rect 322846 431704 322902 431760
rect 318798 423272 318854 423328
rect 322846 423272 322902 423328
rect 350446 431704 350502 431760
rect 350446 423136 350502 423192
rect 352654 419464 352710 419520
rect 378046 431704 378102 431760
rect 378046 423272 378102 423328
rect 260378 414432 260434 414488
rect 234710 404232 234766 404288
rect 234710 395936 234766 395992
rect 262218 404232 262274 404288
rect 266266 404232 266322 404288
rect 266266 395936 266322 395992
rect 262218 395664 262274 395720
rect 291198 404232 291254 404288
rect 291198 395800 291254 395856
rect 361946 414432 362002 414488
rect 318798 404232 318854 404288
rect 318798 395936 318854 395992
rect 344650 391856 344706 391912
rect 346398 404232 346454 404288
rect 350446 404232 350502 404288
rect 350446 395936 350502 395992
rect 346398 395664 346454 395720
rect 375378 404232 375434 404288
rect 378046 404232 378102 404288
rect 375378 395800 375434 395856
rect 378046 395800 378102 395856
rect 234710 377712 234766 377768
rect 238666 377712 238722 377768
rect 234710 369280 234766 369336
rect 238666 369280 238722 369336
rect 262218 377712 262274 377768
rect 266266 377712 266322 377768
rect 291198 377712 291254 377768
rect 293866 377712 293922 377768
rect 291198 369280 291254 369336
rect 293866 369280 293922 369336
rect 318798 377712 318854 377768
rect 322846 377712 322902 377768
rect 346398 377712 346454 377768
rect 350446 377712 350502 377768
rect 346398 369280 346454 369336
rect 350446 369280 350502 369336
rect 352654 365608 352710 365664
rect 375378 377712 375434 377768
rect 378046 377712 378102 377768
rect 260378 360440 260434 360496
rect 234710 350240 234766 350296
rect 234710 341944 234766 342000
rect 262218 350240 262274 350296
rect 266266 350240 266322 350296
rect 266266 341944 266322 342000
rect 262218 341672 262274 341728
rect 291198 350240 291254 350296
rect 291198 341808 291254 341864
rect 361946 360440 362002 360496
rect 318798 350240 318854 350296
rect 318798 341944 318854 342000
rect 346398 350240 346454 350296
rect 350446 350240 350502 350296
rect 350446 341944 350502 342000
rect 346398 341672 346454 341728
rect 344650 338000 344706 338056
rect 375378 350240 375434 350296
rect 378046 350240 378102 350296
rect 375378 341808 375434 341864
rect 378046 341808 378102 341864
rect 234710 323720 234766 323776
rect 238666 323720 238722 323776
rect 234710 315288 234766 315344
rect 238666 315288 238722 315344
rect 262218 323720 262274 323776
rect 266266 323720 266322 323776
rect 291198 323720 291254 323776
rect 293866 323720 293922 323776
rect 291198 315288 291254 315344
rect 293866 315288 293922 315344
rect 318798 323720 318854 323776
rect 322846 323720 322902 323776
rect 346398 323720 346454 323776
rect 350446 323720 350502 323776
rect 346398 315288 346454 315344
rect 350446 315288 350502 315344
rect 352654 311752 352710 311808
rect 375378 323720 375434 323776
rect 378046 323720 378102 323776
rect 260378 306448 260434 306504
rect 234710 296248 234766 296304
rect 238666 296248 238722 296304
rect 234710 287952 234766 288008
rect 238666 287680 238722 287736
rect 262218 296248 262274 296304
rect 266266 296248 266322 296304
rect 266266 287952 266322 288008
rect 262218 287816 262274 287872
rect 361946 306448 362002 306504
rect 318798 296248 318854 296304
rect 322846 296248 322902 296304
rect 318798 287952 318854 288008
rect 322846 287952 322902 288008
rect 346398 296248 346454 296304
rect 350446 296248 350502 296304
rect 346398 287816 346454 287872
rect 350446 287816 350502 287872
rect 378046 296248 378102 296304
rect 378046 287952 378102 288008
rect 344650 284144 344706 284200
rect 234710 278024 234766 278080
rect 238666 278024 238722 278080
rect 234710 269728 234766 269784
rect 238666 269728 238722 269784
rect 262218 269728 262274 269784
rect 266266 269728 266322 269784
rect 278226 279792 278282 279848
rect 291198 278024 291254 278080
rect 293866 278024 293922 278080
rect 291198 269728 291254 269784
rect 293866 269728 293922 269784
rect 318798 269728 318854 269784
rect 322846 269728 322902 269784
rect 240322 256536 240378 256592
rect 346398 278024 346454 278080
rect 350446 278024 350502 278080
rect 346398 269728 346454 269784
rect 350446 269728 350502 269784
rect 375378 269728 375434 269784
rect 378046 269728 378102 269784
rect 352654 256536 352710 256592
rect 260378 252592 260434 252648
rect 234710 242256 234766 242312
rect 238666 242256 238722 242312
rect 234710 233960 234766 234016
rect 238666 233960 238722 234016
rect 262218 242256 262274 242312
rect 266266 242256 266322 242312
rect 291198 242256 291254 242312
rect 293866 242256 293922 242312
rect 291198 233960 291254 234016
rect 293866 233960 293922 234016
rect 361946 252592 362002 252648
rect 318798 242256 318854 242312
rect 322846 242256 322902 242312
rect 346398 242256 346454 242312
rect 350446 242256 350502 242312
rect 346398 233960 346454 234016
rect 350446 233960 350502 234016
rect 344650 230424 344706 230480
rect 375378 242256 375434 242312
rect 378046 242256 378102 242312
rect 238666 224304 238722 224360
rect 234710 224032 234766 224088
rect 234710 215736 234766 215792
rect 238666 215736 238722 215792
rect 266266 224032 266322 224088
rect 266266 215736 266322 215792
rect 293866 215736 293922 215792
rect 318798 224032 318854 224088
rect 318798 215736 318854 215792
rect 322846 215736 322902 215792
rect 346398 215736 346454 215792
rect 350446 224032 350502 224088
rect 350446 215736 350502 215792
rect 378046 224168 378102 224224
rect 375378 215736 375434 215792
rect 378046 215736 378102 215792
rect 260378 198464 260434 198520
rect 234710 196696 234766 196752
rect 238666 196696 238722 196752
rect 234710 188264 234766 188320
rect 238666 188264 238722 188320
rect 262218 188264 262274 188320
rect 266266 188264 266322 188320
rect 291198 196696 291254 196752
rect 293866 196696 293922 196752
rect 291198 188264 291254 188320
rect 293866 188264 293922 188320
rect 361946 198464 362002 198520
rect 318798 188264 318854 188320
rect 322846 188264 322902 188320
rect 346398 196696 346454 196752
rect 350446 196696 350502 196752
rect 346398 188264 346454 188320
rect 350446 188264 350502 188320
rect 375378 188264 375434 188320
rect 378046 188264 378102 188320
rect 344650 176568 344706 176624
rect 234710 170040 234766 170096
rect 234710 161744 234766 161800
rect 238666 161744 238722 161800
rect 262218 161744 262274 161800
rect 266266 170040 266322 170096
rect 266266 161744 266322 161800
rect 293866 170176 293922 170232
rect 291198 161744 291254 161800
rect 293866 161744 293922 161800
rect 322846 170312 322902 170368
rect 318798 170040 318854 170096
rect 318798 161744 318854 161800
rect 322846 161744 322902 161800
rect 350446 170040 350502 170096
rect 350446 161744 350502 161800
rect 378046 170176 378102 170232
rect 378046 161744 378102 161800
rect 234710 134272 234766 134328
rect 238666 134272 238722 134328
rect 262218 142704 262274 142760
rect 262218 134272 262274 134328
rect 266266 142704 266322 142760
rect 266266 134272 266322 134328
rect 291198 134272 291254 134328
rect 293866 134272 293922 134328
rect 361946 144472 362002 144528
rect 318798 142704 318854 142760
rect 322846 142704 322902 142760
rect 318798 134272 318854 134328
rect 322846 134272 322902 134328
rect 346398 134272 346454 134328
rect 350446 134272 350502 134328
rect 375378 142704 375434 142760
rect 378046 142704 378102 142760
rect 375378 134272 375434 134328
rect 378046 134272 378102 134328
rect 344650 122712 344706 122768
rect 234710 116320 234766 116376
rect 234710 107752 234766 107808
rect 238666 107752 238722 107808
rect 266266 116048 266322 116104
rect 266266 107752 266322 107808
rect 291198 107752 291254 107808
rect 293866 107752 293922 107808
rect 318798 116048 318854 116104
rect 324226 117272 324282 117328
rect 318798 107752 318854 107808
rect 322846 107752 322902 107808
rect 306930 95104 306986 95160
rect 346398 107752 346454 107808
rect 350446 116048 350502 116104
rect 350446 107752 350502 107808
rect 378046 116184 378102 116240
rect 375378 107752 375434 107808
rect 378046 107752 378102 107808
rect 238666 88848 238722 88904
rect 234710 88712 234766 88768
rect 234710 80280 234766 80336
rect 238666 80280 238722 80336
rect 266266 88712 266322 88768
rect 262218 80280 262274 80336
rect 266266 80280 266322 80336
rect 322846 88984 322902 89040
rect 318798 88712 318854 88768
rect 318798 80280 318854 80336
rect 322846 80280 322902 80336
rect 346398 88848 346454 88904
rect 350446 88712 350502 88768
rect 346398 80280 346454 80336
rect 350446 80280 350502 80336
rect 378046 88848 378102 88904
rect 378046 80280 378102 80336
rect 234710 53760 234766 53816
rect 238666 53760 238722 53816
rect 234710 45328 234766 45384
rect 238666 45056 238722 45112
rect 266266 53760 266322 53816
rect 266266 45328 266322 45384
rect 293866 53760 293922 53816
rect 293866 45192 293922 45248
rect 318798 53760 318854 53816
rect 322846 53760 322902 53816
rect 318798 45328 318854 45384
rect 322846 45056 322902 45112
rect 350446 53760 350502 53816
rect 350446 45328 350502 45384
rect 378046 53760 378102 53816
rect 378046 45192 378102 45248
rect 250074 36488 250130 36544
rect 234618 34856 234674 34912
rect 234618 26288 234674 26344
rect 262218 34720 262274 34776
rect 266266 34720 266322 34776
rect 262218 26288 262274 26344
rect 266266 26288 266322 26344
rect 291198 34856 291254 34912
rect 291198 26288 291254 26344
rect 318798 34720 318854 34776
rect 318798 26288 318854 26344
rect 346398 34992 346454 35048
rect 350446 34720 350502 34776
rect 346398 26288 346454 26344
rect 350446 26288 350502 26344
rect 375378 34856 375434 34912
rect 378046 34856 378102 34912
rect 375378 26288 375434 26344
rect 378046 26288 378102 26344
rect 402978 674192 403034 674248
rect 405646 674192 405702 674248
rect 402978 665896 403034 665952
rect 405646 665896 405702 665952
rect 428646 662360 428702 662416
rect 390834 657328 390890 657384
rect 402978 655968 403034 656024
rect 402978 647672 403034 647728
rect 408130 655968 408186 656024
rect 408130 648216 408186 648272
rect 402978 620200 403034 620256
rect 405646 620200 405702 620256
rect 402978 611904 403034 611960
rect 405646 611904 405702 611960
rect 428646 608504 428702 608560
rect 390834 603336 390890 603392
rect 402978 602112 403034 602168
rect 405646 602112 405702 602168
rect 402978 593680 403034 593736
rect 405646 593680 405702 593736
rect 402978 574640 403034 574696
rect 405646 574640 405702 574696
rect 402978 566208 403034 566264
rect 405646 566208 405702 566264
rect 428646 554648 428702 554704
rect 390834 549344 390890 549400
rect 402978 547984 403034 548040
rect 402978 539688 403034 539744
rect 402978 520784 403034 520840
rect 402978 512216 403034 512272
rect 428646 500792 428702 500848
rect 390834 495488 390890 495544
rect 402978 485696 403034 485752
rect 402978 477264 403034 477320
rect 402978 466792 403034 466848
rect 402978 458224 403034 458280
rect 418342 445576 418398 445632
rect 428646 445440 428702 445496
rect 390834 441632 390890 441688
rect 402978 431704 403034 431760
rect 405646 431704 405702 431760
rect 402978 423136 403034 423192
rect 405646 423136 405702 423192
rect 402978 404232 403034 404288
rect 402978 395936 403034 395992
rect 418342 391856 418398 391912
rect 428646 391720 428702 391776
rect 390834 387368 390890 387424
rect 402978 377712 403034 377768
rect 405646 377712 405702 377768
rect 402978 369280 403034 369336
rect 405646 369280 405702 369336
rect 402978 350240 403034 350296
rect 402978 341944 403034 342000
rect 428646 338000 428702 338056
rect 390834 333240 390890 333296
rect 402978 323720 403034 323776
rect 405646 323720 405702 323776
rect 402978 315288 403034 315344
rect 405646 315288 405702 315344
rect 402978 296248 403034 296304
rect 402978 287816 403034 287872
rect 428646 284144 428702 284200
rect 390834 279248 390890 279304
rect 402978 278024 403034 278080
rect 405646 278024 405702 278080
rect 402978 269728 403034 269784
rect 405646 269728 405702 269784
rect 402978 242256 403034 242312
rect 405646 242256 405702 242312
rect 402978 233960 403034 234016
rect 405646 233960 405702 234016
rect 428646 230424 428702 230480
rect 402978 224032 403034 224088
rect 402978 215736 403034 215792
rect 405646 215736 405702 215792
rect 402978 196696 403034 196752
rect 405646 196696 405702 196752
rect 402978 188264 403034 188320
rect 405646 188264 405702 188320
rect 428646 176568 428702 176624
rect 402978 170040 403034 170096
rect 402978 161744 403034 161800
rect 402978 134272 403034 134328
rect 405646 134272 405702 134328
rect 428646 122712 428702 122768
rect 402978 116048 403034 116104
rect 402978 107752 403034 107808
rect 402978 88712 403034 88768
rect 402978 80280 403034 80336
rect 405646 80280 405702 80336
rect 402978 53760 403034 53816
rect 405646 53760 405702 53816
rect 402978 45328 403034 45384
rect 405646 45328 405702 45384
rect 402978 34720 403034 34776
rect 402978 26288 403034 26344
rect 446034 684528 446090 684584
rect 430578 674192 430634 674248
rect 434626 674192 434682 674248
rect 462226 674192 462282 674248
rect 458178 673784 458234 673840
rect 458178 665896 458234 665952
rect 462226 665896 462282 665952
rect 487158 674192 487214 674248
rect 489826 674192 489882 674248
rect 514758 674192 514814 674248
rect 514758 665896 514814 665952
rect 430578 647672 430634 647728
rect 434626 647672 434682 647728
rect 436650 634752 436706 634808
rect 474278 657328 474334 657384
rect 464158 655968 464214 656024
rect 464158 648216 464214 648272
rect 487158 647672 487214 647728
rect 489826 647672 489882 647728
rect 502614 634752 502670 634808
rect 514758 655968 514814 656024
rect 514758 647672 514814 647728
rect 446034 630400 446090 630456
rect 430578 620200 430634 620256
rect 434626 620200 434682 620256
rect 458178 620200 458234 620256
rect 462226 620200 462282 620256
rect 458178 611904 458234 611960
rect 462226 611904 462282 611960
rect 487158 620200 487214 620256
rect 489826 620200 489882 620256
rect 514758 620200 514814 620256
rect 514758 611904 514814 611960
rect 434626 602248 434682 602304
rect 430578 601976 430634 602032
rect 430578 593680 430634 593736
rect 434626 593680 434682 593736
rect 462226 601976 462282 602032
rect 462226 593680 462282 593736
rect 514758 601976 514814 602032
rect 514758 593680 514814 593736
rect 446034 576408 446090 576464
rect 430578 566208 430634 566264
rect 434626 566208 434682 566264
rect 458178 574640 458234 574696
rect 462226 574640 462282 574696
rect 458178 566208 458234 566264
rect 462226 566208 462282 566264
rect 487158 566208 487214 566264
rect 489826 566208 489882 566264
rect 514758 574640 514814 574696
rect 514758 566208 514814 566264
rect 430578 548120 430634 548176
rect 434626 548120 434682 548176
rect 430578 539688 430634 539744
rect 434626 539688 434682 539744
rect 458178 547984 458234 548040
rect 462226 547984 462282 548040
rect 458178 539688 458234 539744
rect 462226 539688 462282 539744
rect 489826 548120 489882 548176
rect 489826 539688 489882 539744
rect 514758 547984 514814 548040
rect 514758 539688 514814 539744
rect 446034 522416 446090 522472
rect 434626 520920 434682 520976
rect 430578 520648 430634 520704
rect 430578 512216 430634 512272
rect 434626 512216 434682 512272
rect 458178 520784 458234 520840
rect 463882 520648 463938 520704
rect 458178 512216 458234 512272
rect 462226 512216 462282 512272
rect 514758 520648 514814 520704
rect 514758 512216 514814 512272
rect 430578 485696 430634 485752
rect 434626 485696 434682 485752
rect 430578 477128 430634 477184
rect 434626 477128 434682 477184
rect 458178 485696 458234 485752
rect 462226 485696 462282 485752
rect 458178 477264 458234 477320
rect 462226 477264 462282 477320
rect 489826 485696 489882 485752
rect 489826 477128 489882 477184
rect 514758 485696 514814 485752
rect 514758 477264 514814 477320
rect 446034 468424 446090 468480
rect 456338 468424 456394 468480
rect 430578 466656 430634 466712
rect 430578 458224 430634 458280
rect 458178 466928 458234 466984
rect 462226 466656 462282 466712
rect 458178 458224 458234 458280
rect 462226 458224 462282 458280
rect 487158 466792 487214 466848
rect 487158 458224 487214 458280
rect 514758 466656 514814 466712
rect 514758 458224 514814 458280
rect 430578 431704 430634 431760
rect 434626 431704 434682 431760
rect 430578 423272 430634 423328
rect 434626 423000 434682 423056
rect 462226 431704 462282 431760
rect 462226 423272 462282 423328
rect 514758 431704 514814 431760
rect 514758 423272 514814 423328
rect 446034 414432 446090 414488
rect 456338 414432 456394 414488
rect 430578 404232 430634 404288
rect 430578 395800 430634 395856
rect 458178 404232 458234 404288
rect 462226 404232 462282 404288
rect 458178 395936 458234 395992
rect 462226 395936 462282 395992
rect 487158 404232 487214 404288
rect 487158 395800 487214 395856
rect 514758 404232 514814 404288
rect 514758 395936 514814 395992
rect 430578 377712 430634 377768
rect 434626 377712 434682 377768
rect 462226 377712 462282 377768
rect 462226 369280 462282 369336
rect 487158 377712 487214 377768
rect 489826 377712 489882 377768
rect 514758 377712 514814 377768
rect 514758 369280 514814 369336
rect 446034 360440 446090 360496
rect 430578 350240 430634 350296
rect 430578 341808 430634 341864
rect 458178 350240 458234 350296
rect 462226 350240 462282 350296
rect 458178 341944 458234 342000
rect 462226 341944 462282 342000
rect 487158 350240 487214 350296
rect 487158 341808 487214 341864
rect 514758 350240 514814 350296
rect 514758 341944 514814 342000
rect 430578 323720 430634 323776
rect 434626 323720 434682 323776
rect 462226 323720 462282 323776
rect 462226 315288 462282 315344
rect 487158 323720 487214 323776
rect 489826 323720 489882 323776
rect 514758 323720 514814 323776
rect 514758 315288 514814 315344
rect 446034 306448 446090 306504
rect 430578 296248 430634 296304
rect 434626 296248 434682 296304
rect 430578 287952 430634 288008
rect 434626 287680 434682 287736
rect 458178 296248 458234 296304
rect 462226 296248 462282 296304
rect 462226 287952 462282 288008
rect 458178 287816 458234 287872
rect 514758 296248 514814 296304
rect 514758 287952 514814 288008
rect 430578 269728 430634 269784
rect 434626 269728 434682 269784
rect 462226 278024 462282 278080
rect 462226 269728 462282 269784
rect 474278 279248 474334 279304
rect 487158 269728 487214 269784
rect 489826 269728 489882 269784
rect 436650 256536 436706 256592
rect 514758 278024 514814 278080
rect 514758 269728 514814 269784
rect 502614 256536 502670 256592
rect 446034 252592 446090 252648
rect 430578 242256 430634 242312
rect 434626 242256 434682 242312
rect 458178 242256 458234 242312
rect 462226 242256 462282 242312
rect 458178 233960 458234 234016
rect 462226 233960 462282 234016
rect 487158 242256 487214 242312
rect 489826 242256 489882 242312
rect 514758 242256 514814 242312
rect 514758 233960 514814 234016
rect 430578 224168 430634 224224
rect 430578 215736 430634 215792
rect 434626 215736 434682 215792
rect 458178 215736 458234 215792
rect 462226 224032 462282 224088
rect 462226 215736 462282 215792
rect 487158 215736 487214 215792
rect 514758 224032 514814 224088
rect 514758 215736 514814 215792
rect 446034 198464 446090 198520
rect 430578 188264 430634 188320
rect 434626 188264 434682 188320
rect 458178 196696 458234 196752
rect 462226 196696 462282 196752
rect 458178 188264 458234 188320
rect 462226 188264 462282 188320
rect 487158 188264 487214 188320
rect 489826 188264 489882 188320
rect 514758 196696 514814 196752
rect 514758 188264 514814 188320
rect 430578 170176 430634 170232
rect 430578 161744 430634 161800
rect 434626 161744 434682 161800
rect 458178 170040 458234 170096
rect 458178 161744 458234 161800
rect 462226 161744 462282 161800
rect 489826 170176 489882 170232
rect 487158 161744 487214 161800
rect 489826 161744 489882 161800
rect 514758 161744 514814 161800
rect 446034 144472 446090 144528
rect 430578 142704 430634 142760
rect 434626 142704 434682 142760
rect 430578 134272 430634 134328
rect 434626 134272 434682 134328
rect 458178 134272 458234 134328
rect 462226 134272 462282 134328
rect 487158 142704 487214 142760
rect 489826 142704 489882 142760
rect 487158 134272 487214 134328
rect 489826 134272 489882 134328
rect 514758 134272 514814 134328
rect 430578 116184 430634 116240
rect 430578 107752 430634 107808
rect 434626 107752 434682 107808
rect 458178 116048 458234 116104
rect 458178 108296 458234 108352
rect 462226 116048 462282 116104
rect 462226 107752 462282 107808
rect 489826 116184 489882 116240
rect 487158 107752 487214 107808
rect 489826 107752 489882 107808
rect 514758 116048 514814 116104
rect 514758 107752 514814 107808
rect 430578 88848 430634 88904
rect 434626 88848 434682 88904
rect 430578 80280 430634 80336
rect 434626 80280 434682 80336
rect 458178 80280 458234 80336
rect 462226 88712 462282 88768
rect 462226 80280 462282 80336
rect 489826 80280 489882 80336
rect 514758 88712 514814 88768
rect 514758 80280 514814 80336
rect 430578 53760 430634 53816
rect 434626 53760 434682 53816
rect 430578 45192 430634 45248
rect 434626 45192 434682 45248
rect 462226 53760 462282 53816
rect 462226 45328 462282 45384
rect 489826 53760 489882 53816
rect 514758 53760 514814 53816
rect 514758 45328 514814 45384
rect 456338 36488 456394 36544
rect 430578 34856 430634 34912
rect 430578 26288 430634 26344
rect 418342 13368 418398 13424
rect 458178 34720 458234 34776
rect 462226 34720 462282 34776
rect 458178 26832 458234 26888
rect 462226 26288 462282 26344
rect 487158 34856 487214 34912
rect 487158 26288 487214 26344
rect 514758 34720 514814 34776
rect 514758 26288 514814 26344
rect 557998 684528 558054 684584
rect 518806 674192 518862 674248
rect 518806 665896 518862 665952
rect 540610 662360 540666 662416
rect 542358 674192 542414 674248
rect 545762 674192 545818 674248
rect 520186 657192 520242 657248
rect 518806 655968 518862 656024
rect 518806 647672 518862 647728
rect 542358 647672 542414 647728
rect 518806 620200 518862 620256
rect 518806 611904 518862 611960
rect 540610 608504 540666 608560
rect 542358 620200 542414 620256
rect 542358 602112 542414 602168
rect 542358 593680 542414 593736
rect 518806 574640 518862 574696
rect 518806 566208 518862 566264
rect 540610 554648 540666 554704
rect 542358 566208 542414 566264
rect 540610 500792 540666 500848
rect 542358 520784 542414 520840
rect 542358 512216 542414 512272
rect 540610 445576 540666 445632
rect 542358 466792 542414 466848
rect 542358 458224 542414 458280
rect 542358 431704 542414 431760
rect 542358 423136 542414 423192
rect 540610 391856 540666 391912
rect 542358 404232 542414 404288
rect 542358 395800 542414 395856
rect 518806 377712 518862 377768
rect 518806 369280 518862 369336
rect 542358 377712 542414 377768
rect 540610 338000 540666 338056
rect 542358 350240 542414 350296
rect 542358 341808 542414 341864
rect 518806 323720 518862 323776
rect 518806 315288 518862 315344
rect 542358 323720 542414 323776
rect 540610 284144 540666 284200
rect 542358 296248 542414 296304
rect 542358 287816 542414 287872
rect 520186 279248 520242 279304
rect 518806 278024 518862 278080
rect 518806 269728 518862 269784
rect 542358 269728 542414 269784
rect 518806 242256 518862 242312
rect 518806 233960 518862 234016
rect 540610 230424 540666 230480
rect 542358 242256 542414 242312
rect 542358 224168 542414 224224
rect 542358 215736 542414 215792
rect 518806 196696 518862 196752
rect 518806 188264 518862 188320
rect 542358 188264 542414 188320
rect 518806 134272 518862 134328
rect 542358 142704 542414 142760
rect 542358 134272 542414 134328
rect 542358 80280 542414 80336
rect 542358 53760 542414 53816
rect 571338 674192 571394 674248
rect 571338 665896 571394 665952
rect 546406 647672 546462 647728
rect 546406 620200 546462 620256
rect 557998 630400 558054 630456
rect 571338 620200 571394 620256
rect 580262 617480 580318 617536
rect 571338 611904 571394 611960
rect 546406 593680 546462 593736
rect 546406 566208 546462 566264
rect 557998 576408 558054 576464
rect 571338 601976 571394 602032
rect 571338 593680 571394 593736
rect 571338 574640 571394 574696
rect 571338 566208 571394 566264
rect 546406 539688 546462 539744
rect 546406 512216 546462 512272
rect 557998 522416 558054 522472
rect 571338 547984 571394 548040
rect 571338 539688 571394 539744
rect 568946 520648 569002 520704
rect 568946 512760 569002 512816
rect 546406 485696 546462 485752
rect 546406 458224 546462 458280
rect 557998 468424 558054 468480
rect 571338 485696 571394 485752
rect 571338 477264 571394 477320
rect 579986 471416 580042 471472
rect 571338 466656 571394 466712
rect 571338 458224 571394 458280
rect 546406 431704 546462 431760
rect 546406 404232 546462 404288
rect 557998 414432 558054 414488
rect 571338 431704 571394 431760
rect 571338 423272 571394 423328
rect 571338 404232 571394 404288
rect 571338 395936 571394 395992
rect 546406 377712 546462 377768
rect 546406 350240 546462 350296
rect 557998 360440 558054 360496
rect 579802 378392 579858 378448
rect 546406 323720 546462 323776
rect 546406 296248 546462 296304
rect 557998 306448 558054 306504
rect 546406 269728 546462 269784
rect 546406 242256 546462 242312
rect 557998 252592 558054 252648
rect 546406 215736 546462 215792
rect 546406 188264 546462 188320
rect 546406 161744 546462 161800
rect 546406 134272 546462 134328
rect 546406 107752 546462 107808
rect 546406 80280 546462 80336
rect 546406 53216 546462 53272
rect 542358 34856 542414 34912
rect 542358 26288 542414 26344
rect 546406 26288 546462 26344
rect 557998 36488 558054 36544
rect 580170 351872 580226 351928
rect 571338 350240 571394 350296
rect 571338 341944 571394 342000
rect 580078 325216 580134 325272
rect 571338 296248 571394 296304
rect 571338 287952 571394 288008
rect 571338 242256 571394 242312
rect 571338 233960 571394 234016
rect 571338 224032 571394 224088
rect 571338 215736 571394 215792
rect 571338 196696 571394 196752
rect 571338 188264 571394 188320
rect 571338 170040 571394 170096
rect 571338 161744 571394 161800
rect 571338 134272 571394 134328
rect 571338 116048 571394 116104
rect 571338 107752 571394 107808
rect 571338 88712 571394 88768
rect 571338 80280 571394 80336
rect 571338 53760 571394 53816
rect 571338 45328 571394 45384
rect 540610 13368 540666 13424
rect 571338 34720 571394 34776
rect 571338 26288 571394 26344
rect 578882 272176 578938 272232
rect 580078 232328 580134 232384
rect 580078 192480 580134 192536
rect 580078 152632 580134 152688
rect 580078 112784 580134 112840
rect 580078 72936 580134 72992
rect 580354 590960 580410 591016
rect 580446 564304 580502 564360
rect 580538 537784 580594 537840
rect 580630 511264 580686 511320
rect 580722 484608 580778 484664
rect 580814 431568 580870 431624
rect 580906 404912 580962 404968
rect 580906 33088 580962 33144
<< metal3 >>
rect -960 697220 480 697460
rect 580206 697172 580212 697236
rect 580276 697234 580282 697236
rect 583520 697234 584960 697324
rect 580276 697174 584960 697234
rect 580276 697172 580282 697174
rect 583520 697084 584960 697174
rect 165654 684524 165660 684588
rect 165724 684586 165730 684588
rect 165981 684586 166047 684589
rect 165724 684584 166047 684586
rect 165724 684528 165986 684584
rect 166042 684528 166047 684584
rect 165724 684526 166047 684528
rect 165724 684524 165730 684526
rect 165981 684523 166047 684526
rect 259494 684524 259500 684588
rect 259564 684586 259570 684588
rect 260373 684586 260439 684589
rect 259564 684584 260439 684586
rect 259564 684528 260378 684584
rect 260434 684528 260439 684584
rect 259564 684526 260439 684528
rect 259564 684524 259570 684526
rect 260373 684523 260439 684526
rect 361614 684524 361620 684588
rect 361684 684586 361690 684588
rect 361941 684586 362007 684589
rect 361684 684584 362007 684586
rect 361684 684528 361946 684584
rect 362002 684528 362007 684584
rect 361684 684526 362007 684528
rect 361684 684524 361690 684526
rect 361941 684523 362007 684526
rect 445702 684524 445708 684588
rect 445772 684586 445778 684588
rect 446029 684586 446095 684589
rect 445772 684584 446095 684586
rect 445772 684528 446034 684584
rect 446090 684528 446095 684584
rect 445772 684526 446095 684528
rect 445772 684524 445778 684526
rect 446029 684523 446095 684526
rect 557574 684524 557580 684588
rect 557644 684586 557650 684588
rect 557993 684586 558059 684589
rect 557644 684584 558059 684586
rect 557644 684528 557998 684584
rect 558054 684528 558059 684584
rect 557644 684526 558059 684528
rect 557644 684524 557650 684526
rect 557993 684523 558059 684526
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 583520 683756 584960 683996
rect 13629 674250 13695 674253
rect 38653 674250 38719 674253
rect 13629 674248 16100 674250
rect 13629 674192 13634 674248
rect 13690 674192 16100 674248
rect 13629 674190 16100 674192
rect 36892 674248 38719 674250
rect 36892 674192 38658 674248
rect 38714 674192 38719 674248
rect 36892 674190 38719 674192
rect 13629 674187 13695 674190
rect 38653 674187 38719 674190
rect 42701 674250 42767 674253
rect 66253 674250 66319 674253
rect 95233 674250 95299 674253
rect 42701 674248 44068 674250
rect 42701 674192 42706 674248
rect 42762 674192 44068 674248
rect 42701 674190 44068 674192
rect 64860 674248 66319 674250
rect 64860 674192 66258 674248
rect 66314 674192 66319 674248
rect 92828 674248 95299 674250
rect 64860 674190 66319 674192
rect 42701 674187 42767 674190
rect 66253 674187 66319 674190
rect 70301 673842 70367 673845
rect 72006 673842 72066 674220
rect 92828 674192 95238 674248
rect 95294 674192 95299 674248
rect 92828 674190 95299 674192
rect 95233 674187 95299 674190
rect 97901 674250 97967 674253
rect 122833 674250 122899 674253
rect 97901 674248 100188 674250
rect 97901 674192 97906 674248
rect 97962 674192 100188 674248
rect 97901 674190 100188 674192
rect 120796 674248 122899 674250
rect 120796 674192 122838 674248
rect 122894 674192 122899 674248
rect 120796 674190 122899 674192
rect 97901 674187 97967 674190
rect 122833 674187 122899 674190
rect 126881 674250 126947 674253
rect 150433 674250 150499 674253
rect 126881 674248 128156 674250
rect 126881 674192 126886 674248
rect 126942 674192 128156 674248
rect 126881 674190 128156 674192
rect 148948 674248 150499 674250
rect 148948 674192 150438 674248
rect 150494 674192 150499 674248
rect 148948 674190 150499 674192
rect 126881 674187 126947 674190
rect 150433 674187 150499 674190
rect 154481 674250 154547 674253
rect 178033 674250 178099 674253
rect 154481 674248 156124 674250
rect 154481 674192 154486 674248
rect 154542 674192 156124 674248
rect 154481 674190 156124 674192
rect 176916 674248 178099 674250
rect 176916 674192 178038 674248
rect 178094 674192 178099 674248
rect 176916 674190 178099 674192
rect 154481 674187 154547 674190
rect 178033 674187 178099 674190
rect 182081 674250 182147 674253
rect 207013 674250 207079 674253
rect 182081 674248 184092 674250
rect 182081 674192 182086 674248
rect 182142 674192 184092 674248
rect 182081 674190 184092 674192
rect 204884 674248 207079 674250
rect 204884 674192 207018 674248
rect 207074 674192 207079 674248
rect 204884 674190 207079 674192
rect 182081 674187 182147 674190
rect 207013 674187 207079 674190
rect 209681 674250 209747 674253
rect 234705 674250 234771 674253
rect 209681 674248 212060 674250
rect 209681 674192 209686 674248
rect 209742 674192 212060 674248
rect 209681 674190 212060 674192
rect 232852 674248 234771 674250
rect 232852 674192 234710 674248
rect 234766 674192 234771 674248
rect 232852 674190 234771 674192
rect 209681 674187 209747 674190
rect 234705 674187 234771 674190
rect 238661 674250 238727 674253
rect 262213 674250 262279 674253
rect 238661 674248 240212 674250
rect 238661 674192 238666 674248
rect 238722 674192 240212 674248
rect 238661 674190 240212 674192
rect 260820 674248 262279 674250
rect 260820 674192 262218 674248
rect 262274 674192 262279 674248
rect 260820 674190 262279 674192
rect 238661 674187 238727 674190
rect 262213 674187 262279 674190
rect 266261 674250 266327 674253
rect 291193 674250 291259 674253
rect 266261 674248 268180 674250
rect 266261 674192 266266 674248
rect 266322 674192 268180 674248
rect 266261 674190 268180 674192
rect 288788 674248 291259 674250
rect 288788 674192 291198 674248
rect 291254 674192 291259 674248
rect 288788 674190 291259 674192
rect 266261 674187 266327 674190
rect 291193 674187 291259 674190
rect 293861 674250 293927 674253
rect 318793 674250 318859 674253
rect 293861 674248 296148 674250
rect 293861 674192 293866 674248
rect 293922 674192 296148 674248
rect 293861 674190 296148 674192
rect 316940 674248 318859 674250
rect 316940 674192 318798 674248
rect 318854 674192 318859 674248
rect 316940 674190 318859 674192
rect 293861 674187 293927 674190
rect 318793 674187 318859 674190
rect 322841 674250 322907 674253
rect 346393 674250 346459 674253
rect 322841 674248 324116 674250
rect 322841 674192 322846 674248
rect 322902 674192 324116 674248
rect 322841 674190 324116 674192
rect 344908 674248 346459 674250
rect 344908 674192 346398 674248
rect 346454 674192 346459 674248
rect 344908 674190 346459 674192
rect 322841 674187 322907 674190
rect 346393 674187 346459 674190
rect 350441 674250 350507 674253
rect 375373 674250 375439 674253
rect 350441 674248 352084 674250
rect 350441 674192 350446 674248
rect 350502 674192 352084 674248
rect 350441 674190 352084 674192
rect 372876 674248 375439 674250
rect 372876 674192 375378 674248
rect 375434 674192 375439 674248
rect 372876 674190 375439 674192
rect 350441 674187 350507 674190
rect 375373 674187 375439 674190
rect 378041 674250 378107 674253
rect 402973 674250 403039 674253
rect 378041 674248 380052 674250
rect 378041 674192 378046 674248
rect 378102 674192 380052 674248
rect 378041 674190 380052 674192
rect 400844 674248 403039 674250
rect 400844 674192 402978 674248
rect 403034 674192 403039 674248
rect 400844 674190 403039 674192
rect 378041 674187 378107 674190
rect 402973 674187 403039 674190
rect 405641 674250 405707 674253
rect 430573 674250 430639 674253
rect 405641 674248 408204 674250
rect 405641 674192 405646 674248
rect 405702 674192 408204 674248
rect 405641 674190 408204 674192
rect 428812 674248 430639 674250
rect 428812 674192 430578 674248
rect 430634 674192 430639 674248
rect 428812 674190 430639 674192
rect 405641 674187 405707 674190
rect 430573 674187 430639 674190
rect 434621 674250 434687 674253
rect 462221 674250 462287 674253
rect 487153 674250 487219 674253
rect 434621 674248 436172 674250
rect 434621 674192 434626 674248
rect 434682 674192 436172 674248
rect 462221 674248 464140 674250
rect 434621 674190 436172 674192
rect 434621 674187 434687 674190
rect 70301 673840 72066 673842
rect 70301 673784 70306 673840
rect 70362 673784 72066 673840
rect 70301 673782 72066 673784
rect 456934 673842 456994 674220
rect 462221 674192 462226 674248
rect 462282 674192 464140 674248
rect 462221 674190 464140 674192
rect 484932 674248 487219 674250
rect 484932 674192 487158 674248
rect 487214 674192 487219 674248
rect 484932 674190 487219 674192
rect 462221 674187 462287 674190
rect 487153 674187 487219 674190
rect 489821 674250 489887 674253
rect 514753 674250 514819 674253
rect 489821 674248 492108 674250
rect 489821 674192 489826 674248
rect 489882 674192 492108 674248
rect 489821 674190 492108 674192
rect 512900 674248 514819 674250
rect 512900 674192 514758 674248
rect 514814 674192 514819 674248
rect 512900 674190 514819 674192
rect 489821 674187 489887 674190
rect 514753 674187 514819 674190
rect 518801 674250 518867 674253
rect 542353 674250 542419 674253
rect 518801 674248 520076 674250
rect 518801 674192 518806 674248
rect 518862 674192 520076 674248
rect 518801 674190 520076 674192
rect 540868 674248 542419 674250
rect 540868 674192 542358 674248
rect 542414 674192 542419 674248
rect 540868 674190 542419 674192
rect 518801 674187 518867 674190
rect 542353 674187 542419 674190
rect 545757 674250 545823 674253
rect 571333 674250 571399 674253
rect 545757 674248 548044 674250
rect 545757 674192 545762 674248
rect 545818 674192 548044 674248
rect 545757 674190 548044 674192
rect 568836 674248 571399 674250
rect 568836 674192 571338 674248
rect 571394 674192 571399 674248
rect 568836 674190 571399 674192
rect 545757 674187 545823 674190
rect 571333 674187 571399 674190
rect 458173 673842 458239 673845
rect 456934 673840 458239 673842
rect 456934 673784 458178 673840
rect 458234 673784 458239 673840
rect 456934 673782 458239 673784
rect 70301 673779 70367 673782
rect 458173 673779 458239 673782
rect -960 671108 480 671348
rect 580390 670652 580396 670716
rect 580460 670714 580466 670716
rect 583520 670714 584960 670804
rect 580460 670654 584960 670714
rect 580460 670652 580466 670654
rect 583520 670564 584960 670654
rect 13629 665954 13695 665957
rect 66253 665954 66319 665957
rect 13629 665952 66319 665954
rect 13629 665896 13634 665952
rect 13690 665896 66258 665952
rect 66314 665896 66319 665952
rect 13629 665894 66319 665896
rect 13629 665891 13695 665894
rect 66253 665891 66319 665894
rect 70301 665954 70367 665957
rect 122833 665954 122899 665957
rect 70301 665952 122899 665954
rect 70301 665896 70306 665952
rect 70362 665896 122838 665952
rect 122894 665896 122899 665952
rect 70301 665894 122899 665896
rect 70301 665891 70367 665894
rect 122833 665891 122899 665894
rect 126881 665954 126947 665957
rect 178033 665954 178099 665957
rect 126881 665952 178099 665954
rect 126881 665896 126886 665952
rect 126942 665896 178038 665952
rect 178094 665896 178099 665952
rect 126881 665894 178099 665896
rect 126881 665891 126947 665894
rect 178033 665891 178099 665894
rect 182081 665954 182147 665957
rect 234705 665954 234771 665957
rect 182081 665952 234771 665954
rect 182081 665896 182086 665952
rect 182142 665896 234710 665952
rect 234766 665896 234771 665952
rect 182081 665894 234771 665896
rect 182081 665891 182147 665894
rect 234705 665891 234771 665894
rect 238661 665954 238727 665957
rect 291193 665954 291259 665957
rect 238661 665952 291259 665954
rect 238661 665896 238666 665952
rect 238722 665896 291198 665952
rect 291254 665896 291259 665952
rect 238661 665894 291259 665896
rect 238661 665891 238727 665894
rect 291193 665891 291259 665894
rect 293861 665954 293927 665957
rect 346393 665954 346459 665957
rect 293861 665952 346459 665954
rect 293861 665896 293866 665952
rect 293922 665896 346398 665952
rect 346454 665896 346459 665952
rect 293861 665894 346459 665896
rect 293861 665891 293927 665894
rect 346393 665891 346459 665894
rect 350441 665954 350507 665957
rect 402973 665954 403039 665957
rect 350441 665952 403039 665954
rect 350441 665896 350446 665952
rect 350502 665896 402978 665952
rect 403034 665896 403039 665952
rect 350441 665894 403039 665896
rect 350441 665891 350507 665894
rect 402973 665891 403039 665894
rect 405641 665954 405707 665957
rect 458173 665954 458239 665957
rect 405641 665952 458239 665954
rect 405641 665896 405646 665952
rect 405702 665896 458178 665952
rect 458234 665896 458239 665952
rect 405641 665894 458239 665896
rect 405641 665891 405707 665894
rect 458173 665891 458239 665894
rect 462221 665954 462287 665957
rect 514753 665954 514819 665957
rect 462221 665952 514819 665954
rect 462221 665896 462226 665952
rect 462282 665896 514758 665952
rect 514814 665896 514819 665952
rect 462221 665894 514819 665896
rect 462221 665891 462287 665894
rect 514753 665891 514819 665894
rect 518801 665954 518867 665957
rect 571333 665954 571399 665957
rect 518801 665952 571399 665954
rect 518801 665896 518806 665952
rect 518862 665896 571338 665952
rect 571394 665896 571399 665952
rect 518801 665894 571399 665896
rect 518801 665891 518867 665894
rect 571333 665891 571399 665894
rect 148685 662418 148751 662421
rect 165654 662418 165660 662420
rect 148685 662416 165660 662418
rect 148685 662360 148690 662416
rect 148746 662360 165660 662416
rect 148685 662358 165660 662360
rect 148685 662355 148751 662358
rect 165654 662356 165660 662358
rect 165724 662356 165730 662420
rect 222653 662418 222719 662421
rect 259494 662418 259500 662420
rect 222653 662416 259500 662418
rect 222653 662360 222658 662416
rect 222714 662360 259500 662416
rect 222653 662358 259500 662360
rect 222653 662355 222719 662358
rect 259494 662356 259500 662358
rect 259564 662356 259570 662420
rect 344921 662418 344987 662421
rect 361614 662418 361620 662420
rect 344921 662416 361620 662418
rect 344921 662360 344926 662416
rect 344982 662360 361620 662416
rect 344921 662358 361620 662360
rect 344921 662355 344987 662358
rect 361614 662356 361620 662358
rect 361684 662356 361690 662420
rect 428641 662418 428707 662421
rect 445702 662418 445708 662420
rect 428641 662416 445708 662418
rect 428641 662360 428646 662416
rect 428702 662360 445708 662416
rect 428641 662358 445708 662360
rect 428641 662355 428707 662358
rect 445702 662356 445708 662358
rect 445772 662356 445778 662420
rect 540605 662418 540671 662421
rect 557574 662418 557580 662420
rect 540605 662416 557580 662418
rect 540605 662360 540610 662416
rect 540666 662360 557580 662416
rect 540605 662358 557580 662360
rect 540605 662355 540671 662358
rect 557574 662356 557580 662358
rect 557644 662356 557650 662420
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 81382 657324 81388 657388
rect 81452 657386 81458 657388
rect 82261 657386 82327 657389
rect 81452 657384 82327 657386
rect 81452 657328 82266 657384
rect 82322 657328 82327 657384
rect 81452 657326 82327 657328
rect 81452 657324 81458 657326
rect 82261 657323 82327 657326
rect 128302 657324 128308 657388
rect 128372 657386 128378 657388
rect 128445 657386 128511 657389
rect 194777 657388 194843 657389
rect 194726 657386 194732 657388
rect 128372 657384 128511 657386
rect 128372 657328 128450 657384
rect 128506 657328 128511 657384
rect 128372 657326 128511 657328
rect 194686 657326 194732 657386
rect 194796 657384 194843 657388
rect 194838 657328 194843 657384
rect 128372 657324 128378 657326
rect 128445 657323 128511 657326
rect 194726 657324 194732 657326
rect 194796 657324 194843 657328
rect 277526 657324 277532 657388
rect 277596 657386 277602 657388
rect 278221 657386 278287 657389
rect 277596 657384 278287 657386
rect 277596 657328 278226 657384
rect 278282 657328 278287 657384
rect 277596 657326 278287 657328
rect 277596 657324 277602 657326
rect 194777 657323 194843 657324
rect 278221 657323 278287 657326
rect 390829 657388 390895 657389
rect 390829 657384 390876 657388
rect 390940 657386 390946 657388
rect 390829 657328 390834 657384
rect 390829 657324 390876 657328
rect 390940 657326 390986 657386
rect 390940 657324 390946 657326
rect 473486 657324 473492 657388
rect 473556 657386 473562 657388
rect 474273 657386 474339 657389
rect 473556 657384 474339 657386
rect 473556 657328 474278 657384
rect 474334 657328 474339 657384
rect 473556 657326 474339 657328
rect 473556 657324 473562 657326
rect 390829 657323 390895 657324
rect 474273 657323 474339 657326
rect 520181 657252 520247 657253
rect 520181 657248 520228 657252
rect 520292 657250 520298 657252
rect 520181 657192 520186 657248
rect 520181 657188 520228 657192
rect 520292 657190 520338 657250
rect 583520 657236 584960 657476
rect 520292 657188 520298 657190
rect 520181 657187 520247 657188
rect 13721 656026 13787 656029
rect 66253 656026 66319 656029
rect 13721 656024 66319 656026
rect 13721 655968 13726 656024
rect 13782 655968 66258 656024
rect 66314 655968 66319 656024
rect 13721 655966 66319 655968
rect 13721 655963 13787 655966
rect 66253 655963 66319 655966
rect 70301 656026 70367 656029
rect 122833 656026 122899 656029
rect 70301 656024 122899 656026
rect 70301 655968 70306 656024
rect 70362 655968 122838 656024
rect 122894 655968 122899 656024
rect 70301 655966 122899 655968
rect 70301 655963 70367 655966
rect 122833 655963 122899 655966
rect 126881 656026 126947 656029
rect 176326 656026 176332 656028
rect 126881 656024 176332 656026
rect 126881 655968 126886 656024
rect 126942 655968 176332 656024
rect 126881 655966 176332 655968
rect 126881 655963 126947 655966
rect 176326 655964 176332 655966
rect 176396 655964 176402 656028
rect 184197 656026 184263 656029
rect 234705 656026 234771 656029
rect 184197 656024 234771 656026
rect 184197 655968 184202 656024
rect 184258 655968 234710 656024
rect 234766 655968 234771 656024
rect 184197 655966 234771 655968
rect 184197 655963 184263 655966
rect 234705 655963 234771 655966
rect 238661 656026 238727 656029
rect 291193 656026 291259 656029
rect 238661 656024 291259 656026
rect 238661 655968 238666 656024
rect 238722 655968 291198 656024
rect 291254 655968 291259 656024
rect 238661 655966 291259 655968
rect 238661 655963 238727 655966
rect 291193 655963 291259 655966
rect 293861 656026 293927 656029
rect 346393 656026 346459 656029
rect 293861 656024 346459 656026
rect 293861 655968 293866 656024
rect 293922 655968 346398 656024
rect 346454 655968 346459 656024
rect 293861 655966 346459 655968
rect 293861 655963 293927 655966
rect 346393 655963 346459 655966
rect 350441 656026 350507 656029
rect 402973 656026 403039 656029
rect 350441 656024 403039 656026
rect 350441 655968 350446 656024
rect 350502 655968 402978 656024
rect 403034 655968 403039 656024
rect 350441 655966 403039 655968
rect 350441 655963 350507 655966
rect 402973 655963 403039 655966
rect 408125 656026 408191 656029
rect 456374 656026 456380 656028
rect 408125 656024 456380 656026
rect 408125 655968 408130 656024
rect 408186 655968 456380 656024
rect 408125 655966 456380 655968
rect 408125 655963 408191 655966
rect 456374 655964 456380 655966
rect 456444 655964 456450 656028
rect 464153 656026 464219 656029
rect 514753 656026 514819 656029
rect 464153 656024 514819 656026
rect 464153 655968 464158 656024
rect 464214 655968 514758 656024
rect 514814 655968 514819 656024
rect 464153 655966 514819 655968
rect 464153 655963 464219 655966
rect 514753 655963 514819 655966
rect 518801 656026 518867 656029
rect 568430 656026 568436 656028
rect 518801 656024 568436 656026
rect 518801 655968 518806 656024
rect 518862 655968 568436 656024
rect 518801 655966 568436 655968
rect 518801 655963 518867 655966
rect 568430 655964 568436 655966
rect 568500 655964 568506 656028
rect 176326 648212 176332 648276
rect 176396 648212 176402 648276
rect 184197 648274 184263 648277
rect 408125 648274 408191 648277
rect 184197 648272 184306 648274
rect 184197 648216 184202 648272
rect 184258 648216 184306 648272
rect 13721 647730 13787 647733
rect 38653 647730 38719 647733
rect 13721 647728 16100 647730
rect 13721 647672 13726 647728
rect 13782 647672 16100 647728
rect 13721 647670 16100 647672
rect 36892 647728 38719 647730
rect 36892 647672 38658 647728
rect 38714 647672 38719 647728
rect 36892 647670 38719 647672
rect 13721 647667 13787 647670
rect 38653 647667 38719 647670
rect 42701 647730 42767 647733
rect 66253 647730 66319 647733
rect 42701 647728 44068 647730
rect 42701 647672 42706 647728
rect 42762 647672 44068 647728
rect 42701 647670 44068 647672
rect 64860 647728 66319 647730
rect 64860 647672 66258 647728
rect 66314 647672 66319 647728
rect 64860 647670 66319 647672
rect 42701 647667 42767 647670
rect 66253 647667 66319 647670
rect 70301 647730 70367 647733
rect 95233 647730 95299 647733
rect 70301 647728 72036 647730
rect 70301 647672 70306 647728
rect 70362 647672 72036 647728
rect 70301 647670 72036 647672
rect 92828 647728 95299 647730
rect 92828 647672 95238 647728
rect 95294 647672 95299 647728
rect 92828 647670 95299 647672
rect 70301 647667 70367 647670
rect 95233 647667 95299 647670
rect 97901 647730 97967 647733
rect 122833 647730 122899 647733
rect 97901 647728 100188 647730
rect 97901 647672 97906 647728
rect 97962 647672 100188 647728
rect 97901 647670 100188 647672
rect 120796 647728 122899 647730
rect 120796 647672 122838 647728
rect 122894 647672 122899 647728
rect 120796 647670 122899 647672
rect 97901 647667 97967 647670
rect 122833 647667 122899 647670
rect 126881 647730 126947 647733
rect 150433 647730 150499 647733
rect 126881 647728 128156 647730
rect 126881 647672 126886 647728
rect 126942 647672 128156 647728
rect 126881 647670 128156 647672
rect 148948 647728 150499 647730
rect 148948 647672 150438 647728
rect 150494 647672 150499 647728
rect 148948 647670 150499 647672
rect 126881 647667 126947 647670
rect 150433 647667 150499 647670
rect 154481 647730 154547 647733
rect 154481 647728 156124 647730
rect 154481 647672 154486 647728
rect 154542 647672 156124 647728
rect 176334 647700 176394 648212
rect 184197 648211 184306 648216
rect 408125 648272 408234 648274
rect 408125 648216 408130 648272
rect 408186 648216 408234 648272
rect 408125 648211 408234 648216
rect 456374 648212 456380 648276
rect 456444 648212 456450 648276
rect 464153 648274 464219 648277
rect 464110 648272 464219 648274
rect 464110 648216 464158 648272
rect 464214 648216 464219 648272
rect 184246 647700 184306 648211
rect 207013 647730 207079 647733
rect 204884 647728 207079 647730
rect 154481 647670 156124 647672
rect 204884 647672 207018 647728
rect 207074 647672 207079 647728
rect 204884 647670 207079 647672
rect 154481 647667 154547 647670
rect 207013 647667 207079 647670
rect 209681 647730 209747 647733
rect 234705 647730 234771 647733
rect 209681 647728 212060 647730
rect 209681 647672 209686 647728
rect 209742 647672 212060 647728
rect 209681 647670 212060 647672
rect 232852 647728 234771 647730
rect 232852 647672 234710 647728
rect 234766 647672 234771 647728
rect 232852 647670 234771 647672
rect 209681 647667 209747 647670
rect 234705 647667 234771 647670
rect 238661 647730 238727 647733
rect 262213 647730 262279 647733
rect 238661 647728 240212 647730
rect 238661 647672 238666 647728
rect 238722 647672 240212 647728
rect 238661 647670 240212 647672
rect 260820 647728 262279 647730
rect 260820 647672 262218 647728
rect 262274 647672 262279 647728
rect 260820 647670 262279 647672
rect 238661 647667 238727 647670
rect 262213 647667 262279 647670
rect 266261 647730 266327 647733
rect 291193 647730 291259 647733
rect 266261 647728 268180 647730
rect 266261 647672 266266 647728
rect 266322 647672 268180 647728
rect 266261 647670 268180 647672
rect 288788 647728 291259 647730
rect 288788 647672 291198 647728
rect 291254 647672 291259 647728
rect 288788 647670 291259 647672
rect 266261 647667 266327 647670
rect 291193 647667 291259 647670
rect 293861 647730 293927 647733
rect 318793 647730 318859 647733
rect 293861 647728 296148 647730
rect 293861 647672 293866 647728
rect 293922 647672 296148 647728
rect 293861 647670 296148 647672
rect 316940 647728 318859 647730
rect 316940 647672 318798 647728
rect 318854 647672 318859 647728
rect 316940 647670 318859 647672
rect 293861 647667 293927 647670
rect 318793 647667 318859 647670
rect 322841 647730 322907 647733
rect 346393 647730 346459 647733
rect 322841 647728 324116 647730
rect 322841 647672 322846 647728
rect 322902 647672 324116 647728
rect 322841 647670 324116 647672
rect 344908 647728 346459 647730
rect 344908 647672 346398 647728
rect 346454 647672 346459 647728
rect 344908 647670 346459 647672
rect 322841 647667 322907 647670
rect 346393 647667 346459 647670
rect 350441 647730 350507 647733
rect 375373 647730 375439 647733
rect 350441 647728 352084 647730
rect 350441 647672 350446 647728
rect 350502 647672 352084 647728
rect 350441 647670 352084 647672
rect 372876 647728 375439 647730
rect 372876 647672 375378 647728
rect 375434 647672 375439 647728
rect 372876 647670 375439 647672
rect 350441 647667 350507 647670
rect 375373 647667 375439 647670
rect 378041 647730 378107 647733
rect 402973 647730 403039 647733
rect 378041 647728 380052 647730
rect 378041 647672 378046 647728
rect 378102 647672 380052 647728
rect 378041 647670 380052 647672
rect 400844 647728 403039 647730
rect 400844 647672 402978 647728
rect 403034 647672 403039 647728
rect 408174 647700 408234 648211
rect 430573 647730 430639 647733
rect 428812 647728 430639 647730
rect 400844 647670 403039 647672
rect 428812 647672 430578 647728
rect 430634 647672 430639 647728
rect 428812 647670 430639 647672
rect 378041 647667 378107 647670
rect 402973 647667 403039 647670
rect 430573 647667 430639 647670
rect 434621 647730 434687 647733
rect 434621 647728 436172 647730
rect 434621 647672 434626 647728
rect 434682 647672 436172 647728
rect 456382 647700 456442 648212
rect 464110 648211 464219 648216
rect 568430 648212 568436 648276
rect 568500 648212 568506 648276
rect 464110 647700 464170 648211
rect 487153 647730 487219 647733
rect 484932 647728 487219 647730
rect 434621 647670 436172 647672
rect 484932 647672 487158 647728
rect 487214 647672 487219 647728
rect 484932 647670 487219 647672
rect 434621 647667 434687 647670
rect 487153 647667 487219 647670
rect 489821 647730 489887 647733
rect 514753 647730 514819 647733
rect 489821 647728 492108 647730
rect 489821 647672 489826 647728
rect 489882 647672 492108 647728
rect 489821 647670 492108 647672
rect 512900 647728 514819 647730
rect 512900 647672 514758 647728
rect 514814 647672 514819 647728
rect 512900 647670 514819 647672
rect 489821 647667 489887 647670
rect 514753 647667 514819 647670
rect 518801 647730 518867 647733
rect 542353 647730 542419 647733
rect 518801 647728 520076 647730
rect 518801 647672 518806 647728
rect 518862 647672 520076 647728
rect 518801 647670 520076 647672
rect 540868 647728 542419 647730
rect 540868 647672 542358 647728
rect 542414 647672 542419 647728
rect 540868 647670 542419 647672
rect 518801 647667 518867 647670
rect 542353 647667 542419 647670
rect 546401 647730 546467 647733
rect 546401 647728 548044 647730
rect 546401 647672 546406 647728
rect 546462 647672 548044 647728
rect 568438 647700 568498 648212
rect 546401 647670 548044 647672
rect 546401 647667 546467 647670
rect -960 644996 480 645236
rect 580574 643996 580580 644060
rect 580644 644058 580650 644060
rect 583520 644058 584960 644148
rect 580644 643998 584960 644058
rect 580644 643996 580650 643998
rect 583520 643908 584960 643998
rect 44633 634810 44699 634813
rect 81382 634810 81388 634812
rect 44633 634808 81388 634810
rect 44633 634752 44638 634808
rect 44694 634752 81388 634808
rect 44633 634750 81388 634752
rect 44633 634747 44699 634750
rect 81382 634748 81388 634750
rect 81452 634748 81458 634812
rect 110597 634810 110663 634813
rect 128302 634810 128308 634812
rect 110597 634808 128308 634810
rect 110597 634752 110602 634808
rect 110658 634752 128308 634808
rect 110597 634750 128308 634752
rect 110597 634747 110663 634750
rect 128302 634748 128308 634750
rect 128372 634748 128378 634812
rect 156321 634810 156387 634813
rect 194726 634810 194732 634812
rect 156321 634808 194732 634810
rect 156321 634752 156326 634808
rect 156382 634752 194732 634808
rect 156321 634750 194732 634752
rect 156321 634747 156387 634750
rect 194726 634748 194732 634750
rect 194796 634748 194802 634812
rect 240317 634810 240383 634813
rect 277158 634810 277164 634812
rect 240317 634808 277164 634810
rect 240317 634752 240322 634808
rect 240378 634752 277164 634808
rect 240317 634750 277164 634752
rect 240317 634747 240383 634750
rect 277158 634748 277164 634750
rect 277228 634748 277234 634812
rect 352649 634810 352715 634813
rect 390870 634810 390876 634812
rect 352649 634808 390876 634810
rect 352649 634752 352654 634808
rect 352710 634752 390876 634808
rect 352649 634750 390876 634752
rect 352649 634747 352715 634750
rect 390870 634748 390876 634750
rect 390940 634748 390946 634812
rect 436645 634810 436711 634813
rect 473486 634810 473492 634812
rect 436645 634808 473492 634810
rect 436645 634752 436650 634808
rect 436706 634752 473492 634808
rect 436645 634750 473492 634752
rect 436645 634747 436711 634750
rect 473486 634748 473492 634750
rect 473556 634748 473562 634812
rect 502609 634810 502675 634813
rect 520222 634810 520228 634812
rect 502609 634808 520228 634810
rect 502609 634752 502614 634808
rect 502670 634752 520228 634808
rect 502609 634750 520228 634752
rect 502609 634747 502675 634750
rect 520222 634748 520228 634750
rect 520292 634748 520298 634812
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 583520 630716 584960 630956
rect 165654 630396 165660 630460
rect 165724 630458 165730 630460
rect 165981 630458 166047 630461
rect 165724 630456 166047 630458
rect 165724 630400 165986 630456
rect 166042 630400 166047 630456
rect 165724 630398 166047 630400
rect 165724 630396 165730 630398
rect 165981 630395 166047 630398
rect 259494 630396 259500 630460
rect 259564 630458 259570 630460
rect 260373 630458 260439 630461
rect 259564 630456 260439 630458
rect 259564 630400 260378 630456
rect 260434 630400 260439 630456
rect 259564 630398 260439 630400
rect 259564 630396 259570 630398
rect 260373 630395 260439 630398
rect 361614 630396 361620 630460
rect 361684 630458 361690 630460
rect 361941 630458 362007 630461
rect 361684 630456 362007 630458
rect 361684 630400 361946 630456
rect 362002 630400 362007 630456
rect 361684 630398 362007 630400
rect 361684 630396 361690 630398
rect 361941 630395 362007 630398
rect 445702 630396 445708 630460
rect 445772 630458 445778 630460
rect 446029 630458 446095 630461
rect 445772 630456 446095 630458
rect 445772 630400 446034 630456
rect 446090 630400 446095 630456
rect 445772 630398 446095 630400
rect 445772 630396 445778 630398
rect 446029 630395 446095 630398
rect 557574 630396 557580 630460
rect 557644 630458 557650 630460
rect 557993 630458 558059 630461
rect 557644 630456 558059 630458
rect 557644 630400 557998 630456
rect 558054 630400 558059 630456
rect 557644 630398 558059 630400
rect 557644 630396 557650 630398
rect 557993 630395 558059 630398
rect 13537 620258 13603 620261
rect 38653 620258 38719 620261
rect 13537 620256 16100 620258
rect 13537 620200 13542 620256
rect 13598 620200 16100 620256
rect 13537 620198 16100 620200
rect 36892 620256 38719 620258
rect 36892 620200 38658 620256
rect 38714 620200 38719 620256
rect 36892 620198 38719 620200
rect 13537 620195 13603 620198
rect 38653 620195 38719 620198
rect 42701 620258 42767 620261
rect 66253 620258 66319 620261
rect 42701 620256 44068 620258
rect 42701 620200 42706 620256
rect 42762 620200 44068 620256
rect 42701 620198 44068 620200
rect 64860 620256 66319 620258
rect 64860 620200 66258 620256
rect 66314 620200 66319 620256
rect 64860 620198 66319 620200
rect 42701 620195 42767 620198
rect 66253 620195 66319 620198
rect 70301 620258 70367 620261
rect 95233 620258 95299 620261
rect 70301 620256 72036 620258
rect 70301 620200 70306 620256
rect 70362 620200 72036 620256
rect 70301 620198 72036 620200
rect 92828 620256 95299 620258
rect 92828 620200 95238 620256
rect 95294 620200 95299 620256
rect 92828 620198 95299 620200
rect 70301 620195 70367 620198
rect 95233 620195 95299 620198
rect 97901 620258 97967 620261
rect 122833 620258 122899 620261
rect 97901 620256 100188 620258
rect 97901 620200 97906 620256
rect 97962 620200 100188 620256
rect 97901 620198 100188 620200
rect 120796 620256 122899 620258
rect 120796 620200 122838 620256
rect 122894 620200 122899 620256
rect 120796 620198 122899 620200
rect 97901 620195 97967 620198
rect 122833 620195 122899 620198
rect 126881 620258 126947 620261
rect 150433 620258 150499 620261
rect 126881 620256 128156 620258
rect 126881 620200 126886 620256
rect 126942 620200 128156 620256
rect 126881 620198 128156 620200
rect 148948 620256 150499 620258
rect 148948 620200 150438 620256
rect 150494 620200 150499 620256
rect 148948 620198 150499 620200
rect 126881 620195 126947 620198
rect 150433 620195 150499 620198
rect 154481 620258 154547 620261
rect 178033 620258 178099 620261
rect 154481 620256 156124 620258
rect 154481 620200 154486 620256
rect 154542 620200 156124 620256
rect 154481 620198 156124 620200
rect 176916 620256 178099 620258
rect 176916 620200 178038 620256
rect 178094 620200 178099 620256
rect 176916 620198 178099 620200
rect 154481 620195 154547 620198
rect 178033 620195 178099 620198
rect 182081 620258 182147 620261
rect 207013 620258 207079 620261
rect 182081 620256 184092 620258
rect 182081 620200 182086 620256
rect 182142 620200 184092 620256
rect 182081 620198 184092 620200
rect 204884 620256 207079 620258
rect 204884 620200 207018 620256
rect 207074 620200 207079 620256
rect 204884 620198 207079 620200
rect 182081 620195 182147 620198
rect 207013 620195 207079 620198
rect 209681 620258 209747 620261
rect 234705 620258 234771 620261
rect 209681 620256 212060 620258
rect 209681 620200 209686 620256
rect 209742 620200 212060 620256
rect 209681 620198 212060 620200
rect 232852 620256 234771 620258
rect 232852 620200 234710 620256
rect 234766 620200 234771 620256
rect 232852 620198 234771 620200
rect 209681 620195 209747 620198
rect 234705 620195 234771 620198
rect 238661 620258 238727 620261
rect 262213 620258 262279 620261
rect 238661 620256 240212 620258
rect 238661 620200 238666 620256
rect 238722 620200 240212 620256
rect 238661 620198 240212 620200
rect 260820 620256 262279 620258
rect 260820 620200 262218 620256
rect 262274 620200 262279 620256
rect 260820 620198 262279 620200
rect 238661 620195 238727 620198
rect 262213 620195 262279 620198
rect 266261 620258 266327 620261
rect 291193 620258 291259 620261
rect 266261 620256 268180 620258
rect 266261 620200 266266 620256
rect 266322 620200 268180 620256
rect 266261 620198 268180 620200
rect 288788 620256 291259 620258
rect 288788 620200 291198 620256
rect 291254 620200 291259 620256
rect 288788 620198 291259 620200
rect 266261 620195 266327 620198
rect 291193 620195 291259 620198
rect 293861 620258 293927 620261
rect 318793 620258 318859 620261
rect 293861 620256 296148 620258
rect 293861 620200 293866 620256
rect 293922 620200 296148 620256
rect 293861 620198 296148 620200
rect 316940 620256 318859 620258
rect 316940 620200 318798 620256
rect 318854 620200 318859 620256
rect 316940 620198 318859 620200
rect 293861 620195 293927 620198
rect 318793 620195 318859 620198
rect 322841 620258 322907 620261
rect 346393 620258 346459 620261
rect 322841 620256 324116 620258
rect 322841 620200 322846 620256
rect 322902 620200 324116 620256
rect 322841 620198 324116 620200
rect 344908 620256 346459 620258
rect 344908 620200 346398 620256
rect 346454 620200 346459 620256
rect 344908 620198 346459 620200
rect 322841 620195 322907 620198
rect 346393 620195 346459 620198
rect 350441 620258 350507 620261
rect 375373 620258 375439 620261
rect 350441 620256 352084 620258
rect 350441 620200 350446 620256
rect 350502 620200 352084 620256
rect 350441 620198 352084 620200
rect 372876 620256 375439 620258
rect 372876 620200 375378 620256
rect 375434 620200 375439 620256
rect 372876 620198 375439 620200
rect 350441 620195 350507 620198
rect 375373 620195 375439 620198
rect 378041 620258 378107 620261
rect 402973 620258 403039 620261
rect 378041 620256 380052 620258
rect 378041 620200 378046 620256
rect 378102 620200 380052 620256
rect 378041 620198 380052 620200
rect 400844 620256 403039 620258
rect 400844 620200 402978 620256
rect 403034 620200 403039 620256
rect 400844 620198 403039 620200
rect 378041 620195 378107 620198
rect 402973 620195 403039 620198
rect 405641 620258 405707 620261
rect 430573 620258 430639 620261
rect 405641 620256 408204 620258
rect 405641 620200 405646 620256
rect 405702 620200 408204 620256
rect 405641 620198 408204 620200
rect 428812 620256 430639 620258
rect 428812 620200 430578 620256
rect 430634 620200 430639 620256
rect 428812 620198 430639 620200
rect 405641 620195 405707 620198
rect 430573 620195 430639 620198
rect 434621 620258 434687 620261
rect 458173 620258 458239 620261
rect 434621 620256 436172 620258
rect 434621 620200 434626 620256
rect 434682 620200 436172 620256
rect 434621 620198 436172 620200
rect 456964 620256 458239 620258
rect 456964 620200 458178 620256
rect 458234 620200 458239 620256
rect 456964 620198 458239 620200
rect 434621 620195 434687 620198
rect 458173 620195 458239 620198
rect 462221 620258 462287 620261
rect 487153 620258 487219 620261
rect 462221 620256 464140 620258
rect 462221 620200 462226 620256
rect 462282 620200 464140 620256
rect 462221 620198 464140 620200
rect 484932 620256 487219 620258
rect 484932 620200 487158 620256
rect 487214 620200 487219 620256
rect 484932 620198 487219 620200
rect 462221 620195 462287 620198
rect 487153 620195 487219 620198
rect 489821 620258 489887 620261
rect 514753 620258 514819 620261
rect 489821 620256 492108 620258
rect 489821 620200 489826 620256
rect 489882 620200 492108 620256
rect 489821 620198 492108 620200
rect 512900 620256 514819 620258
rect 512900 620200 514758 620256
rect 514814 620200 514819 620256
rect 512900 620198 514819 620200
rect 489821 620195 489887 620198
rect 514753 620195 514819 620198
rect 518801 620258 518867 620261
rect 542353 620258 542419 620261
rect 518801 620256 520076 620258
rect 518801 620200 518806 620256
rect 518862 620200 520076 620256
rect 518801 620198 520076 620200
rect 540868 620256 542419 620258
rect 540868 620200 542358 620256
rect 542414 620200 542419 620256
rect 540868 620198 542419 620200
rect 518801 620195 518867 620198
rect 542353 620195 542419 620198
rect 546401 620258 546467 620261
rect 571333 620258 571399 620261
rect 546401 620256 548044 620258
rect 546401 620200 546406 620256
rect 546462 620200 548044 620256
rect 546401 620198 548044 620200
rect 568836 620256 571399 620258
rect 568836 620200 571338 620256
rect 571394 620200 571399 620256
rect 568836 620198 571399 620200
rect 546401 620195 546467 620198
rect 571333 620195 571399 620198
rect -960 619020 480 619260
rect 580257 617538 580323 617541
rect 583520 617538 584960 617628
rect 580257 617536 584960 617538
rect 580257 617480 580262 617536
rect 580318 617480 584960 617536
rect 580257 617478 584960 617480
rect 580257 617475 580323 617478
rect 583520 617388 584960 617478
rect 13537 611962 13603 611965
rect 66253 611962 66319 611965
rect 13537 611960 66319 611962
rect 13537 611904 13542 611960
rect 13598 611904 66258 611960
rect 66314 611904 66319 611960
rect 13537 611902 66319 611904
rect 13537 611899 13603 611902
rect 66253 611899 66319 611902
rect 70301 611962 70367 611965
rect 122833 611962 122899 611965
rect 70301 611960 122899 611962
rect 70301 611904 70306 611960
rect 70362 611904 122838 611960
rect 122894 611904 122899 611960
rect 70301 611902 122899 611904
rect 70301 611899 70367 611902
rect 122833 611899 122899 611902
rect 126881 611962 126947 611965
rect 178033 611962 178099 611965
rect 126881 611960 178099 611962
rect 126881 611904 126886 611960
rect 126942 611904 178038 611960
rect 178094 611904 178099 611960
rect 126881 611902 178099 611904
rect 126881 611899 126947 611902
rect 178033 611899 178099 611902
rect 182081 611962 182147 611965
rect 234705 611962 234771 611965
rect 182081 611960 234771 611962
rect 182081 611904 182086 611960
rect 182142 611904 234710 611960
rect 234766 611904 234771 611960
rect 182081 611902 234771 611904
rect 182081 611899 182147 611902
rect 234705 611899 234771 611902
rect 238661 611962 238727 611965
rect 291193 611962 291259 611965
rect 238661 611960 291259 611962
rect 238661 611904 238666 611960
rect 238722 611904 291198 611960
rect 291254 611904 291259 611960
rect 238661 611902 291259 611904
rect 238661 611899 238727 611902
rect 291193 611899 291259 611902
rect 293861 611962 293927 611965
rect 346393 611962 346459 611965
rect 293861 611960 346459 611962
rect 293861 611904 293866 611960
rect 293922 611904 346398 611960
rect 346454 611904 346459 611960
rect 293861 611902 346459 611904
rect 293861 611899 293927 611902
rect 346393 611899 346459 611902
rect 350441 611962 350507 611965
rect 402973 611962 403039 611965
rect 350441 611960 403039 611962
rect 350441 611904 350446 611960
rect 350502 611904 402978 611960
rect 403034 611904 403039 611960
rect 350441 611902 403039 611904
rect 350441 611899 350507 611902
rect 402973 611899 403039 611902
rect 405641 611962 405707 611965
rect 458173 611962 458239 611965
rect 405641 611960 458239 611962
rect 405641 611904 405646 611960
rect 405702 611904 458178 611960
rect 458234 611904 458239 611960
rect 405641 611902 458239 611904
rect 405641 611899 405707 611902
rect 458173 611899 458239 611902
rect 462221 611962 462287 611965
rect 514753 611962 514819 611965
rect 462221 611960 514819 611962
rect 462221 611904 462226 611960
rect 462282 611904 514758 611960
rect 514814 611904 514819 611960
rect 462221 611902 514819 611904
rect 462221 611899 462287 611902
rect 514753 611899 514819 611902
rect 518801 611962 518867 611965
rect 571333 611962 571399 611965
rect 518801 611960 571399 611962
rect 518801 611904 518806 611960
rect 518862 611904 571338 611960
rect 571394 611904 571399 611960
rect 518801 611902 571399 611904
rect 518801 611899 518867 611902
rect 571333 611899 571399 611902
rect 148593 608562 148659 608565
rect 165654 608562 165660 608564
rect 148593 608560 165660 608562
rect 148593 608504 148598 608560
rect 148654 608504 165660 608560
rect 148593 608502 165660 608504
rect 148593 608499 148659 608502
rect 165654 608500 165660 608502
rect 165724 608500 165730 608564
rect 222653 608562 222719 608565
rect 259494 608562 259500 608564
rect 222653 608560 259500 608562
rect 222653 608504 222658 608560
rect 222714 608504 259500 608560
rect 222653 608502 259500 608504
rect 222653 608499 222719 608502
rect 259494 608500 259500 608502
rect 259564 608500 259570 608564
rect 344645 608562 344711 608565
rect 361614 608562 361620 608564
rect 344645 608560 361620 608562
rect 344645 608504 344650 608560
rect 344706 608504 361620 608560
rect 344645 608502 361620 608504
rect 344645 608499 344711 608502
rect 361614 608500 361620 608502
rect 361684 608500 361690 608564
rect 428641 608562 428707 608565
rect 445702 608562 445708 608564
rect 428641 608560 445708 608562
rect 428641 608504 428646 608560
rect 428702 608504 445708 608560
rect 428641 608502 445708 608504
rect 428641 608499 428707 608502
rect 445702 608500 445708 608502
rect 445772 608500 445778 608564
rect 540605 608562 540671 608565
rect 557574 608562 557580 608564
rect 540605 608560 557580 608562
rect 540605 608504 540610 608560
rect 540666 608504 557580 608560
rect 540605 608502 557580 608504
rect 540605 608499 540671 608502
rect 557574 608500 557580 608502
rect 557644 608500 557650 608564
rect -960 606114 480 606204
rect 2773 606114 2839 606117
rect -960 606112 2839 606114
rect -960 606056 2778 606112
rect 2834 606056 2839 606112
rect -960 606054 2839 606056
rect -960 605964 480 606054
rect 2773 606051 2839 606054
rect 583520 604060 584960 604300
rect 128302 603332 128308 603396
rect 128372 603394 128378 603396
rect 128445 603394 128511 603397
rect 194777 603396 194843 603397
rect 194726 603394 194732 603396
rect 128372 603392 128511 603394
rect 128372 603336 128450 603392
rect 128506 603336 128511 603392
rect 128372 603334 128511 603336
rect 194686 603334 194732 603394
rect 194796 603392 194843 603396
rect 194838 603336 194843 603392
rect 128372 603332 128378 603334
rect 128445 603331 128511 603334
rect 194726 603332 194732 603334
rect 194796 603332 194843 603336
rect 194777 603331 194843 603332
rect 390829 603396 390895 603397
rect 390829 603392 390876 603396
rect 390940 603394 390946 603396
rect 390829 603336 390834 603392
rect 390829 603332 390876 603336
rect 390940 603334 390986 603394
rect 390940 603332 390946 603334
rect 390829 603331 390895 603332
rect 238661 602306 238727 602309
rect 288382 602306 288388 602308
rect 238661 602304 288388 602306
rect 238661 602248 238666 602304
rect 238722 602248 288388 602304
rect 238661 602246 288388 602248
rect 238661 602243 238727 602246
rect 288382 602244 288388 602246
rect 288452 602244 288458 602308
rect 434621 602306 434687 602309
rect 484342 602306 484348 602308
rect 434621 602304 484348 602306
rect 434621 602248 434626 602304
rect 434682 602248 484348 602304
rect 434621 602246 484348 602248
rect 434621 602243 434687 602246
rect 484342 602244 484348 602246
rect 484412 602244 484418 602308
rect 42701 602170 42767 602173
rect 92422 602170 92428 602172
rect 42701 602168 92428 602170
rect 42701 602112 42706 602168
rect 42762 602112 92428 602168
rect 42701 602110 92428 602112
rect 42701 602107 42767 602110
rect 92422 602108 92428 602110
rect 92492 602108 92498 602172
rect 97901 602170 97967 602173
rect 148358 602170 148364 602172
rect 97901 602168 148364 602170
rect 97901 602112 97906 602168
rect 97962 602112 148364 602168
rect 97901 602110 148364 602112
rect 97901 602107 97967 602110
rect 148358 602108 148364 602110
rect 148428 602108 148434 602172
rect 154481 602170 154547 602173
rect 207013 602170 207079 602173
rect 154481 602168 207079 602170
rect 154481 602112 154486 602168
rect 154542 602112 207018 602168
rect 207074 602112 207079 602168
rect 154481 602110 207079 602112
rect 154481 602107 154547 602110
rect 207013 602107 207079 602110
rect 209681 602170 209747 602173
rect 260414 602170 260420 602172
rect 209681 602168 260420 602170
rect 209681 602112 209686 602168
rect 209742 602112 260420 602168
rect 209681 602110 260420 602112
rect 209681 602107 209747 602110
rect 260414 602108 260420 602110
rect 260484 602108 260490 602172
rect 293861 602170 293927 602173
rect 344318 602170 344324 602172
rect 293861 602168 344324 602170
rect 293861 602112 293866 602168
rect 293922 602112 344324 602168
rect 293861 602110 344324 602112
rect 293861 602107 293927 602110
rect 344318 602108 344324 602110
rect 344388 602108 344394 602172
rect 350441 602170 350507 602173
rect 402973 602170 403039 602173
rect 350441 602168 403039 602170
rect 350441 602112 350446 602168
rect 350502 602112 402978 602168
rect 403034 602112 403039 602168
rect 350441 602110 403039 602112
rect 350441 602107 350507 602110
rect 402973 602107 403039 602110
rect 405641 602170 405707 602173
rect 456374 602170 456380 602172
rect 405641 602168 456380 602170
rect 405641 602112 405646 602168
rect 405702 602112 456380 602168
rect 405641 602110 456380 602112
rect 405641 602107 405707 602110
rect 456374 602108 456380 602110
rect 456444 602108 456450 602172
rect 492806 602108 492812 602172
rect 492876 602170 492882 602172
rect 542353 602170 542419 602173
rect 492876 602168 542419 602170
rect 492876 602112 542358 602168
rect 542414 602112 542419 602168
rect 492876 602110 542419 602112
rect 492876 602108 492882 602110
rect 542353 602107 542419 602110
rect 13537 602034 13603 602037
rect 64454 602034 64460 602036
rect 13537 602032 64460 602034
rect 13537 601976 13542 602032
rect 13598 601976 64460 602032
rect 13537 601974 64460 601976
rect 13537 601971 13603 601974
rect 64454 601972 64460 601974
rect 64524 601972 64530 602036
rect 70301 602034 70367 602037
rect 122833 602034 122899 602037
rect 70301 602032 122899 602034
rect 70301 601976 70306 602032
rect 70362 601976 122838 602032
rect 122894 601976 122899 602032
rect 70301 601974 122899 601976
rect 70301 601971 70367 601974
rect 122833 601971 122899 601974
rect 126881 602034 126947 602037
rect 176326 602034 176332 602036
rect 126881 602032 176332 602034
rect 126881 601976 126886 602032
rect 126942 601976 176332 602032
rect 126881 601974 176332 601976
rect 126881 601971 126947 601974
rect 176326 601972 176332 601974
rect 176396 601972 176402 602036
rect 182081 602034 182147 602037
rect 234705 602034 234771 602037
rect 182081 602032 234771 602034
rect 182081 601976 182086 602032
rect 182142 601976 234710 602032
rect 234766 601976 234771 602032
rect 182081 601974 234771 601976
rect 182081 601971 182147 601974
rect 234705 601971 234771 601974
rect 266261 602034 266327 602037
rect 318793 602034 318859 602037
rect 266261 602032 318859 602034
rect 266261 601976 266266 602032
rect 266322 601976 318798 602032
rect 318854 601976 318859 602032
rect 266261 601974 318859 601976
rect 266261 601971 266327 601974
rect 318793 601971 318859 601974
rect 322841 602034 322907 602037
rect 372286 602034 372292 602036
rect 322841 602032 372292 602034
rect 322841 601976 322846 602032
rect 322902 601976 372292 602032
rect 322841 601974 372292 601976
rect 322841 601971 322907 601974
rect 372286 601972 372292 601974
rect 372356 601972 372362 602036
rect 378041 602034 378107 602037
rect 430573 602034 430639 602037
rect 378041 602032 430639 602034
rect 378041 601976 378046 602032
rect 378102 601976 430578 602032
rect 430634 601976 430639 602032
rect 378041 601974 430639 601976
rect 378041 601971 378107 601974
rect 430573 601971 430639 601974
rect 462221 602034 462287 602037
rect 514753 602034 514819 602037
rect 462221 602032 514819 602034
rect 462221 601976 462226 602032
rect 462282 601976 514758 602032
rect 514814 601976 514819 602032
rect 462221 601974 514819 601976
rect 462221 601971 462287 601974
rect 514753 601971 514819 601974
rect 520590 601972 520596 602036
rect 520660 602034 520666 602036
rect 571333 602034 571399 602037
rect 520660 602032 571399 602034
rect 520660 601976 571338 602032
rect 571394 601976 571399 602032
rect 520660 601974 571399 601976
rect 520660 601972 520666 601974
rect 571333 601971 571399 601974
rect 64454 594220 64460 594284
rect 64524 594220 64530 594284
rect 92422 594220 92428 594284
rect 92492 594220 92498 594284
rect 148358 594220 148364 594284
rect 148428 594220 148434 594284
rect 176326 594220 176332 594284
rect 176396 594220 176402 594284
rect 260414 594220 260420 594284
rect 260484 594220 260490 594284
rect 288382 594220 288388 594284
rect 288452 594220 288458 594284
rect 344318 594220 344324 594284
rect 344388 594220 344394 594284
rect 372286 594220 372292 594284
rect 372356 594220 372362 594284
rect 456374 594220 456380 594284
rect 456444 594220 456450 594284
rect 484342 594220 484348 594284
rect 484412 594220 484418 594284
rect 492622 594220 492628 594284
rect 492692 594220 492698 594284
rect 520590 594220 520596 594284
rect 520660 594220 520666 594284
rect 13537 593738 13603 593741
rect 38653 593738 38719 593741
rect 13537 593736 16100 593738
rect 13537 593680 13542 593736
rect 13598 593680 16100 593736
rect 13537 593678 16100 593680
rect 36892 593736 38719 593738
rect 36892 593680 38658 593736
rect 38714 593680 38719 593736
rect 36892 593678 38719 593680
rect 13537 593675 13603 593678
rect 38653 593675 38719 593678
rect 42701 593738 42767 593741
rect 42701 593736 44068 593738
rect 42701 593680 42706 593736
rect 42762 593680 44068 593736
rect 64462 593708 64522 594220
rect 70301 593738 70367 593741
rect 70301 593736 72036 593738
rect 42701 593678 44068 593680
rect 70301 593680 70306 593736
rect 70362 593680 72036 593736
rect 92430 593708 92490 594220
rect 97901 593738 97967 593741
rect 122833 593738 122899 593741
rect 97901 593736 100188 593738
rect 70301 593678 72036 593680
rect 97901 593680 97906 593736
rect 97962 593680 100188 593736
rect 97901 593678 100188 593680
rect 120796 593736 122899 593738
rect 120796 593680 122838 593736
rect 122894 593680 122899 593736
rect 120796 593678 122899 593680
rect 42701 593675 42767 593678
rect 70301 593675 70367 593678
rect 97901 593675 97967 593678
rect 122833 593675 122899 593678
rect 126881 593738 126947 593741
rect 126881 593736 128156 593738
rect 126881 593680 126886 593736
rect 126942 593680 128156 593736
rect 148366 593708 148426 594220
rect 154481 593738 154547 593741
rect 154481 593736 156124 593738
rect 126881 593678 128156 593680
rect 154481 593680 154486 593736
rect 154542 593680 156124 593736
rect 176334 593708 176394 594220
rect 182081 593738 182147 593741
rect 207013 593738 207079 593741
rect 182081 593736 184092 593738
rect 154481 593678 156124 593680
rect 182081 593680 182086 593736
rect 182142 593680 184092 593736
rect 182081 593678 184092 593680
rect 204884 593736 207079 593738
rect 204884 593680 207018 593736
rect 207074 593680 207079 593736
rect 204884 593678 207079 593680
rect 126881 593675 126947 593678
rect 154481 593675 154547 593678
rect 182081 593675 182147 593678
rect 207013 593675 207079 593678
rect 209681 593738 209747 593741
rect 234705 593738 234771 593741
rect 209681 593736 212060 593738
rect 209681 593680 209686 593736
rect 209742 593680 212060 593736
rect 209681 593678 212060 593680
rect 232852 593736 234771 593738
rect 232852 593680 234710 593736
rect 234766 593680 234771 593736
rect 232852 593678 234771 593680
rect 209681 593675 209747 593678
rect 234705 593675 234771 593678
rect 238661 593738 238727 593741
rect 238661 593736 240212 593738
rect 238661 593680 238666 593736
rect 238722 593680 240212 593736
rect 260422 593708 260482 594220
rect 266261 593738 266327 593741
rect 266261 593736 268180 593738
rect 238661 593678 240212 593680
rect 266261 593680 266266 593736
rect 266322 593680 268180 593736
rect 288390 593708 288450 594220
rect 293861 593738 293927 593741
rect 318793 593738 318859 593741
rect 293861 593736 296148 593738
rect 266261 593678 268180 593680
rect 293861 593680 293866 593736
rect 293922 593680 296148 593736
rect 293861 593678 296148 593680
rect 316940 593736 318859 593738
rect 316940 593680 318798 593736
rect 318854 593680 318859 593736
rect 316940 593678 318859 593680
rect 238661 593675 238727 593678
rect 266261 593675 266327 593678
rect 293861 593675 293927 593678
rect 318793 593675 318859 593678
rect 322841 593738 322907 593741
rect 322841 593736 324116 593738
rect 322841 593680 322846 593736
rect 322902 593680 324116 593736
rect 344326 593708 344386 594220
rect 350441 593738 350507 593741
rect 350441 593736 352084 593738
rect 322841 593678 324116 593680
rect 350441 593680 350446 593736
rect 350502 593680 352084 593736
rect 372294 593708 372354 594220
rect 378041 593738 378107 593741
rect 402973 593738 403039 593741
rect 378041 593736 380052 593738
rect 350441 593678 352084 593680
rect 378041 593680 378046 593736
rect 378102 593680 380052 593736
rect 378041 593678 380052 593680
rect 400844 593736 403039 593738
rect 400844 593680 402978 593736
rect 403034 593680 403039 593736
rect 400844 593678 403039 593680
rect 322841 593675 322907 593678
rect 350441 593675 350507 593678
rect 378041 593675 378107 593678
rect 402973 593675 403039 593678
rect 405641 593738 405707 593741
rect 430573 593738 430639 593741
rect 405641 593736 408204 593738
rect 405641 593680 405646 593736
rect 405702 593680 408204 593736
rect 405641 593678 408204 593680
rect 428812 593736 430639 593738
rect 428812 593680 430578 593736
rect 430634 593680 430639 593736
rect 428812 593678 430639 593680
rect 405641 593675 405707 593678
rect 430573 593675 430639 593678
rect 434621 593738 434687 593741
rect 434621 593736 436172 593738
rect 434621 593680 434626 593736
rect 434682 593680 436172 593736
rect 456382 593708 456442 594220
rect 462221 593738 462287 593741
rect 462221 593736 464140 593738
rect 434621 593678 436172 593680
rect 462221 593680 462226 593736
rect 462282 593680 464140 593736
rect 484350 593708 484410 594220
rect 492630 593708 492690 594220
rect 514753 593738 514819 593741
rect 512900 593736 514819 593738
rect 462221 593678 464140 593680
rect 512900 593680 514758 593736
rect 514814 593680 514819 593736
rect 520598 593708 520658 594220
rect 542353 593738 542419 593741
rect 540868 593736 542419 593738
rect 512900 593678 514819 593680
rect 540868 593680 542358 593736
rect 542414 593680 542419 593736
rect 540868 593678 542419 593680
rect 434621 593675 434687 593678
rect 462221 593675 462287 593678
rect 514753 593675 514819 593678
rect 542353 593675 542419 593678
rect 546401 593738 546467 593741
rect 571333 593738 571399 593741
rect 546401 593736 548044 593738
rect 546401 593680 546406 593736
rect 546462 593680 548044 593736
rect 546401 593678 548044 593680
rect 568836 593736 571399 593738
rect 568836 593680 571338 593736
rect 571394 593680 571399 593736
rect 568836 593678 571399 593680
rect 546401 593675 546467 593678
rect 571333 593675 571399 593678
rect -960 592908 480 593148
rect 580349 591018 580415 591021
rect 583520 591018 584960 591108
rect 580349 591016 584960 591018
rect 580349 590960 580354 591016
rect 580410 590960 584960 591016
rect 580349 590958 584960 590960
rect 580349 590955 580415 590958
rect 583520 590868 584960 590958
rect 110597 580954 110663 580957
rect 128118 580954 128124 580956
rect 110597 580952 128124 580954
rect 110597 580896 110602 580952
rect 110658 580896 128124 580952
rect 110597 580894 128124 580896
rect 110597 580891 110663 580894
rect 128118 580892 128124 580894
rect 128188 580892 128194 580956
rect 156321 580954 156387 580957
rect 194726 580954 194732 580956
rect 156321 580952 194732 580954
rect 156321 580896 156326 580952
rect 156382 580896 194732 580952
rect 156321 580894 194732 580896
rect 156321 580891 156387 580894
rect 194726 580892 194732 580894
rect 194796 580892 194802 580956
rect 352649 580954 352715 580957
rect 390870 580954 390876 580956
rect 352649 580952 390876 580954
rect 352649 580896 352654 580952
rect 352710 580896 390876 580952
rect 352649 580894 390876 580896
rect 352649 580891 352715 580894
rect 390870 580892 390876 580894
rect 390940 580892 390946 580956
rect -960 580002 480 580092
rect 3509 580002 3575 580005
rect -960 580000 3575 580002
rect -960 579944 3514 580000
rect 3570 579944 3575 580000
rect -960 579942 3575 579944
rect -960 579852 480 579942
rect 3509 579939 3575 579942
rect 583520 577540 584960 577780
rect 165654 576404 165660 576468
rect 165724 576466 165730 576468
rect 165981 576466 166047 576469
rect 165724 576464 166047 576466
rect 165724 576408 165986 576464
rect 166042 576408 166047 576464
rect 165724 576406 166047 576408
rect 165724 576404 165730 576406
rect 165981 576403 166047 576406
rect 259494 576404 259500 576468
rect 259564 576466 259570 576468
rect 260373 576466 260439 576469
rect 259564 576464 260439 576466
rect 259564 576408 260378 576464
rect 260434 576408 260439 576464
rect 259564 576406 260439 576408
rect 259564 576404 259570 576406
rect 260373 576403 260439 576406
rect 361614 576404 361620 576468
rect 361684 576466 361690 576468
rect 361941 576466 362007 576469
rect 361684 576464 362007 576466
rect 361684 576408 361946 576464
rect 362002 576408 362007 576464
rect 361684 576406 362007 576408
rect 361684 576404 361690 576406
rect 361941 576403 362007 576406
rect 445702 576404 445708 576468
rect 445772 576466 445778 576468
rect 446029 576466 446095 576469
rect 445772 576464 446095 576466
rect 445772 576408 446034 576464
rect 446090 576408 446095 576464
rect 445772 576406 446095 576408
rect 445772 576404 445778 576406
rect 446029 576403 446095 576406
rect 557574 576404 557580 576468
rect 557644 576466 557650 576468
rect 557993 576466 558059 576469
rect 557644 576464 558059 576466
rect 557644 576408 557998 576464
rect 558054 576408 558059 576464
rect 557644 576406 558059 576408
rect 557644 576404 557650 576406
rect 557993 576403 558059 576406
rect 13537 574698 13603 574701
rect 66253 574698 66319 574701
rect 13537 574696 66319 574698
rect 13537 574640 13542 574696
rect 13598 574640 66258 574696
rect 66314 574640 66319 574696
rect 13537 574638 66319 574640
rect 13537 574635 13603 574638
rect 66253 574635 66319 574638
rect 70301 574698 70367 574701
rect 122833 574698 122899 574701
rect 70301 574696 122899 574698
rect 70301 574640 70306 574696
rect 70362 574640 122838 574696
rect 122894 574640 122899 574696
rect 70301 574638 122899 574640
rect 70301 574635 70367 574638
rect 122833 574635 122899 574638
rect 126881 574698 126947 574701
rect 178033 574698 178099 574701
rect 126881 574696 178099 574698
rect 126881 574640 126886 574696
rect 126942 574640 178038 574696
rect 178094 574640 178099 574696
rect 126881 574638 178099 574640
rect 126881 574635 126947 574638
rect 178033 574635 178099 574638
rect 182081 574698 182147 574701
rect 234705 574698 234771 574701
rect 182081 574696 234771 574698
rect 182081 574640 182086 574696
rect 182142 574640 234710 574696
rect 234766 574640 234771 574696
rect 182081 574638 234771 574640
rect 182081 574635 182147 574638
rect 234705 574635 234771 574638
rect 238661 574698 238727 574701
rect 291193 574698 291259 574701
rect 238661 574696 291259 574698
rect 238661 574640 238666 574696
rect 238722 574640 291198 574696
rect 291254 574640 291259 574696
rect 238661 574638 291259 574640
rect 238661 574635 238727 574638
rect 291193 574635 291259 574638
rect 293861 574698 293927 574701
rect 346393 574698 346459 574701
rect 293861 574696 346459 574698
rect 293861 574640 293866 574696
rect 293922 574640 346398 574696
rect 346454 574640 346459 574696
rect 293861 574638 346459 574640
rect 293861 574635 293927 574638
rect 346393 574635 346459 574638
rect 350441 574698 350507 574701
rect 402973 574698 403039 574701
rect 350441 574696 403039 574698
rect 350441 574640 350446 574696
rect 350502 574640 402978 574696
rect 403034 574640 403039 574696
rect 350441 574638 403039 574640
rect 350441 574635 350507 574638
rect 402973 574635 403039 574638
rect 405641 574698 405707 574701
rect 458173 574698 458239 574701
rect 405641 574696 458239 574698
rect 405641 574640 405646 574696
rect 405702 574640 458178 574696
rect 458234 574640 458239 574696
rect 405641 574638 458239 574640
rect 405641 574635 405707 574638
rect 458173 574635 458239 574638
rect 462221 574698 462287 574701
rect 514753 574698 514819 574701
rect 462221 574696 514819 574698
rect 462221 574640 462226 574696
rect 462282 574640 514758 574696
rect 514814 574640 514819 574696
rect 462221 574638 514819 574640
rect 462221 574635 462287 574638
rect 514753 574635 514819 574638
rect 518801 574698 518867 574701
rect 571333 574698 571399 574701
rect 518801 574696 571399 574698
rect 518801 574640 518806 574696
rect 518862 574640 571338 574696
rect 571394 574640 571399 574696
rect 518801 574638 571399 574640
rect 518801 574635 518867 574638
rect 571333 574635 571399 574638
rect -960 566796 480 567036
rect 13537 566266 13603 566269
rect 38653 566266 38719 566269
rect 13537 566264 16100 566266
rect 13537 566208 13542 566264
rect 13598 566208 16100 566264
rect 13537 566206 16100 566208
rect 36892 566264 38719 566266
rect 36892 566208 38658 566264
rect 38714 566208 38719 566264
rect 36892 566206 38719 566208
rect 13537 566203 13603 566206
rect 38653 566203 38719 566206
rect 42701 566266 42767 566269
rect 66253 566266 66319 566269
rect 42701 566264 44068 566266
rect 42701 566208 42706 566264
rect 42762 566208 44068 566264
rect 42701 566206 44068 566208
rect 64860 566264 66319 566266
rect 64860 566208 66258 566264
rect 66314 566208 66319 566264
rect 64860 566206 66319 566208
rect 42701 566203 42767 566206
rect 66253 566203 66319 566206
rect 70301 566266 70367 566269
rect 95233 566266 95299 566269
rect 70301 566264 72036 566266
rect 70301 566208 70306 566264
rect 70362 566208 72036 566264
rect 70301 566206 72036 566208
rect 92828 566264 95299 566266
rect 92828 566208 95238 566264
rect 95294 566208 95299 566264
rect 92828 566206 95299 566208
rect 70301 566203 70367 566206
rect 95233 566203 95299 566206
rect 97901 566266 97967 566269
rect 122833 566266 122899 566269
rect 97901 566264 100188 566266
rect 97901 566208 97906 566264
rect 97962 566208 100188 566264
rect 97901 566206 100188 566208
rect 120796 566264 122899 566266
rect 120796 566208 122838 566264
rect 122894 566208 122899 566264
rect 120796 566206 122899 566208
rect 97901 566203 97967 566206
rect 122833 566203 122899 566206
rect 126881 566266 126947 566269
rect 150433 566266 150499 566269
rect 126881 566264 128156 566266
rect 126881 566208 126886 566264
rect 126942 566208 128156 566264
rect 126881 566206 128156 566208
rect 148948 566264 150499 566266
rect 148948 566208 150438 566264
rect 150494 566208 150499 566264
rect 148948 566206 150499 566208
rect 126881 566203 126947 566206
rect 150433 566203 150499 566206
rect 154481 566266 154547 566269
rect 178033 566266 178099 566269
rect 154481 566264 156124 566266
rect 154481 566208 154486 566264
rect 154542 566208 156124 566264
rect 154481 566206 156124 566208
rect 176916 566264 178099 566266
rect 176916 566208 178038 566264
rect 178094 566208 178099 566264
rect 176916 566206 178099 566208
rect 154481 566203 154547 566206
rect 178033 566203 178099 566206
rect 182081 566266 182147 566269
rect 207013 566266 207079 566269
rect 182081 566264 184092 566266
rect 182081 566208 182086 566264
rect 182142 566208 184092 566264
rect 182081 566206 184092 566208
rect 204884 566264 207079 566266
rect 204884 566208 207018 566264
rect 207074 566208 207079 566264
rect 204884 566206 207079 566208
rect 182081 566203 182147 566206
rect 207013 566203 207079 566206
rect 209681 566266 209747 566269
rect 234705 566266 234771 566269
rect 209681 566264 212060 566266
rect 209681 566208 209686 566264
rect 209742 566208 212060 566264
rect 209681 566206 212060 566208
rect 232852 566264 234771 566266
rect 232852 566208 234710 566264
rect 234766 566208 234771 566264
rect 232852 566206 234771 566208
rect 209681 566203 209747 566206
rect 234705 566203 234771 566206
rect 238661 566266 238727 566269
rect 262213 566266 262279 566269
rect 238661 566264 240212 566266
rect 238661 566208 238666 566264
rect 238722 566208 240212 566264
rect 238661 566206 240212 566208
rect 260820 566264 262279 566266
rect 260820 566208 262218 566264
rect 262274 566208 262279 566264
rect 260820 566206 262279 566208
rect 238661 566203 238727 566206
rect 262213 566203 262279 566206
rect 266261 566266 266327 566269
rect 291193 566266 291259 566269
rect 266261 566264 268180 566266
rect 266261 566208 266266 566264
rect 266322 566208 268180 566264
rect 266261 566206 268180 566208
rect 288788 566264 291259 566266
rect 288788 566208 291198 566264
rect 291254 566208 291259 566264
rect 288788 566206 291259 566208
rect 266261 566203 266327 566206
rect 291193 566203 291259 566206
rect 293861 566266 293927 566269
rect 318793 566266 318859 566269
rect 293861 566264 296148 566266
rect 293861 566208 293866 566264
rect 293922 566208 296148 566264
rect 293861 566206 296148 566208
rect 316940 566264 318859 566266
rect 316940 566208 318798 566264
rect 318854 566208 318859 566264
rect 316940 566206 318859 566208
rect 293861 566203 293927 566206
rect 318793 566203 318859 566206
rect 322841 566266 322907 566269
rect 346393 566266 346459 566269
rect 322841 566264 324116 566266
rect 322841 566208 322846 566264
rect 322902 566208 324116 566264
rect 322841 566206 324116 566208
rect 344908 566264 346459 566266
rect 344908 566208 346398 566264
rect 346454 566208 346459 566264
rect 344908 566206 346459 566208
rect 322841 566203 322907 566206
rect 346393 566203 346459 566206
rect 350441 566266 350507 566269
rect 375373 566266 375439 566269
rect 350441 566264 352084 566266
rect 350441 566208 350446 566264
rect 350502 566208 352084 566264
rect 350441 566206 352084 566208
rect 372876 566264 375439 566266
rect 372876 566208 375378 566264
rect 375434 566208 375439 566264
rect 372876 566206 375439 566208
rect 350441 566203 350507 566206
rect 375373 566203 375439 566206
rect 378041 566266 378107 566269
rect 402973 566266 403039 566269
rect 378041 566264 380052 566266
rect 378041 566208 378046 566264
rect 378102 566208 380052 566264
rect 378041 566206 380052 566208
rect 400844 566264 403039 566266
rect 400844 566208 402978 566264
rect 403034 566208 403039 566264
rect 400844 566206 403039 566208
rect 378041 566203 378107 566206
rect 402973 566203 403039 566206
rect 405641 566266 405707 566269
rect 430573 566266 430639 566269
rect 405641 566264 408204 566266
rect 405641 566208 405646 566264
rect 405702 566208 408204 566264
rect 405641 566206 408204 566208
rect 428812 566264 430639 566266
rect 428812 566208 430578 566264
rect 430634 566208 430639 566264
rect 428812 566206 430639 566208
rect 405641 566203 405707 566206
rect 430573 566203 430639 566206
rect 434621 566266 434687 566269
rect 458173 566266 458239 566269
rect 434621 566264 436172 566266
rect 434621 566208 434626 566264
rect 434682 566208 436172 566264
rect 434621 566206 436172 566208
rect 456964 566264 458239 566266
rect 456964 566208 458178 566264
rect 458234 566208 458239 566264
rect 456964 566206 458239 566208
rect 434621 566203 434687 566206
rect 458173 566203 458239 566206
rect 462221 566266 462287 566269
rect 487153 566266 487219 566269
rect 462221 566264 464140 566266
rect 462221 566208 462226 566264
rect 462282 566208 464140 566264
rect 462221 566206 464140 566208
rect 484932 566264 487219 566266
rect 484932 566208 487158 566264
rect 487214 566208 487219 566264
rect 484932 566206 487219 566208
rect 462221 566203 462287 566206
rect 487153 566203 487219 566206
rect 489821 566266 489887 566269
rect 514753 566266 514819 566269
rect 489821 566264 492108 566266
rect 489821 566208 489826 566264
rect 489882 566208 492108 566264
rect 489821 566206 492108 566208
rect 512900 566264 514819 566266
rect 512900 566208 514758 566264
rect 514814 566208 514819 566264
rect 512900 566206 514819 566208
rect 489821 566203 489887 566206
rect 514753 566203 514819 566206
rect 518801 566266 518867 566269
rect 542353 566266 542419 566269
rect 518801 566264 520076 566266
rect 518801 566208 518806 566264
rect 518862 566208 520076 566264
rect 518801 566206 520076 566208
rect 540868 566264 542419 566266
rect 540868 566208 542358 566264
rect 542414 566208 542419 566264
rect 540868 566206 542419 566208
rect 518801 566203 518867 566206
rect 542353 566203 542419 566206
rect 546401 566266 546467 566269
rect 571333 566266 571399 566269
rect 546401 566264 548044 566266
rect 546401 566208 546406 566264
rect 546462 566208 548044 566264
rect 546401 566206 548044 566208
rect 568836 566264 571399 566266
rect 568836 566208 571338 566264
rect 571394 566208 571399 566264
rect 568836 566206 571399 566208
rect 546401 566203 546467 566206
rect 571333 566203 571399 566206
rect 580441 564362 580507 564365
rect 583520 564362 584960 564452
rect 580441 564360 584960 564362
rect 580441 564304 580446 564360
rect 580502 564304 584960 564360
rect 580441 564302 584960 564304
rect 580441 564299 580507 564302
rect 583520 564212 584960 564302
rect 148593 554706 148659 554709
rect 165654 554706 165660 554708
rect 148593 554704 165660 554706
rect 148593 554648 148598 554704
rect 148654 554648 165660 554704
rect 148593 554646 165660 554648
rect 148593 554643 148659 554646
rect 165654 554644 165660 554646
rect 165724 554644 165730 554708
rect 222653 554706 222719 554709
rect 259494 554706 259500 554708
rect 222653 554704 259500 554706
rect 222653 554648 222658 554704
rect 222714 554648 259500 554704
rect 222653 554646 259500 554648
rect 222653 554643 222719 554646
rect 259494 554644 259500 554646
rect 259564 554644 259570 554708
rect 344645 554706 344711 554709
rect 361614 554706 361620 554708
rect 344645 554704 361620 554706
rect 344645 554648 344650 554704
rect 344706 554648 361620 554704
rect 344645 554646 361620 554648
rect 344645 554643 344711 554646
rect 361614 554644 361620 554646
rect 361684 554644 361690 554708
rect 428641 554706 428707 554709
rect 445702 554706 445708 554708
rect 428641 554704 445708 554706
rect 428641 554648 428646 554704
rect 428702 554648 445708 554704
rect 428641 554646 445708 554648
rect 428641 554643 428707 554646
rect 445702 554644 445708 554646
rect 445772 554644 445778 554708
rect 540605 554706 540671 554709
rect 557574 554706 557580 554708
rect 540605 554704 557580 554706
rect 540605 554648 540610 554704
rect 540666 554648 557580 554704
rect 540605 554646 557580 554648
rect 540605 554643 540671 554646
rect 557574 554644 557580 554646
rect 557644 554644 557650 554708
rect -960 553890 480 553980
rect 3601 553890 3667 553893
rect -960 553888 3667 553890
rect -960 553832 3606 553888
rect 3662 553832 3667 553888
rect -960 553830 3667 553832
rect -960 553740 480 553830
rect 3601 553827 3667 553830
rect 583520 551020 584960 551260
rect 128302 549340 128308 549404
rect 128372 549402 128378 549404
rect 128445 549402 128511 549405
rect 194777 549404 194843 549405
rect 194726 549402 194732 549404
rect 128372 549400 128511 549402
rect 128372 549344 128450 549400
rect 128506 549344 128511 549400
rect 128372 549342 128511 549344
rect 194686 549342 194732 549402
rect 194796 549400 194843 549404
rect 194838 549344 194843 549400
rect 128372 549340 128378 549342
rect 128445 549339 128511 549342
rect 194726 549340 194732 549342
rect 194796 549340 194843 549344
rect 194777 549339 194843 549340
rect 390829 549404 390895 549405
rect 390829 549400 390876 549404
rect 390940 549402 390946 549404
rect 390829 549344 390834 549400
rect 390829 549340 390876 549344
rect 390940 549342 390986 549402
rect 390940 549340 390946 549342
rect 390829 549339 390895 549340
rect 238661 548314 238727 548317
rect 288382 548314 288388 548316
rect 238661 548312 288388 548314
rect 238661 548256 238666 548312
rect 238722 548256 288388 548312
rect 238661 548254 288388 548256
rect 238661 548251 238727 548254
rect 288382 548252 288388 548254
rect 288452 548252 288458 548316
rect 322841 548314 322907 548317
rect 372286 548314 372292 548316
rect 322841 548312 372292 548314
rect 322841 548256 322846 548312
rect 322902 548256 372292 548312
rect 322841 548254 372292 548256
rect 322841 548251 322907 548254
rect 372286 548252 372292 548254
rect 372356 548252 372362 548316
rect 42701 548178 42767 548181
rect 92422 548178 92428 548180
rect 42701 548176 92428 548178
rect 42701 548120 42706 548176
rect 42762 548120 92428 548176
rect 42701 548118 92428 548120
rect 42701 548115 42767 548118
rect 92422 548116 92428 548118
rect 92492 548116 92498 548180
rect 97901 548178 97967 548181
rect 148358 548178 148364 548180
rect 97901 548176 148364 548178
rect 97901 548120 97906 548176
rect 97962 548120 148364 548176
rect 97901 548118 148364 548120
rect 97901 548115 97967 548118
rect 148358 548116 148364 548118
rect 148428 548116 148434 548180
rect 154481 548178 154547 548181
rect 207013 548178 207079 548181
rect 154481 548176 207079 548178
rect 154481 548120 154486 548176
rect 154542 548120 207018 548176
rect 207074 548120 207079 548176
rect 154481 548118 207079 548120
rect 154481 548115 154547 548118
rect 207013 548115 207079 548118
rect 212574 548116 212580 548180
rect 212644 548178 212650 548180
rect 262213 548178 262279 548181
rect 212644 548176 262279 548178
rect 212644 548120 262218 548176
rect 262274 548120 262279 548176
rect 212644 548118 262279 548120
rect 212644 548116 212650 548118
rect 262213 548115 262279 548118
rect 296846 548116 296852 548180
rect 296916 548178 296922 548180
rect 346393 548178 346459 548181
rect 296916 548176 346459 548178
rect 296916 548120 346398 548176
rect 346454 548120 346459 548176
rect 296916 548118 346459 548120
rect 296916 548116 296922 548118
rect 346393 548115 346459 548118
rect 378041 548178 378107 548181
rect 430573 548178 430639 548181
rect 378041 548176 430639 548178
rect 378041 548120 378046 548176
rect 378102 548120 430578 548176
rect 430634 548120 430639 548176
rect 378041 548118 430639 548120
rect 378041 548115 378107 548118
rect 430573 548115 430639 548118
rect 434621 548178 434687 548181
rect 484342 548178 484348 548180
rect 434621 548176 484348 548178
rect 434621 548120 434626 548176
rect 434682 548120 484348 548176
rect 434621 548118 484348 548120
rect 434621 548115 434687 548118
rect 484342 548116 484348 548118
rect 484412 548116 484418 548180
rect 489821 548178 489887 548181
rect 540462 548178 540468 548180
rect 489821 548176 540468 548178
rect 489821 548120 489826 548176
rect 489882 548120 540468 548176
rect 489821 548118 540468 548120
rect 489821 548115 489887 548118
rect 540462 548116 540468 548118
rect 540532 548116 540538 548180
rect 13537 548042 13603 548045
rect 64454 548042 64460 548044
rect 13537 548040 64460 548042
rect 13537 547984 13542 548040
rect 13598 547984 64460 548040
rect 13537 547982 64460 547984
rect 13537 547979 13603 547982
rect 64454 547980 64460 547982
rect 64524 547980 64530 548044
rect 70301 548042 70367 548045
rect 122833 548042 122899 548045
rect 70301 548040 122899 548042
rect 70301 547984 70306 548040
rect 70362 547984 122838 548040
rect 122894 547984 122899 548040
rect 70301 547982 122899 547984
rect 70301 547979 70367 547982
rect 122833 547979 122899 547982
rect 126881 548042 126947 548045
rect 176326 548042 176332 548044
rect 126881 548040 176332 548042
rect 126881 547984 126886 548040
rect 126942 547984 176332 548040
rect 126881 547982 176332 547984
rect 126881 547979 126947 547982
rect 176326 547980 176332 547982
rect 176396 547980 176402 548044
rect 182081 548042 182147 548045
rect 234705 548042 234771 548045
rect 182081 548040 234771 548042
rect 182081 547984 182086 548040
rect 182142 547984 234710 548040
rect 234766 547984 234771 548040
rect 182081 547982 234771 547984
rect 182081 547979 182147 547982
rect 234705 547979 234771 547982
rect 266261 548042 266327 548045
rect 318793 548042 318859 548045
rect 266261 548040 318859 548042
rect 266261 547984 266266 548040
rect 266322 547984 318798 548040
rect 318854 547984 318859 548040
rect 266261 547982 318859 547984
rect 266261 547979 266327 547982
rect 318793 547979 318859 547982
rect 350441 548042 350507 548045
rect 402973 548042 403039 548045
rect 350441 548040 403039 548042
rect 350441 547984 350446 548040
rect 350502 547984 402978 548040
rect 403034 547984 403039 548040
rect 350441 547982 403039 547984
rect 350441 547979 350507 547982
rect 402973 547979 403039 547982
rect 408534 547980 408540 548044
rect 408604 548042 408610 548044
rect 458173 548042 458239 548045
rect 408604 548040 458239 548042
rect 408604 547984 458178 548040
rect 458234 547984 458239 548040
rect 408604 547982 458239 547984
rect 408604 547980 408610 547982
rect 458173 547979 458239 547982
rect 462221 548042 462287 548045
rect 514753 548042 514819 548045
rect 462221 548040 514819 548042
rect 462221 547984 462226 548040
rect 462282 547984 514758 548040
rect 514814 547984 514819 548040
rect 462221 547982 514819 547984
rect 462221 547979 462287 547982
rect 514753 547979 514819 547982
rect 520590 547980 520596 548044
rect 520660 548042 520666 548044
rect 571333 548042 571399 548045
rect 520660 548040 571399 548042
rect 520660 547984 571338 548040
rect 571394 547984 571399 548040
rect 520660 547982 571399 547984
rect 520660 547980 520666 547982
rect 571333 547979 571399 547982
rect -960 540684 480 540924
rect 64454 540228 64460 540292
rect 64524 540228 64530 540292
rect 92422 540228 92428 540292
rect 92492 540228 92498 540292
rect 148358 540228 148364 540292
rect 148428 540228 148434 540292
rect 176326 540228 176332 540292
rect 176396 540228 176402 540292
rect 212574 540228 212580 540292
rect 212644 540228 212650 540292
rect 288382 540228 288388 540292
rect 288452 540228 288458 540292
rect 296478 540228 296484 540292
rect 296548 540228 296554 540292
rect 372286 540228 372292 540292
rect 372356 540228 372362 540292
rect 408534 540228 408540 540292
rect 408604 540228 408610 540292
rect 484342 540228 484348 540292
rect 484412 540228 484418 540292
rect 520590 540228 520596 540292
rect 520660 540228 520666 540292
rect 540462 540228 540468 540292
rect 540532 540228 540538 540292
rect 13537 539746 13603 539749
rect 38653 539746 38719 539749
rect 13537 539744 16100 539746
rect 13537 539688 13542 539744
rect 13598 539688 16100 539744
rect 13537 539686 16100 539688
rect 36892 539744 38719 539746
rect 36892 539688 38658 539744
rect 38714 539688 38719 539744
rect 36892 539686 38719 539688
rect 13537 539683 13603 539686
rect 38653 539683 38719 539686
rect 42701 539746 42767 539749
rect 42701 539744 44068 539746
rect 42701 539688 42706 539744
rect 42762 539688 44068 539744
rect 64462 539716 64522 540228
rect 70301 539746 70367 539749
rect 70301 539744 72036 539746
rect 42701 539686 44068 539688
rect 70301 539688 70306 539744
rect 70362 539688 72036 539744
rect 92430 539716 92490 540228
rect 97901 539746 97967 539749
rect 122833 539746 122899 539749
rect 97901 539744 100188 539746
rect 70301 539686 72036 539688
rect 97901 539688 97906 539744
rect 97962 539688 100188 539744
rect 97901 539686 100188 539688
rect 120796 539744 122899 539746
rect 120796 539688 122838 539744
rect 122894 539688 122899 539744
rect 120796 539686 122899 539688
rect 42701 539683 42767 539686
rect 70301 539683 70367 539686
rect 97901 539683 97967 539686
rect 122833 539683 122899 539686
rect 126881 539746 126947 539749
rect 126881 539744 128156 539746
rect 126881 539688 126886 539744
rect 126942 539688 128156 539744
rect 148366 539716 148426 540228
rect 154481 539746 154547 539749
rect 154481 539744 156124 539746
rect 126881 539686 128156 539688
rect 154481 539688 154486 539744
rect 154542 539688 156124 539744
rect 176334 539716 176394 540228
rect 182081 539746 182147 539749
rect 207013 539746 207079 539749
rect 182081 539744 184092 539746
rect 154481 539686 156124 539688
rect 182081 539688 182086 539744
rect 182142 539688 184092 539744
rect 182081 539686 184092 539688
rect 204884 539744 207079 539746
rect 204884 539688 207018 539744
rect 207074 539688 207079 539744
rect 212582 539716 212642 540228
rect 234705 539746 234771 539749
rect 232852 539744 234771 539746
rect 204884 539686 207079 539688
rect 232852 539688 234710 539744
rect 234766 539688 234771 539744
rect 232852 539686 234771 539688
rect 126881 539683 126947 539686
rect 154481 539683 154547 539686
rect 182081 539683 182147 539686
rect 207013 539683 207079 539686
rect 234705 539683 234771 539686
rect 238661 539746 238727 539749
rect 262213 539746 262279 539749
rect 238661 539744 240212 539746
rect 238661 539688 238666 539744
rect 238722 539688 240212 539744
rect 238661 539686 240212 539688
rect 260820 539744 262279 539746
rect 260820 539688 262218 539744
rect 262274 539688 262279 539744
rect 260820 539686 262279 539688
rect 238661 539683 238727 539686
rect 262213 539683 262279 539686
rect 266261 539746 266327 539749
rect 266261 539744 268180 539746
rect 266261 539688 266266 539744
rect 266322 539688 268180 539744
rect 288390 539716 288450 540228
rect 296486 539716 296546 540228
rect 318793 539746 318859 539749
rect 316940 539744 318859 539746
rect 266261 539686 268180 539688
rect 316940 539688 318798 539744
rect 318854 539688 318859 539744
rect 316940 539686 318859 539688
rect 266261 539683 266327 539686
rect 318793 539683 318859 539686
rect 322841 539746 322907 539749
rect 346393 539746 346459 539749
rect 322841 539744 324116 539746
rect 322841 539688 322846 539744
rect 322902 539688 324116 539744
rect 322841 539686 324116 539688
rect 344908 539744 346459 539746
rect 344908 539688 346398 539744
rect 346454 539688 346459 539744
rect 344908 539686 346459 539688
rect 322841 539683 322907 539686
rect 346393 539683 346459 539686
rect 350441 539746 350507 539749
rect 350441 539744 352084 539746
rect 350441 539688 350446 539744
rect 350502 539688 352084 539744
rect 372294 539716 372354 540228
rect 378041 539746 378107 539749
rect 402973 539746 403039 539749
rect 378041 539744 380052 539746
rect 350441 539686 352084 539688
rect 378041 539688 378046 539744
rect 378102 539688 380052 539744
rect 378041 539686 380052 539688
rect 400844 539744 403039 539746
rect 400844 539688 402978 539744
rect 403034 539688 403039 539744
rect 408542 539716 408602 540228
rect 430573 539746 430639 539749
rect 428812 539744 430639 539746
rect 400844 539686 403039 539688
rect 428812 539688 430578 539744
rect 430634 539688 430639 539744
rect 428812 539686 430639 539688
rect 350441 539683 350507 539686
rect 378041 539683 378107 539686
rect 402973 539683 403039 539686
rect 430573 539683 430639 539686
rect 434621 539746 434687 539749
rect 458173 539746 458239 539749
rect 434621 539744 436172 539746
rect 434621 539688 434626 539744
rect 434682 539688 436172 539744
rect 434621 539686 436172 539688
rect 456964 539744 458239 539746
rect 456964 539688 458178 539744
rect 458234 539688 458239 539744
rect 456964 539686 458239 539688
rect 434621 539683 434687 539686
rect 458173 539683 458239 539686
rect 462221 539746 462287 539749
rect 462221 539744 464140 539746
rect 462221 539688 462226 539744
rect 462282 539688 464140 539744
rect 484350 539716 484410 540228
rect 489821 539746 489887 539749
rect 514753 539746 514819 539749
rect 489821 539744 492108 539746
rect 462221 539686 464140 539688
rect 489821 539688 489826 539744
rect 489882 539688 492108 539744
rect 489821 539686 492108 539688
rect 512900 539744 514819 539746
rect 512900 539688 514758 539744
rect 514814 539688 514819 539744
rect 520598 539716 520658 540228
rect 540470 539716 540530 540228
rect 546401 539746 546467 539749
rect 571333 539746 571399 539749
rect 546401 539744 548044 539746
rect 512900 539686 514819 539688
rect 462221 539683 462287 539686
rect 489821 539683 489887 539686
rect 514753 539683 514819 539686
rect 546401 539688 546406 539744
rect 546462 539688 548044 539744
rect 546401 539686 548044 539688
rect 568836 539744 571399 539746
rect 568836 539688 571338 539744
rect 571394 539688 571399 539744
rect 568836 539686 571399 539688
rect 546401 539683 546467 539686
rect 571333 539683 571399 539686
rect 580533 537842 580599 537845
rect 583520 537842 584960 537932
rect 580533 537840 584960 537842
rect 580533 537784 580538 537840
rect 580594 537784 584960 537840
rect 580533 537782 584960 537784
rect 580533 537779 580599 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 110597 527098 110663 527101
rect 128302 527098 128308 527100
rect 110597 527096 128308 527098
rect 110597 527040 110602 527096
rect 110658 527040 128308 527096
rect 110597 527038 128308 527040
rect 110597 527035 110663 527038
rect 128302 527036 128308 527038
rect 128372 527036 128378 527100
rect 156321 527098 156387 527101
rect 194726 527098 194732 527100
rect 156321 527096 194732 527098
rect 156321 527040 156326 527096
rect 156382 527040 194732 527096
rect 156321 527038 194732 527040
rect 156321 527035 156387 527038
rect 194726 527036 194732 527038
rect 194796 527036 194802 527100
rect 352649 527098 352715 527101
rect 390870 527098 390876 527100
rect 352649 527096 390876 527098
rect 352649 527040 352654 527096
rect 352710 527040 390876 527096
rect 352649 527038 390876 527040
rect 352649 527035 352715 527038
rect 390870 527036 390876 527038
rect 390940 527036 390946 527100
rect 583520 524364 584960 524604
rect 165654 522412 165660 522476
rect 165724 522474 165730 522476
rect 165981 522474 166047 522477
rect 165724 522472 166047 522474
rect 165724 522416 165986 522472
rect 166042 522416 166047 522472
rect 165724 522414 166047 522416
rect 165724 522412 165730 522414
rect 165981 522411 166047 522414
rect 259494 522412 259500 522476
rect 259564 522474 259570 522476
rect 260373 522474 260439 522477
rect 259564 522472 260439 522474
rect 259564 522416 260378 522472
rect 260434 522416 260439 522472
rect 259564 522414 260439 522416
rect 259564 522412 259570 522414
rect 260373 522411 260439 522414
rect 361614 522412 361620 522476
rect 361684 522474 361690 522476
rect 361941 522474 362007 522477
rect 361684 522472 362007 522474
rect 361684 522416 361946 522472
rect 362002 522416 362007 522472
rect 361684 522414 362007 522416
rect 361684 522412 361690 522414
rect 361941 522411 362007 522414
rect 445702 522412 445708 522476
rect 445772 522474 445778 522476
rect 446029 522474 446095 522477
rect 445772 522472 446095 522474
rect 445772 522416 446034 522472
rect 446090 522416 446095 522472
rect 445772 522414 446095 522416
rect 445772 522412 445778 522414
rect 446029 522411 446095 522414
rect 557574 522412 557580 522476
rect 557644 522474 557650 522476
rect 557993 522474 558059 522477
rect 557644 522472 558059 522474
rect 557644 522416 557998 522472
rect 558054 522416 558059 522472
rect 557644 522414 558059 522416
rect 557644 522412 557650 522414
rect 557993 522411 558059 522414
rect 44582 520916 44588 520980
rect 44652 520978 44658 520980
rect 95233 520978 95299 520981
rect 44652 520976 95299 520978
rect 44652 520920 95238 520976
rect 95294 520920 95299 520976
rect 44652 520918 95299 520920
rect 44652 520916 44658 520918
rect 95233 520915 95299 520918
rect 126881 520978 126947 520981
rect 176326 520978 176332 520980
rect 126881 520976 176332 520978
rect 126881 520920 126886 520976
rect 126942 520920 176332 520976
rect 126881 520918 176332 520920
rect 126881 520915 126947 520918
rect 176326 520916 176332 520918
rect 176396 520916 176402 520980
rect 238661 520978 238727 520981
rect 288382 520978 288388 520980
rect 238661 520976 288388 520978
rect 238661 520920 238666 520976
rect 238722 520920 288388 520976
rect 238661 520918 288388 520920
rect 238661 520915 238727 520918
rect 288382 520916 288388 520918
rect 288452 520916 288458 520980
rect 434621 520978 434687 520981
rect 484342 520978 484348 520980
rect 434621 520976 484348 520978
rect 434621 520920 434626 520976
rect 434682 520920 484348 520976
rect 434621 520918 484348 520920
rect 434621 520915 434687 520918
rect 484342 520916 484348 520918
rect 484412 520916 484418 520980
rect 70301 520842 70367 520845
rect 122833 520842 122899 520845
rect 70301 520840 122899 520842
rect 70301 520784 70306 520840
rect 70362 520784 122838 520840
rect 122894 520784 122899 520840
rect 70301 520782 122899 520784
rect 70301 520779 70367 520782
rect 122833 520779 122899 520782
rect 155861 520842 155927 520845
rect 207013 520842 207079 520845
rect 155861 520840 207079 520842
rect 155861 520784 155866 520840
rect 155922 520784 207018 520840
rect 207074 520784 207079 520840
rect 155861 520782 207079 520784
rect 155861 520779 155927 520782
rect 207013 520779 207079 520782
rect 212574 520780 212580 520844
rect 212644 520842 212650 520844
rect 262213 520842 262279 520845
rect 212644 520840 262279 520842
rect 212644 520784 262218 520840
rect 262274 520784 262279 520840
rect 212644 520782 262279 520784
rect 212644 520780 212650 520782
rect 262213 520779 262279 520782
rect 296846 520780 296852 520844
rect 296916 520842 296922 520844
rect 346393 520842 346459 520845
rect 296916 520840 346459 520842
rect 296916 520784 346398 520840
rect 346454 520784 346459 520840
rect 296916 520782 346459 520784
rect 296916 520780 296922 520782
rect 346393 520779 346459 520782
rect 350441 520842 350507 520845
rect 402973 520842 403039 520845
rect 350441 520840 403039 520842
rect 350441 520784 350446 520840
rect 350502 520784 402978 520840
rect 403034 520784 403039 520840
rect 350441 520782 403039 520784
rect 350441 520779 350507 520782
rect 402973 520779 403039 520782
rect 408534 520780 408540 520844
rect 408604 520842 408610 520844
rect 458173 520842 458239 520845
rect 408604 520840 458239 520842
rect 408604 520784 458178 520840
rect 458234 520784 458239 520840
rect 408604 520782 458239 520784
rect 408604 520780 408610 520782
rect 458173 520779 458239 520782
rect 492806 520780 492812 520844
rect 492876 520842 492882 520844
rect 542353 520842 542419 520845
rect 492876 520840 542419 520842
rect 492876 520784 542358 520840
rect 542414 520784 542419 520840
rect 492876 520782 542419 520784
rect 492876 520780 492882 520782
rect 542353 520779 542419 520782
rect 13721 520706 13787 520709
rect 66253 520706 66319 520709
rect 13721 520704 66319 520706
rect 13721 520648 13726 520704
rect 13782 520648 66258 520704
rect 66314 520648 66319 520704
rect 13721 520646 66319 520648
rect 13721 520643 13787 520646
rect 66253 520643 66319 520646
rect 97901 520706 97967 520709
rect 150433 520706 150499 520709
rect 97901 520704 150499 520706
rect 97901 520648 97906 520704
rect 97962 520648 150438 520704
rect 150494 520648 150499 520704
rect 97901 520646 150499 520648
rect 97901 520643 97967 520646
rect 150433 520643 150499 520646
rect 182081 520706 182147 520709
rect 234705 520706 234771 520709
rect 182081 520704 234771 520706
rect 182081 520648 182086 520704
rect 182142 520648 234710 520704
rect 234766 520648 234771 520704
rect 182081 520646 234771 520648
rect 182081 520643 182147 520646
rect 234705 520643 234771 520646
rect 266261 520706 266327 520709
rect 317045 520706 317111 520709
rect 266261 520704 317111 520706
rect 266261 520648 266266 520704
rect 266322 520648 317050 520704
rect 317106 520648 317111 520704
rect 266261 520646 317111 520648
rect 266261 520643 266327 520646
rect 317045 520643 317111 520646
rect 322841 520706 322907 520709
rect 372286 520706 372292 520708
rect 322841 520704 372292 520706
rect 322841 520648 322846 520704
rect 322902 520648 372292 520704
rect 322841 520646 372292 520648
rect 322841 520643 322907 520646
rect 372286 520644 372292 520646
rect 372356 520644 372362 520708
rect 378041 520706 378107 520709
rect 430573 520706 430639 520709
rect 378041 520704 430639 520706
rect 378041 520648 378046 520704
rect 378102 520648 430578 520704
rect 430634 520648 430639 520704
rect 378041 520646 430639 520648
rect 378041 520643 378107 520646
rect 430573 520643 430639 520646
rect 463877 520706 463943 520709
rect 514753 520706 514819 520709
rect 463877 520704 514819 520706
rect 463877 520648 463882 520704
rect 463938 520648 514758 520704
rect 514814 520648 514819 520704
rect 463877 520646 514819 520648
rect 463877 520643 463943 520646
rect 514753 520643 514819 520646
rect 520590 520644 520596 520708
rect 520660 520706 520666 520708
rect 568941 520706 569007 520709
rect 520660 520704 569007 520706
rect 520660 520648 568946 520704
rect 569002 520648 569007 520704
rect 520660 520646 569007 520648
rect 520660 520644 520666 520646
rect 568941 520643 569007 520646
rect -960 514708 480 514948
rect 44582 512756 44588 512820
rect 44652 512756 44658 512820
rect 176326 512756 176332 512820
rect 176396 512756 176402 512820
rect 212574 512756 212580 512820
rect 212644 512756 212650 512820
rect 288382 512756 288388 512820
rect 288452 512756 288458 512820
rect 296478 512756 296484 512820
rect 296548 512756 296554 512820
rect 317045 512818 317111 512821
rect 316910 512816 317111 512818
rect 316910 512760 317050 512816
rect 317106 512760 317111 512816
rect 316910 512758 317111 512760
rect 13721 512274 13787 512277
rect 38653 512274 38719 512277
rect 13721 512272 16100 512274
rect 13721 512216 13726 512272
rect 13782 512216 16100 512272
rect 13721 512214 16100 512216
rect 36892 512272 38719 512274
rect 36892 512216 38658 512272
rect 38714 512216 38719 512272
rect 44590 512244 44650 512756
rect 66253 512274 66319 512277
rect 64860 512272 66319 512274
rect 36892 512214 38719 512216
rect 64860 512216 66258 512272
rect 66314 512216 66319 512272
rect 64860 512214 66319 512216
rect 13721 512211 13787 512214
rect 38653 512211 38719 512214
rect 66253 512211 66319 512214
rect 70301 512274 70367 512277
rect 95233 512274 95299 512277
rect 70301 512272 72036 512274
rect 70301 512216 70306 512272
rect 70362 512216 72036 512272
rect 70301 512214 72036 512216
rect 92828 512272 95299 512274
rect 92828 512216 95238 512272
rect 95294 512216 95299 512272
rect 92828 512214 95299 512216
rect 70301 512211 70367 512214
rect 95233 512211 95299 512214
rect 97901 512274 97967 512277
rect 122833 512274 122899 512277
rect 97901 512272 100188 512274
rect 97901 512216 97906 512272
rect 97962 512216 100188 512272
rect 97901 512214 100188 512216
rect 120796 512272 122899 512274
rect 120796 512216 122838 512272
rect 122894 512216 122899 512272
rect 120796 512214 122899 512216
rect 97901 512211 97967 512214
rect 122833 512211 122899 512214
rect 126881 512274 126947 512277
rect 150433 512274 150499 512277
rect 126881 512272 128156 512274
rect 126881 512216 126886 512272
rect 126942 512216 128156 512272
rect 126881 512214 128156 512216
rect 148948 512272 150499 512274
rect 148948 512216 150438 512272
rect 150494 512216 150499 512272
rect 148948 512214 150499 512216
rect 126881 512211 126947 512214
rect 150433 512211 150499 512214
rect 154481 512274 154547 512277
rect 154481 512272 156124 512274
rect 154481 512216 154486 512272
rect 154542 512216 156124 512272
rect 176334 512244 176394 512756
rect 182081 512274 182147 512277
rect 207013 512274 207079 512277
rect 182081 512272 184092 512274
rect 154481 512214 156124 512216
rect 182081 512216 182086 512272
rect 182142 512216 184092 512272
rect 182081 512214 184092 512216
rect 204884 512272 207079 512274
rect 204884 512216 207018 512272
rect 207074 512216 207079 512272
rect 212582 512244 212642 512756
rect 234705 512274 234771 512277
rect 232852 512272 234771 512274
rect 204884 512214 207079 512216
rect 232852 512216 234710 512272
rect 234766 512216 234771 512272
rect 232852 512214 234771 512216
rect 154481 512211 154547 512214
rect 182081 512211 182147 512214
rect 207013 512211 207079 512214
rect 234705 512211 234771 512214
rect 238661 512274 238727 512277
rect 262213 512274 262279 512277
rect 238661 512272 240212 512274
rect 238661 512216 238666 512272
rect 238722 512216 240212 512272
rect 238661 512214 240212 512216
rect 260820 512272 262279 512274
rect 260820 512216 262218 512272
rect 262274 512216 262279 512272
rect 260820 512214 262279 512216
rect 238661 512211 238727 512214
rect 262213 512211 262279 512214
rect 266261 512274 266327 512277
rect 266261 512272 268180 512274
rect 266261 512216 266266 512272
rect 266322 512216 268180 512272
rect 288390 512244 288450 512756
rect 296486 512244 296546 512756
rect 316910 512244 316970 512758
rect 317045 512755 317111 512758
rect 372286 512756 372292 512820
rect 372356 512756 372362 512820
rect 408534 512756 408540 512820
rect 408604 512756 408610 512820
rect 484342 512756 484348 512820
rect 484412 512756 484418 512820
rect 492622 512756 492628 512820
rect 492692 512756 492698 512820
rect 520590 512756 520596 512820
rect 520660 512756 520666 512820
rect 568941 512818 569007 512821
rect 568806 512816 569007 512818
rect 568806 512760 568946 512816
rect 569002 512760 569007 512816
rect 568806 512758 569007 512760
rect 322841 512274 322907 512277
rect 346393 512274 346459 512277
rect 322841 512272 324116 512274
rect 266261 512214 268180 512216
rect 322841 512216 322846 512272
rect 322902 512216 324116 512272
rect 322841 512214 324116 512216
rect 344908 512272 346459 512274
rect 344908 512216 346398 512272
rect 346454 512216 346459 512272
rect 344908 512214 346459 512216
rect 266261 512211 266327 512214
rect 322841 512211 322907 512214
rect 346393 512211 346459 512214
rect 350441 512274 350507 512277
rect 350441 512272 352084 512274
rect 350441 512216 350446 512272
rect 350502 512216 352084 512272
rect 372294 512244 372354 512756
rect 378041 512274 378107 512277
rect 402973 512274 403039 512277
rect 378041 512272 380052 512274
rect 350441 512214 352084 512216
rect 378041 512216 378046 512272
rect 378102 512216 380052 512272
rect 378041 512214 380052 512216
rect 400844 512272 403039 512274
rect 400844 512216 402978 512272
rect 403034 512216 403039 512272
rect 408542 512244 408602 512756
rect 430573 512274 430639 512277
rect 428812 512272 430639 512274
rect 400844 512214 403039 512216
rect 428812 512216 430578 512272
rect 430634 512216 430639 512272
rect 428812 512214 430639 512216
rect 350441 512211 350507 512214
rect 378041 512211 378107 512214
rect 402973 512211 403039 512214
rect 430573 512211 430639 512214
rect 434621 512274 434687 512277
rect 458173 512274 458239 512277
rect 434621 512272 436172 512274
rect 434621 512216 434626 512272
rect 434682 512216 436172 512272
rect 434621 512214 436172 512216
rect 456964 512272 458239 512274
rect 456964 512216 458178 512272
rect 458234 512216 458239 512272
rect 456964 512214 458239 512216
rect 434621 512211 434687 512214
rect 458173 512211 458239 512214
rect 462221 512274 462287 512277
rect 462221 512272 464140 512274
rect 462221 512216 462226 512272
rect 462282 512216 464140 512272
rect 484350 512244 484410 512756
rect 492630 512244 492690 512756
rect 514753 512274 514819 512277
rect 512900 512272 514819 512274
rect 462221 512214 464140 512216
rect 512900 512216 514758 512272
rect 514814 512216 514819 512272
rect 520598 512244 520658 512756
rect 542353 512274 542419 512277
rect 540868 512272 542419 512274
rect 512900 512214 514819 512216
rect 540868 512216 542358 512272
rect 542414 512216 542419 512272
rect 540868 512214 542419 512216
rect 462221 512211 462287 512214
rect 514753 512211 514819 512214
rect 542353 512211 542419 512214
rect 546401 512274 546467 512277
rect 546401 512272 548044 512274
rect 546401 512216 546406 512272
rect 546462 512216 548044 512272
rect 568806 512244 568866 512758
rect 568941 512755 569007 512758
rect 546401 512214 548044 512216
rect 546401 512211 546467 512214
rect 580625 511322 580691 511325
rect 583520 511322 584960 511412
rect 580625 511320 584960 511322
rect 580625 511264 580630 511320
rect 580686 511264 584960 511320
rect 580625 511262 584960 511264
rect 580625 511259 580691 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3601 501802 3667 501805
rect -960 501800 3667 501802
rect -960 501744 3606 501800
rect 3662 501744 3667 501800
rect -960 501742 3667 501744
rect -960 501652 480 501742
rect 3601 501739 3667 501742
rect 148593 500850 148659 500853
rect 165654 500850 165660 500852
rect 148593 500848 165660 500850
rect 148593 500792 148598 500848
rect 148654 500792 165660 500848
rect 148593 500790 165660 500792
rect 148593 500787 148659 500790
rect 165654 500788 165660 500790
rect 165724 500788 165730 500852
rect 222653 500850 222719 500853
rect 259494 500850 259500 500852
rect 222653 500848 259500 500850
rect 222653 500792 222658 500848
rect 222714 500792 259500 500848
rect 222653 500790 259500 500792
rect 222653 500787 222719 500790
rect 259494 500788 259500 500790
rect 259564 500788 259570 500852
rect 344645 500850 344711 500853
rect 361614 500850 361620 500852
rect 344645 500848 361620 500850
rect 344645 500792 344650 500848
rect 344706 500792 361620 500848
rect 344645 500790 361620 500792
rect 344645 500787 344711 500790
rect 361614 500788 361620 500790
rect 361684 500788 361690 500852
rect 428641 500850 428707 500853
rect 445702 500850 445708 500852
rect 428641 500848 445708 500850
rect 428641 500792 428646 500848
rect 428702 500792 445708 500848
rect 428641 500790 445708 500792
rect 428641 500787 428707 500790
rect 445702 500788 445708 500790
rect 445772 500788 445778 500852
rect 540605 500850 540671 500853
rect 557574 500850 557580 500852
rect 540605 500848 557580 500850
rect 540605 500792 540610 500848
rect 540666 500792 557580 500848
rect 540605 500790 557580 500792
rect 540605 500787 540671 500790
rect 557574 500788 557580 500790
rect 557644 500788 557650 500852
rect 583520 497844 584960 498084
rect 194777 495548 194843 495549
rect 194726 495546 194732 495548
rect 194686 495486 194732 495546
rect 194796 495544 194843 495548
rect 194838 495488 194843 495544
rect 194726 495484 194732 495486
rect 194796 495484 194843 495488
rect 194777 495483 194843 495484
rect 390829 495548 390895 495549
rect 390829 495544 390876 495548
rect 390940 495546 390946 495548
rect 390829 495488 390834 495544
rect 390829 495484 390876 495488
rect 390940 495486 390986 495546
rect 390940 495484 390946 495486
rect 390829 495483 390895 495484
rect 128169 495274 128235 495277
rect 128302 495274 128308 495276
rect 128169 495272 128308 495274
rect 128169 495216 128174 495272
rect 128230 495216 128308 495272
rect 128169 495214 128308 495216
rect 128169 495211 128235 495214
rect 128302 495212 128308 495214
rect 128372 495212 128378 495276
rect -960 488596 480 488836
rect 13537 485754 13603 485757
rect 38653 485754 38719 485757
rect 13537 485752 16100 485754
rect 13537 485696 13542 485752
rect 13598 485696 16100 485752
rect 13537 485694 16100 485696
rect 36892 485752 38719 485754
rect 36892 485696 38658 485752
rect 38714 485696 38719 485752
rect 36892 485694 38719 485696
rect 13537 485691 13603 485694
rect 38653 485691 38719 485694
rect 42701 485754 42767 485757
rect 70301 485754 70367 485757
rect 97901 485754 97967 485757
rect 122833 485754 122899 485757
rect 42701 485752 44068 485754
rect 42701 485696 42706 485752
rect 42762 485696 44068 485752
rect 70301 485752 72036 485754
rect 42701 485694 44068 485696
rect 42701 485691 42767 485694
rect 64462 485212 64522 485724
rect 70301 485696 70306 485752
rect 70362 485696 72036 485752
rect 97901 485752 100188 485754
rect 70301 485694 72036 485696
rect 70301 485691 70367 485694
rect 92430 485212 92490 485724
rect 97901 485696 97906 485752
rect 97962 485696 100188 485752
rect 97901 485694 100188 485696
rect 120796 485752 122899 485754
rect 120796 485696 122838 485752
rect 122894 485696 122899 485752
rect 120796 485694 122899 485696
rect 97901 485691 97967 485694
rect 122833 485691 122899 485694
rect 126881 485754 126947 485757
rect 154481 485754 154547 485757
rect 182081 485754 182147 485757
rect 207013 485754 207079 485757
rect 234705 485754 234771 485757
rect 126881 485752 128156 485754
rect 126881 485696 126886 485752
rect 126942 485696 128156 485752
rect 154481 485752 156124 485754
rect 126881 485694 128156 485696
rect 126881 485691 126947 485694
rect 148366 485212 148426 485724
rect 154481 485696 154486 485752
rect 154542 485696 156124 485752
rect 182081 485752 184092 485754
rect 154481 485694 156124 485696
rect 154481 485691 154547 485694
rect 176334 485212 176394 485724
rect 182081 485696 182086 485752
rect 182142 485696 184092 485752
rect 182081 485694 184092 485696
rect 204884 485752 207079 485754
rect 204884 485696 207018 485752
rect 207074 485696 207079 485752
rect 232852 485752 234771 485754
rect 204884 485694 207079 485696
rect 182081 485691 182147 485694
rect 207013 485691 207079 485694
rect 212582 485212 212642 485724
rect 232852 485696 234710 485752
rect 234766 485696 234771 485752
rect 232852 485694 234771 485696
rect 234705 485691 234771 485694
rect 238661 485754 238727 485757
rect 262213 485754 262279 485757
rect 238661 485752 240212 485754
rect 238661 485696 238666 485752
rect 238722 485696 240212 485752
rect 238661 485694 240212 485696
rect 260820 485752 262279 485754
rect 260820 485696 262218 485752
rect 262274 485696 262279 485752
rect 260820 485694 262279 485696
rect 238661 485691 238727 485694
rect 262213 485691 262279 485694
rect 266261 485754 266327 485757
rect 318793 485754 318859 485757
rect 266261 485752 268180 485754
rect 266261 485696 266266 485752
rect 266322 485696 268180 485752
rect 316940 485752 318859 485754
rect 266261 485694 268180 485696
rect 266261 485691 266327 485694
rect 288390 485212 288450 485724
rect 296486 485212 296546 485724
rect 316940 485696 318798 485752
rect 318854 485696 318859 485752
rect 316940 485694 318859 485696
rect 318793 485691 318859 485694
rect 322841 485754 322907 485757
rect 346393 485754 346459 485757
rect 322841 485752 324116 485754
rect 322841 485696 322846 485752
rect 322902 485696 324116 485752
rect 322841 485694 324116 485696
rect 344908 485752 346459 485754
rect 344908 485696 346398 485752
rect 346454 485696 346459 485752
rect 344908 485694 346459 485696
rect 322841 485691 322907 485694
rect 346393 485691 346459 485694
rect 350441 485754 350507 485757
rect 378041 485754 378107 485757
rect 402973 485754 403039 485757
rect 430573 485754 430639 485757
rect 350441 485752 352084 485754
rect 350441 485696 350446 485752
rect 350502 485696 352084 485752
rect 378041 485752 380052 485754
rect 350441 485694 352084 485696
rect 350441 485691 350507 485694
rect 372294 485212 372354 485724
rect 378041 485696 378046 485752
rect 378102 485696 380052 485752
rect 378041 485694 380052 485696
rect 400844 485752 403039 485754
rect 400844 485696 402978 485752
rect 403034 485696 403039 485752
rect 428812 485752 430639 485754
rect 400844 485694 403039 485696
rect 378041 485691 378107 485694
rect 402973 485691 403039 485694
rect 408542 485212 408602 485724
rect 428812 485696 430578 485752
rect 430634 485696 430639 485752
rect 428812 485694 430639 485696
rect 430573 485691 430639 485694
rect 434621 485754 434687 485757
rect 458173 485754 458239 485757
rect 434621 485752 436172 485754
rect 434621 485696 434626 485752
rect 434682 485696 436172 485752
rect 434621 485694 436172 485696
rect 456964 485752 458239 485754
rect 456964 485696 458178 485752
rect 458234 485696 458239 485752
rect 456964 485694 458239 485696
rect 434621 485691 434687 485694
rect 458173 485691 458239 485694
rect 462221 485754 462287 485757
rect 489821 485754 489887 485757
rect 514753 485754 514819 485757
rect 462221 485752 464140 485754
rect 462221 485696 462226 485752
rect 462282 485696 464140 485752
rect 489821 485752 492108 485754
rect 462221 485694 464140 485696
rect 462221 485691 462287 485694
rect 484350 485212 484410 485724
rect 489821 485696 489826 485752
rect 489882 485696 492108 485752
rect 489821 485694 492108 485696
rect 512900 485752 514819 485754
rect 512900 485696 514758 485752
rect 514814 485696 514819 485752
rect 546401 485754 546467 485757
rect 571333 485754 571399 485757
rect 546401 485752 548044 485754
rect 512900 485694 514819 485696
rect 489821 485691 489887 485694
rect 514753 485691 514819 485694
rect 520598 485212 520658 485724
rect 540470 485212 540530 485724
rect 546401 485696 546406 485752
rect 546462 485696 548044 485752
rect 546401 485694 548044 485696
rect 568836 485752 571399 485754
rect 568836 485696 571338 485752
rect 571394 485696 571399 485752
rect 568836 485694 571399 485696
rect 546401 485691 546467 485694
rect 571333 485691 571399 485694
rect 64454 485148 64460 485212
rect 64524 485148 64530 485212
rect 92422 485148 92428 485212
rect 92492 485148 92498 485212
rect 148358 485148 148364 485212
rect 148428 485148 148434 485212
rect 176326 485148 176332 485212
rect 176396 485148 176402 485212
rect 212574 485148 212580 485212
rect 212644 485148 212650 485212
rect 288382 485148 288388 485212
rect 288452 485148 288458 485212
rect 296478 485148 296484 485212
rect 296548 485148 296554 485212
rect 372286 485148 372292 485212
rect 372356 485148 372362 485212
rect 408534 485148 408540 485212
rect 408604 485148 408610 485212
rect 484342 485148 484348 485212
rect 484412 485148 484418 485212
rect 520590 485148 520596 485212
rect 520660 485148 520666 485212
rect 540462 485148 540468 485212
rect 540532 485148 540538 485212
rect 580717 484666 580783 484669
rect 583520 484666 584960 484756
rect 580717 484664 584960 484666
rect 580717 484608 580722 484664
rect 580778 484608 584960 484664
rect 580717 484606 584960 484608
rect 580717 484603 580783 484606
rect 583520 484516 584960 484606
rect 13537 477322 13603 477325
rect 64454 477322 64460 477324
rect 13537 477320 64460 477322
rect 13537 477264 13542 477320
rect 13598 477264 64460 477320
rect 13537 477262 64460 477264
rect 13537 477259 13603 477262
rect 64454 477260 64460 477262
rect 64524 477260 64530 477324
rect 70301 477322 70367 477325
rect 122833 477322 122899 477325
rect 70301 477320 122899 477322
rect 70301 477264 70306 477320
rect 70362 477264 122838 477320
rect 122894 477264 122899 477320
rect 70301 477262 122899 477264
rect 70301 477259 70367 477262
rect 122833 477259 122899 477262
rect 126881 477322 126947 477325
rect 176326 477322 176332 477324
rect 126881 477320 176332 477322
rect 126881 477264 126886 477320
rect 126942 477264 176332 477320
rect 126881 477262 176332 477264
rect 126881 477259 126947 477262
rect 176326 477260 176332 477262
rect 176396 477260 176402 477324
rect 182081 477322 182147 477325
rect 234705 477322 234771 477325
rect 182081 477320 234771 477322
rect 182081 477264 182086 477320
rect 182142 477264 234710 477320
rect 234766 477264 234771 477320
rect 182081 477262 234771 477264
rect 182081 477259 182147 477262
rect 234705 477259 234771 477262
rect 266261 477322 266327 477325
rect 318793 477322 318859 477325
rect 266261 477320 318859 477322
rect 266261 477264 266266 477320
rect 266322 477264 318798 477320
rect 318854 477264 318859 477320
rect 266261 477262 318859 477264
rect 266261 477259 266327 477262
rect 318793 477259 318859 477262
rect 350441 477322 350507 477325
rect 402973 477322 403039 477325
rect 350441 477320 403039 477322
rect 350441 477264 350446 477320
rect 350502 477264 402978 477320
rect 403034 477264 403039 477320
rect 350441 477262 403039 477264
rect 350441 477259 350507 477262
rect 402973 477259 403039 477262
rect 408534 477260 408540 477324
rect 408604 477322 408610 477324
rect 458173 477322 458239 477325
rect 408604 477320 458239 477322
rect 408604 477264 458178 477320
rect 458234 477264 458239 477320
rect 408604 477262 458239 477264
rect 408604 477260 408610 477262
rect 458173 477259 458239 477262
rect 462221 477322 462287 477325
rect 514753 477322 514819 477325
rect 462221 477320 514819 477322
rect 462221 477264 462226 477320
rect 462282 477264 514758 477320
rect 514814 477264 514819 477320
rect 462221 477262 514819 477264
rect 462221 477259 462287 477262
rect 514753 477259 514819 477262
rect 520590 477260 520596 477324
rect 520660 477322 520666 477324
rect 571333 477322 571399 477325
rect 520660 477320 571399 477322
rect 520660 477264 571338 477320
rect 571394 477264 571399 477320
rect 520660 477262 571399 477264
rect 520660 477260 520666 477262
rect 571333 477259 571399 477262
rect 42701 477186 42767 477189
rect 92422 477186 92428 477188
rect 42701 477184 92428 477186
rect 42701 477128 42706 477184
rect 42762 477128 92428 477184
rect 42701 477126 92428 477128
rect 42701 477123 42767 477126
rect 92422 477124 92428 477126
rect 92492 477124 92498 477188
rect 97901 477186 97967 477189
rect 148358 477186 148364 477188
rect 97901 477184 148364 477186
rect 97901 477128 97906 477184
rect 97962 477128 148364 477184
rect 97901 477126 148364 477128
rect 97901 477123 97967 477126
rect 148358 477124 148364 477126
rect 148428 477124 148434 477188
rect 154481 477186 154547 477189
rect 207013 477186 207079 477189
rect 154481 477184 207079 477186
rect 154481 477128 154486 477184
rect 154542 477128 207018 477184
rect 207074 477128 207079 477184
rect 154481 477126 207079 477128
rect 154481 477123 154547 477126
rect 207013 477123 207079 477126
rect 212574 477124 212580 477188
rect 212644 477186 212650 477188
rect 262213 477186 262279 477189
rect 212644 477184 262279 477186
rect 212644 477128 262218 477184
rect 262274 477128 262279 477184
rect 212644 477126 262279 477128
rect 212644 477124 212650 477126
rect 262213 477123 262279 477126
rect 296846 477124 296852 477188
rect 296916 477186 296922 477188
rect 346393 477186 346459 477189
rect 296916 477184 346459 477186
rect 296916 477128 346398 477184
rect 346454 477128 346459 477184
rect 296916 477126 346459 477128
rect 296916 477124 296922 477126
rect 346393 477123 346459 477126
rect 378041 477186 378107 477189
rect 430573 477186 430639 477189
rect 378041 477184 430639 477186
rect 378041 477128 378046 477184
rect 378102 477128 430578 477184
rect 430634 477128 430639 477184
rect 378041 477126 430639 477128
rect 378041 477123 378107 477126
rect 430573 477123 430639 477126
rect 434621 477186 434687 477189
rect 484342 477186 484348 477188
rect 434621 477184 484348 477186
rect 434621 477128 434626 477184
rect 434682 477128 484348 477184
rect 434621 477126 484348 477128
rect 434621 477123 434687 477126
rect 484342 477124 484348 477126
rect 484412 477124 484418 477188
rect 489821 477186 489887 477189
rect 540462 477186 540468 477188
rect 489821 477184 540468 477186
rect 489821 477128 489826 477184
rect 489882 477128 540468 477184
rect 489821 477126 540468 477128
rect 489821 477123 489887 477126
rect 540462 477124 540468 477126
rect 540532 477124 540538 477188
rect 238661 477050 238727 477053
rect 288382 477050 288388 477052
rect 238661 477048 288388 477050
rect 238661 476992 238666 477048
rect 238722 476992 288388 477048
rect 238661 476990 288388 476992
rect 238661 476987 238727 476990
rect 288382 476988 288388 476990
rect 288452 476988 288458 477052
rect 322841 477050 322907 477053
rect 372286 477050 372292 477052
rect 322841 477048 372292 477050
rect 322841 476992 322846 477048
rect 322902 476992 372292 477048
rect 322841 476990 372292 476992
rect 322841 476987 322907 476990
rect 372286 476988 372292 476990
rect 372356 476988 372362 477052
rect -960 475690 480 475780
rect 3693 475690 3759 475693
rect -960 475688 3759 475690
rect -960 475632 3698 475688
rect 3754 475632 3759 475688
rect -960 475630 3759 475632
rect -960 475540 480 475630
rect 3693 475627 3759 475630
rect 110597 473242 110663 473245
rect 128302 473242 128308 473244
rect 110597 473240 128308 473242
rect 110597 473184 110602 473240
rect 110658 473184 128308 473240
rect 110597 473182 128308 473184
rect 110597 473179 110663 473182
rect 128302 473180 128308 473182
rect 128372 473180 128378 473244
rect 156321 473242 156387 473245
rect 194726 473242 194732 473244
rect 156321 473240 194732 473242
rect 156321 473184 156326 473240
rect 156382 473184 194732 473240
rect 156321 473182 194732 473184
rect 156321 473179 156387 473182
rect 194726 473180 194732 473182
rect 194796 473180 194802 473244
rect 352649 473242 352715 473245
rect 390870 473242 390876 473244
rect 352649 473240 390876 473242
rect 352649 473184 352654 473240
rect 352710 473184 390876 473240
rect 352649 473182 390876 473184
rect 352649 473179 352715 473182
rect 390870 473180 390876 473182
rect 390940 473180 390946 473244
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect 81382 468420 81388 468484
rect 81452 468482 81458 468484
rect 81985 468482 82051 468485
rect 81452 468480 82051 468482
rect 81452 468424 81990 468480
rect 82046 468424 82051 468480
rect 81452 468422 82051 468424
rect 81452 468420 81458 468422
rect 81985 468419 82051 468422
rect 165654 468420 165660 468484
rect 165724 468482 165730 468484
rect 165981 468482 166047 468485
rect 165724 468480 166047 468482
rect 165724 468424 165986 468480
rect 166042 468424 166047 468480
rect 165724 468422 166047 468424
rect 165724 468420 165730 468422
rect 165981 468419 166047 468422
rect 259494 468420 259500 468484
rect 259564 468482 259570 468484
rect 260373 468482 260439 468485
rect 259564 468480 260439 468482
rect 259564 468424 260378 468480
rect 260434 468424 260439 468480
rect 259564 468422 260439 468424
rect 259564 468420 259570 468422
rect 260373 468419 260439 468422
rect 361614 468420 361620 468484
rect 361684 468482 361690 468484
rect 361941 468482 362007 468485
rect 361684 468480 362007 468482
rect 361684 468424 361946 468480
rect 362002 468424 362007 468480
rect 361684 468422 362007 468424
rect 361684 468420 361690 468422
rect 361941 468419 362007 468422
rect 445702 468420 445708 468484
rect 445772 468482 445778 468484
rect 446029 468482 446095 468485
rect 445772 468480 446095 468482
rect 445772 468424 446034 468480
rect 446090 468424 446095 468480
rect 445772 468422 446095 468424
rect 445772 468420 445778 468422
rect 446029 468419 446095 468422
rect 455454 468420 455460 468484
rect 455524 468482 455530 468484
rect 456333 468482 456399 468485
rect 455524 468480 456399 468482
rect 455524 468424 456338 468480
rect 456394 468424 456399 468480
rect 455524 468422 456399 468424
rect 455524 468420 455530 468422
rect 456333 468419 456399 468422
rect 557574 468420 557580 468484
rect 557644 468482 557650 468484
rect 557993 468482 558059 468485
rect 557644 468480 558059 468482
rect 557644 468424 557998 468480
rect 558054 468424 558059 468480
rect 557644 468422 558059 468424
rect 557644 468420 557650 468422
rect 557993 468419 558059 468422
rect 212574 466924 212580 466988
rect 212644 466986 212650 466988
rect 262213 466986 262279 466989
rect 212644 466984 262279 466986
rect 212644 466928 262218 466984
rect 262274 466928 262279 466984
rect 212644 466926 262279 466928
rect 212644 466924 212650 466926
rect 262213 466923 262279 466926
rect 408534 466924 408540 466988
rect 408604 466986 408610 466988
rect 458173 466986 458239 466989
rect 408604 466984 458239 466986
rect 408604 466928 458178 466984
rect 458234 466928 458239 466984
rect 408604 466926 458239 466928
rect 408604 466924 408610 466926
rect 458173 466923 458239 466926
rect 44582 466788 44588 466852
rect 44652 466850 44658 466852
rect 95233 466850 95299 466853
rect 44652 466848 95299 466850
rect 44652 466792 95238 466848
rect 95294 466792 95299 466848
rect 44652 466790 95299 466792
rect 44652 466788 44658 466790
rect 95233 466787 95299 466790
rect 97901 466850 97967 466853
rect 150433 466850 150499 466853
rect 97901 466848 150499 466850
rect 97901 466792 97906 466848
rect 97962 466792 150438 466848
rect 150494 466792 150499 466848
rect 97901 466790 150499 466792
rect 97901 466787 97967 466790
rect 150433 466787 150499 466790
rect 154481 466850 154547 466853
rect 207013 466850 207079 466853
rect 154481 466848 207079 466850
rect 154481 466792 154486 466848
rect 154542 466792 207018 466848
rect 207074 466792 207079 466848
rect 154481 466790 207079 466792
rect 154481 466787 154547 466790
rect 207013 466787 207079 466790
rect 240542 466788 240548 466852
rect 240612 466850 240618 466852
rect 291193 466850 291259 466853
rect 240612 466848 291259 466850
rect 240612 466792 291198 466848
rect 291254 466792 291259 466848
rect 240612 466790 291259 466792
rect 240612 466788 240618 466790
rect 291193 466787 291259 466790
rect 296846 466788 296852 466852
rect 296916 466850 296922 466852
rect 346393 466850 346459 466853
rect 296916 466848 346459 466850
rect 296916 466792 346398 466848
rect 346454 466792 346459 466848
rect 296916 466790 346459 466792
rect 296916 466788 296922 466790
rect 346393 466787 346459 466790
rect 350441 466850 350507 466853
rect 402973 466850 403039 466853
rect 350441 466848 403039 466850
rect 350441 466792 350446 466848
rect 350502 466792 402978 466848
rect 403034 466792 403039 466848
rect 350441 466790 403039 466792
rect 350441 466787 350507 466790
rect 402973 466787 403039 466790
rect 436502 466788 436508 466852
rect 436572 466850 436578 466852
rect 487153 466850 487219 466853
rect 436572 466848 487219 466850
rect 436572 466792 487158 466848
rect 487214 466792 487219 466848
rect 436572 466790 487219 466792
rect 436572 466788 436578 466790
rect 487153 466787 487219 466790
rect 492806 466788 492812 466852
rect 492876 466850 492882 466852
rect 542353 466850 542419 466853
rect 492876 466848 542419 466850
rect 492876 466792 542358 466848
rect 542414 466792 542419 466848
rect 492876 466790 542419 466792
rect 492876 466788 492882 466790
rect 542353 466787 542419 466790
rect 13537 466714 13603 466717
rect 66253 466714 66319 466717
rect 13537 466712 66319 466714
rect 13537 466656 13542 466712
rect 13598 466656 66258 466712
rect 66314 466656 66319 466712
rect 13537 466654 66319 466656
rect 13537 466651 13603 466654
rect 66253 466651 66319 466654
rect 70301 466714 70367 466717
rect 122833 466714 122899 466717
rect 70301 466712 122899 466714
rect 70301 466656 70306 466712
rect 70362 466656 122838 466712
rect 122894 466656 122899 466712
rect 70301 466654 122899 466656
rect 70301 466651 70367 466654
rect 122833 466651 122899 466654
rect 128486 466652 128492 466716
rect 128556 466714 128562 466716
rect 178033 466714 178099 466717
rect 128556 466712 178099 466714
rect 128556 466656 178038 466712
rect 178094 466656 178099 466712
rect 128556 466654 178099 466656
rect 128556 466652 128562 466654
rect 178033 466651 178099 466654
rect 182081 466714 182147 466717
rect 234705 466714 234771 466717
rect 182081 466712 234771 466714
rect 182081 466656 182086 466712
rect 182142 466656 234710 466712
rect 234766 466656 234771 466712
rect 182081 466654 234771 466656
rect 182081 466651 182147 466654
rect 234705 466651 234771 466654
rect 266261 466714 266327 466717
rect 318793 466714 318859 466717
rect 266261 466712 318859 466714
rect 266261 466656 266266 466712
rect 266322 466656 318798 466712
rect 318854 466656 318859 466712
rect 266261 466654 318859 466656
rect 266261 466651 266327 466654
rect 318793 466651 318859 466654
rect 324630 466652 324636 466716
rect 324700 466714 324706 466716
rect 375373 466714 375439 466717
rect 324700 466712 375439 466714
rect 324700 466656 375378 466712
rect 375434 466656 375439 466712
rect 324700 466654 375439 466656
rect 324700 466652 324706 466654
rect 375373 466651 375439 466654
rect 378041 466714 378107 466717
rect 430573 466714 430639 466717
rect 378041 466712 430639 466714
rect 378041 466656 378046 466712
rect 378102 466656 430578 466712
rect 430634 466656 430639 466712
rect 378041 466654 430639 466656
rect 378041 466651 378107 466654
rect 430573 466651 430639 466654
rect 462221 466714 462287 466717
rect 514753 466714 514819 466717
rect 462221 466712 514819 466714
rect 462221 466656 462226 466712
rect 462282 466656 514758 466712
rect 514814 466656 514819 466712
rect 462221 466654 514819 466656
rect 462221 466651 462287 466654
rect 514753 466651 514819 466654
rect 520590 466652 520596 466716
rect 520660 466714 520666 466716
rect 571333 466714 571399 466717
rect 520660 466712 571399 466714
rect 520660 466656 571338 466712
rect 571394 466656 571399 466712
rect 520660 466654 571399 466656
rect 520660 466652 520666 466654
rect 571333 466651 571399 466654
rect -960 462484 480 462724
rect 44582 458764 44588 458828
rect 44652 458764 44658 458828
rect 128486 458764 128492 458828
rect 128556 458764 128562 458828
rect 212574 458764 212580 458828
rect 212644 458764 212650 458828
rect 240542 458764 240548 458828
rect 240612 458764 240618 458828
rect 296478 458764 296484 458828
rect 296548 458764 296554 458828
rect 324630 458764 324636 458828
rect 324700 458764 324706 458828
rect 408534 458764 408540 458828
rect 408604 458764 408610 458828
rect 436502 458764 436508 458828
rect 436572 458764 436578 458828
rect 492622 458764 492628 458828
rect 492692 458764 492698 458828
rect 520590 458764 520596 458828
rect 520660 458764 520666 458828
rect 13537 458282 13603 458285
rect 38653 458282 38719 458285
rect 13537 458280 16100 458282
rect 13537 458224 13542 458280
rect 13598 458224 16100 458280
rect 13537 458222 16100 458224
rect 36892 458280 38719 458282
rect 36892 458224 38658 458280
rect 38714 458224 38719 458280
rect 44590 458252 44650 458764
rect 66253 458282 66319 458285
rect 64860 458280 66319 458282
rect 36892 458222 38719 458224
rect 64860 458224 66258 458280
rect 66314 458224 66319 458280
rect 64860 458222 66319 458224
rect 13537 458219 13603 458222
rect 38653 458219 38719 458222
rect 66253 458219 66319 458222
rect 70301 458282 70367 458285
rect 95233 458282 95299 458285
rect 70301 458280 72036 458282
rect 70301 458224 70306 458280
rect 70362 458224 72036 458280
rect 70301 458222 72036 458224
rect 92828 458280 95299 458282
rect 92828 458224 95238 458280
rect 95294 458224 95299 458280
rect 92828 458222 95299 458224
rect 70301 458219 70367 458222
rect 95233 458219 95299 458222
rect 97901 458282 97967 458285
rect 122833 458282 122899 458285
rect 97901 458280 100188 458282
rect 97901 458224 97906 458280
rect 97962 458224 100188 458280
rect 97901 458222 100188 458224
rect 120796 458280 122899 458282
rect 120796 458224 122838 458280
rect 122894 458224 122899 458280
rect 128494 458252 128554 458764
rect 150433 458282 150499 458285
rect 148948 458280 150499 458282
rect 120796 458222 122899 458224
rect 148948 458224 150438 458280
rect 150494 458224 150499 458280
rect 148948 458222 150499 458224
rect 97901 458219 97967 458222
rect 122833 458219 122899 458222
rect 150433 458219 150499 458222
rect 154481 458282 154547 458285
rect 178033 458282 178099 458285
rect 154481 458280 156124 458282
rect 154481 458224 154486 458280
rect 154542 458224 156124 458280
rect 154481 458222 156124 458224
rect 176916 458280 178099 458282
rect 176916 458224 178038 458280
rect 178094 458224 178099 458280
rect 176916 458222 178099 458224
rect 154481 458219 154547 458222
rect 178033 458219 178099 458222
rect 182081 458282 182147 458285
rect 207013 458282 207079 458285
rect 182081 458280 184092 458282
rect 182081 458224 182086 458280
rect 182142 458224 184092 458280
rect 182081 458222 184092 458224
rect 204884 458280 207079 458282
rect 204884 458224 207018 458280
rect 207074 458224 207079 458280
rect 212582 458252 212642 458764
rect 234705 458282 234771 458285
rect 232852 458280 234771 458282
rect 204884 458222 207079 458224
rect 232852 458224 234710 458280
rect 234766 458224 234771 458280
rect 240550 458252 240610 458764
rect 262213 458282 262279 458285
rect 260820 458280 262279 458282
rect 232852 458222 234771 458224
rect 260820 458224 262218 458280
rect 262274 458224 262279 458280
rect 260820 458222 262279 458224
rect 182081 458219 182147 458222
rect 207013 458219 207079 458222
rect 234705 458219 234771 458222
rect 262213 458219 262279 458222
rect 266261 458282 266327 458285
rect 291193 458282 291259 458285
rect 266261 458280 268180 458282
rect 266261 458224 266266 458280
rect 266322 458224 268180 458280
rect 266261 458222 268180 458224
rect 288788 458280 291259 458282
rect 288788 458224 291198 458280
rect 291254 458224 291259 458280
rect 296486 458252 296546 458764
rect 318793 458282 318859 458285
rect 316940 458280 318859 458282
rect 288788 458222 291259 458224
rect 316940 458224 318798 458280
rect 318854 458224 318859 458280
rect 324638 458252 324698 458764
rect 346393 458282 346459 458285
rect 344908 458280 346459 458282
rect 316940 458222 318859 458224
rect 344908 458224 346398 458280
rect 346454 458224 346459 458280
rect 344908 458222 346459 458224
rect 266261 458219 266327 458222
rect 291193 458219 291259 458222
rect 318793 458219 318859 458222
rect 346393 458219 346459 458222
rect 350441 458282 350507 458285
rect 375373 458282 375439 458285
rect 350441 458280 352084 458282
rect 350441 458224 350446 458280
rect 350502 458224 352084 458280
rect 350441 458222 352084 458224
rect 372876 458280 375439 458282
rect 372876 458224 375378 458280
rect 375434 458224 375439 458280
rect 372876 458222 375439 458224
rect 350441 458219 350507 458222
rect 375373 458219 375439 458222
rect 378041 458282 378107 458285
rect 402973 458282 403039 458285
rect 378041 458280 380052 458282
rect 378041 458224 378046 458280
rect 378102 458224 380052 458280
rect 378041 458222 380052 458224
rect 400844 458280 403039 458282
rect 400844 458224 402978 458280
rect 403034 458224 403039 458280
rect 408542 458252 408602 458764
rect 430573 458282 430639 458285
rect 428812 458280 430639 458282
rect 400844 458222 403039 458224
rect 428812 458224 430578 458280
rect 430634 458224 430639 458280
rect 436510 458252 436570 458764
rect 458173 458282 458239 458285
rect 456964 458280 458239 458282
rect 428812 458222 430639 458224
rect 456964 458224 458178 458280
rect 458234 458224 458239 458280
rect 456964 458222 458239 458224
rect 378041 458219 378107 458222
rect 402973 458219 403039 458222
rect 430573 458219 430639 458222
rect 458173 458219 458239 458222
rect 462221 458282 462287 458285
rect 487153 458282 487219 458285
rect 462221 458280 464140 458282
rect 462221 458224 462226 458280
rect 462282 458224 464140 458280
rect 462221 458222 464140 458224
rect 484932 458280 487219 458282
rect 484932 458224 487158 458280
rect 487214 458224 487219 458280
rect 492630 458252 492690 458764
rect 514753 458282 514819 458285
rect 512900 458280 514819 458282
rect 484932 458222 487219 458224
rect 512900 458224 514758 458280
rect 514814 458224 514819 458280
rect 520598 458252 520658 458764
rect 542353 458282 542419 458285
rect 540868 458280 542419 458282
rect 512900 458222 514819 458224
rect 540868 458224 542358 458280
rect 542414 458224 542419 458280
rect 540868 458222 542419 458224
rect 462221 458219 462287 458222
rect 487153 458219 487219 458222
rect 514753 458219 514819 458222
rect 542353 458219 542419 458222
rect 546401 458282 546467 458285
rect 571333 458282 571399 458285
rect 546401 458280 548044 458282
rect 546401 458224 546406 458280
rect 546462 458224 548044 458280
rect 546401 458222 548044 458224
rect 568836 458280 571399 458282
rect 568836 458224 571338 458280
rect 571394 458224 571399 458280
rect 568836 458222 571399 458224
rect 546401 458219 546467 458222
rect 571333 458219 571399 458222
rect 583520 457996 584960 458236
rect -960 449578 480 449668
rect 2773 449578 2839 449581
rect -960 449576 2839 449578
rect -960 449520 2778 449576
rect 2834 449520 2839 449576
rect -960 449518 2839 449520
rect -960 449428 480 449518
rect 2773 449515 2839 449518
rect 64597 445634 64663 445637
rect 81382 445634 81388 445636
rect 64597 445632 81388 445634
rect 64597 445576 64602 445632
rect 64658 445576 81388 445632
rect 64597 445574 81388 445576
rect 64597 445571 64663 445574
rect 81382 445572 81388 445574
rect 81452 445572 81458 445636
rect 148593 445634 148659 445637
rect 165654 445634 165660 445636
rect 148593 445632 165660 445634
rect 148593 445576 148598 445632
rect 148654 445576 165660 445632
rect 148593 445574 165660 445576
rect 148593 445571 148659 445574
rect 165654 445572 165660 445574
rect 165724 445572 165730 445636
rect 222653 445634 222719 445637
rect 259494 445634 259500 445636
rect 222653 445632 259500 445634
rect 222653 445576 222658 445632
rect 222714 445576 259500 445632
rect 222653 445574 259500 445576
rect 222653 445571 222719 445574
rect 259494 445572 259500 445574
rect 259564 445572 259570 445636
rect 344645 445634 344711 445637
rect 361614 445634 361620 445636
rect 344645 445632 361620 445634
rect 344645 445576 344650 445632
rect 344706 445576 361620 445632
rect 344645 445574 361620 445576
rect 344645 445571 344711 445574
rect 361614 445572 361620 445574
rect 361684 445572 361690 445636
rect 418337 445634 418403 445637
rect 455454 445634 455460 445636
rect 418337 445632 455460 445634
rect 418337 445576 418342 445632
rect 418398 445576 455460 445632
rect 418337 445574 455460 445576
rect 418337 445571 418403 445574
rect 455454 445572 455460 445574
rect 455524 445572 455530 445636
rect 540605 445634 540671 445637
rect 557574 445634 557580 445636
rect 540605 445632 557580 445634
rect 540605 445576 540610 445632
rect 540666 445576 557580 445632
rect 540605 445574 557580 445576
rect 540605 445571 540671 445574
rect 557574 445572 557580 445574
rect 557644 445572 557650 445636
rect 428641 445498 428707 445501
rect 445702 445498 445708 445500
rect 428641 445496 445708 445498
rect 428641 445440 428646 445496
rect 428702 445440 445708 445496
rect 428641 445438 445708 445440
rect 428641 445435 428707 445438
rect 445702 445436 445708 445438
rect 445772 445436 445778 445500
rect 583520 444668 584960 444908
rect 128302 441628 128308 441692
rect 128372 441690 128378 441692
rect 128445 441690 128511 441693
rect 194777 441692 194843 441693
rect 194726 441690 194732 441692
rect 128372 441688 128511 441690
rect 128372 441632 128450 441688
rect 128506 441632 128511 441688
rect 128372 441630 128511 441632
rect 194686 441630 194732 441690
rect 194796 441688 194843 441692
rect 194838 441632 194843 441688
rect 128372 441628 128378 441630
rect 128445 441627 128511 441630
rect 194726 441628 194732 441630
rect 194796 441628 194843 441632
rect 194777 441627 194843 441628
rect 390829 441692 390895 441693
rect 390829 441688 390876 441692
rect 390940 441690 390946 441692
rect 390829 441632 390834 441688
rect 390829 441628 390876 441632
rect 390940 441630 390986 441690
rect 390940 441628 390946 441630
rect 390829 441627 390895 441628
rect -960 436508 480 436748
rect 13721 431762 13787 431765
rect 38653 431762 38719 431765
rect 13721 431760 16100 431762
rect 13721 431704 13726 431760
rect 13782 431704 16100 431760
rect 13721 431702 16100 431704
rect 36892 431760 38719 431762
rect 36892 431704 38658 431760
rect 38714 431704 38719 431760
rect 36892 431702 38719 431704
rect 13721 431699 13787 431702
rect 38653 431699 38719 431702
rect 42701 431762 42767 431765
rect 70301 431762 70367 431765
rect 97901 431762 97967 431765
rect 122833 431762 122899 431765
rect 42701 431760 44068 431762
rect 42701 431704 42706 431760
rect 42762 431704 44068 431760
rect 70301 431760 72036 431762
rect 42701 431702 44068 431704
rect 42701 431699 42767 431702
rect 64462 431220 64522 431732
rect 70301 431704 70306 431760
rect 70362 431704 72036 431760
rect 97901 431760 100188 431762
rect 70301 431702 72036 431704
rect 70301 431699 70367 431702
rect 92430 431220 92490 431732
rect 97901 431704 97906 431760
rect 97962 431704 100188 431760
rect 97901 431702 100188 431704
rect 120796 431760 122899 431762
rect 120796 431704 122838 431760
rect 122894 431704 122899 431760
rect 120796 431702 122899 431704
rect 97901 431699 97967 431702
rect 122833 431699 122899 431702
rect 126881 431762 126947 431765
rect 154481 431762 154547 431765
rect 182081 431762 182147 431765
rect 207013 431762 207079 431765
rect 126881 431760 128156 431762
rect 126881 431704 126886 431760
rect 126942 431704 128156 431760
rect 154481 431760 156124 431762
rect 126881 431702 128156 431704
rect 126881 431699 126947 431702
rect 148366 431220 148426 431732
rect 154481 431704 154486 431760
rect 154542 431704 156124 431760
rect 182081 431760 184092 431762
rect 154481 431702 156124 431704
rect 154481 431699 154547 431702
rect 176334 431220 176394 431732
rect 182081 431704 182086 431760
rect 182142 431704 184092 431760
rect 182081 431702 184092 431704
rect 204884 431760 207079 431762
rect 204884 431704 207018 431760
rect 207074 431704 207079 431760
rect 204884 431702 207079 431704
rect 182081 431699 182147 431702
rect 207013 431699 207079 431702
rect 209681 431762 209747 431765
rect 234705 431762 234771 431765
rect 209681 431760 212060 431762
rect 209681 431704 209686 431760
rect 209742 431704 212060 431760
rect 209681 431702 212060 431704
rect 232852 431760 234771 431762
rect 232852 431704 234710 431760
rect 234766 431704 234771 431760
rect 232852 431702 234771 431704
rect 209681 431699 209747 431702
rect 234705 431699 234771 431702
rect 238661 431762 238727 431765
rect 266261 431762 266327 431765
rect 293861 431762 293927 431765
rect 318793 431762 318859 431765
rect 238661 431760 240212 431762
rect 238661 431704 238666 431760
rect 238722 431704 240212 431760
rect 266261 431760 268180 431762
rect 238661 431702 240212 431704
rect 238661 431699 238727 431702
rect 260422 431220 260482 431732
rect 266261 431704 266266 431760
rect 266322 431704 268180 431760
rect 293861 431760 296148 431762
rect 266261 431702 268180 431704
rect 266261 431699 266327 431702
rect 288390 431220 288450 431732
rect 293861 431704 293866 431760
rect 293922 431704 296148 431760
rect 293861 431702 296148 431704
rect 316940 431760 318859 431762
rect 316940 431704 318798 431760
rect 318854 431704 318859 431760
rect 316940 431702 318859 431704
rect 293861 431699 293927 431702
rect 318793 431699 318859 431702
rect 322841 431762 322907 431765
rect 350441 431762 350507 431765
rect 378041 431762 378107 431765
rect 402973 431762 403039 431765
rect 322841 431760 324116 431762
rect 322841 431704 322846 431760
rect 322902 431704 324116 431760
rect 350441 431760 352084 431762
rect 322841 431702 324116 431704
rect 322841 431699 322907 431702
rect 344326 431220 344386 431732
rect 350441 431704 350446 431760
rect 350502 431704 352084 431760
rect 378041 431760 380052 431762
rect 350441 431702 352084 431704
rect 350441 431699 350507 431702
rect 372294 431220 372354 431732
rect 378041 431704 378046 431760
rect 378102 431704 380052 431760
rect 378041 431702 380052 431704
rect 400844 431760 403039 431762
rect 400844 431704 402978 431760
rect 403034 431704 403039 431760
rect 400844 431702 403039 431704
rect 378041 431699 378107 431702
rect 402973 431699 403039 431702
rect 405641 431762 405707 431765
rect 430573 431762 430639 431765
rect 405641 431760 408204 431762
rect 405641 431704 405646 431760
rect 405702 431704 408204 431760
rect 405641 431702 408204 431704
rect 428812 431760 430639 431762
rect 428812 431704 430578 431760
rect 430634 431704 430639 431760
rect 428812 431702 430639 431704
rect 405641 431699 405707 431702
rect 430573 431699 430639 431702
rect 434621 431762 434687 431765
rect 462221 431762 462287 431765
rect 514753 431762 514819 431765
rect 542353 431762 542419 431765
rect 434621 431760 436172 431762
rect 434621 431704 434626 431760
rect 434682 431704 436172 431760
rect 462221 431760 464140 431762
rect 434621 431702 436172 431704
rect 434621 431699 434687 431702
rect 456382 431220 456442 431732
rect 462221 431704 462226 431760
rect 462282 431704 464140 431760
rect 512900 431760 514819 431762
rect 462221 431702 464140 431704
rect 462221 431699 462287 431702
rect 484350 431220 484410 431732
rect 492630 431220 492690 431732
rect 512900 431704 514758 431760
rect 514814 431704 514819 431760
rect 540868 431760 542419 431762
rect 512900 431702 514819 431704
rect 514753 431699 514819 431702
rect 520598 431220 520658 431732
rect 540868 431704 542358 431760
rect 542414 431704 542419 431760
rect 540868 431702 542419 431704
rect 542353 431699 542419 431702
rect 546401 431762 546467 431765
rect 571333 431762 571399 431765
rect 546401 431760 548044 431762
rect 546401 431704 546406 431760
rect 546462 431704 548044 431760
rect 546401 431702 548044 431704
rect 568836 431760 571399 431762
rect 568836 431704 571338 431760
rect 571394 431704 571399 431760
rect 568836 431702 571399 431704
rect 546401 431699 546467 431702
rect 571333 431699 571399 431702
rect 580809 431626 580875 431629
rect 583520 431626 584960 431716
rect 580809 431624 584960 431626
rect 580809 431568 580814 431624
rect 580870 431568 584960 431624
rect 580809 431566 584960 431568
rect 580809 431563 580875 431566
rect 583520 431476 584960 431566
rect 64454 431156 64460 431220
rect 64524 431156 64530 431220
rect 92422 431156 92428 431220
rect 92492 431156 92498 431220
rect 148358 431156 148364 431220
rect 148428 431156 148434 431220
rect 176326 431156 176332 431220
rect 176396 431156 176402 431220
rect 260414 431156 260420 431220
rect 260484 431156 260490 431220
rect 288382 431156 288388 431220
rect 288452 431156 288458 431220
rect 344318 431156 344324 431220
rect 344388 431156 344394 431220
rect 372286 431156 372292 431220
rect 372356 431156 372362 431220
rect 456374 431156 456380 431220
rect 456444 431156 456450 431220
rect 484342 431156 484348 431220
rect 484412 431156 484418 431220
rect 492622 431156 492628 431220
rect 492692 431156 492698 431220
rect 520590 431156 520596 431220
rect 520660 431156 520666 431220
rect -960 423452 480 423692
rect 13721 423330 13787 423333
rect 64454 423330 64460 423332
rect 13721 423328 64460 423330
rect 13721 423272 13726 423328
rect 13782 423272 64460 423328
rect 13721 423270 64460 423272
rect 13721 423267 13787 423270
rect 64454 423268 64460 423270
rect 64524 423268 64530 423332
rect 70301 423330 70367 423333
rect 122833 423330 122899 423333
rect 70301 423328 122899 423330
rect 70301 423272 70306 423328
rect 70362 423272 122838 423328
rect 122894 423272 122899 423328
rect 70301 423270 122899 423272
rect 70301 423267 70367 423270
rect 122833 423267 122899 423270
rect 126881 423330 126947 423333
rect 176326 423330 176332 423332
rect 126881 423328 176332 423330
rect 126881 423272 126886 423328
rect 126942 423272 176332 423328
rect 126881 423270 176332 423272
rect 126881 423267 126947 423270
rect 176326 423268 176332 423270
rect 176396 423268 176402 423332
rect 182081 423330 182147 423333
rect 234705 423330 234771 423333
rect 182081 423328 234771 423330
rect 182081 423272 182086 423328
rect 182142 423272 234710 423328
rect 234766 423272 234771 423328
rect 182081 423270 234771 423272
rect 182081 423267 182147 423270
rect 234705 423267 234771 423270
rect 266261 423330 266327 423333
rect 318793 423330 318859 423333
rect 266261 423328 318859 423330
rect 266261 423272 266266 423328
rect 266322 423272 318798 423328
rect 318854 423272 318859 423328
rect 266261 423270 318859 423272
rect 266261 423267 266327 423270
rect 318793 423267 318859 423270
rect 322841 423330 322907 423333
rect 372286 423330 372292 423332
rect 322841 423328 372292 423330
rect 322841 423272 322846 423328
rect 322902 423272 372292 423328
rect 322841 423270 372292 423272
rect 322841 423267 322907 423270
rect 372286 423268 372292 423270
rect 372356 423268 372362 423332
rect 378041 423330 378107 423333
rect 430573 423330 430639 423333
rect 378041 423328 430639 423330
rect 378041 423272 378046 423328
rect 378102 423272 430578 423328
rect 430634 423272 430639 423328
rect 378041 423270 430639 423272
rect 378041 423267 378107 423270
rect 430573 423267 430639 423270
rect 462221 423330 462287 423333
rect 514753 423330 514819 423333
rect 462221 423328 514819 423330
rect 462221 423272 462226 423328
rect 462282 423272 514758 423328
rect 514814 423272 514819 423328
rect 462221 423270 514819 423272
rect 462221 423267 462287 423270
rect 514753 423267 514819 423270
rect 520590 423268 520596 423332
rect 520660 423330 520666 423332
rect 571333 423330 571399 423333
rect 520660 423328 571399 423330
rect 520660 423272 571338 423328
rect 571394 423272 571399 423328
rect 520660 423270 571399 423272
rect 520660 423268 520666 423270
rect 571333 423267 571399 423270
rect 42701 423194 42767 423197
rect 92422 423194 92428 423196
rect 42701 423192 92428 423194
rect 42701 423136 42706 423192
rect 42762 423136 92428 423192
rect 42701 423134 92428 423136
rect 42701 423131 42767 423134
rect 92422 423132 92428 423134
rect 92492 423132 92498 423196
rect 97901 423194 97967 423197
rect 148358 423194 148364 423196
rect 97901 423192 148364 423194
rect 97901 423136 97906 423192
rect 97962 423136 148364 423192
rect 97901 423134 148364 423136
rect 97901 423131 97967 423134
rect 148358 423132 148364 423134
rect 148428 423132 148434 423196
rect 154481 423194 154547 423197
rect 207013 423194 207079 423197
rect 154481 423192 207079 423194
rect 154481 423136 154486 423192
rect 154542 423136 207018 423192
rect 207074 423136 207079 423192
rect 154481 423134 207079 423136
rect 154481 423131 154547 423134
rect 207013 423131 207079 423134
rect 209681 423194 209747 423197
rect 260414 423194 260420 423196
rect 209681 423192 260420 423194
rect 209681 423136 209686 423192
rect 209742 423136 260420 423192
rect 209681 423134 260420 423136
rect 209681 423131 209747 423134
rect 260414 423132 260420 423134
rect 260484 423132 260490 423196
rect 293861 423194 293927 423197
rect 344318 423194 344324 423196
rect 293861 423192 344324 423194
rect 293861 423136 293866 423192
rect 293922 423136 344324 423192
rect 293861 423134 344324 423136
rect 293861 423131 293927 423134
rect 344318 423132 344324 423134
rect 344388 423132 344394 423196
rect 350441 423194 350507 423197
rect 402973 423194 403039 423197
rect 350441 423192 403039 423194
rect 350441 423136 350446 423192
rect 350502 423136 402978 423192
rect 403034 423136 403039 423192
rect 350441 423134 403039 423136
rect 350441 423131 350507 423134
rect 402973 423131 403039 423134
rect 405641 423194 405707 423197
rect 456374 423194 456380 423196
rect 405641 423192 456380 423194
rect 405641 423136 405646 423192
rect 405702 423136 456380 423192
rect 405641 423134 456380 423136
rect 405641 423131 405707 423134
rect 456374 423132 456380 423134
rect 456444 423132 456450 423196
rect 492622 423132 492628 423196
rect 492692 423194 492698 423196
rect 542353 423194 542419 423197
rect 492692 423192 542419 423194
rect 492692 423136 542358 423192
rect 542414 423136 542419 423192
rect 492692 423134 542419 423136
rect 492692 423132 492698 423134
rect 542353 423131 542419 423134
rect 238661 423058 238727 423061
rect 288382 423058 288388 423060
rect 238661 423056 288388 423058
rect 238661 423000 238666 423056
rect 238722 423000 288388 423056
rect 238661 422998 288388 423000
rect 238661 422995 238727 422998
rect 288382 422996 288388 422998
rect 288452 422996 288458 423060
rect 434621 423058 434687 423061
rect 484342 423058 484348 423060
rect 434621 423056 484348 423058
rect 434621 423000 434626 423056
rect 434682 423000 484348 423056
rect 434621 422998 484348 423000
rect 434621 422995 434687 422998
rect 484342 422996 484348 422998
rect 484412 422996 484418 423060
rect 110597 419522 110663 419525
rect 128302 419522 128308 419524
rect 110597 419520 128308 419522
rect 110597 419464 110602 419520
rect 110658 419464 128308 419520
rect 110597 419462 128308 419464
rect 110597 419459 110663 419462
rect 128302 419460 128308 419462
rect 128372 419460 128378 419524
rect 156321 419522 156387 419525
rect 194726 419522 194732 419524
rect 156321 419520 194732 419522
rect 156321 419464 156326 419520
rect 156382 419464 194732 419520
rect 156321 419462 194732 419464
rect 156321 419459 156387 419462
rect 194726 419460 194732 419462
rect 194796 419460 194802 419524
rect 352649 419522 352715 419525
rect 390870 419522 390876 419524
rect 352649 419520 390876 419522
rect 352649 419464 352654 419520
rect 352710 419464 390876 419520
rect 352649 419462 390876 419464
rect 352649 419459 352715 419462
rect 390870 419460 390876 419462
rect 390940 419460 390946 419524
rect 583520 418148 584960 418388
rect 81382 414428 81388 414492
rect 81452 414490 81458 414492
rect 81985 414490 82051 414493
rect 81452 414488 82051 414490
rect 81452 414432 81990 414488
rect 82046 414432 82051 414488
rect 81452 414430 82051 414432
rect 81452 414428 81458 414430
rect 81985 414427 82051 414430
rect 165654 414428 165660 414492
rect 165724 414490 165730 414492
rect 165981 414490 166047 414493
rect 165724 414488 166047 414490
rect 165724 414432 165986 414488
rect 166042 414432 166047 414488
rect 165724 414430 166047 414432
rect 165724 414428 165730 414430
rect 165981 414427 166047 414430
rect 259494 414428 259500 414492
rect 259564 414490 259570 414492
rect 260373 414490 260439 414493
rect 259564 414488 260439 414490
rect 259564 414432 260378 414488
rect 260434 414432 260439 414488
rect 259564 414430 260439 414432
rect 259564 414428 259570 414430
rect 260373 414427 260439 414430
rect 361614 414428 361620 414492
rect 361684 414490 361690 414492
rect 361941 414490 362007 414493
rect 361684 414488 362007 414490
rect 361684 414432 361946 414488
rect 362002 414432 362007 414488
rect 361684 414430 362007 414432
rect 361684 414428 361690 414430
rect 361941 414427 362007 414430
rect 445702 414428 445708 414492
rect 445772 414490 445778 414492
rect 446029 414490 446095 414493
rect 445772 414488 446095 414490
rect 445772 414432 446034 414488
rect 446090 414432 446095 414488
rect 445772 414430 446095 414432
rect 445772 414428 445778 414430
rect 446029 414427 446095 414430
rect 455454 414428 455460 414492
rect 455524 414490 455530 414492
rect 456333 414490 456399 414493
rect 455524 414488 456399 414490
rect 455524 414432 456338 414488
rect 456394 414432 456399 414488
rect 455524 414430 456399 414432
rect 455524 414428 455530 414430
rect 456333 414427 456399 414430
rect 557574 414428 557580 414492
rect 557644 414490 557650 414492
rect 557993 414490 558059 414493
rect 557644 414488 558059 414490
rect 557644 414432 557998 414488
rect 558054 414432 558059 414488
rect 557644 414430 558059 414432
rect 557644 414428 557650 414430
rect 557993 414427 558059 414430
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 580901 404970 580967 404973
rect 583520 404970 584960 405060
rect 580901 404968 584960 404970
rect 580901 404912 580906 404968
rect 580962 404912 584960 404968
rect 580901 404910 584960 404912
rect 580901 404907 580967 404910
rect 583520 404820 584960 404910
rect 13537 404290 13603 404293
rect 38653 404290 38719 404293
rect 66253 404290 66319 404293
rect 13537 404288 16100 404290
rect 13537 404232 13542 404288
rect 13598 404232 16100 404288
rect 13537 404230 16100 404232
rect 36892 404288 38719 404290
rect 36892 404232 38658 404288
rect 38714 404232 38719 404288
rect 64860 404288 66319 404290
rect 36892 404230 38719 404232
rect 13537 404227 13603 404230
rect 38653 404227 38719 404230
rect 44590 403748 44650 404260
rect 64860 404232 66258 404288
rect 66314 404232 66319 404288
rect 64860 404230 66319 404232
rect 66253 404227 66319 404230
rect 70301 404290 70367 404293
rect 95233 404290 95299 404293
rect 70301 404288 72036 404290
rect 70301 404232 70306 404288
rect 70362 404232 72036 404288
rect 70301 404230 72036 404232
rect 92828 404288 95299 404290
rect 92828 404232 95238 404288
rect 95294 404232 95299 404288
rect 92828 404230 95299 404232
rect 70301 404227 70367 404230
rect 95233 404227 95299 404230
rect 97901 404290 97967 404293
rect 122833 404290 122899 404293
rect 150433 404290 150499 404293
rect 97901 404288 100188 404290
rect 97901 404232 97906 404288
rect 97962 404232 100188 404288
rect 97901 404230 100188 404232
rect 120796 404288 122899 404290
rect 120796 404232 122838 404288
rect 122894 404232 122899 404288
rect 148948 404288 150499 404290
rect 120796 404230 122899 404232
rect 97901 404227 97967 404230
rect 122833 404227 122899 404230
rect 128494 403748 128554 404260
rect 148948 404232 150438 404288
rect 150494 404232 150499 404288
rect 148948 404230 150499 404232
rect 150433 404227 150499 404230
rect 154481 404290 154547 404293
rect 178033 404290 178099 404293
rect 154481 404288 156124 404290
rect 154481 404232 154486 404288
rect 154542 404232 156124 404288
rect 154481 404230 156124 404232
rect 176916 404288 178099 404290
rect 176916 404232 178038 404288
rect 178094 404232 178099 404288
rect 176916 404230 178099 404232
rect 154481 404227 154547 404230
rect 178033 404227 178099 404230
rect 182081 404290 182147 404293
rect 207013 404290 207079 404293
rect 234705 404290 234771 404293
rect 262213 404290 262279 404293
rect 182081 404288 184092 404290
rect 182081 404232 182086 404288
rect 182142 404232 184092 404288
rect 182081 404230 184092 404232
rect 204884 404288 207079 404290
rect 204884 404232 207018 404288
rect 207074 404232 207079 404288
rect 232852 404288 234771 404290
rect 204884 404230 207079 404232
rect 182081 404227 182147 404230
rect 207013 404227 207079 404230
rect 212582 403748 212642 404260
rect 232852 404232 234710 404288
rect 234766 404232 234771 404288
rect 260820 404288 262279 404290
rect 232852 404230 234771 404232
rect 234705 404227 234771 404230
rect 240550 403748 240610 404260
rect 260820 404232 262218 404288
rect 262274 404232 262279 404288
rect 260820 404230 262279 404232
rect 262213 404227 262279 404230
rect 266261 404290 266327 404293
rect 291193 404290 291259 404293
rect 318793 404290 318859 404293
rect 346393 404290 346459 404293
rect 266261 404288 268180 404290
rect 266261 404232 266266 404288
rect 266322 404232 268180 404288
rect 266261 404230 268180 404232
rect 288788 404288 291259 404290
rect 288788 404232 291198 404288
rect 291254 404232 291259 404288
rect 316940 404288 318859 404290
rect 288788 404230 291259 404232
rect 266261 404227 266327 404230
rect 291193 404227 291259 404230
rect 296486 403748 296546 404260
rect 316940 404232 318798 404288
rect 318854 404232 318859 404288
rect 344908 404288 346459 404290
rect 316940 404230 318859 404232
rect 318793 404227 318859 404230
rect 324638 403748 324698 404260
rect 344908 404232 346398 404288
rect 346454 404232 346459 404288
rect 344908 404230 346459 404232
rect 346393 404227 346459 404230
rect 350441 404290 350507 404293
rect 375373 404290 375439 404293
rect 350441 404288 352084 404290
rect 350441 404232 350446 404288
rect 350502 404232 352084 404288
rect 350441 404230 352084 404232
rect 372876 404288 375439 404290
rect 372876 404232 375378 404288
rect 375434 404232 375439 404288
rect 372876 404230 375439 404232
rect 350441 404227 350507 404230
rect 375373 404227 375439 404230
rect 378041 404290 378107 404293
rect 402973 404290 403039 404293
rect 430573 404290 430639 404293
rect 458173 404290 458239 404293
rect 378041 404288 380052 404290
rect 378041 404232 378046 404288
rect 378102 404232 380052 404288
rect 378041 404230 380052 404232
rect 400844 404288 403039 404290
rect 400844 404232 402978 404288
rect 403034 404232 403039 404288
rect 428812 404288 430639 404290
rect 400844 404230 403039 404232
rect 378041 404227 378107 404230
rect 402973 404227 403039 404230
rect 408542 403748 408602 404260
rect 428812 404232 430578 404288
rect 430634 404232 430639 404288
rect 456964 404288 458239 404290
rect 428812 404230 430639 404232
rect 430573 404227 430639 404230
rect 436510 403748 436570 404260
rect 456964 404232 458178 404288
rect 458234 404232 458239 404288
rect 456964 404230 458239 404232
rect 458173 404227 458239 404230
rect 462221 404290 462287 404293
rect 487153 404290 487219 404293
rect 514753 404290 514819 404293
rect 542353 404290 542419 404293
rect 462221 404288 464140 404290
rect 462221 404232 462226 404288
rect 462282 404232 464140 404288
rect 462221 404230 464140 404232
rect 484932 404288 487219 404290
rect 484932 404232 487158 404288
rect 487214 404232 487219 404288
rect 512900 404288 514819 404290
rect 484932 404230 487219 404232
rect 462221 404227 462287 404230
rect 487153 404227 487219 404230
rect 492630 403748 492690 404260
rect 512900 404232 514758 404288
rect 514814 404232 514819 404288
rect 540868 404288 542419 404290
rect 512900 404230 514819 404232
rect 514753 404227 514819 404230
rect 520598 403748 520658 404260
rect 540868 404232 542358 404288
rect 542414 404232 542419 404288
rect 540868 404230 542419 404232
rect 542353 404227 542419 404230
rect 546401 404290 546467 404293
rect 571333 404290 571399 404293
rect 546401 404288 548044 404290
rect 546401 404232 546406 404288
rect 546462 404232 548044 404288
rect 546401 404230 548044 404232
rect 568836 404288 571399 404290
rect 568836 404232 571338 404288
rect 571394 404232 571399 404288
rect 568836 404230 571399 404232
rect 546401 404227 546467 404230
rect 571333 404227 571399 404230
rect 44582 403684 44588 403748
rect 44652 403684 44658 403748
rect 128486 403684 128492 403748
rect 128556 403684 128562 403748
rect 212574 403684 212580 403748
rect 212644 403684 212650 403748
rect 240542 403684 240548 403748
rect 240612 403684 240618 403748
rect 296478 403684 296484 403748
rect 296548 403684 296554 403748
rect 324630 403684 324636 403748
rect 324700 403684 324706 403748
rect 408534 403684 408540 403748
rect 408604 403684 408610 403748
rect 436502 403684 436508 403748
rect 436572 403684 436578 403748
rect 492622 403684 492628 403748
rect 492692 403684 492698 403748
rect 520590 403684 520596 403748
rect 520660 403684 520666 403748
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 13537 395994 13603 395997
rect 66253 395994 66319 395997
rect 13537 395992 66319 395994
rect 13537 395936 13542 395992
rect 13598 395936 66258 395992
rect 66314 395936 66319 395992
rect 13537 395934 66319 395936
rect 13537 395931 13603 395934
rect 66253 395931 66319 395934
rect 70301 395994 70367 395997
rect 122833 395994 122899 395997
rect 70301 395992 122899 395994
rect 70301 395936 70306 395992
rect 70362 395936 122838 395992
rect 122894 395936 122899 395992
rect 70301 395934 122899 395936
rect 70301 395931 70367 395934
rect 122833 395931 122899 395934
rect 128486 395932 128492 395996
rect 128556 395994 128562 395996
rect 178033 395994 178099 395997
rect 128556 395992 178099 395994
rect 128556 395936 178038 395992
rect 178094 395936 178099 395992
rect 128556 395934 178099 395936
rect 128556 395932 128562 395934
rect 178033 395931 178099 395934
rect 182081 395994 182147 395997
rect 234705 395994 234771 395997
rect 182081 395992 234771 395994
rect 182081 395936 182086 395992
rect 182142 395936 234710 395992
rect 234766 395936 234771 395992
rect 182081 395934 234771 395936
rect 182081 395931 182147 395934
rect 234705 395931 234771 395934
rect 266261 395994 266327 395997
rect 318793 395994 318859 395997
rect 266261 395992 318859 395994
rect 266261 395936 266266 395992
rect 266322 395936 318798 395992
rect 318854 395936 318859 395992
rect 266261 395934 318859 395936
rect 266261 395931 266327 395934
rect 318793 395931 318859 395934
rect 350441 395994 350507 395997
rect 402973 395994 403039 395997
rect 350441 395992 403039 395994
rect 350441 395936 350446 395992
rect 350502 395936 402978 395992
rect 403034 395936 403039 395992
rect 350441 395934 403039 395936
rect 350441 395931 350507 395934
rect 402973 395931 403039 395934
rect 408534 395932 408540 395996
rect 408604 395994 408610 395996
rect 458173 395994 458239 395997
rect 408604 395992 458239 395994
rect 408604 395936 458178 395992
rect 458234 395936 458239 395992
rect 408604 395934 458239 395936
rect 408604 395932 408610 395934
rect 458173 395931 458239 395934
rect 462221 395994 462287 395997
rect 514753 395994 514819 395997
rect 462221 395992 514819 395994
rect 462221 395936 462226 395992
rect 462282 395936 514758 395992
rect 514814 395936 514819 395992
rect 462221 395934 514819 395936
rect 462221 395931 462287 395934
rect 514753 395931 514819 395934
rect 520590 395932 520596 395996
rect 520660 395994 520666 395996
rect 571333 395994 571399 395997
rect 520660 395992 571399 395994
rect 520660 395936 571338 395992
rect 571394 395936 571399 395992
rect 520660 395934 571399 395936
rect 520660 395932 520666 395934
rect 571333 395931 571399 395934
rect 44582 395796 44588 395860
rect 44652 395858 44658 395860
rect 95233 395858 95299 395861
rect 44652 395856 95299 395858
rect 44652 395800 95238 395856
rect 95294 395800 95299 395856
rect 44652 395798 95299 395800
rect 44652 395796 44658 395798
rect 95233 395795 95299 395798
rect 97901 395858 97967 395861
rect 150433 395858 150499 395861
rect 97901 395856 150499 395858
rect 97901 395800 97906 395856
rect 97962 395800 150438 395856
rect 150494 395800 150499 395856
rect 97901 395798 150499 395800
rect 97901 395795 97967 395798
rect 150433 395795 150499 395798
rect 154481 395858 154547 395861
rect 207013 395858 207079 395861
rect 154481 395856 207079 395858
rect 154481 395800 154486 395856
rect 154542 395800 207018 395856
rect 207074 395800 207079 395856
rect 154481 395798 207079 395800
rect 154481 395795 154547 395798
rect 207013 395795 207079 395798
rect 240542 395796 240548 395860
rect 240612 395858 240618 395860
rect 291193 395858 291259 395861
rect 240612 395856 291259 395858
rect 240612 395800 291198 395856
rect 291254 395800 291259 395856
rect 240612 395798 291259 395800
rect 240612 395796 240618 395798
rect 291193 395795 291259 395798
rect 324630 395796 324636 395860
rect 324700 395858 324706 395860
rect 375373 395858 375439 395861
rect 324700 395856 375439 395858
rect 324700 395800 375378 395856
rect 375434 395800 375439 395856
rect 324700 395798 375439 395800
rect 324700 395796 324706 395798
rect 375373 395795 375439 395798
rect 378041 395858 378107 395861
rect 430573 395858 430639 395861
rect 378041 395856 430639 395858
rect 378041 395800 378046 395856
rect 378102 395800 430578 395856
rect 430634 395800 430639 395856
rect 378041 395798 430639 395800
rect 378041 395795 378107 395798
rect 430573 395795 430639 395798
rect 436502 395796 436508 395860
rect 436572 395858 436578 395860
rect 487153 395858 487219 395861
rect 436572 395856 487219 395858
rect 436572 395800 487158 395856
rect 487214 395800 487219 395856
rect 436572 395798 487219 395800
rect 436572 395796 436578 395798
rect 487153 395795 487219 395798
rect 492622 395796 492628 395860
rect 492692 395858 492698 395860
rect 542353 395858 542419 395861
rect 492692 395856 542419 395858
rect 492692 395800 542358 395856
rect 542414 395800 542419 395856
rect 492692 395798 542419 395800
rect 492692 395796 492698 395798
rect 542353 395795 542419 395798
rect 212574 395660 212580 395724
rect 212644 395722 212650 395724
rect 262213 395722 262279 395725
rect 212644 395720 262279 395722
rect 212644 395664 262218 395720
rect 262274 395664 262279 395720
rect 212644 395662 262279 395664
rect 212644 395660 212650 395662
rect 262213 395659 262279 395662
rect 296846 395660 296852 395724
rect 296916 395722 296922 395724
rect 346393 395722 346459 395725
rect 296916 395720 346459 395722
rect 296916 395664 346398 395720
rect 346454 395664 346459 395720
rect 296916 395662 346459 395664
rect 296916 395660 296922 395662
rect 346393 395659 346459 395662
rect 64597 391914 64663 391917
rect 81382 391914 81388 391916
rect 64597 391912 81388 391914
rect 64597 391856 64602 391912
rect 64658 391856 81388 391912
rect 64597 391854 81388 391856
rect 64597 391851 64663 391854
rect 81382 391852 81388 391854
rect 81452 391852 81458 391916
rect 148593 391914 148659 391917
rect 165654 391914 165660 391916
rect 148593 391912 165660 391914
rect 148593 391856 148598 391912
rect 148654 391856 165660 391912
rect 148593 391854 165660 391856
rect 148593 391851 148659 391854
rect 165654 391852 165660 391854
rect 165724 391852 165730 391916
rect 222653 391914 222719 391917
rect 259494 391914 259500 391916
rect 222653 391912 259500 391914
rect 222653 391856 222658 391912
rect 222714 391856 259500 391912
rect 222653 391854 259500 391856
rect 222653 391851 222719 391854
rect 259494 391852 259500 391854
rect 259564 391852 259570 391916
rect 344645 391914 344711 391917
rect 361614 391914 361620 391916
rect 344645 391912 361620 391914
rect 344645 391856 344650 391912
rect 344706 391856 361620 391912
rect 344645 391854 361620 391856
rect 344645 391851 344711 391854
rect 361614 391852 361620 391854
rect 361684 391852 361690 391916
rect 418337 391914 418403 391917
rect 455454 391914 455460 391916
rect 418337 391912 455460 391914
rect 418337 391856 418342 391912
rect 418398 391856 455460 391912
rect 418337 391854 455460 391856
rect 418337 391851 418403 391854
rect 455454 391852 455460 391854
rect 455524 391852 455530 391916
rect 540605 391914 540671 391917
rect 557574 391914 557580 391916
rect 540605 391912 557580 391914
rect 540605 391856 540610 391912
rect 540666 391856 557580 391912
rect 540605 391854 557580 391856
rect 540605 391851 540671 391854
rect 557574 391852 557580 391854
rect 557644 391852 557650 391916
rect 428641 391778 428707 391781
rect 445702 391778 445708 391780
rect 428641 391776 445708 391778
rect 428641 391720 428646 391776
rect 428702 391720 445708 391776
rect 428641 391718 445708 391720
rect 428641 391715 428707 391718
rect 445702 391716 445708 391718
rect 445772 391716 445778 391780
rect 583520 391628 584960 391868
rect 128302 387364 128308 387428
rect 128372 387426 128378 387428
rect 128445 387426 128511 387429
rect 194777 387428 194843 387429
rect 194726 387426 194732 387428
rect 128372 387424 128511 387426
rect 128372 387368 128450 387424
rect 128506 387368 128511 387424
rect 128372 387366 128511 387368
rect 194686 387366 194732 387426
rect 194796 387424 194843 387428
rect 194838 387368 194843 387424
rect 128372 387364 128378 387366
rect 128445 387363 128511 387366
rect 194726 387364 194732 387366
rect 194796 387364 194843 387368
rect 194777 387363 194843 387364
rect 390829 387428 390895 387429
rect 390829 387424 390876 387428
rect 390940 387426 390946 387428
rect 390829 387368 390834 387424
rect 390829 387364 390876 387368
rect 390940 387366 390986 387426
rect 390940 387364 390946 387366
rect 390829 387363 390895 387364
rect -960 384284 480 384524
rect 579797 378450 579863 378453
rect 583520 378450 584960 378540
rect 579797 378448 584960 378450
rect 579797 378392 579802 378448
rect 579858 378392 584960 378448
rect 579797 378390 584960 378392
rect 579797 378387 579863 378390
rect 583520 378300 584960 378390
rect 13537 377770 13603 377773
rect 38653 377770 38719 377773
rect 13537 377768 16100 377770
rect 13537 377712 13542 377768
rect 13598 377712 16100 377768
rect 13537 377710 16100 377712
rect 36892 377768 38719 377770
rect 36892 377712 38658 377768
rect 38714 377712 38719 377768
rect 36892 377710 38719 377712
rect 13537 377707 13603 377710
rect 38653 377707 38719 377710
rect 42701 377770 42767 377773
rect 66253 377770 66319 377773
rect 42701 377768 44068 377770
rect 42701 377712 42706 377768
rect 42762 377712 44068 377768
rect 42701 377710 44068 377712
rect 64860 377768 66319 377770
rect 64860 377712 66258 377768
rect 66314 377712 66319 377768
rect 64860 377710 66319 377712
rect 42701 377707 42767 377710
rect 66253 377707 66319 377710
rect 70301 377770 70367 377773
rect 95233 377770 95299 377773
rect 70301 377768 72036 377770
rect 70301 377712 70306 377768
rect 70362 377712 72036 377768
rect 70301 377710 72036 377712
rect 92828 377768 95299 377770
rect 92828 377712 95238 377768
rect 95294 377712 95299 377768
rect 92828 377710 95299 377712
rect 70301 377707 70367 377710
rect 95233 377707 95299 377710
rect 97901 377770 97967 377773
rect 122833 377770 122899 377773
rect 97901 377768 100188 377770
rect 97901 377712 97906 377768
rect 97962 377712 100188 377768
rect 97901 377710 100188 377712
rect 120796 377768 122899 377770
rect 120796 377712 122838 377768
rect 122894 377712 122899 377768
rect 120796 377710 122899 377712
rect 97901 377707 97967 377710
rect 122833 377707 122899 377710
rect 126881 377770 126947 377773
rect 150433 377770 150499 377773
rect 126881 377768 128156 377770
rect 126881 377712 126886 377768
rect 126942 377712 128156 377768
rect 126881 377710 128156 377712
rect 148948 377768 150499 377770
rect 148948 377712 150438 377768
rect 150494 377712 150499 377768
rect 148948 377710 150499 377712
rect 126881 377707 126947 377710
rect 150433 377707 150499 377710
rect 154481 377770 154547 377773
rect 182081 377770 182147 377773
rect 207013 377770 207079 377773
rect 154481 377768 156124 377770
rect 154481 377712 154486 377768
rect 154542 377712 156124 377768
rect 182081 377768 184092 377770
rect 154481 377710 156124 377712
rect 154481 377707 154547 377710
rect 176334 377228 176394 377740
rect 182081 377712 182086 377768
rect 182142 377712 184092 377768
rect 182081 377710 184092 377712
rect 204884 377768 207079 377770
rect 204884 377712 207018 377768
rect 207074 377712 207079 377768
rect 204884 377710 207079 377712
rect 182081 377707 182147 377710
rect 207013 377707 207079 377710
rect 209681 377770 209747 377773
rect 234705 377770 234771 377773
rect 209681 377768 212060 377770
rect 209681 377712 209686 377768
rect 209742 377712 212060 377768
rect 209681 377710 212060 377712
rect 232852 377768 234771 377770
rect 232852 377712 234710 377768
rect 234766 377712 234771 377768
rect 232852 377710 234771 377712
rect 209681 377707 209747 377710
rect 234705 377707 234771 377710
rect 238661 377770 238727 377773
rect 262213 377770 262279 377773
rect 238661 377768 240212 377770
rect 238661 377712 238666 377768
rect 238722 377712 240212 377768
rect 238661 377710 240212 377712
rect 260820 377768 262279 377770
rect 260820 377712 262218 377768
rect 262274 377712 262279 377768
rect 260820 377710 262279 377712
rect 238661 377707 238727 377710
rect 262213 377707 262279 377710
rect 266261 377770 266327 377773
rect 291193 377770 291259 377773
rect 266261 377768 268180 377770
rect 266261 377712 266266 377768
rect 266322 377712 268180 377768
rect 266261 377710 268180 377712
rect 288788 377768 291259 377770
rect 288788 377712 291198 377768
rect 291254 377712 291259 377768
rect 288788 377710 291259 377712
rect 266261 377707 266327 377710
rect 291193 377707 291259 377710
rect 293861 377770 293927 377773
rect 318793 377770 318859 377773
rect 293861 377768 296148 377770
rect 293861 377712 293866 377768
rect 293922 377712 296148 377768
rect 293861 377710 296148 377712
rect 316940 377768 318859 377770
rect 316940 377712 318798 377768
rect 318854 377712 318859 377768
rect 316940 377710 318859 377712
rect 293861 377707 293927 377710
rect 318793 377707 318859 377710
rect 322841 377770 322907 377773
rect 346393 377770 346459 377773
rect 322841 377768 324116 377770
rect 322841 377712 322846 377768
rect 322902 377712 324116 377768
rect 322841 377710 324116 377712
rect 344908 377768 346459 377770
rect 344908 377712 346398 377768
rect 346454 377712 346459 377768
rect 344908 377710 346459 377712
rect 322841 377707 322907 377710
rect 346393 377707 346459 377710
rect 350441 377770 350507 377773
rect 375373 377770 375439 377773
rect 350441 377768 352084 377770
rect 350441 377712 350446 377768
rect 350502 377712 352084 377768
rect 350441 377710 352084 377712
rect 372876 377768 375439 377770
rect 372876 377712 375378 377768
rect 375434 377712 375439 377768
rect 372876 377710 375439 377712
rect 350441 377707 350507 377710
rect 375373 377707 375439 377710
rect 378041 377770 378107 377773
rect 402973 377770 403039 377773
rect 378041 377768 380052 377770
rect 378041 377712 378046 377768
rect 378102 377712 380052 377768
rect 378041 377710 380052 377712
rect 400844 377768 403039 377770
rect 400844 377712 402978 377768
rect 403034 377712 403039 377768
rect 400844 377710 403039 377712
rect 378041 377707 378107 377710
rect 402973 377707 403039 377710
rect 405641 377770 405707 377773
rect 430573 377770 430639 377773
rect 405641 377768 408204 377770
rect 405641 377712 405646 377768
rect 405702 377712 408204 377768
rect 405641 377710 408204 377712
rect 428812 377768 430639 377770
rect 428812 377712 430578 377768
rect 430634 377712 430639 377768
rect 428812 377710 430639 377712
rect 405641 377707 405707 377710
rect 430573 377707 430639 377710
rect 434621 377770 434687 377773
rect 462221 377770 462287 377773
rect 487153 377770 487219 377773
rect 434621 377768 436172 377770
rect 434621 377712 434626 377768
rect 434682 377712 436172 377768
rect 462221 377768 464140 377770
rect 434621 377710 436172 377712
rect 434621 377707 434687 377710
rect 456382 377228 456442 377740
rect 462221 377712 462226 377768
rect 462282 377712 464140 377768
rect 462221 377710 464140 377712
rect 484932 377768 487219 377770
rect 484932 377712 487158 377768
rect 487214 377712 487219 377768
rect 484932 377710 487219 377712
rect 462221 377707 462287 377710
rect 487153 377707 487219 377710
rect 489821 377770 489887 377773
rect 514753 377770 514819 377773
rect 489821 377768 492108 377770
rect 489821 377712 489826 377768
rect 489882 377712 492108 377768
rect 489821 377710 492108 377712
rect 512900 377768 514819 377770
rect 512900 377712 514758 377768
rect 514814 377712 514819 377768
rect 512900 377710 514819 377712
rect 489821 377707 489887 377710
rect 514753 377707 514819 377710
rect 518801 377770 518867 377773
rect 542353 377770 542419 377773
rect 518801 377768 520076 377770
rect 518801 377712 518806 377768
rect 518862 377712 520076 377768
rect 518801 377710 520076 377712
rect 540868 377768 542419 377770
rect 540868 377712 542358 377768
rect 542414 377712 542419 377768
rect 540868 377710 542419 377712
rect 518801 377707 518867 377710
rect 542353 377707 542419 377710
rect 546401 377770 546467 377773
rect 546401 377768 548044 377770
rect 546401 377712 546406 377768
rect 546462 377712 548044 377768
rect 546401 377710 548044 377712
rect 546401 377707 546467 377710
rect 568438 377228 568498 377740
rect 176326 377164 176332 377228
rect 176396 377164 176402 377228
rect 456374 377164 456380 377228
rect 456444 377164 456450 377228
rect 568430 377164 568436 377228
rect 568500 377164 568506 377228
rect -960 371228 480 371468
rect 13537 369338 13603 369341
rect 66253 369338 66319 369341
rect 13537 369336 66319 369338
rect 13537 369280 13542 369336
rect 13598 369280 66258 369336
rect 66314 369280 66319 369336
rect 13537 369278 66319 369280
rect 13537 369275 13603 369278
rect 66253 369275 66319 369278
rect 70301 369338 70367 369341
rect 122833 369338 122899 369341
rect 70301 369336 122899 369338
rect 70301 369280 70306 369336
rect 70362 369280 122838 369336
rect 122894 369280 122899 369336
rect 70301 369278 122899 369280
rect 70301 369275 70367 369278
rect 122833 369275 122899 369278
rect 126881 369338 126947 369341
rect 175222 369338 175228 369340
rect 126881 369336 175228 369338
rect 126881 369280 126886 369336
rect 126942 369280 175228 369336
rect 126881 369278 175228 369280
rect 126881 369275 126947 369278
rect 175222 369276 175228 369278
rect 175292 369276 175298 369340
rect 182081 369338 182147 369341
rect 234705 369338 234771 369341
rect 182081 369336 234771 369338
rect 182081 369280 182086 369336
rect 182142 369280 234710 369336
rect 234766 369280 234771 369336
rect 182081 369278 234771 369280
rect 182081 369275 182147 369278
rect 234705 369275 234771 369278
rect 238661 369338 238727 369341
rect 291193 369338 291259 369341
rect 238661 369336 291259 369338
rect 238661 369280 238666 369336
rect 238722 369280 291198 369336
rect 291254 369280 291259 369336
rect 238661 369278 291259 369280
rect 238661 369275 238727 369278
rect 291193 369275 291259 369278
rect 293861 369338 293927 369341
rect 346393 369338 346459 369341
rect 293861 369336 346459 369338
rect 293861 369280 293866 369336
rect 293922 369280 346398 369336
rect 346454 369280 346459 369336
rect 293861 369278 346459 369280
rect 293861 369275 293927 369278
rect 346393 369275 346459 369278
rect 350441 369338 350507 369341
rect 402973 369338 403039 369341
rect 350441 369336 403039 369338
rect 350441 369280 350446 369336
rect 350502 369280 402978 369336
rect 403034 369280 403039 369336
rect 350441 369278 403039 369280
rect 350441 369275 350507 369278
rect 402973 369275 403039 369278
rect 405641 369338 405707 369341
rect 455454 369338 455460 369340
rect 405641 369336 455460 369338
rect 405641 369280 405646 369336
rect 405702 369280 455460 369336
rect 405641 369278 455460 369280
rect 405641 369275 405707 369278
rect 455454 369276 455460 369278
rect 455524 369276 455530 369340
rect 462221 369338 462287 369341
rect 514753 369338 514819 369341
rect 462221 369336 514819 369338
rect 462221 369280 462226 369336
rect 462282 369280 514758 369336
rect 514814 369280 514819 369336
rect 462221 369278 514819 369280
rect 462221 369275 462287 369278
rect 514753 369275 514819 369278
rect 518801 369338 518867 369341
rect 566958 369338 566964 369340
rect 518801 369336 566964 369338
rect 518801 369280 518806 369336
rect 518862 369280 566964 369336
rect 518801 369278 566964 369280
rect 518801 369275 518867 369278
rect 566958 369276 566964 369278
rect 567028 369276 567034 369340
rect 110597 365666 110663 365669
rect 128302 365666 128308 365668
rect 110597 365664 128308 365666
rect 110597 365608 110602 365664
rect 110658 365608 128308 365664
rect 110597 365606 128308 365608
rect 110597 365603 110663 365606
rect 128302 365604 128308 365606
rect 128372 365604 128378 365668
rect 156321 365666 156387 365669
rect 194726 365666 194732 365668
rect 156321 365664 194732 365666
rect 156321 365608 156326 365664
rect 156382 365608 194732 365664
rect 156321 365606 194732 365608
rect 156321 365603 156387 365606
rect 194726 365604 194732 365606
rect 194796 365604 194802 365668
rect 352649 365666 352715 365669
rect 390870 365666 390876 365668
rect 352649 365664 390876 365666
rect 352649 365608 352654 365664
rect 352710 365608 390876 365664
rect 352649 365606 390876 365608
rect 352649 365603 352715 365606
rect 390870 365604 390876 365606
rect 390940 365604 390946 365668
rect 583520 364972 584960 365212
rect 165654 360436 165660 360500
rect 165724 360498 165730 360500
rect 165981 360498 166047 360501
rect 165724 360496 166047 360498
rect 165724 360440 165986 360496
rect 166042 360440 166047 360496
rect 165724 360438 166047 360440
rect 165724 360436 165730 360438
rect 165981 360435 166047 360438
rect 259494 360436 259500 360500
rect 259564 360498 259570 360500
rect 260373 360498 260439 360501
rect 259564 360496 260439 360498
rect 259564 360440 260378 360496
rect 260434 360440 260439 360496
rect 259564 360438 260439 360440
rect 259564 360436 259570 360438
rect 260373 360435 260439 360438
rect 361614 360436 361620 360500
rect 361684 360498 361690 360500
rect 361941 360498 362007 360501
rect 361684 360496 362007 360498
rect 361684 360440 361946 360496
rect 362002 360440 362007 360496
rect 361684 360438 362007 360440
rect 361684 360436 361690 360438
rect 361941 360435 362007 360438
rect 445702 360436 445708 360500
rect 445772 360498 445778 360500
rect 446029 360498 446095 360501
rect 445772 360496 446095 360498
rect 445772 360440 446034 360496
rect 446090 360440 446095 360496
rect 445772 360438 446095 360440
rect 445772 360436 445778 360438
rect 446029 360435 446095 360438
rect 557574 360436 557580 360500
rect 557644 360498 557650 360500
rect 557993 360498 558059 360501
rect 557644 360496 558059 360498
rect 557644 360440 557998 360496
rect 558054 360440 558059 360496
rect 557644 360438 558059 360440
rect 557644 360436 557650 360438
rect 557993 360435 558059 360438
rect -960 358458 480 358548
rect 3785 358458 3851 358461
rect -960 358456 3851 358458
rect -960 358400 3790 358456
rect 3846 358400 3851 358456
rect -960 358398 3851 358400
rect -960 358308 480 358398
rect 3785 358395 3851 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 13537 350298 13603 350301
rect 38653 350298 38719 350301
rect 66253 350298 66319 350301
rect 13537 350296 16100 350298
rect 13537 350240 13542 350296
rect 13598 350240 16100 350296
rect 13537 350238 16100 350240
rect 36892 350296 38719 350298
rect 36892 350240 38658 350296
rect 38714 350240 38719 350296
rect 64860 350296 66319 350298
rect 36892 350238 38719 350240
rect 13537 350235 13603 350238
rect 38653 350235 38719 350238
rect 44590 349756 44650 350268
rect 64860 350240 66258 350296
rect 66314 350240 66319 350296
rect 64860 350238 66319 350240
rect 66253 350235 66319 350238
rect 70301 350298 70367 350301
rect 95233 350298 95299 350301
rect 70301 350296 72036 350298
rect 70301 350240 70306 350296
rect 70362 350240 72036 350296
rect 70301 350238 72036 350240
rect 92828 350296 95299 350298
rect 92828 350240 95238 350296
rect 95294 350240 95299 350296
rect 92828 350238 95299 350240
rect 70301 350235 70367 350238
rect 95233 350235 95299 350238
rect 97901 350298 97967 350301
rect 122833 350298 122899 350301
rect 150433 350298 150499 350301
rect 97901 350296 100188 350298
rect 97901 350240 97906 350296
rect 97962 350240 100188 350296
rect 97901 350238 100188 350240
rect 120796 350296 122899 350298
rect 120796 350240 122838 350296
rect 122894 350240 122899 350296
rect 148948 350296 150499 350298
rect 120796 350238 122899 350240
rect 97901 350235 97967 350238
rect 122833 350235 122899 350238
rect 128494 349756 128554 350268
rect 148948 350240 150438 350296
rect 150494 350240 150499 350296
rect 148948 350238 150499 350240
rect 150433 350235 150499 350238
rect 154481 350298 154547 350301
rect 178033 350298 178099 350301
rect 154481 350296 156124 350298
rect 154481 350240 154486 350296
rect 154542 350240 156124 350296
rect 154481 350238 156124 350240
rect 176916 350296 178099 350298
rect 176916 350240 178038 350296
rect 178094 350240 178099 350296
rect 176916 350238 178099 350240
rect 154481 350235 154547 350238
rect 178033 350235 178099 350238
rect 182081 350298 182147 350301
rect 207013 350298 207079 350301
rect 234705 350298 234771 350301
rect 262213 350298 262279 350301
rect 182081 350296 184092 350298
rect 182081 350240 182086 350296
rect 182142 350240 184092 350296
rect 182081 350238 184092 350240
rect 204884 350296 207079 350298
rect 204884 350240 207018 350296
rect 207074 350240 207079 350296
rect 232852 350296 234771 350298
rect 204884 350238 207079 350240
rect 182081 350235 182147 350238
rect 207013 350235 207079 350238
rect 212582 349756 212642 350268
rect 232852 350240 234710 350296
rect 234766 350240 234771 350296
rect 260820 350296 262279 350298
rect 232852 350238 234771 350240
rect 234705 350235 234771 350238
rect 240550 349756 240610 350268
rect 260820 350240 262218 350296
rect 262274 350240 262279 350296
rect 260820 350238 262279 350240
rect 262213 350235 262279 350238
rect 266261 350298 266327 350301
rect 291193 350298 291259 350301
rect 318793 350298 318859 350301
rect 346393 350298 346459 350301
rect 266261 350296 268180 350298
rect 266261 350240 266266 350296
rect 266322 350240 268180 350296
rect 266261 350238 268180 350240
rect 288788 350296 291259 350298
rect 288788 350240 291198 350296
rect 291254 350240 291259 350296
rect 316940 350296 318859 350298
rect 288788 350238 291259 350240
rect 266261 350235 266327 350238
rect 291193 350235 291259 350238
rect 296486 349756 296546 350268
rect 316940 350240 318798 350296
rect 318854 350240 318859 350296
rect 344908 350296 346459 350298
rect 316940 350238 318859 350240
rect 318793 350235 318859 350238
rect 324638 349756 324698 350268
rect 344908 350240 346398 350296
rect 346454 350240 346459 350296
rect 344908 350238 346459 350240
rect 346393 350235 346459 350238
rect 350441 350298 350507 350301
rect 375373 350298 375439 350301
rect 350441 350296 352084 350298
rect 350441 350240 350446 350296
rect 350502 350240 352084 350296
rect 350441 350238 352084 350240
rect 372876 350296 375439 350298
rect 372876 350240 375378 350296
rect 375434 350240 375439 350296
rect 372876 350238 375439 350240
rect 350441 350235 350507 350238
rect 375373 350235 375439 350238
rect 378041 350298 378107 350301
rect 402973 350298 403039 350301
rect 430573 350298 430639 350301
rect 458173 350298 458239 350301
rect 378041 350296 380052 350298
rect 378041 350240 378046 350296
rect 378102 350240 380052 350296
rect 378041 350238 380052 350240
rect 400844 350296 403039 350298
rect 400844 350240 402978 350296
rect 403034 350240 403039 350296
rect 428812 350296 430639 350298
rect 400844 350238 403039 350240
rect 378041 350235 378107 350238
rect 402973 350235 403039 350238
rect 408542 349756 408602 350268
rect 428812 350240 430578 350296
rect 430634 350240 430639 350296
rect 456964 350296 458239 350298
rect 428812 350238 430639 350240
rect 430573 350235 430639 350238
rect 436510 349756 436570 350268
rect 456964 350240 458178 350296
rect 458234 350240 458239 350296
rect 456964 350238 458239 350240
rect 458173 350235 458239 350238
rect 462221 350298 462287 350301
rect 487153 350298 487219 350301
rect 514753 350298 514819 350301
rect 542353 350298 542419 350301
rect 462221 350296 464140 350298
rect 462221 350240 462226 350296
rect 462282 350240 464140 350296
rect 462221 350238 464140 350240
rect 484932 350296 487219 350298
rect 484932 350240 487158 350296
rect 487214 350240 487219 350296
rect 512900 350296 514819 350298
rect 484932 350238 487219 350240
rect 462221 350235 462287 350238
rect 487153 350235 487219 350238
rect 492630 349756 492690 350268
rect 512900 350240 514758 350296
rect 514814 350240 514819 350296
rect 540868 350296 542419 350298
rect 512900 350238 514819 350240
rect 514753 350235 514819 350238
rect 520598 349756 520658 350268
rect 540868 350240 542358 350296
rect 542414 350240 542419 350296
rect 540868 350238 542419 350240
rect 542353 350235 542419 350238
rect 546401 350298 546467 350301
rect 571333 350298 571399 350301
rect 546401 350296 548044 350298
rect 546401 350240 546406 350296
rect 546462 350240 548044 350296
rect 546401 350238 548044 350240
rect 568836 350296 571399 350298
rect 568836 350240 571338 350296
rect 571394 350240 571399 350296
rect 568836 350238 571399 350240
rect 546401 350235 546467 350238
rect 571333 350235 571399 350238
rect 44582 349692 44588 349756
rect 44652 349692 44658 349756
rect 128486 349692 128492 349756
rect 128556 349692 128562 349756
rect 212574 349692 212580 349756
rect 212644 349692 212650 349756
rect 240542 349692 240548 349756
rect 240612 349692 240618 349756
rect 296478 349692 296484 349756
rect 296548 349692 296554 349756
rect 324630 349692 324636 349756
rect 324700 349692 324706 349756
rect 408534 349692 408540 349756
rect 408604 349692 408610 349756
rect 436502 349692 436508 349756
rect 436572 349692 436578 349756
rect 492622 349692 492628 349756
rect 492692 349692 492698 349756
rect 520590 349692 520596 349756
rect 520660 349692 520666 349756
rect -960 345402 480 345492
rect 2773 345402 2839 345405
rect -960 345400 2839 345402
rect -960 345344 2778 345400
rect 2834 345344 2839 345400
rect -960 345342 2839 345344
rect -960 345252 480 345342
rect 2773 345339 2839 345342
rect 13537 342002 13603 342005
rect 66253 342002 66319 342005
rect 13537 342000 66319 342002
rect 13537 341944 13542 342000
rect 13598 341944 66258 342000
rect 66314 341944 66319 342000
rect 13537 341942 66319 341944
rect 13537 341939 13603 341942
rect 66253 341939 66319 341942
rect 97901 342002 97967 342005
rect 150433 342002 150499 342005
rect 97901 342000 150499 342002
rect 97901 341944 97906 342000
rect 97962 341944 150438 342000
rect 150494 341944 150499 342000
rect 97901 341942 150499 341944
rect 97901 341939 97967 341942
rect 150433 341939 150499 341942
rect 182081 342002 182147 342005
rect 234705 342002 234771 342005
rect 182081 342000 234771 342002
rect 182081 341944 182086 342000
rect 182142 341944 234710 342000
rect 234766 341944 234771 342000
rect 182081 341942 234771 341944
rect 182081 341939 182147 341942
rect 234705 341939 234771 341942
rect 266261 342002 266327 342005
rect 318793 342002 318859 342005
rect 266261 342000 318859 342002
rect 266261 341944 266266 342000
rect 266322 341944 318798 342000
rect 318854 341944 318859 342000
rect 266261 341942 318859 341944
rect 266261 341939 266327 341942
rect 318793 341939 318859 341942
rect 350441 342002 350507 342005
rect 402973 342002 403039 342005
rect 350441 342000 403039 342002
rect 350441 341944 350446 342000
rect 350502 341944 402978 342000
rect 403034 341944 403039 342000
rect 350441 341942 403039 341944
rect 350441 341939 350507 341942
rect 402973 341939 403039 341942
rect 408534 341940 408540 342004
rect 408604 342002 408610 342004
rect 458173 342002 458239 342005
rect 408604 342000 458239 342002
rect 408604 341944 458178 342000
rect 458234 341944 458239 342000
rect 408604 341942 458239 341944
rect 408604 341940 408610 341942
rect 458173 341939 458239 341942
rect 462221 342002 462287 342005
rect 514753 342002 514819 342005
rect 462221 342000 514819 342002
rect 462221 341944 462226 342000
rect 462282 341944 514758 342000
rect 514814 341944 514819 342000
rect 462221 341942 514819 341944
rect 462221 341939 462287 341942
rect 514753 341939 514819 341942
rect 520590 341940 520596 342004
rect 520660 342002 520666 342004
rect 571333 342002 571399 342005
rect 520660 342000 571399 342002
rect 520660 341944 571338 342000
rect 571394 341944 571399 342000
rect 520660 341942 571399 341944
rect 520660 341940 520666 341942
rect 571333 341939 571399 341942
rect 70301 341866 70367 341869
rect 122833 341866 122899 341869
rect 70301 341864 122899 341866
rect 70301 341808 70306 341864
rect 70362 341808 122838 341864
rect 122894 341808 122899 341864
rect 70301 341806 122899 341808
rect 70301 341803 70367 341806
rect 122833 341803 122899 341806
rect 154481 341866 154547 341869
rect 207013 341866 207079 341869
rect 154481 341864 207079 341866
rect 154481 341808 154486 341864
rect 154542 341808 207018 341864
rect 207074 341808 207079 341864
rect 154481 341806 207079 341808
rect 154481 341803 154547 341806
rect 207013 341803 207079 341806
rect 240542 341804 240548 341868
rect 240612 341866 240618 341868
rect 291193 341866 291259 341869
rect 240612 341864 291259 341866
rect 240612 341808 291198 341864
rect 291254 341808 291259 341864
rect 240612 341806 291259 341808
rect 240612 341804 240618 341806
rect 291193 341803 291259 341806
rect 324630 341804 324636 341868
rect 324700 341866 324706 341868
rect 375373 341866 375439 341869
rect 324700 341864 375439 341866
rect 324700 341808 375378 341864
rect 375434 341808 375439 341864
rect 324700 341806 375439 341808
rect 324700 341804 324706 341806
rect 375373 341803 375439 341806
rect 378041 341866 378107 341869
rect 430573 341866 430639 341869
rect 378041 341864 430639 341866
rect 378041 341808 378046 341864
rect 378102 341808 430578 341864
rect 430634 341808 430639 341864
rect 378041 341806 430639 341808
rect 378041 341803 378107 341806
rect 430573 341803 430639 341806
rect 436502 341804 436508 341868
rect 436572 341866 436578 341868
rect 487153 341866 487219 341869
rect 436572 341864 487219 341866
rect 436572 341808 487158 341864
rect 487214 341808 487219 341864
rect 436572 341806 487219 341808
rect 436572 341804 436578 341806
rect 487153 341803 487219 341806
rect 492622 341804 492628 341868
rect 492692 341866 492698 341868
rect 542353 341866 542419 341869
rect 492692 341864 542419 341866
rect 492692 341808 542358 341864
rect 542414 341808 542419 341864
rect 492692 341806 542419 341808
rect 492692 341804 492698 341806
rect 542353 341803 542419 341806
rect 44582 341668 44588 341732
rect 44652 341730 44658 341732
rect 95233 341730 95299 341733
rect 44652 341728 95299 341730
rect 44652 341672 95238 341728
rect 95294 341672 95299 341728
rect 44652 341670 95299 341672
rect 44652 341668 44658 341670
rect 95233 341667 95299 341670
rect 128486 341668 128492 341732
rect 128556 341730 128562 341732
rect 178033 341730 178099 341733
rect 128556 341728 178099 341730
rect 128556 341672 178038 341728
rect 178094 341672 178099 341728
rect 128556 341670 178099 341672
rect 128556 341668 128562 341670
rect 178033 341667 178099 341670
rect 212574 341668 212580 341732
rect 212644 341730 212650 341732
rect 262213 341730 262279 341733
rect 212644 341728 262279 341730
rect 212644 341672 262218 341728
rect 262274 341672 262279 341728
rect 212644 341670 262279 341672
rect 212644 341668 212650 341670
rect 262213 341667 262279 341670
rect 296846 341668 296852 341732
rect 296916 341730 296922 341732
rect 346393 341730 346459 341733
rect 296916 341728 346459 341730
rect 296916 341672 346398 341728
rect 346454 341672 346459 341728
rect 296916 341670 346459 341672
rect 296916 341668 296922 341670
rect 346393 341667 346459 341670
rect 583520 338452 584960 338692
rect 148593 338058 148659 338061
rect 165654 338058 165660 338060
rect 148593 338056 165660 338058
rect 148593 338000 148598 338056
rect 148654 338000 165660 338056
rect 148593 337998 165660 338000
rect 148593 337995 148659 337998
rect 165654 337996 165660 337998
rect 165724 337996 165730 338060
rect 222653 338058 222719 338061
rect 259494 338058 259500 338060
rect 222653 338056 259500 338058
rect 222653 338000 222658 338056
rect 222714 338000 259500 338056
rect 222653 337998 259500 338000
rect 222653 337995 222719 337998
rect 259494 337996 259500 337998
rect 259564 337996 259570 338060
rect 344645 338058 344711 338061
rect 361614 338058 361620 338060
rect 344645 338056 361620 338058
rect 344645 338000 344650 338056
rect 344706 338000 361620 338056
rect 344645 337998 361620 338000
rect 344645 337995 344711 337998
rect 361614 337996 361620 337998
rect 361684 337996 361690 338060
rect 428641 338058 428707 338061
rect 445702 338058 445708 338060
rect 428641 338056 445708 338058
rect 428641 338000 428646 338056
rect 428702 338000 445708 338056
rect 428641 337998 445708 338000
rect 428641 337995 428707 337998
rect 445702 337996 445708 337998
rect 445772 337996 445778 338060
rect 540605 338058 540671 338061
rect 557574 338058 557580 338060
rect 540605 338056 557580 338058
rect 540605 338000 540610 338056
rect 540666 338000 557580 338056
rect 540605 337998 557580 338000
rect 540605 337995 540671 337998
rect 557574 337996 557580 337998
rect 557644 337996 557650 338060
rect 128302 333236 128308 333300
rect 128372 333298 128378 333300
rect 128445 333298 128511 333301
rect 194777 333300 194843 333301
rect 194726 333298 194732 333300
rect 128372 333296 128511 333298
rect 128372 333240 128450 333296
rect 128506 333240 128511 333296
rect 128372 333238 128511 333240
rect 194686 333238 194732 333298
rect 194796 333296 194843 333300
rect 194838 333240 194843 333296
rect 128372 333236 128378 333238
rect 128445 333235 128511 333238
rect 194726 333236 194732 333238
rect 194796 333236 194843 333240
rect 194777 333235 194843 333236
rect 390829 333300 390895 333301
rect 390829 333296 390876 333300
rect 390940 333298 390946 333300
rect 390829 333240 390834 333296
rect 390829 333236 390876 333240
rect 390940 333238 390986 333298
rect 390940 333236 390946 333238
rect 390829 333235 390895 333236
rect -960 332196 480 332436
rect 580073 325274 580139 325277
rect 583520 325274 584960 325364
rect 580073 325272 584960 325274
rect 580073 325216 580078 325272
rect 580134 325216 584960 325272
rect 580073 325214 584960 325216
rect 580073 325211 580139 325214
rect 583520 325124 584960 325214
rect 13537 323778 13603 323781
rect 38653 323778 38719 323781
rect 13537 323776 16100 323778
rect 13537 323720 13542 323776
rect 13598 323720 16100 323776
rect 13537 323718 16100 323720
rect 36892 323776 38719 323778
rect 36892 323720 38658 323776
rect 38714 323720 38719 323776
rect 36892 323718 38719 323720
rect 13537 323715 13603 323718
rect 38653 323715 38719 323718
rect 42701 323778 42767 323781
rect 66253 323778 66319 323781
rect 42701 323776 44068 323778
rect 42701 323720 42706 323776
rect 42762 323720 44068 323776
rect 42701 323718 44068 323720
rect 64860 323776 66319 323778
rect 64860 323720 66258 323776
rect 66314 323720 66319 323776
rect 64860 323718 66319 323720
rect 42701 323715 42767 323718
rect 66253 323715 66319 323718
rect 70301 323778 70367 323781
rect 95233 323778 95299 323781
rect 70301 323776 72036 323778
rect 70301 323720 70306 323776
rect 70362 323720 72036 323776
rect 70301 323718 72036 323720
rect 92828 323776 95299 323778
rect 92828 323720 95238 323776
rect 95294 323720 95299 323776
rect 92828 323718 95299 323720
rect 70301 323715 70367 323718
rect 95233 323715 95299 323718
rect 97901 323778 97967 323781
rect 122833 323778 122899 323781
rect 97901 323776 100188 323778
rect 97901 323720 97906 323776
rect 97962 323720 100188 323776
rect 97901 323718 100188 323720
rect 120796 323776 122899 323778
rect 120796 323720 122838 323776
rect 122894 323720 122899 323776
rect 120796 323718 122899 323720
rect 97901 323715 97967 323718
rect 122833 323715 122899 323718
rect 126881 323778 126947 323781
rect 150433 323778 150499 323781
rect 126881 323776 128156 323778
rect 126881 323720 126886 323776
rect 126942 323720 128156 323776
rect 126881 323718 128156 323720
rect 148948 323776 150499 323778
rect 148948 323720 150438 323776
rect 150494 323720 150499 323776
rect 148948 323718 150499 323720
rect 126881 323715 126947 323718
rect 150433 323715 150499 323718
rect 154481 323778 154547 323781
rect 182081 323778 182147 323781
rect 207013 323778 207079 323781
rect 154481 323776 156124 323778
rect 154481 323720 154486 323776
rect 154542 323720 156124 323776
rect 182081 323776 184092 323778
rect 154481 323718 156124 323720
rect 154481 323715 154547 323718
rect 176334 323236 176394 323748
rect 182081 323720 182086 323776
rect 182142 323720 184092 323776
rect 182081 323718 184092 323720
rect 204884 323776 207079 323778
rect 204884 323720 207018 323776
rect 207074 323720 207079 323776
rect 204884 323718 207079 323720
rect 182081 323715 182147 323718
rect 207013 323715 207079 323718
rect 209681 323778 209747 323781
rect 234705 323778 234771 323781
rect 209681 323776 212060 323778
rect 209681 323720 209686 323776
rect 209742 323720 212060 323776
rect 209681 323718 212060 323720
rect 232852 323776 234771 323778
rect 232852 323720 234710 323776
rect 234766 323720 234771 323776
rect 232852 323718 234771 323720
rect 209681 323715 209747 323718
rect 234705 323715 234771 323718
rect 238661 323778 238727 323781
rect 262213 323778 262279 323781
rect 238661 323776 240212 323778
rect 238661 323720 238666 323776
rect 238722 323720 240212 323776
rect 238661 323718 240212 323720
rect 260820 323776 262279 323778
rect 260820 323720 262218 323776
rect 262274 323720 262279 323776
rect 260820 323718 262279 323720
rect 238661 323715 238727 323718
rect 262213 323715 262279 323718
rect 266261 323778 266327 323781
rect 291193 323778 291259 323781
rect 266261 323776 268180 323778
rect 266261 323720 266266 323776
rect 266322 323720 268180 323776
rect 266261 323718 268180 323720
rect 288788 323776 291259 323778
rect 288788 323720 291198 323776
rect 291254 323720 291259 323776
rect 288788 323718 291259 323720
rect 266261 323715 266327 323718
rect 291193 323715 291259 323718
rect 293861 323778 293927 323781
rect 318793 323778 318859 323781
rect 293861 323776 296148 323778
rect 293861 323720 293866 323776
rect 293922 323720 296148 323776
rect 293861 323718 296148 323720
rect 316940 323776 318859 323778
rect 316940 323720 318798 323776
rect 318854 323720 318859 323776
rect 316940 323718 318859 323720
rect 293861 323715 293927 323718
rect 318793 323715 318859 323718
rect 322841 323778 322907 323781
rect 346393 323778 346459 323781
rect 322841 323776 324116 323778
rect 322841 323720 322846 323776
rect 322902 323720 324116 323776
rect 322841 323718 324116 323720
rect 344908 323776 346459 323778
rect 344908 323720 346398 323776
rect 346454 323720 346459 323776
rect 344908 323718 346459 323720
rect 322841 323715 322907 323718
rect 346393 323715 346459 323718
rect 350441 323778 350507 323781
rect 375373 323778 375439 323781
rect 350441 323776 352084 323778
rect 350441 323720 350446 323776
rect 350502 323720 352084 323776
rect 350441 323718 352084 323720
rect 372876 323776 375439 323778
rect 372876 323720 375378 323776
rect 375434 323720 375439 323776
rect 372876 323718 375439 323720
rect 350441 323715 350507 323718
rect 375373 323715 375439 323718
rect 378041 323778 378107 323781
rect 402973 323778 403039 323781
rect 378041 323776 380052 323778
rect 378041 323720 378046 323776
rect 378102 323720 380052 323776
rect 378041 323718 380052 323720
rect 400844 323776 403039 323778
rect 400844 323720 402978 323776
rect 403034 323720 403039 323776
rect 400844 323718 403039 323720
rect 378041 323715 378107 323718
rect 402973 323715 403039 323718
rect 405641 323778 405707 323781
rect 430573 323778 430639 323781
rect 405641 323776 408204 323778
rect 405641 323720 405646 323776
rect 405702 323720 408204 323776
rect 405641 323718 408204 323720
rect 428812 323776 430639 323778
rect 428812 323720 430578 323776
rect 430634 323720 430639 323776
rect 428812 323718 430639 323720
rect 405641 323715 405707 323718
rect 430573 323715 430639 323718
rect 434621 323778 434687 323781
rect 462221 323778 462287 323781
rect 487153 323778 487219 323781
rect 434621 323776 436172 323778
rect 434621 323720 434626 323776
rect 434682 323720 436172 323776
rect 462221 323776 464140 323778
rect 434621 323718 436172 323720
rect 434621 323715 434687 323718
rect 456382 323236 456442 323748
rect 462221 323720 462226 323776
rect 462282 323720 464140 323776
rect 462221 323718 464140 323720
rect 484932 323776 487219 323778
rect 484932 323720 487158 323776
rect 487214 323720 487219 323776
rect 484932 323718 487219 323720
rect 462221 323715 462287 323718
rect 487153 323715 487219 323718
rect 489821 323778 489887 323781
rect 514753 323778 514819 323781
rect 489821 323776 492108 323778
rect 489821 323720 489826 323776
rect 489882 323720 492108 323776
rect 489821 323718 492108 323720
rect 512900 323776 514819 323778
rect 512900 323720 514758 323776
rect 514814 323720 514819 323776
rect 512900 323718 514819 323720
rect 489821 323715 489887 323718
rect 514753 323715 514819 323718
rect 518801 323778 518867 323781
rect 542353 323778 542419 323781
rect 518801 323776 520076 323778
rect 518801 323720 518806 323776
rect 518862 323720 520076 323776
rect 518801 323718 520076 323720
rect 540868 323776 542419 323778
rect 540868 323720 542358 323776
rect 542414 323720 542419 323776
rect 540868 323718 542419 323720
rect 518801 323715 518867 323718
rect 542353 323715 542419 323718
rect 546401 323778 546467 323781
rect 546401 323776 548044 323778
rect 546401 323720 546406 323776
rect 546462 323720 548044 323776
rect 546401 323718 548044 323720
rect 546401 323715 546467 323718
rect 568438 323372 568498 323748
rect 568430 323308 568436 323372
rect 568500 323308 568506 323372
rect 176326 323172 176332 323236
rect 176396 323172 176402 323236
rect 456374 323172 456380 323236
rect 456444 323172 456450 323236
rect -960 319140 480 319380
rect 13537 315346 13603 315349
rect 66253 315346 66319 315349
rect 13537 315344 66319 315346
rect 13537 315288 13542 315344
rect 13598 315288 66258 315344
rect 66314 315288 66319 315344
rect 13537 315286 66319 315288
rect 13537 315283 13603 315286
rect 66253 315283 66319 315286
rect 70301 315346 70367 315349
rect 122833 315346 122899 315349
rect 70301 315344 122899 315346
rect 70301 315288 70306 315344
rect 70362 315288 122838 315344
rect 122894 315288 122899 315344
rect 70301 315286 122899 315288
rect 70301 315283 70367 315286
rect 122833 315283 122899 315286
rect 126881 315346 126947 315349
rect 175222 315346 175228 315348
rect 126881 315344 175228 315346
rect 126881 315288 126886 315344
rect 126942 315288 175228 315344
rect 126881 315286 175228 315288
rect 126881 315283 126947 315286
rect 175222 315284 175228 315286
rect 175292 315284 175298 315348
rect 182081 315346 182147 315349
rect 234705 315346 234771 315349
rect 182081 315344 234771 315346
rect 182081 315288 182086 315344
rect 182142 315288 234710 315344
rect 234766 315288 234771 315344
rect 182081 315286 234771 315288
rect 182081 315283 182147 315286
rect 234705 315283 234771 315286
rect 238661 315346 238727 315349
rect 291193 315346 291259 315349
rect 238661 315344 291259 315346
rect 238661 315288 238666 315344
rect 238722 315288 291198 315344
rect 291254 315288 291259 315344
rect 238661 315286 291259 315288
rect 238661 315283 238727 315286
rect 291193 315283 291259 315286
rect 293861 315346 293927 315349
rect 346393 315346 346459 315349
rect 293861 315344 346459 315346
rect 293861 315288 293866 315344
rect 293922 315288 346398 315344
rect 346454 315288 346459 315344
rect 293861 315286 346459 315288
rect 293861 315283 293927 315286
rect 346393 315283 346459 315286
rect 350441 315346 350507 315349
rect 402973 315346 403039 315349
rect 350441 315344 403039 315346
rect 350441 315288 350446 315344
rect 350502 315288 402978 315344
rect 403034 315288 403039 315344
rect 350441 315286 403039 315288
rect 350441 315283 350507 315286
rect 402973 315283 403039 315286
rect 405641 315346 405707 315349
rect 455454 315346 455460 315348
rect 405641 315344 455460 315346
rect 405641 315288 405646 315344
rect 405702 315288 455460 315344
rect 405641 315286 455460 315288
rect 405641 315283 405707 315286
rect 455454 315284 455460 315286
rect 455524 315284 455530 315348
rect 462221 315346 462287 315349
rect 514753 315346 514819 315349
rect 462221 315344 514819 315346
rect 462221 315288 462226 315344
rect 462282 315288 514758 315344
rect 514814 315288 514819 315344
rect 462221 315286 514819 315288
rect 462221 315283 462287 315286
rect 514753 315283 514819 315286
rect 518801 315346 518867 315349
rect 566958 315346 566964 315348
rect 518801 315344 566964 315346
rect 518801 315288 518806 315344
rect 518862 315288 566964 315344
rect 518801 315286 566964 315288
rect 518801 315283 518867 315286
rect 566958 315284 566964 315286
rect 567028 315284 567034 315348
rect 583520 311932 584960 312172
rect 110597 311810 110663 311813
rect 128302 311810 128308 311812
rect 110597 311808 128308 311810
rect 110597 311752 110602 311808
rect 110658 311752 128308 311808
rect 110597 311750 128308 311752
rect 110597 311747 110663 311750
rect 128302 311748 128308 311750
rect 128372 311748 128378 311812
rect 156321 311810 156387 311813
rect 194726 311810 194732 311812
rect 156321 311808 194732 311810
rect 156321 311752 156326 311808
rect 156382 311752 194732 311808
rect 156321 311750 194732 311752
rect 156321 311747 156387 311750
rect 194726 311748 194732 311750
rect 194796 311748 194802 311812
rect 352649 311810 352715 311813
rect 390870 311810 390876 311812
rect 352649 311808 390876 311810
rect 352649 311752 352654 311808
rect 352710 311752 390876 311808
rect 352649 311750 390876 311752
rect 352649 311747 352715 311750
rect 390870 311748 390876 311750
rect 390940 311748 390946 311812
rect 165654 306444 165660 306508
rect 165724 306506 165730 306508
rect 165981 306506 166047 306509
rect 165724 306504 166047 306506
rect 165724 306448 165986 306504
rect 166042 306448 166047 306504
rect 165724 306446 166047 306448
rect 165724 306444 165730 306446
rect 165981 306443 166047 306446
rect 259494 306444 259500 306508
rect 259564 306506 259570 306508
rect 260373 306506 260439 306509
rect 259564 306504 260439 306506
rect 259564 306448 260378 306504
rect 260434 306448 260439 306504
rect 259564 306446 260439 306448
rect 259564 306444 259570 306446
rect 260373 306443 260439 306446
rect 361614 306444 361620 306508
rect 361684 306506 361690 306508
rect 361941 306506 362007 306509
rect 361684 306504 362007 306506
rect 361684 306448 361946 306504
rect 362002 306448 362007 306504
rect 361684 306446 362007 306448
rect 361684 306444 361690 306446
rect 361941 306443 362007 306446
rect 445702 306444 445708 306508
rect 445772 306506 445778 306508
rect 446029 306506 446095 306509
rect 445772 306504 446095 306506
rect 445772 306448 446034 306504
rect 446090 306448 446095 306504
rect 445772 306446 446095 306448
rect 445772 306444 445778 306446
rect 446029 306443 446095 306446
rect 557574 306444 557580 306508
rect 557644 306506 557650 306508
rect 557993 306506 558059 306509
rect 557644 306504 558059 306506
rect 557644 306448 557998 306504
rect 558054 306448 558059 306504
rect 557644 306446 558059 306448
rect 557644 306444 557650 306446
rect 557993 306443 558059 306446
rect -960 306234 480 306324
rect 3877 306234 3943 306237
rect -960 306232 3943 306234
rect -960 306176 3882 306232
rect 3938 306176 3943 306232
rect -960 306174 3943 306176
rect -960 306084 480 306174
rect 3877 306171 3943 306174
rect 583520 298604 584960 298844
rect 13721 296306 13787 296309
rect 38653 296306 38719 296309
rect 66253 296306 66319 296309
rect 13721 296304 16100 296306
rect 13721 296248 13726 296304
rect 13782 296248 16100 296304
rect 13721 296246 16100 296248
rect 36892 296304 38719 296306
rect 36892 296248 38658 296304
rect 38714 296248 38719 296304
rect 64860 296304 66319 296306
rect 36892 296246 38719 296248
rect 13721 296243 13787 296246
rect 38653 296243 38719 296246
rect 44590 295764 44650 296276
rect 64860 296248 66258 296304
rect 66314 296248 66319 296304
rect 64860 296246 66319 296248
rect 66253 296243 66319 296246
rect 70301 296306 70367 296309
rect 95233 296306 95299 296309
rect 70301 296304 72036 296306
rect 70301 296248 70306 296304
rect 70362 296248 72036 296304
rect 70301 296246 72036 296248
rect 92828 296304 95299 296306
rect 92828 296248 95238 296304
rect 95294 296248 95299 296304
rect 92828 296246 95299 296248
rect 70301 296243 70367 296246
rect 95233 296243 95299 296246
rect 97901 296306 97967 296309
rect 122833 296306 122899 296309
rect 97901 296304 100188 296306
rect 97901 296248 97906 296304
rect 97962 296248 100188 296304
rect 97901 296246 100188 296248
rect 120796 296304 122899 296306
rect 120796 296248 122838 296304
rect 122894 296248 122899 296304
rect 120796 296246 122899 296248
rect 97901 296243 97967 296246
rect 122833 296243 122899 296246
rect 126881 296306 126947 296309
rect 150433 296306 150499 296309
rect 126881 296304 128156 296306
rect 126881 296248 126886 296304
rect 126942 296248 128156 296304
rect 126881 296246 128156 296248
rect 148948 296304 150499 296306
rect 148948 296248 150438 296304
rect 150494 296248 150499 296304
rect 148948 296246 150499 296248
rect 126881 296243 126947 296246
rect 150433 296243 150499 296246
rect 154481 296306 154547 296309
rect 182081 296306 182147 296309
rect 207013 296306 207079 296309
rect 234705 296306 234771 296309
rect 154481 296304 156124 296306
rect 154481 296248 154486 296304
rect 154542 296248 156124 296304
rect 182081 296304 184092 296306
rect 154481 296246 156124 296248
rect 154481 296243 154547 296246
rect 176334 295764 176394 296276
rect 182081 296248 182086 296304
rect 182142 296248 184092 296304
rect 182081 296246 184092 296248
rect 204884 296304 207079 296306
rect 204884 296248 207018 296304
rect 207074 296248 207079 296304
rect 232852 296304 234771 296306
rect 204884 296246 207079 296248
rect 182081 296243 182147 296246
rect 207013 296243 207079 296246
rect 212582 295764 212642 296276
rect 232852 296248 234710 296304
rect 234766 296248 234771 296304
rect 232852 296246 234771 296248
rect 234705 296243 234771 296246
rect 238661 296306 238727 296309
rect 262213 296306 262279 296309
rect 238661 296304 240212 296306
rect 238661 296248 238666 296304
rect 238722 296248 240212 296304
rect 238661 296246 240212 296248
rect 260820 296304 262279 296306
rect 260820 296248 262218 296304
rect 262274 296248 262279 296304
rect 260820 296246 262279 296248
rect 238661 296243 238727 296246
rect 262213 296243 262279 296246
rect 266261 296306 266327 296309
rect 318793 296306 318859 296309
rect 266261 296304 268180 296306
rect 266261 296248 266266 296304
rect 266322 296248 268180 296304
rect 316940 296304 318859 296306
rect 266261 296246 268180 296248
rect 266261 296243 266327 296246
rect 288390 295764 288450 296276
rect 296486 295764 296546 296276
rect 316940 296248 318798 296304
rect 318854 296248 318859 296304
rect 316940 296246 318859 296248
rect 318793 296243 318859 296246
rect 322841 296306 322907 296309
rect 346393 296306 346459 296309
rect 322841 296304 324116 296306
rect 322841 296248 322846 296304
rect 322902 296248 324116 296304
rect 322841 296246 324116 296248
rect 344908 296304 346459 296306
rect 344908 296248 346398 296304
rect 346454 296248 346459 296304
rect 344908 296246 346459 296248
rect 322841 296243 322907 296246
rect 346393 296243 346459 296246
rect 350441 296306 350507 296309
rect 378041 296306 378107 296309
rect 402973 296306 403039 296309
rect 430573 296306 430639 296309
rect 350441 296304 352084 296306
rect 350441 296248 350446 296304
rect 350502 296248 352084 296304
rect 378041 296304 380052 296306
rect 350441 296246 352084 296248
rect 350441 296243 350507 296246
rect 372294 295764 372354 296276
rect 378041 296248 378046 296304
rect 378102 296248 380052 296304
rect 378041 296246 380052 296248
rect 400844 296304 403039 296306
rect 400844 296248 402978 296304
rect 403034 296248 403039 296304
rect 428812 296304 430639 296306
rect 400844 296246 403039 296248
rect 378041 296243 378107 296246
rect 402973 296243 403039 296246
rect 408542 295764 408602 296276
rect 428812 296248 430578 296304
rect 430634 296248 430639 296304
rect 428812 296246 430639 296248
rect 430573 296243 430639 296246
rect 434621 296306 434687 296309
rect 458173 296306 458239 296309
rect 434621 296304 436172 296306
rect 434621 296248 434626 296304
rect 434682 296248 436172 296304
rect 434621 296246 436172 296248
rect 456964 296304 458239 296306
rect 456964 296248 458178 296304
rect 458234 296248 458239 296304
rect 456964 296246 458239 296248
rect 434621 296243 434687 296246
rect 458173 296243 458239 296246
rect 462221 296306 462287 296309
rect 514753 296306 514819 296309
rect 542353 296306 542419 296309
rect 462221 296304 464140 296306
rect 462221 296248 462226 296304
rect 462282 296248 464140 296304
rect 512900 296304 514819 296306
rect 462221 296246 464140 296248
rect 462221 296243 462287 296246
rect 484350 295764 484410 296276
rect 492630 295764 492690 296276
rect 512900 296248 514758 296304
rect 514814 296248 514819 296304
rect 540868 296304 542419 296306
rect 512900 296246 514819 296248
rect 514753 296243 514819 296246
rect 520598 295764 520658 296276
rect 540868 296248 542358 296304
rect 542414 296248 542419 296304
rect 540868 296246 542419 296248
rect 542353 296243 542419 296246
rect 546401 296306 546467 296309
rect 571333 296306 571399 296309
rect 546401 296304 548044 296306
rect 546401 296248 546406 296304
rect 546462 296248 548044 296304
rect 546401 296246 548044 296248
rect 568836 296304 571399 296306
rect 568836 296248 571338 296304
rect 571394 296248 571399 296304
rect 568836 296246 571399 296248
rect 546401 296243 546467 296246
rect 571333 296243 571399 296246
rect 44582 295700 44588 295764
rect 44652 295700 44658 295764
rect 176326 295700 176332 295764
rect 176396 295700 176402 295764
rect 212574 295700 212580 295764
rect 212644 295700 212650 295764
rect 288382 295700 288388 295764
rect 288452 295700 288458 295764
rect 296478 295700 296484 295764
rect 296548 295700 296554 295764
rect 372286 295700 372292 295764
rect 372356 295700 372362 295764
rect 408534 295700 408540 295764
rect 408604 295700 408610 295764
rect 484342 295700 484348 295764
rect 484412 295700 484418 295764
rect 492622 295700 492628 295764
rect 492692 295700 492698 295764
rect 520590 295700 520596 295764
rect 520660 295700 520666 295764
rect -960 293178 480 293268
rect 3141 293178 3207 293181
rect -960 293176 3207 293178
rect -960 293120 3146 293176
rect 3202 293120 3207 293176
rect -960 293118 3207 293120
rect -960 293028 480 293118
rect 3141 293115 3207 293118
rect 13721 288010 13787 288013
rect 66253 288010 66319 288013
rect 13721 288008 66319 288010
rect 13721 287952 13726 288008
rect 13782 287952 66258 288008
rect 66314 287952 66319 288008
rect 13721 287950 66319 287952
rect 13721 287947 13787 287950
rect 66253 287947 66319 287950
rect 70301 288010 70367 288013
rect 122833 288010 122899 288013
rect 70301 288008 122899 288010
rect 70301 287952 70306 288008
rect 70362 287952 122838 288008
rect 122894 287952 122899 288008
rect 70301 287950 122899 287952
rect 70301 287947 70367 287950
rect 122833 287947 122899 287950
rect 126881 288010 126947 288013
rect 176326 288010 176332 288012
rect 126881 288008 176332 288010
rect 126881 287952 126886 288008
rect 126942 287952 176332 288008
rect 126881 287950 176332 287952
rect 126881 287947 126947 287950
rect 176326 287948 176332 287950
rect 176396 287948 176402 288012
rect 182081 288010 182147 288013
rect 234705 288010 234771 288013
rect 182081 288008 234771 288010
rect 182081 287952 182086 288008
rect 182142 287952 234710 288008
rect 234766 287952 234771 288008
rect 182081 287950 234771 287952
rect 182081 287947 182147 287950
rect 234705 287947 234771 287950
rect 266261 288010 266327 288013
rect 318793 288010 318859 288013
rect 266261 288008 318859 288010
rect 266261 287952 266266 288008
rect 266322 287952 318798 288008
rect 318854 287952 318859 288008
rect 266261 287950 318859 287952
rect 266261 287947 266327 287950
rect 318793 287947 318859 287950
rect 322841 288010 322907 288013
rect 372286 288010 372292 288012
rect 322841 288008 372292 288010
rect 322841 287952 322846 288008
rect 322902 287952 372292 288008
rect 322841 287950 372292 287952
rect 322841 287947 322907 287950
rect 372286 287948 372292 287950
rect 372356 287948 372362 288012
rect 378041 288010 378107 288013
rect 430573 288010 430639 288013
rect 378041 288008 430639 288010
rect 378041 287952 378046 288008
rect 378102 287952 430578 288008
rect 430634 287952 430639 288008
rect 378041 287950 430639 287952
rect 378041 287947 378107 287950
rect 430573 287947 430639 287950
rect 462221 288010 462287 288013
rect 514753 288010 514819 288013
rect 462221 288008 514819 288010
rect 462221 287952 462226 288008
rect 462282 287952 514758 288008
rect 514814 287952 514819 288008
rect 462221 287950 514819 287952
rect 462221 287947 462287 287950
rect 514753 287947 514819 287950
rect 520590 287948 520596 288012
rect 520660 288010 520666 288012
rect 571333 288010 571399 288013
rect 520660 288008 571399 288010
rect 520660 287952 571338 288008
rect 571394 287952 571399 288008
rect 520660 287950 571399 287952
rect 520660 287948 520666 287950
rect 571333 287947 571399 287950
rect 44582 287812 44588 287876
rect 44652 287874 44658 287876
rect 95233 287874 95299 287877
rect 44652 287872 95299 287874
rect 44652 287816 95238 287872
rect 95294 287816 95299 287872
rect 44652 287814 95299 287816
rect 44652 287812 44658 287814
rect 95233 287811 95299 287814
rect 97901 287874 97967 287877
rect 150433 287874 150499 287877
rect 97901 287872 150499 287874
rect 97901 287816 97906 287872
rect 97962 287816 150438 287872
rect 150494 287816 150499 287872
rect 97901 287814 150499 287816
rect 97901 287811 97967 287814
rect 150433 287811 150499 287814
rect 154481 287874 154547 287877
rect 207013 287874 207079 287877
rect 154481 287872 207079 287874
rect 154481 287816 154486 287872
rect 154542 287816 207018 287872
rect 207074 287816 207079 287872
rect 154481 287814 207079 287816
rect 154481 287811 154547 287814
rect 207013 287811 207079 287814
rect 212574 287812 212580 287876
rect 212644 287874 212650 287876
rect 262213 287874 262279 287877
rect 212644 287872 262279 287874
rect 212644 287816 262218 287872
rect 262274 287816 262279 287872
rect 212644 287814 262279 287816
rect 212644 287812 212650 287814
rect 262213 287811 262279 287814
rect 296846 287812 296852 287876
rect 296916 287874 296922 287876
rect 346393 287874 346459 287877
rect 296916 287872 346459 287874
rect 296916 287816 346398 287872
rect 346454 287816 346459 287872
rect 296916 287814 346459 287816
rect 296916 287812 296922 287814
rect 346393 287811 346459 287814
rect 350441 287874 350507 287877
rect 402973 287874 403039 287877
rect 350441 287872 403039 287874
rect 350441 287816 350446 287872
rect 350502 287816 402978 287872
rect 403034 287816 403039 287872
rect 350441 287814 403039 287816
rect 350441 287811 350507 287814
rect 402973 287811 403039 287814
rect 408534 287812 408540 287876
rect 408604 287874 408610 287876
rect 458173 287874 458239 287877
rect 408604 287872 458239 287874
rect 408604 287816 458178 287872
rect 458234 287816 458239 287872
rect 408604 287814 458239 287816
rect 408604 287812 408610 287814
rect 458173 287811 458239 287814
rect 492622 287812 492628 287876
rect 492692 287874 492698 287876
rect 542353 287874 542419 287877
rect 492692 287872 542419 287874
rect 492692 287816 542358 287872
rect 542414 287816 542419 287872
rect 492692 287814 542419 287816
rect 492692 287812 492698 287814
rect 542353 287811 542419 287814
rect 238661 287738 238727 287741
rect 288382 287738 288388 287740
rect 238661 287736 288388 287738
rect 238661 287680 238666 287736
rect 238722 287680 288388 287736
rect 238661 287678 288388 287680
rect 238661 287675 238727 287678
rect 288382 287676 288388 287678
rect 288452 287676 288458 287740
rect 434621 287738 434687 287741
rect 484342 287738 484348 287740
rect 434621 287736 484348 287738
rect 434621 287680 434626 287736
rect 434682 287680 484348 287736
rect 434621 287678 484348 287680
rect 434621 287675 434687 287678
rect 484342 287676 484348 287678
rect 484412 287676 484418 287740
rect 583520 285276 584960 285516
rect 148593 284202 148659 284205
rect 165654 284202 165660 284204
rect 148593 284200 165660 284202
rect 148593 284144 148598 284200
rect 148654 284144 165660 284200
rect 148593 284142 165660 284144
rect 148593 284139 148659 284142
rect 165654 284140 165660 284142
rect 165724 284140 165730 284204
rect 222653 284202 222719 284205
rect 259494 284202 259500 284204
rect 222653 284200 259500 284202
rect 222653 284144 222658 284200
rect 222714 284144 259500 284200
rect 222653 284142 259500 284144
rect 222653 284139 222719 284142
rect 259494 284140 259500 284142
rect 259564 284140 259570 284204
rect 344645 284202 344711 284205
rect 361614 284202 361620 284204
rect 344645 284200 361620 284202
rect 344645 284144 344650 284200
rect 344706 284144 361620 284200
rect 344645 284142 361620 284144
rect 344645 284139 344711 284142
rect 361614 284140 361620 284142
rect 361684 284140 361690 284204
rect 428641 284202 428707 284205
rect 445702 284202 445708 284204
rect 428641 284200 445708 284202
rect 428641 284144 428646 284200
rect 428702 284144 445708 284200
rect 428641 284142 445708 284144
rect 428641 284139 428707 284142
rect 445702 284140 445708 284142
rect 445772 284140 445778 284204
rect 540605 284202 540671 284205
rect 557574 284202 557580 284204
rect 540605 284200 557580 284202
rect 540605 284144 540610 284200
rect 540666 284144 557580 284200
rect 540605 284142 557580 284144
rect 540605 284139 540671 284142
rect 557574 284140 557580 284142
rect 557644 284140 557650 284204
rect -960 279972 480 280212
rect 277342 279788 277348 279852
rect 277412 279850 277418 279852
rect 278221 279850 278287 279853
rect 277412 279848 278287 279850
rect 277412 279792 278226 279848
rect 278282 279792 278287 279848
rect 277412 279790 278287 279792
rect 277412 279788 277418 279790
rect 278221 279787 278287 279790
rect 81382 279244 81388 279308
rect 81452 279306 81458 279308
rect 82261 279306 82327 279309
rect 81452 279304 82327 279306
rect 81452 279248 82266 279304
rect 82322 279248 82327 279304
rect 81452 279246 82327 279248
rect 81452 279244 81458 279246
rect 82261 279243 82327 279246
rect 128302 279244 128308 279308
rect 128372 279306 128378 279308
rect 128445 279306 128511 279309
rect 194777 279308 194843 279309
rect 194726 279306 194732 279308
rect 128372 279304 128511 279306
rect 128372 279248 128450 279304
rect 128506 279248 128511 279304
rect 128372 279246 128511 279248
rect 194686 279246 194732 279306
rect 194796 279304 194843 279308
rect 194838 279248 194843 279304
rect 128372 279244 128378 279246
rect 128445 279243 128511 279246
rect 194726 279244 194732 279246
rect 194796 279244 194843 279248
rect 194777 279243 194843 279244
rect 390829 279308 390895 279309
rect 390829 279304 390876 279308
rect 390940 279306 390946 279308
rect 390829 279248 390834 279304
rect 390829 279244 390876 279248
rect 390940 279246 390986 279306
rect 390940 279244 390946 279246
rect 473486 279244 473492 279308
rect 473556 279306 473562 279308
rect 474273 279306 474339 279309
rect 473556 279304 474339 279306
rect 473556 279248 474278 279304
rect 474334 279248 474339 279304
rect 473556 279246 474339 279248
rect 473556 279244 473562 279246
rect 390829 279243 390895 279244
rect 474273 279243 474339 279246
rect 520181 279308 520247 279309
rect 520181 279304 520228 279308
rect 520292 279306 520298 279308
rect 520181 279248 520186 279304
rect 520181 279244 520228 279248
rect 520292 279246 520338 279306
rect 520292 279244 520298 279246
rect 520181 279243 520247 279244
rect 13537 278082 13603 278085
rect 66253 278082 66319 278085
rect 13537 278080 66319 278082
rect 13537 278024 13542 278080
rect 13598 278024 66258 278080
rect 66314 278024 66319 278080
rect 13537 278022 66319 278024
rect 13537 278019 13603 278022
rect 66253 278019 66319 278022
rect 70301 278082 70367 278085
rect 122833 278082 122899 278085
rect 70301 278080 122899 278082
rect 70301 278024 70306 278080
rect 70362 278024 122838 278080
rect 122894 278024 122899 278080
rect 70301 278022 122899 278024
rect 70301 278019 70367 278022
rect 122833 278019 122899 278022
rect 126881 278082 126947 278085
rect 176326 278082 176332 278084
rect 126881 278080 176332 278082
rect 126881 278024 126886 278080
rect 126942 278024 176332 278080
rect 126881 278022 176332 278024
rect 126881 278019 126947 278022
rect 176326 278020 176332 278022
rect 176396 278020 176402 278084
rect 182081 278082 182147 278085
rect 234705 278082 234771 278085
rect 182081 278080 234771 278082
rect 182081 278024 182086 278080
rect 182142 278024 234710 278080
rect 234766 278024 234771 278080
rect 182081 278022 234771 278024
rect 182081 278019 182147 278022
rect 234705 278019 234771 278022
rect 238661 278082 238727 278085
rect 291193 278082 291259 278085
rect 238661 278080 291259 278082
rect 238661 278024 238666 278080
rect 238722 278024 291198 278080
rect 291254 278024 291259 278080
rect 238661 278022 291259 278024
rect 238661 278019 238727 278022
rect 291193 278019 291259 278022
rect 293861 278082 293927 278085
rect 346393 278082 346459 278085
rect 293861 278080 346459 278082
rect 293861 278024 293866 278080
rect 293922 278024 346398 278080
rect 346454 278024 346459 278080
rect 293861 278022 346459 278024
rect 293861 278019 293927 278022
rect 346393 278019 346459 278022
rect 350441 278082 350507 278085
rect 402973 278082 403039 278085
rect 350441 278080 403039 278082
rect 350441 278024 350446 278080
rect 350502 278024 402978 278080
rect 403034 278024 403039 278080
rect 350441 278022 403039 278024
rect 350441 278019 350507 278022
rect 402973 278019 403039 278022
rect 405641 278082 405707 278085
rect 456374 278082 456380 278084
rect 405641 278080 456380 278082
rect 405641 278024 405646 278080
rect 405702 278024 456380 278080
rect 405641 278022 456380 278024
rect 405641 278019 405707 278022
rect 456374 278020 456380 278022
rect 456444 278020 456450 278084
rect 462221 278082 462287 278085
rect 514753 278082 514819 278085
rect 462221 278080 514819 278082
rect 462221 278024 462226 278080
rect 462282 278024 514758 278080
rect 514814 278024 514819 278080
rect 462221 278022 514819 278024
rect 462221 278019 462287 278022
rect 514753 278019 514819 278022
rect 518801 278082 518867 278085
rect 566958 278082 566964 278084
rect 518801 278080 566964 278082
rect 518801 278024 518806 278080
rect 518862 278024 566964 278080
rect 518801 278022 566964 278024
rect 518801 278019 518867 278022
rect 566958 278020 566964 278022
rect 567028 278020 567034 278084
rect 578877 272234 578943 272237
rect 583520 272234 584960 272324
rect 578877 272232 584960 272234
rect 578877 272176 578882 272232
rect 578938 272176 584960 272232
rect 578877 272174 584960 272176
rect 578877 272171 578943 272174
rect 583520 272084 584960 272174
rect 176326 270268 176332 270332
rect 176396 270268 176402 270332
rect 456374 270268 456380 270332
rect 456444 270268 456450 270332
rect 13537 269786 13603 269789
rect 38653 269786 38719 269789
rect 13537 269784 16100 269786
rect 13537 269728 13542 269784
rect 13598 269728 16100 269784
rect 13537 269726 16100 269728
rect 36892 269784 38719 269786
rect 36892 269728 38658 269784
rect 38714 269728 38719 269784
rect 36892 269726 38719 269728
rect 13537 269723 13603 269726
rect 38653 269723 38719 269726
rect 42701 269786 42767 269789
rect 66253 269786 66319 269789
rect 42701 269784 44068 269786
rect 42701 269728 42706 269784
rect 42762 269728 44068 269784
rect 42701 269726 44068 269728
rect 64860 269784 66319 269786
rect 64860 269728 66258 269784
rect 66314 269728 66319 269784
rect 64860 269726 66319 269728
rect 42701 269723 42767 269726
rect 66253 269723 66319 269726
rect 70301 269786 70367 269789
rect 95233 269786 95299 269789
rect 70301 269784 72036 269786
rect 70301 269728 70306 269784
rect 70362 269728 72036 269784
rect 70301 269726 72036 269728
rect 92828 269784 95299 269786
rect 92828 269728 95238 269784
rect 95294 269728 95299 269784
rect 92828 269726 95299 269728
rect 70301 269723 70367 269726
rect 95233 269723 95299 269726
rect 97901 269786 97967 269789
rect 122833 269786 122899 269789
rect 97901 269784 100188 269786
rect 97901 269728 97906 269784
rect 97962 269728 100188 269784
rect 97901 269726 100188 269728
rect 120796 269784 122899 269786
rect 120796 269728 122838 269784
rect 122894 269728 122899 269784
rect 120796 269726 122899 269728
rect 97901 269723 97967 269726
rect 122833 269723 122899 269726
rect 126881 269786 126947 269789
rect 150433 269786 150499 269789
rect 126881 269784 128156 269786
rect 126881 269728 126886 269784
rect 126942 269728 128156 269784
rect 126881 269726 128156 269728
rect 148948 269784 150499 269786
rect 148948 269728 150438 269784
rect 150494 269728 150499 269784
rect 148948 269726 150499 269728
rect 126881 269723 126947 269726
rect 150433 269723 150499 269726
rect 154481 269786 154547 269789
rect 154481 269784 156124 269786
rect 154481 269728 154486 269784
rect 154542 269728 156124 269784
rect 176334 269756 176394 270268
rect 182081 269786 182147 269789
rect 207013 269786 207079 269789
rect 182081 269784 184092 269786
rect 154481 269726 156124 269728
rect 182081 269728 182086 269784
rect 182142 269728 184092 269784
rect 182081 269726 184092 269728
rect 204884 269784 207079 269786
rect 204884 269728 207018 269784
rect 207074 269728 207079 269784
rect 204884 269726 207079 269728
rect 154481 269723 154547 269726
rect 182081 269723 182147 269726
rect 207013 269723 207079 269726
rect 209681 269786 209747 269789
rect 234705 269786 234771 269789
rect 209681 269784 212060 269786
rect 209681 269728 209686 269784
rect 209742 269728 212060 269784
rect 209681 269726 212060 269728
rect 232852 269784 234771 269786
rect 232852 269728 234710 269784
rect 234766 269728 234771 269784
rect 232852 269726 234771 269728
rect 209681 269723 209747 269726
rect 234705 269723 234771 269726
rect 238661 269786 238727 269789
rect 262213 269786 262279 269789
rect 238661 269784 240212 269786
rect 238661 269728 238666 269784
rect 238722 269728 240212 269784
rect 238661 269726 240212 269728
rect 260820 269784 262279 269786
rect 260820 269728 262218 269784
rect 262274 269728 262279 269784
rect 260820 269726 262279 269728
rect 238661 269723 238727 269726
rect 262213 269723 262279 269726
rect 266261 269786 266327 269789
rect 291193 269786 291259 269789
rect 266261 269784 268180 269786
rect 266261 269728 266266 269784
rect 266322 269728 268180 269784
rect 266261 269726 268180 269728
rect 288788 269784 291259 269786
rect 288788 269728 291198 269784
rect 291254 269728 291259 269784
rect 288788 269726 291259 269728
rect 266261 269723 266327 269726
rect 291193 269723 291259 269726
rect 293861 269786 293927 269789
rect 318793 269786 318859 269789
rect 293861 269784 296148 269786
rect 293861 269728 293866 269784
rect 293922 269728 296148 269784
rect 293861 269726 296148 269728
rect 316940 269784 318859 269786
rect 316940 269728 318798 269784
rect 318854 269728 318859 269784
rect 316940 269726 318859 269728
rect 293861 269723 293927 269726
rect 318793 269723 318859 269726
rect 322841 269786 322907 269789
rect 346393 269786 346459 269789
rect 322841 269784 324116 269786
rect 322841 269728 322846 269784
rect 322902 269728 324116 269784
rect 322841 269726 324116 269728
rect 344908 269784 346459 269786
rect 344908 269728 346398 269784
rect 346454 269728 346459 269784
rect 344908 269726 346459 269728
rect 322841 269723 322907 269726
rect 346393 269723 346459 269726
rect 350441 269786 350507 269789
rect 375373 269786 375439 269789
rect 350441 269784 352084 269786
rect 350441 269728 350446 269784
rect 350502 269728 352084 269784
rect 350441 269726 352084 269728
rect 372876 269784 375439 269786
rect 372876 269728 375378 269784
rect 375434 269728 375439 269784
rect 372876 269726 375439 269728
rect 350441 269723 350507 269726
rect 375373 269723 375439 269726
rect 378041 269786 378107 269789
rect 402973 269786 403039 269789
rect 378041 269784 380052 269786
rect 378041 269728 378046 269784
rect 378102 269728 380052 269784
rect 378041 269726 380052 269728
rect 400844 269784 403039 269786
rect 400844 269728 402978 269784
rect 403034 269728 403039 269784
rect 400844 269726 403039 269728
rect 378041 269723 378107 269726
rect 402973 269723 403039 269726
rect 405641 269786 405707 269789
rect 430573 269786 430639 269789
rect 405641 269784 408204 269786
rect 405641 269728 405646 269784
rect 405702 269728 408204 269784
rect 405641 269726 408204 269728
rect 428812 269784 430639 269786
rect 428812 269728 430578 269784
rect 430634 269728 430639 269784
rect 428812 269726 430639 269728
rect 405641 269723 405707 269726
rect 430573 269723 430639 269726
rect 434621 269786 434687 269789
rect 434621 269784 436172 269786
rect 434621 269728 434626 269784
rect 434682 269728 436172 269784
rect 456382 269756 456442 270268
rect 568430 270132 568436 270196
rect 568500 270132 568506 270196
rect 462221 269786 462287 269789
rect 487153 269786 487219 269789
rect 462221 269784 464140 269786
rect 434621 269726 436172 269728
rect 462221 269728 462226 269784
rect 462282 269728 464140 269784
rect 462221 269726 464140 269728
rect 484932 269784 487219 269786
rect 484932 269728 487158 269784
rect 487214 269728 487219 269784
rect 484932 269726 487219 269728
rect 434621 269723 434687 269726
rect 462221 269723 462287 269726
rect 487153 269723 487219 269726
rect 489821 269786 489887 269789
rect 514753 269786 514819 269789
rect 489821 269784 492108 269786
rect 489821 269728 489826 269784
rect 489882 269728 492108 269784
rect 489821 269726 492108 269728
rect 512900 269784 514819 269786
rect 512900 269728 514758 269784
rect 514814 269728 514819 269784
rect 512900 269726 514819 269728
rect 489821 269723 489887 269726
rect 514753 269723 514819 269726
rect 518801 269786 518867 269789
rect 542353 269786 542419 269789
rect 518801 269784 520076 269786
rect 518801 269728 518806 269784
rect 518862 269728 520076 269784
rect 518801 269726 520076 269728
rect 540868 269784 542419 269786
rect 540868 269728 542358 269784
rect 542414 269728 542419 269784
rect 540868 269726 542419 269728
rect 518801 269723 518867 269726
rect 542353 269723 542419 269726
rect 546401 269786 546467 269789
rect 546401 269784 548044 269786
rect 546401 269728 546406 269784
rect 546462 269728 548044 269784
rect 568438 269756 568498 270132
rect 546401 269726 548044 269728
rect 546401 269723 546467 269726
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect 44633 256594 44699 256597
rect 81382 256594 81388 256596
rect 44633 256592 81388 256594
rect 44633 256536 44638 256592
rect 44694 256536 81388 256592
rect 44633 256534 81388 256536
rect 44633 256531 44699 256534
rect 81382 256532 81388 256534
rect 81452 256532 81458 256596
rect 110597 256594 110663 256597
rect 128302 256594 128308 256596
rect 110597 256592 128308 256594
rect 110597 256536 110602 256592
rect 110658 256536 128308 256592
rect 110597 256534 128308 256536
rect 110597 256531 110663 256534
rect 128302 256532 128308 256534
rect 128372 256532 128378 256596
rect 156321 256594 156387 256597
rect 194726 256594 194732 256596
rect 156321 256592 194732 256594
rect 156321 256536 156326 256592
rect 156382 256536 194732 256592
rect 156321 256534 194732 256536
rect 156321 256531 156387 256534
rect 194726 256532 194732 256534
rect 194796 256532 194802 256596
rect 240317 256594 240383 256597
rect 277158 256594 277164 256596
rect 240317 256592 277164 256594
rect 240317 256536 240322 256592
rect 240378 256536 277164 256592
rect 240317 256534 277164 256536
rect 240317 256531 240383 256534
rect 277158 256532 277164 256534
rect 277228 256532 277234 256596
rect 352649 256594 352715 256597
rect 390870 256594 390876 256596
rect 352649 256592 390876 256594
rect 352649 256536 352654 256592
rect 352710 256536 390876 256592
rect 352649 256534 390876 256536
rect 352649 256531 352715 256534
rect 390870 256532 390876 256534
rect 390940 256532 390946 256596
rect 436645 256594 436711 256597
rect 473486 256594 473492 256596
rect 436645 256592 473492 256594
rect 436645 256536 436650 256592
rect 436706 256536 473492 256592
rect 436645 256534 473492 256536
rect 436645 256531 436711 256534
rect 473486 256532 473492 256534
rect 473556 256532 473562 256596
rect 502609 256594 502675 256597
rect 520222 256594 520228 256596
rect 502609 256592 520228 256594
rect 502609 256536 502614 256592
rect 502670 256536 520228 256592
rect 502609 256534 520228 256536
rect 502609 256531 502675 256534
rect 520222 256532 520228 256534
rect 520292 256532 520298 256596
rect -960 254146 480 254236
rect 3969 254146 4035 254149
rect -960 254144 4035 254146
rect -960 254088 3974 254144
rect 4030 254088 4035 254144
rect -960 254086 4035 254088
rect -960 253996 480 254086
rect 3969 254083 4035 254086
rect 165654 252588 165660 252652
rect 165724 252650 165730 252652
rect 165981 252650 166047 252653
rect 165724 252648 166047 252650
rect 165724 252592 165986 252648
rect 166042 252592 166047 252648
rect 165724 252590 166047 252592
rect 165724 252588 165730 252590
rect 165981 252587 166047 252590
rect 259494 252588 259500 252652
rect 259564 252650 259570 252652
rect 260373 252650 260439 252653
rect 259564 252648 260439 252650
rect 259564 252592 260378 252648
rect 260434 252592 260439 252648
rect 259564 252590 260439 252592
rect 259564 252588 259570 252590
rect 260373 252587 260439 252590
rect 361614 252588 361620 252652
rect 361684 252650 361690 252652
rect 361941 252650 362007 252653
rect 361684 252648 362007 252650
rect 361684 252592 361946 252648
rect 362002 252592 362007 252648
rect 361684 252590 362007 252592
rect 361684 252588 361690 252590
rect 361941 252587 362007 252590
rect 445702 252588 445708 252652
rect 445772 252650 445778 252652
rect 446029 252650 446095 252653
rect 445772 252648 446095 252650
rect 445772 252592 446034 252648
rect 446090 252592 446095 252648
rect 445772 252590 446095 252592
rect 445772 252588 445778 252590
rect 446029 252587 446095 252590
rect 557574 252588 557580 252652
rect 557644 252650 557650 252652
rect 557993 252650 558059 252653
rect 557644 252648 558059 252650
rect 557644 252592 557998 252648
rect 558054 252592 558059 252648
rect 557644 252590 558059 252592
rect 557644 252588 557650 252590
rect 557993 252587 558059 252590
rect 583520 245428 584960 245668
rect 13537 242314 13603 242317
rect 38653 242314 38719 242317
rect 13537 242312 16100 242314
rect 13537 242256 13542 242312
rect 13598 242256 16100 242312
rect 13537 242254 16100 242256
rect 36892 242312 38719 242314
rect 36892 242256 38658 242312
rect 38714 242256 38719 242312
rect 36892 242254 38719 242256
rect 13537 242251 13603 242254
rect 38653 242251 38719 242254
rect 42701 242314 42767 242317
rect 66253 242314 66319 242317
rect 42701 242312 44068 242314
rect 42701 242256 42706 242312
rect 42762 242256 44068 242312
rect 42701 242254 44068 242256
rect 64860 242312 66319 242314
rect 64860 242256 66258 242312
rect 66314 242256 66319 242312
rect 64860 242254 66319 242256
rect 42701 242251 42767 242254
rect 66253 242251 66319 242254
rect 70301 242314 70367 242317
rect 95233 242314 95299 242317
rect 70301 242312 72036 242314
rect 70301 242256 70306 242312
rect 70362 242256 72036 242312
rect 70301 242254 72036 242256
rect 92828 242312 95299 242314
rect 92828 242256 95238 242312
rect 95294 242256 95299 242312
rect 92828 242254 95299 242256
rect 70301 242251 70367 242254
rect 95233 242251 95299 242254
rect 97901 242314 97967 242317
rect 122833 242314 122899 242317
rect 97901 242312 100188 242314
rect 97901 242256 97906 242312
rect 97962 242256 100188 242312
rect 97901 242254 100188 242256
rect 120796 242312 122899 242314
rect 120796 242256 122838 242312
rect 122894 242256 122899 242312
rect 120796 242254 122899 242256
rect 97901 242251 97967 242254
rect 122833 242251 122899 242254
rect 126881 242314 126947 242317
rect 150433 242314 150499 242317
rect 126881 242312 128156 242314
rect 126881 242256 126886 242312
rect 126942 242256 128156 242312
rect 126881 242254 128156 242256
rect 148948 242312 150499 242314
rect 148948 242256 150438 242312
rect 150494 242256 150499 242312
rect 148948 242254 150499 242256
rect 126881 242251 126947 242254
rect 150433 242251 150499 242254
rect 154481 242314 154547 242317
rect 178033 242314 178099 242317
rect 154481 242312 156124 242314
rect 154481 242256 154486 242312
rect 154542 242256 156124 242312
rect 154481 242254 156124 242256
rect 176916 242312 178099 242314
rect 176916 242256 178038 242312
rect 178094 242256 178099 242312
rect 176916 242254 178099 242256
rect 154481 242251 154547 242254
rect 178033 242251 178099 242254
rect 182081 242314 182147 242317
rect 207013 242314 207079 242317
rect 182081 242312 184092 242314
rect 182081 242256 182086 242312
rect 182142 242256 184092 242312
rect 182081 242254 184092 242256
rect 204884 242312 207079 242314
rect 204884 242256 207018 242312
rect 207074 242256 207079 242312
rect 204884 242254 207079 242256
rect 182081 242251 182147 242254
rect 207013 242251 207079 242254
rect 209681 242314 209747 242317
rect 234705 242314 234771 242317
rect 209681 242312 212060 242314
rect 209681 242256 209686 242312
rect 209742 242256 212060 242312
rect 209681 242254 212060 242256
rect 232852 242312 234771 242314
rect 232852 242256 234710 242312
rect 234766 242256 234771 242312
rect 232852 242254 234771 242256
rect 209681 242251 209747 242254
rect 234705 242251 234771 242254
rect 238661 242314 238727 242317
rect 262213 242314 262279 242317
rect 238661 242312 240212 242314
rect 238661 242256 238666 242312
rect 238722 242256 240212 242312
rect 238661 242254 240212 242256
rect 260820 242312 262279 242314
rect 260820 242256 262218 242312
rect 262274 242256 262279 242312
rect 260820 242254 262279 242256
rect 238661 242251 238727 242254
rect 262213 242251 262279 242254
rect 266261 242314 266327 242317
rect 291193 242314 291259 242317
rect 266261 242312 268180 242314
rect 266261 242256 266266 242312
rect 266322 242256 268180 242312
rect 266261 242254 268180 242256
rect 288788 242312 291259 242314
rect 288788 242256 291198 242312
rect 291254 242256 291259 242312
rect 288788 242254 291259 242256
rect 266261 242251 266327 242254
rect 291193 242251 291259 242254
rect 293861 242314 293927 242317
rect 318793 242314 318859 242317
rect 293861 242312 296148 242314
rect 293861 242256 293866 242312
rect 293922 242256 296148 242312
rect 293861 242254 296148 242256
rect 316940 242312 318859 242314
rect 316940 242256 318798 242312
rect 318854 242256 318859 242312
rect 316940 242254 318859 242256
rect 293861 242251 293927 242254
rect 318793 242251 318859 242254
rect 322841 242314 322907 242317
rect 346393 242314 346459 242317
rect 322841 242312 324116 242314
rect 322841 242256 322846 242312
rect 322902 242256 324116 242312
rect 322841 242254 324116 242256
rect 344908 242312 346459 242314
rect 344908 242256 346398 242312
rect 346454 242256 346459 242312
rect 344908 242254 346459 242256
rect 322841 242251 322907 242254
rect 346393 242251 346459 242254
rect 350441 242314 350507 242317
rect 375373 242314 375439 242317
rect 350441 242312 352084 242314
rect 350441 242256 350446 242312
rect 350502 242256 352084 242312
rect 350441 242254 352084 242256
rect 372876 242312 375439 242314
rect 372876 242256 375378 242312
rect 375434 242256 375439 242312
rect 372876 242254 375439 242256
rect 350441 242251 350507 242254
rect 375373 242251 375439 242254
rect 378041 242314 378107 242317
rect 402973 242314 403039 242317
rect 378041 242312 380052 242314
rect 378041 242256 378046 242312
rect 378102 242256 380052 242312
rect 378041 242254 380052 242256
rect 400844 242312 403039 242314
rect 400844 242256 402978 242312
rect 403034 242256 403039 242312
rect 400844 242254 403039 242256
rect 378041 242251 378107 242254
rect 402973 242251 403039 242254
rect 405641 242314 405707 242317
rect 430573 242314 430639 242317
rect 405641 242312 408204 242314
rect 405641 242256 405646 242312
rect 405702 242256 408204 242312
rect 405641 242254 408204 242256
rect 428812 242312 430639 242314
rect 428812 242256 430578 242312
rect 430634 242256 430639 242312
rect 428812 242254 430639 242256
rect 405641 242251 405707 242254
rect 430573 242251 430639 242254
rect 434621 242314 434687 242317
rect 458173 242314 458239 242317
rect 434621 242312 436172 242314
rect 434621 242256 434626 242312
rect 434682 242256 436172 242312
rect 434621 242254 436172 242256
rect 456964 242312 458239 242314
rect 456964 242256 458178 242312
rect 458234 242256 458239 242312
rect 456964 242254 458239 242256
rect 434621 242251 434687 242254
rect 458173 242251 458239 242254
rect 462221 242314 462287 242317
rect 487153 242314 487219 242317
rect 462221 242312 464140 242314
rect 462221 242256 462226 242312
rect 462282 242256 464140 242312
rect 462221 242254 464140 242256
rect 484932 242312 487219 242314
rect 484932 242256 487158 242312
rect 487214 242256 487219 242312
rect 484932 242254 487219 242256
rect 462221 242251 462287 242254
rect 487153 242251 487219 242254
rect 489821 242314 489887 242317
rect 514753 242314 514819 242317
rect 489821 242312 492108 242314
rect 489821 242256 489826 242312
rect 489882 242256 492108 242312
rect 489821 242254 492108 242256
rect 512900 242312 514819 242314
rect 512900 242256 514758 242312
rect 514814 242256 514819 242312
rect 512900 242254 514819 242256
rect 489821 242251 489887 242254
rect 514753 242251 514819 242254
rect 518801 242314 518867 242317
rect 542353 242314 542419 242317
rect 518801 242312 520076 242314
rect 518801 242256 518806 242312
rect 518862 242256 520076 242312
rect 518801 242254 520076 242256
rect 540868 242312 542419 242314
rect 540868 242256 542358 242312
rect 542414 242256 542419 242312
rect 540868 242254 542419 242256
rect 518801 242251 518867 242254
rect 542353 242251 542419 242254
rect 546401 242314 546467 242317
rect 571333 242314 571399 242317
rect 546401 242312 548044 242314
rect 546401 242256 546406 242312
rect 546462 242256 548044 242312
rect 546401 242254 548044 242256
rect 568836 242312 571399 242314
rect 568836 242256 571338 242312
rect 571394 242256 571399 242312
rect 568836 242254 571399 242256
rect 546401 242251 546467 242254
rect 571333 242251 571399 242254
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 13537 234018 13603 234021
rect 66253 234018 66319 234021
rect 13537 234016 66319 234018
rect 13537 233960 13542 234016
rect 13598 233960 66258 234016
rect 66314 233960 66319 234016
rect 13537 233958 66319 233960
rect 13537 233955 13603 233958
rect 66253 233955 66319 233958
rect 70301 234018 70367 234021
rect 122833 234018 122899 234021
rect 70301 234016 122899 234018
rect 70301 233960 70306 234016
rect 70362 233960 122838 234016
rect 122894 233960 122899 234016
rect 70301 233958 122899 233960
rect 70301 233955 70367 233958
rect 122833 233955 122899 233958
rect 126881 234018 126947 234021
rect 178033 234018 178099 234021
rect 126881 234016 178099 234018
rect 126881 233960 126886 234016
rect 126942 233960 178038 234016
rect 178094 233960 178099 234016
rect 126881 233958 178099 233960
rect 126881 233955 126947 233958
rect 178033 233955 178099 233958
rect 182081 234018 182147 234021
rect 234705 234018 234771 234021
rect 182081 234016 234771 234018
rect 182081 233960 182086 234016
rect 182142 233960 234710 234016
rect 234766 233960 234771 234016
rect 182081 233958 234771 233960
rect 182081 233955 182147 233958
rect 234705 233955 234771 233958
rect 238661 234018 238727 234021
rect 291193 234018 291259 234021
rect 238661 234016 291259 234018
rect 238661 233960 238666 234016
rect 238722 233960 291198 234016
rect 291254 233960 291259 234016
rect 238661 233958 291259 233960
rect 238661 233955 238727 233958
rect 291193 233955 291259 233958
rect 293861 234018 293927 234021
rect 346393 234018 346459 234021
rect 293861 234016 346459 234018
rect 293861 233960 293866 234016
rect 293922 233960 346398 234016
rect 346454 233960 346459 234016
rect 293861 233958 346459 233960
rect 293861 233955 293927 233958
rect 346393 233955 346459 233958
rect 350441 234018 350507 234021
rect 402973 234018 403039 234021
rect 350441 234016 403039 234018
rect 350441 233960 350446 234016
rect 350502 233960 402978 234016
rect 403034 233960 403039 234016
rect 350441 233958 403039 233960
rect 350441 233955 350507 233958
rect 402973 233955 403039 233958
rect 405641 234018 405707 234021
rect 458173 234018 458239 234021
rect 405641 234016 458239 234018
rect 405641 233960 405646 234016
rect 405702 233960 458178 234016
rect 458234 233960 458239 234016
rect 405641 233958 458239 233960
rect 405641 233955 405707 233958
rect 458173 233955 458239 233958
rect 462221 234018 462287 234021
rect 514753 234018 514819 234021
rect 462221 234016 514819 234018
rect 462221 233960 462226 234016
rect 462282 233960 514758 234016
rect 514814 233960 514819 234016
rect 462221 233958 514819 233960
rect 462221 233955 462287 233958
rect 514753 233955 514819 233958
rect 518801 234018 518867 234021
rect 571333 234018 571399 234021
rect 518801 234016 571399 234018
rect 518801 233960 518806 234016
rect 518862 233960 571338 234016
rect 571394 233960 571399 234016
rect 518801 233958 571399 233960
rect 518801 233955 518867 233958
rect 571333 233955 571399 233958
rect 580073 232386 580139 232389
rect 583520 232386 584960 232476
rect 580073 232384 584960 232386
rect 580073 232328 580078 232384
rect 580134 232328 584960 232384
rect 580073 232326 584960 232328
rect 580073 232323 580139 232326
rect 583520 232236 584960 232326
rect 148593 230482 148659 230485
rect 165654 230482 165660 230484
rect 148593 230480 165660 230482
rect 148593 230424 148598 230480
rect 148654 230424 165660 230480
rect 148593 230422 165660 230424
rect 148593 230419 148659 230422
rect 165654 230420 165660 230422
rect 165724 230420 165730 230484
rect 222653 230482 222719 230485
rect 259494 230482 259500 230484
rect 222653 230480 259500 230482
rect 222653 230424 222658 230480
rect 222714 230424 259500 230480
rect 222653 230422 259500 230424
rect 222653 230419 222719 230422
rect 259494 230420 259500 230422
rect 259564 230420 259570 230484
rect 344645 230482 344711 230485
rect 361614 230482 361620 230484
rect 344645 230480 361620 230482
rect 344645 230424 344650 230480
rect 344706 230424 361620 230480
rect 344645 230422 361620 230424
rect 344645 230419 344711 230422
rect 361614 230420 361620 230422
rect 361684 230420 361690 230484
rect 428641 230482 428707 230485
rect 445702 230482 445708 230484
rect 428641 230480 445708 230482
rect 428641 230424 428646 230480
rect 428702 230424 445708 230480
rect 428641 230422 445708 230424
rect 428641 230419 428707 230422
rect 445702 230420 445708 230422
rect 445772 230420 445778 230484
rect 540605 230482 540671 230485
rect 557574 230482 557580 230484
rect 540605 230480 557580 230482
rect 540605 230424 540610 230480
rect 540666 230424 557580 230480
rect 540605 230422 557580 230424
rect 540605 230419 540671 230422
rect 557574 230420 557580 230422
rect 557644 230420 557650 230484
rect -960 227884 480 228124
rect 128302 225252 128308 225316
rect 128372 225314 128378 225316
rect 128445 225314 128511 225317
rect 194777 225316 194843 225317
rect 194726 225314 194732 225316
rect 128372 225312 128511 225314
rect 128372 225256 128450 225312
rect 128506 225256 128511 225312
rect 128372 225254 128511 225256
rect 194686 225254 194732 225314
rect 194796 225312 194843 225316
rect 194838 225256 194843 225312
rect 128372 225252 128378 225254
rect 128445 225251 128511 225254
rect 194726 225252 194732 225254
rect 194796 225252 194843 225256
rect 194777 225251 194843 225252
rect 238661 224362 238727 224365
rect 288382 224362 288388 224364
rect 238661 224360 288388 224362
rect 238661 224304 238666 224360
rect 238722 224304 288388 224360
rect 238661 224302 288388 224304
rect 238661 224299 238727 224302
rect 288382 224300 288388 224302
rect 288452 224300 288458 224364
rect 42701 224226 42767 224229
rect 92422 224226 92428 224228
rect 42701 224224 92428 224226
rect 42701 224168 42706 224224
rect 42762 224168 92428 224224
rect 42701 224166 92428 224168
rect 42701 224163 42767 224166
rect 92422 224164 92428 224166
rect 92492 224164 92498 224228
rect 97901 224226 97967 224229
rect 148358 224226 148364 224228
rect 97901 224224 148364 224226
rect 97901 224168 97906 224224
rect 97962 224168 148364 224224
rect 97901 224166 148364 224168
rect 97901 224163 97967 224166
rect 148358 224164 148364 224166
rect 148428 224164 148434 224228
rect 154481 224226 154547 224229
rect 207013 224226 207079 224229
rect 154481 224224 207079 224226
rect 154481 224168 154486 224224
rect 154542 224168 207018 224224
rect 207074 224168 207079 224224
rect 154481 224166 207079 224168
rect 154481 224163 154547 224166
rect 207013 224163 207079 224166
rect 209681 224226 209747 224229
rect 260414 224226 260420 224228
rect 209681 224224 260420 224226
rect 209681 224168 209686 224224
rect 209742 224168 260420 224224
rect 209681 224166 260420 224168
rect 209681 224163 209747 224166
rect 260414 224164 260420 224166
rect 260484 224164 260490 224228
rect 378041 224226 378107 224229
rect 430573 224226 430639 224229
rect 378041 224224 430639 224226
rect 378041 224168 378046 224224
rect 378102 224168 430578 224224
rect 430634 224168 430639 224224
rect 378041 224166 430639 224168
rect 378041 224163 378107 224166
rect 430573 224163 430639 224166
rect 492622 224164 492628 224228
rect 492692 224226 492698 224228
rect 542353 224226 542419 224229
rect 492692 224224 542419 224226
rect 492692 224168 542358 224224
rect 542414 224168 542419 224224
rect 492692 224166 542419 224168
rect 492692 224164 492698 224166
rect 542353 224163 542419 224166
rect 13537 224090 13603 224093
rect 64454 224090 64460 224092
rect 13537 224088 64460 224090
rect 13537 224032 13542 224088
rect 13598 224032 64460 224088
rect 13537 224030 64460 224032
rect 13537 224027 13603 224030
rect 64454 224028 64460 224030
rect 64524 224028 64530 224092
rect 70301 224090 70367 224093
rect 122833 224090 122899 224093
rect 70301 224088 122899 224090
rect 70301 224032 70306 224088
rect 70362 224032 122838 224088
rect 122894 224032 122899 224088
rect 70301 224030 122899 224032
rect 70301 224027 70367 224030
rect 122833 224027 122899 224030
rect 126881 224090 126947 224093
rect 176326 224090 176332 224092
rect 126881 224088 176332 224090
rect 126881 224032 126886 224088
rect 126942 224032 176332 224088
rect 126881 224030 176332 224032
rect 126881 224027 126947 224030
rect 176326 224028 176332 224030
rect 176396 224028 176402 224092
rect 182081 224090 182147 224093
rect 234705 224090 234771 224093
rect 182081 224088 234771 224090
rect 182081 224032 182086 224088
rect 182142 224032 234710 224088
rect 234766 224032 234771 224088
rect 182081 224030 234771 224032
rect 182081 224027 182147 224030
rect 234705 224027 234771 224030
rect 266261 224090 266327 224093
rect 318793 224090 318859 224093
rect 266261 224088 318859 224090
rect 266261 224032 266266 224088
rect 266322 224032 318798 224088
rect 318854 224032 318859 224088
rect 266261 224030 318859 224032
rect 266261 224027 266327 224030
rect 318793 224027 318859 224030
rect 350441 224090 350507 224093
rect 402973 224090 403039 224093
rect 350441 224088 403039 224090
rect 350441 224032 350446 224088
rect 350502 224032 402978 224088
rect 403034 224032 403039 224088
rect 350441 224030 403039 224032
rect 350441 224027 350507 224030
rect 402973 224027 403039 224030
rect 462221 224090 462287 224093
rect 514753 224090 514819 224093
rect 462221 224088 514819 224090
rect 462221 224032 462226 224088
rect 462282 224032 514758 224088
rect 514814 224032 514819 224088
rect 462221 224030 514819 224032
rect 462221 224027 462287 224030
rect 514753 224027 514819 224030
rect 520590 224028 520596 224092
rect 520660 224090 520666 224092
rect 571333 224090 571399 224093
rect 520660 224088 571399 224090
rect 520660 224032 571338 224088
rect 571394 224032 571399 224088
rect 520660 224030 571399 224032
rect 520660 224028 520666 224030
rect 571333 224027 571399 224030
rect 583520 218908 584960 219148
rect 64454 216276 64460 216340
rect 64524 216276 64530 216340
rect 92422 216276 92428 216340
rect 92492 216276 92498 216340
rect 148358 216276 148364 216340
rect 148428 216276 148434 216340
rect 176326 216276 176332 216340
rect 176396 216276 176402 216340
rect 260414 216276 260420 216340
rect 260484 216276 260490 216340
rect 288382 216276 288388 216340
rect 288452 216276 288458 216340
rect 492622 216276 492628 216340
rect 492692 216276 492698 216340
rect 520590 216276 520596 216340
rect 520660 216276 520666 216340
rect 13537 215794 13603 215797
rect 38653 215794 38719 215797
rect 13537 215792 16100 215794
rect 13537 215736 13542 215792
rect 13598 215736 16100 215792
rect 13537 215734 16100 215736
rect 36892 215792 38719 215794
rect 36892 215736 38658 215792
rect 38714 215736 38719 215792
rect 36892 215734 38719 215736
rect 13537 215731 13603 215734
rect 38653 215731 38719 215734
rect 42701 215794 42767 215797
rect 42701 215792 44068 215794
rect 42701 215736 42706 215792
rect 42762 215736 44068 215792
rect 64462 215764 64522 216276
rect 70301 215794 70367 215797
rect 70301 215792 72036 215794
rect 42701 215734 44068 215736
rect 70301 215736 70306 215792
rect 70362 215736 72036 215792
rect 92430 215764 92490 216276
rect 97901 215794 97967 215797
rect 122833 215794 122899 215797
rect 97901 215792 100188 215794
rect 70301 215734 72036 215736
rect 97901 215736 97906 215792
rect 97962 215736 100188 215792
rect 97901 215734 100188 215736
rect 120796 215792 122899 215794
rect 120796 215736 122838 215792
rect 122894 215736 122899 215792
rect 120796 215734 122899 215736
rect 42701 215731 42767 215734
rect 70301 215731 70367 215734
rect 97901 215731 97967 215734
rect 122833 215731 122899 215734
rect 126881 215794 126947 215797
rect 126881 215792 128156 215794
rect 126881 215736 126886 215792
rect 126942 215736 128156 215792
rect 148366 215764 148426 216276
rect 154481 215794 154547 215797
rect 154481 215792 156124 215794
rect 126881 215734 128156 215736
rect 154481 215736 154486 215792
rect 154542 215736 156124 215792
rect 176334 215764 176394 216276
rect 182081 215794 182147 215797
rect 207013 215794 207079 215797
rect 182081 215792 184092 215794
rect 154481 215734 156124 215736
rect 182081 215736 182086 215792
rect 182142 215736 184092 215792
rect 182081 215734 184092 215736
rect 204884 215792 207079 215794
rect 204884 215736 207018 215792
rect 207074 215736 207079 215792
rect 204884 215734 207079 215736
rect 126881 215731 126947 215734
rect 154481 215731 154547 215734
rect 182081 215731 182147 215734
rect 207013 215731 207079 215734
rect 209681 215794 209747 215797
rect 234705 215794 234771 215797
rect 209681 215792 212060 215794
rect 209681 215736 209686 215792
rect 209742 215736 212060 215792
rect 209681 215734 212060 215736
rect 232852 215792 234771 215794
rect 232852 215736 234710 215792
rect 234766 215736 234771 215792
rect 232852 215734 234771 215736
rect 209681 215731 209747 215734
rect 234705 215731 234771 215734
rect 238661 215794 238727 215797
rect 238661 215792 240212 215794
rect 238661 215736 238666 215792
rect 238722 215736 240212 215792
rect 260422 215764 260482 216276
rect 266261 215794 266327 215797
rect 266261 215792 268180 215794
rect 238661 215734 240212 215736
rect 266261 215736 266266 215792
rect 266322 215736 268180 215792
rect 288390 215764 288450 216276
rect 293861 215794 293927 215797
rect 318793 215794 318859 215797
rect 293861 215792 296148 215794
rect 266261 215734 268180 215736
rect 293861 215736 293866 215792
rect 293922 215736 296148 215792
rect 293861 215734 296148 215736
rect 316940 215792 318859 215794
rect 316940 215736 318798 215792
rect 318854 215736 318859 215792
rect 316940 215734 318859 215736
rect 238661 215731 238727 215734
rect 266261 215731 266327 215734
rect 293861 215731 293927 215734
rect 318793 215731 318859 215734
rect 322841 215794 322907 215797
rect 346393 215794 346459 215797
rect 322841 215792 324116 215794
rect 322841 215736 322846 215792
rect 322902 215736 324116 215792
rect 322841 215734 324116 215736
rect 344908 215792 346459 215794
rect 344908 215736 346398 215792
rect 346454 215736 346459 215792
rect 344908 215734 346459 215736
rect 322841 215731 322907 215734
rect 346393 215731 346459 215734
rect 350441 215794 350507 215797
rect 375373 215794 375439 215797
rect 350441 215792 352084 215794
rect 350441 215736 350446 215792
rect 350502 215736 352084 215792
rect 350441 215734 352084 215736
rect 372876 215792 375439 215794
rect 372876 215736 375378 215792
rect 375434 215736 375439 215792
rect 372876 215734 375439 215736
rect 350441 215731 350507 215734
rect 375373 215731 375439 215734
rect 378041 215794 378107 215797
rect 402973 215794 403039 215797
rect 378041 215792 380052 215794
rect 378041 215736 378046 215792
rect 378102 215736 380052 215792
rect 378041 215734 380052 215736
rect 400844 215792 403039 215794
rect 400844 215736 402978 215792
rect 403034 215736 403039 215792
rect 400844 215734 403039 215736
rect 378041 215731 378107 215734
rect 402973 215731 403039 215734
rect 405641 215794 405707 215797
rect 430573 215794 430639 215797
rect 405641 215792 408204 215794
rect 405641 215736 405646 215792
rect 405702 215736 408204 215792
rect 405641 215734 408204 215736
rect 428812 215792 430639 215794
rect 428812 215736 430578 215792
rect 430634 215736 430639 215792
rect 428812 215734 430639 215736
rect 405641 215731 405707 215734
rect 430573 215731 430639 215734
rect 434621 215794 434687 215797
rect 458173 215794 458239 215797
rect 434621 215792 436172 215794
rect 434621 215736 434626 215792
rect 434682 215736 436172 215792
rect 434621 215734 436172 215736
rect 456964 215792 458239 215794
rect 456964 215736 458178 215792
rect 458234 215736 458239 215792
rect 456964 215734 458239 215736
rect 434621 215731 434687 215734
rect 458173 215731 458239 215734
rect 462221 215794 462287 215797
rect 487153 215794 487219 215797
rect 462221 215792 464140 215794
rect 462221 215736 462226 215792
rect 462282 215736 464140 215792
rect 462221 215734 464140 215736
rect 484932 215792 487219 215794
rect 484932 215736 487158 215792
rect 487214 215736 487219 215792
rect 492630 215764 492690 216276
rect 514753 215794 514819 215797
rect 512900 215792 514819 215794
rect 484932 215734 487219 215736
rect 512900 215736 514758 215792
rect 514814 215736 514819 215792
rect 520598 215764 520658 216276
rect 542353 215794 542419 215797
rect 540868 215792 542419 215794
rect 512900 215734 514819 215736
rect 540868 215736 542358 215792
rect 542414 215736 542419 215792
rect 540868 215734 542419 215736
rect 462221 215731 462287 215734
rect 487153 215731 487219 215734
rect 514753 215731 514819 215734
rect 542353 215731 542419 215734
rect 546401 215794 546467 215797
rect 571333 215794 571399 215797
rect 546401 215792 548044 215794
rect 546401 215736 546406 215792
rect 546462 215736 548044 215792
rect 546401 215734 548044 215736
rect 568836 215792 571399 215794
rect 568836 215736 571338 215792
rect 571394 215736 571399 215792
rect 568836 215734 571399 215736
rect 546401 215731 546467 215734
rect 571333 215731 571399 215734
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect 110597 202874 110663 202877
rect 128302 202874 128308 202876
rect 110597 202872 128308 202874
rect 110597 202816 110602 202872
rect 110658 202816 128308 202872
rect 110597 202814 128308 202816
rect 110597 202811 110663 202814
rect 128302 202812 128308 202814
rect 128372 202812 128378 202876
rect 156321 202874 156387 202877
rect 194726 202874 194732 202876
rect 156321 202872 194732 202874
rect 156321 202816 156326 202872
rect 156382 202816 194732 202872
rect 156321 202814 194732 202816
rect 156321 202811 156387 202814
rect 194726 202812 194732 202814
rect 194796 202812 194802 202876
rect -960 201922 480 202012
rect -960 201862 6930 201922
rect -960 201772 480 201862
rect 6870 201514 6930 201862
rect 63718 201514 63724 201516
rect 6870 201454 63724 201514
rect 63718 201452 63724 201454
rect 63788 201452 63794 201516
rect 259494 198460 259500 198524
rect 259564 198522 259570 198524
rect 260373 198522 260439 198525
rect 259564 198520 260439 198522
rect 259564 198464 260378 198520
rect 260434 198464 260439 198520
rect 259564 198462 260439 198464
rect 259564 198460 259570 198462
rect 260373 198459 260439 198462
rect 361614 198460 361620 198524
rect 361684 198522 361690 198524
rect 361941 198522 362007 198525
rect 361684 198520 362007 198522
rect 361684 198464 361946 198520
rect 362002 198464 362007 198520
rect 361684 198462 362007 198464
rect 361684 198460 361690 198462
rect 361941 198459 362007 198462
rect 445702 198460 445708 198524
rect 445772 198522 445778 198524
rect 446029 198522 446095 198525
rect 445772 198520 446095 198522
rect 445772 198464 446034 198520
rect 446090 198464 446095 198520
rect 445772 198462 446095 198464
rect 445772 198460 445778 198462
rect 446029 198459 446095 198462
rect 13537 196754 13603 196757
rect 66253 196754 66319 196757
rect 13537 196752 66319 196754
rect 13537 196696 13542 196752
rect 13598 196696 66258 196752
rect 66314 196696 66319 196752
rect 13537 196694 66319 196696
rect 13537 196691 13603 196694
rect 66253 196691 66319 196694
rect 70301 196754 70367 196757
rect 122833 196754 122899 196757
rect 70301 196752 122899 196754
rect 70301 196696 70306 196752
rect 70362 196696 122838 196752
rect 122894 196696 122899 196752
rect 70301 196694 122899 196696
rect 70301 196691 70367 196694
rect 122833 196691 122899 196694
rect 126881 196754 126947 196757
rect 178033 196754 178099 196757
rect 126881 196752 178099 196754
rect 126881 196696 126886 196752
rect 126942 196696 178038 196752
rect 178094 196696 178099 196752
rect 126881 196694 178099 196696
rect 126881 196691 126947 196694
rect 178033 196691 178099 196694
rect 182081 196754 182147 196757
rect 234705 196754 234771 196757
rect 182081 196752 234771 196754
rect 182081 196696 182086 196752
rect 182142 196696 234710 196752
rect 234766 196696 234771 196752
rect 182081 196694 234771 196696
rect 182081 196691 182147 196694
rect 234705 196691 234771 196694
rect 238661 196754 238727 196757
rect 291193 196754 291259 196757
rect 238661 196752 291259 196754
rect 238661 196696 238666 196752
rect 238722 196696 291198 196752
rect 291254 196696 291259 196752
rect 238661 196694 291259 196696
rect 238661 196691 238727 196694
rect 291193 196691 291259 196694
rect 293861 196754 293927 196757
rect 346393 196754 346459 196757
rect 293861 196752 346459 196754
rect 293861 196696 293866 196752
rect 293922 196696 346398 196752
rect 346454 196696 346459 196752
rect 293861 196694 346459 196696
rect 293861 196691 293927 196694
rect 346393 196691 346459 196694
rect 350441 196754 350507 196757
rect 402973 196754 403039 196757
rect 350441 196752 403039 196754
rect 350441 196696 350446 196752
rect 350502 196696 402978 196752
rect 403034 196696 403039 196752
rect 350441 196694 403039 196696
rect 350441 196691 350507 196694
rect 402973 196691 403039 196694
rect 405641 196754 405707 196757
rect 458173 196754 458239 196757
rect 405641 196752 458239 196754
rect 405641 196696 405646 196752
rect 405702 196696 458178 196752
rect 458234 196696 458239 196752
rect 405641 196694 458239 196696
rect 405641 196691 405707 196694
rect 458173 196691 458239 196694
rect 462221 196754 462287 196757
rect 514753 196754 514819 196757
rect 462221 196752 514819 196754
rect 462221 196696 462226 196752
rect 462282 196696 514758 196752
rect 514814 196696 514819 196752
rect 462221 196694 514819 196696
rect 462221 196691 462287 196694
rect 514753 196691 514819 196694
rect 518801 196754 518867 196757
rect 571333 196754 571399 196757
rect 518801 196752 571399 196754
rect 518801 196696 518806 196752
rect 518862 196696 571338 196752
rect 571394 196696 571399 196752
rect 518801 196694 571399 196696
rect 518801 196691 518867 196694
rect 571333 196691 571399 196694
rect 580073 192538 580139 192541
rect 583520 192538 584960 192628
rect 580073 192536 584960 192538
rect 580073 192480 580078 192536
rect 580134 192480 584960 192536
rect 580073 192478 584960 192480
rect 580073 192475 580139 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 2773 188866 2839 188869
rect -960 188864 2839 188866
rect -960 188808 2778 188864
rect 2834 188808 2839 188864
rect -960 188806 2839 188808
rect -960 188716 480 188806
rect 2773 188803 2839 188806
rect 13537 188322 13603 188325
rect 38653 188322 38719 188325
rect 13537 188320 16100 188322
rect 13537 188264 13542 188320
rect 13598 188264 16100 188320
rect 13537 188262 16100 188264
rect 36892 188320 38719 188322
rect 36892 188264 38658 188320
rect 38714 188264 38719 188320
rect 36892 188262 38719 188264
rect 13537 188259 13603 188262
rect 38653 188259 38719 188262
rect 42701 188322 42767 188325
rect 66253 188322 66319 188325
rect 42701 188320 44068 188322
rect 42701 188264 42706 188320
rect 42762 188264 44068 188320
rect 42701 188262 44068 188264
rect 64860 188320 66319 188322
rect 64860 188264 66258 188320
rect 66314 188264 66319 188320
rect 64860 188262 66319 188264
rect 42701 188259 42767 188262
rect 66253 188259 66319 188262
rect 70301 188322 70367 188325
rect 95233 188322 95299 188325
rect 70301 188320 72036 188322
rect 70301 188264 70306 188320
rect 70362 188264 72036 188320
rect 70301 188262 72036 188264
rect 92828 188320 95299 188322
rect 92828 188264 95238 188320
rect 95294 188264 95299 188320
rect 92828 188262 95299 188264
rect 70301 188259 70367 188262
rect 95233 188259 95299 188262
rect 97901 188322 97967 188325
rect 122833 188322 122899 188325
rect 97901 188320 100188 188322
rect 97901 188264 97906 188320
rect 97962 188264 100188 188320
rect 97901 188262 100188 188264
rect 120796 188320 122899 188322
rect 120796 188264 122838 188320
rect 122894 188264 122899 188320
rect 120796 188262 122899 188264
rect 97901 188259 97967 188262
rect 122833 188259 122899 188262
rect 126881 188322 126947 188325
rect 150433 188322 150499 188325
rect 126881 188320 128156 188322
rect 126881 188264 126886 188320
rect 126942 188264 128156 188320
rect 126881 188262 128156 188264
rect 148948 188320 150499 188322
rect 148948 188264 150438 188320
rect 150494 188264 150499 188320
rect 148948 188262 150499 188264
rect 126881 188259 126947 188262
rect 150433 188259 150499 188262
rect 154481 188322 154547 188325
rect 178033 188322 178099 188325
rect 154481 188320 156124 188322
rect 154481 188264 154486 188320
rect 154542 188264 156124 188320
rect 154481 188262 156124 188264
rect 176916 188320 178099 188322
rect 176916 188264 178038 188320
rect 178094 188264 178099 188320
rect 176916 188262 178099 188264
rect 154481 188259 154547 188262
rect 178033 188259 178099 188262
rect 182081 188322 182147 188325
rect 207013 188322 207079 188325
rect 182081 188320 184092 188322
rect 182081 188264 182086 188320
rect 182142 188264 184092 188320
rect 182081 188262 184092 188264
rect 204884 188320 207079 188322
rect 204884 188264 207018 188320
rect 207074 188264 207079 188320
rect 204884 188262 207079 188264
rect 182081 188259 182147 188262
rect 207013 188259 207079 188262
rect 209681 188322 209747 188325
rect 234705 188322 234771 188325
rect 209681 188320 212060 188322
rect 209681 188264 209686 188320
rect 209742 188264 212060 188320
rect 209681 188262 212060 188264
rect 232852 188320 234771 188322
rect 232852 188264 234710 188320
rect 234766 188264 234771 188320
rect 232852 188262 234771 188264
rect 209681 188259 209747 188262
rect 234705 188259 234771 188262
rect 238661 188322 238727 188325
rect 262213 188322 262279 188325
rect 238661 188320 240212 188322
rect 238661 188264 238666 188320
rect 238722 188264 240212 188320
rect 238661 188262 240212 188264
rect 260820 188320 262279 188322
rect 260820 188264 262218 188320
rect 262274 188264 262279 188320
rect 260820 188262 262279 188264
rect 238661 188259 238727 188262
rect 262213 188259 262279 188262
rect 266261 188322 266327 188325
rect 291193 188322 291259 188325
rect 266261 188320 268180 188322
rect 266261 188264 266266 188320
rect 266322 188264 268180 188320
rect 266261 188262 268180 188264
rect 288788 188320 291259 188322
rect 288788 188264 291198 188320
rect 291254 188264 291259 188320
rect 288788 188262 291259 188264
rect 266261 188259 266327 188262
rect 291193 188259 291259 188262
rect 293861 188322 293927 188325
rect 318793 188322 318859 188325
rect 293861 188320 296148 188322
rect 293861 188264 293866 188320
rect 293922 188264 296148 188320
rect 293861 188262 296148 188264
rect 316940 188320 318859 188322
rect 316940 188264 318798 188320
rect 318854 188264 318859 188320
rect 316940 188262 318859 188264
rect 293861 188259 293927 188262
rect 318793 188259 318859 188262
rect 322841 188322 322907 188325
rect 346393 188322 346459 188325
rect 322841 188320 324116 188322
rect 322841 188264 322846 188320
rect 322902 188264 324116 188320
rect 322841 188262 324116 188264
rect 344908 188320 346459 188322
rect 344908 188264 346398 188320
rect 346454 188264 346459 188320
rect 344908 188262 346459 188264
rect 322841 188259 322907 188262
rect 346393 188259 346459 188262
rect 350441 188322 350507 188325
rect 375373 188322 375439 188325
rect 350441 188320 352084 188322
rect 350441 188264 350446 188320
rect 350502 188264 352084 188320
rect 350441 188262 352084 188264
rect 372876 188320 375439 188322
rect 372876 188264 375378 188320
rect 375434 188264 375439 188320
rect 372876 188262 375439 188264
rect 350441 188259 350507 188262
rect 375373 188259 375439 188262
rect 378041 188322 378107 188325
rect 402973 188322 403039 188325
rect 378041 188320 380052 188322
rect 378041 188264 378046 188320
rect 378102 188264 380052 188320
rect 378041 188262 380052 188264
rect 400844 188320 403039 188322
rect 400844 188264 402978 188320
rect 403034 188264 403039 188320
rect 400844 188262 403039 188264
rect 378041 188259 378107 188262
rect 402973 188259 403039 188262
rect 405641 188322 405707 188325
rect 430573 188322 430639 188325
rect 405641 188320 408204 188322
rect 405641 188264 405646 188320
rect 405702 188264 408204 188320
rect 405641 188262 408204 188264
rect 428812 188320 430639 188322
rect 428812 188264 430578 188320
rect 430634 188264 430639 188320
rect 428812 188262 430639 188264
rect 405641 188259 405707 188262
rect 430573 188259 430639 188262
rect 434621 188322 434687 188325
rect 458173 188322 458239 188325
rect 434621 188320 436172 188322
rect 434621 188264 434626 188320
rect 434682 188264 436172 188320
rect 434621 188262 436172 188264
rect 456964 188320 458239 188322
rect 456964 188264 458178 188320
rect 458234 188264 458239 188320
rect 456964 188262 458239 188264
rect 434621 188259 434687 188262
rect 458173 188259 458239 188262
rect 462221 188322 462287 188325
rect 487153 188322 487219 188325
rect 462221 188320 464140 188322
rect 462221 188264 462226 188320
rect 462282 188264 464140 188320
rect 462221 188262 464140 188264
rect 484932 188320 487219 188322
rect 484932 188264 487158 188320
rect 487214 188264 487219 188320
rect 484932 188262 487219 188264
rect 462221 188259 462287 188262
rect 487153 188259 487219 188262
rect 489821 188322 489887 188325
rect 514753 188322 514819 188325
rect 489821 188320 492108 188322
rect 489821 188264 489826 188320
rect 489882 188264 492108 188320
rect 489821 188262 492108 188264
rect 512900 188320 514819 188322
rect 512900 188264 514758 188320
rect 514814 188264 514819 188320
rect 512900 188262 514819 188264
rect 489821 188259 489887 188262
rect 514753 188259 514819 188262
rect 518801 188322 518867 188325
rect 542353 188322 542419 188325
rect 518801 188320 520076 188322
rect 518801 188264 518806 188320
rect 518862 188264 520076 188320
rect 518801 188262 520076 188264
rect 540868 188320 542419 188322
rect 540868 188264 542358 188320
rect 542414 188264 542419 188320
rect 540868 188262 542419 188264
rect 518801 188259 518867 188262
rect 542353 188259 542419 188262
rect 546401 188322 546467 188325
rect 571333 188322 571399 188325
rect 546401 188320 548044 188322
rect 546401 188264 546406 188320
rect 546462 188264 548044 188320
rect 546401 188262 548044 188264
rect 568836 188320 571399 188322
rect 568836 188264 571338 188320
rect 571394 188264 571399 188320
rect 568836 188262 571399 188264
rect 546401 188259 546467 188262
rect 571333 188259 571399 188262
rect 583520 179060 584960 179300
rect 222653 176626 222719 176629
rect 259494 176626 259500 176628
rect 222653 176624 259500 176626
rect 222653 176568 222658 176624
rect 222714 176568 259500 176624
rect 222653 176566 259500 176568
rect 222653 176563 222719 176566
rect 259494 176564 259500 176566
rect 259564 176564 259570 176628
rect 344645 176626 344711 176629
rect 361614 176626 361620 176628
rect 344645 176624 361620 176626
rect 344645 176568 344650 176624
rect 344706 176568 361620 176624
rect 344645 176566 361620 176568
rect 344645 176563 344711 176566
rect 361614 176564 361620 176566
rect 361684 176564 361690 176628
rect 428641 176626 428707 176629
rect 445702 176626 445708 176628
rect 428641 176624 445708 176626
rect 428641 176568 428646 176624
rect 428702 176568 445708 176624
rect 428641 176566 445708 176568
rect 428641 176563 428707 176566
rect 445702 176564 445708 176566
rect 445772 176564 445778 176628
rect -960 175796 480 176036
rect 97901 170642 97967 170645
rect 148358 170642 148364 170644
rect 97901 170640 148364 170642
rect 97901 170584 97906 170640
rect 97962 170584 148364 170640
rect 97901 170582 148364 170584
rect 97901 170579 97967 170582
rect 148358 170580 148364 170582
rect 148428 170580 148434 170644
rect 128486 170308 128492 170372
rect 128556 170370 128562 170372
rect 178033 170370 178099 170373
rect 128556 170368 178099 170370
rect 128556 170312 178038 170368
rect 178094 170312 178099 170368
rect 128556 170310 178099 170312
rect 128556 170308 128562 170310
rect 178033 170307 178099 170310
rect 322841 170370 322907 170373
rect 372286 170370 372292 170372
rect 322841 170368 372292 170370
rect 322841 170312 322846 170368
rect 322902 170312 372292 170368
rect 322841 170310 372292 170312
rect 322841 170307 322907 170310
rect 372286 170308 372292 170310
rect 372356 170308 372362 170372
rect 154481 170234 154547 170237
rect 207013 170234 207079 170237
rect 154481 170232 207079 170234
rect 154481 170176 154486 170232
rect 154542 170176 207018 170232
rect 207074 170176 207079 170232
rect 154481 170174 207079 170176
rect 154481 170171 154547 170174
rect 207013 170171 207079 170174
rect 293861 170234 293927 170237
rect 344318 170234 344324 170236
rect 293861 170232 344324 170234
rect 293861 170176 293866 170232
rect 293922 170176 344324 170232
rect 293861 170174 344324 170176
rect 293861 170171 293927 170174
rect 344318 170172 344324 170174
rect 344388 170172 344394 170236
rect 378041 170234 378107 170237
rect 430573 170234 430639 170237
rect 378041 170232 430639 170234
rect 378041 170176 378046 170232
rect 378102 170176 430578 170232
rect 430634 170176 430639 170232
rect 378041 170174 430639 170176
rect 378041 170171 378107 170174
rect 430573 170171 430639 170174
rect 489821 170234 489887 170237
rect 540462 170234 540468 170236
rect 489821 170232 540468 170234
rect 489821 170176 489826 170232
rect 489882 170176 540468 170232
rect 489821 170174 540468 170176
rect 489821 170171 489887 170174
rect 540462 170172 540468 170174
rect 540532 170172 540538 170236
rect 42701 170098 42767 170101
rect 95233 170098 95299 170101
rect 42701 170096 95299 170098
rect 42701 170040 42706 170096
rect 42762 170040 95238 170096
rect 95294 170040 95299 170096
rect 42701 170038 95299 170040
rect 42701 170035 42767 170038
rect 95233 170035 95299 170038
rect 182081 170098 182147 170101
rect 234705 170098 234771 170101
rect 182081 170096 234771 170098
rect 182081 170040 182086 170096
rect 182142 170040 234710 170096
rect 234766 170040 234771 170096
rect 182081 170038 234771 170040
rect 182081 170035 182147 170038
rect 234705 170035 234771 170038
rect 266261 170098 266327 170101
rect 318793 170098 318859 170101
rect 266261 170096 318859 170098
rect 266261 170040 266266 170096
rect 266322 170040 318798 170096
rect 318854 170040 318859 170096
rect 266261 170038 318859 170040
rect 266261 170035 266327 170038
rect 318793 170035 318859 170038
rect 350441 170098 350507 170101
rect 402973 170098 403039 170101
rect 350441 170096 403039 170098
rect 350441 170040 350446 170096
rect 350502 170040 402978 170096
rect 403034 170040 403039 170096
rect 350441 170038 403039 170040
rect 350441 170035 350507 170038
rect 402973 170035 403039 170038
rect 408534 170036 408540 170100
rect 408604 170098 408610 170100
rect 458173 170098 458239 170101
rect 408604 170096 458239 170098
rect 408604 170040 458178 170096
rect 458234 170040 458239 170096
rect 408604 170038 458239 170040
rect 408604 170036 408610 170038
rect 458173 170035 458239 170038
rect 520590 170036 520596 170100
rect 520660 170098 520666 170100
rect 571333 170098 571399 170101
rect 520660 170096 571399 170098
rect 520660 170040 571338 170096
rect 571394 170040 571399 170096
rect 520660 170038 571399 170040
rect 520660 170036 520666 170038
rect 571333 170035 571399 170038
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 128486 162284 128492 162348
rect 128556 162284 128562 162348
rect 148358 162284 148364 162348
rect 148428 162284 148434 162348
rect 344318 162284 344324 162348
rect 344388 162284 344394 162348
rect 372286 162284 372292 162348
rect 372356 162284 372362 162348
rect 408534 162284 408540 162348
rect 408604 162284 408610 162348
rect 520590 162284 520596 162348
rect 520660 162284 520666 162348
rect 540462 162284 540468 162348
rect 540532 162284 540538 162348
rect 13537 161802 13603 161805
rect 38653 161802 38719 161805
rect 13537 161800 16100 161802
rect 13537 161744 13542 161800
rect 13598 161744 16100 161800
rect 13537 161742 16100 161744
rect 36892 161800 38719 161802
rect 36892 161744 38658 161800
rect 38714 161744 38719 161800
rect 36892 161742 38719 161744
rect 13537 161739 13603 161742
rect 38653 161739 38719 161742
rect 42701 161802 42767 161805
rect 66253 161802 66319 161805
rect 42701 161800 44068 161802
rect 42701 161744 42706 161800
rect 42762 161744 44068 161800
rect 42701 161742 44068 161744
rect 64860 161800 66319 161802
rect 64860 161744 66258 161800
rect 66314 161744 66319 161800
rect 64860 161742 66319 161744
rect 42701 161739 42767 161742
rect 66253 161739 66319 161742
rect 70301 161802 70367 161805
rect 95233 161802 95299 161805
rect 70301 161800 72036 161802
rect 70301 161744 70306 161800
rect 70362 161744 72036 161800
rect 70301 161742 72036 161744
rect 92828 161800 95299 161802
rect 92828 161744 95238 161800
rect 95294 161744 95299 161800
rect 92828 161742 95299 161744
rect 70301 161739 70367 161742
rect 95233 161739 95299 161742
rect 97901 161802 97967 161805
rect 122833 161802 122899 161805
rect 97901 161800 100188 161802
rect 97901 161744 97906 161800
rect 97962 161744 100188 161800
rect 97901 161742 100188 161744
rect 120796 161800 122899 161802
rect 120796 161744 122838 161800
rect 122894 161744 122899 161800
rect 128494 161772 128554 162284
rect 148366 161772 148426 162284
rect 154481 161802 154547 161805
rect 178033 161802 178099 161805
rect 154481 161800 156124 161802
rect 120796 161742 122899 161744
rect 97901 161739 97967 161742
rect 122833 161739 122899 161742
rect 154481 161744 154486 161800
rect 154542 161744 156124 161800
rect 154481 161742 156124 161744
rect 176916 161800 178099 161802
rect 176916 161744 178038 161800
rect 178094 161744 178099 161800
rect 176916 161742 178099 161744
rect 154481 161739 154547 161742
rect 178033 161739 178099 161742
rect 182081 161802 182147 161805
rect 207013 161802 207079 161805
rect 182081 161800 184092 161802
rect 182081 161744 182086 161800
rect 182142 161744 184092 161800
rect 182081 161742 184092 161744
rect 204884 161800 207079 161802
rect 204884 161744 207018 161800
rect 207074 161744 207079 161800
rect 204884 161742 207079 161744
rect 182081 161739 182147 161742
rect 207013 161739 207079 161742
rect 209681 161802 209747 161805
rect 234705 161802 234771 161805
rect 209681 161800 212060 161802
rect 209681 161744 209686 161800
rect 209742 161744 212060 161800
rect 209681 161742 212060 161744
rect 232852 161800 234771 161802
rect 232852 161744 234710 161800
rect 234766 161744 234771 161800
rect 232852 161742 234771 161744
rect 209681 161739 209747 161742
rect 234705 161739 234771 161742
rect 238661 161802 238727 161805
rect 262213 161802 262279 161805
rect 238661 161800 240212 161802
rect 238661 161744 238666 161800
rect 238722 161744 240212 161800
rect 238661 161742 240212 161744
rect 260820 161800 262279 161802
rect 260820 161744 262218 161800
rect 262274 161744 262279 161800
rect 260820 161742 262279 161744
rect 238661 161739 238727 161742
rect 262213 161739 262279 161742
rect 266261 161802 266327 161805
rect 291193 161802 291259 161805
rect 266261 161800 268180 161802
rect 266261 161744 266266 161800
rect 266322 161744 268180 161800
rect 266261 161742 268180 161744
rect 288788 161800 291259 161802
rect 288788 161744 291198 161800
rect 291254 161744 291259 161800
rect 288788 161742 291259 161744
rect 266261 161739 266327 161742
rect 291193 161739 291259 161742
rect 293861 161802 293927 161805
rect 318793 161802 318859 161805
rect 293861 161800 296148 161802
rect 293861 161744 293866 161800
rect 293922 161744 296148 161800
rect 293861 161742 296148 161744
rect 316940 161800 318859 161802
rect 316940 161744 318798 161800
rect 318854 161744 318859 161800
rect 316940 161742 318859 161744
rect 293861 161739 293927 161742
rect 318793 161739 318859 161742
rect 322841 161802 322907 161805
rect 322841 161800 324116 161802
rect 322841 161744 322846 161800
rect 322902 161744 324116 161800
rect 344326 161772 344386 162284
rect 350441 161802 350507 161805
rect 350441 161800 352084 161802
rect 322841 161742 324116 161744
rect 350441 161744 350446 161800
rect 350502 161744 352084 161800
rect 372294 161772 372354 162284
rect 378041 161802 378107 161805
rect 402973 161802 403039 161805
rect 378041 161800 380052 161802
rect 350441 161742 352084 161744
rect 378041 161744 378046 161800
rect 378102 161744 380052 161800
rect 378041 161742 380052 161744
rect 400844 161800 403039 161802
rect 400844 161744 402978 161800
rect 403034 161744 403039 161800
rect 408542 161772 408602 162284
rect 430573 161802 430639 161805
rect 428812 161800 430639 161802
rect 400844 161742 403039 161744
rect 428812 161744 430578 161800
rect 430634 161744 430639 161800
rect 428812 161742 430639 161744
rect 322841 161739 322907 161742
rect 350441 161739 350507 161742
rect 378041 161739 378107 161742
rect 402973 161739 403039 161742
rect 430573 161739 430639 161742
rect 434621 161802 434687 161805
rect 458173 161802 458239 161805
rect 434621 161800 436172 161802
rect 434621 161744 434626 161800
rect 434682 161744 436172 161800
rect 434621 161742 436172 161744
rect 456964 161800 458239 161802
rect 456964 161744 458178 161800
rect 458234 161744 458239 161800
rect 456964 161742 458239 161744
rect 434621 161739 434687 161742
rect 458173 161739 458239 161742
rect 462221 161802 462287 161805
rect 487153 161802 487219 161805
rect 462221 161800 464140 161802
rect 462221 161744 462226 161800
rect 462282 161744 464140 161800
rect 462221 161742 464140 161744
rect 484932 161800 487219 161802
rect 484932 161744 487158 161800
rect 487214 161744 487219 161800
rect 484932 161742 487219 161744
rect 462221 161739 462287 161742
rect 487153 161739 487219 161742
rect 489821 161802 489887 161805
rect 514753 161802 514819 161805
rect 489821 161800 492108 161802
rect 489821 161744 489826 161800
rect 489882 161744 492108 161800
rect 489821 161742 492108 161744
rect 512900 161800 514819 161802
rect 512900 161744 514758 161800
rect 514814 161744 514819 161800
rect 520598 161772 520658 162284
rect 540470 161772 540530 162284
rect 546401 161802 546467 161805
rect 571333 161802 571399 161805
rect 546401 161800 548044 161802
rect 512900 161742 514819 161744
rect 489821 161739 489887 161742
rect 514753 161739 514819 161742
rect 546401 161744 546406 161800
rect 546462 161744 548044 161800
rect 546401 161742 548044 161744
rect 568836 161800 571399 161802
rect 568836 161744 571338 161800
rect 571394 161744 571399 161800
rect 568836 161742 571399 161744
rect 546401 161739 546467 161742
rect 571333 161739 571399 161742
rect 580073 152690 580139 152693
rect 583520 152690 584960 152780
rect 580073 152688 584960 152690
rect 580073 152632 580078 152688
rect 580134 152632 584960 152688
rect 580073 152630 584960 152632
rect 580073 152627 580139 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 2773 149834 2839 149837
rect -960 149832 2839 149834
rect -960 149776 2778 149832
rect 2834 149776 2839 149832
rect -960 149774 2839 149776
rect -960 149684 480 149774
rect 2773 149771 2839 149774
rect 361614 144468 361620 144532
rect 361684 144530 361690 144532
rect 361941 144530 362007 144533
rect 361684 144528 362007 144530
rect 361684 144472 361946 144528
rect 362002 144472 362007 144528
rect 361684 144470 362007 144472
rect 361684 144468 361690 144470
rect 361941 144467 362007 144470
rect 445702 144468 445708 144532
rect 445772 144530 445778 144532
rect 446029 144530 446095 144533
rect 445772 144528 446095 144530
rect 445772 144472 446034 144528
rect 446090 144472 446095 144528
rect 445772 144470 446095 144472
rect 445772 144468 445778 144470
rect 446029 144467 446095 144470
rect 13537 142762 13603 142765
rect 66253 142762 66319 142765
rect 13537 142760 66319 142762
rect 13537 142704 13542 142760
rect 13598 142704 66258 142760
rect 66314 142704 66319 142760
rect 13537 142702 66319 142704
rect 13537 142699 13603 142702
rect 66253 142699 66319 142702
rect 70301 142762 70367 142765
rect 122833 142762 122899 142765
rect 70301 142760 122899 142762
rect 70301 142704 70306 142760
rect 70362 142704 122838 142760
rect 122894 142704 122899 142760
rect 70301 142702 122899 142704
rect 70301 142699 70367 142702
rect 122833 142699 122899 142702
rect 126881 142762 126947 142765
rect 178033 142762 178099 142765
rect 126881 142760 178099 142762
rect 126881 142704 126886 142760
rect 126942 142704 178038 142760
rect 178094 142704 178099 142760
rect 126881 142702 178099 142704
rect 126881 142699 126947 142702
rect 178033 142699 178099 142702
rect 209681 142762 209747 142765
rect 262213 142762 262279 142765
rect 209681 142760 262279 142762
rect 209681 142704 209686 142760
rect 209742 142704 262218 142760
rect 262274 142704 262279 142760
rect 209681 142702 262279 142704
rect 209681 142699 209747 142702
rect 262213 142699 262279 142702
rect 266261 142762 266327 142765
rect 318793 142762 318859 142765
rect 266261 142760 318859 142762
rect 266261 142704 266266 142760
rect 266322 142704 318798 142760
rect 318854 142704 318859 142760
rect 266261 142702 318859 142704
rect 266261 142699 266327 142702
rect 318793 142699 318859 142702
rect 322841 142762 322907 142765
rect 375373 142762 375439 142765
rect 322841 142760 375439 142762
rect 322841 142704 322846 142760
rect 322902 142704 375378 142760
rect 375434 142704 375439 142760
rect 322841 142702 375439 142704
rect 322841 142699 322907 142702
rect 375373 142699 375439 142702
rect 378041 142762 378107 142765
rect 430573 142762 430639 142765
rect 378041 142760 430639 142762
rect 378041 142704 378046 142760
rect 378102 142704 430578 142760
rect 430634 142704 430639 142760
rect 378041 142702 430639 142704
rect 378041 142699 378107 142702
rect 430573 142699 430639 142702
rect 434621 142762 434687 142765
rect 487153 142762 487219 142765
rect 434621 142760 487219 142762
rect 434621 142704 434626 142760
rect 434682 142704 487158 142760
rect 487214 142704 487219 142760
rect 434621 142702 487219 142704
rect 434621 142699 434687 142702
rect 487153 142699 487219 142702
rect 489821 142762 489887 142765
rect 542353 142762 542419 142765
rect 489821 142760 542419 142762
rect 489821 142704 489826 142760
rect 489882 142704 542358 142760
rect 542414 142704 542419 142760
rect 489821 142702 542419 142704
rect 489821 142699 489887 142702
rect 542353 142699 542419 142702
rect 583520 139212 584960 139452
rect -960 136778 480 136868
rect 3325 136778 3391 136781
rect -960 136776 3391 136778
rect -960 136720 3330 136776
rect 3386 136720 3391 136776
rect -960 136718 3391 136720
rect -960 136628 480 136718
rect 3325 136715 3391 136718
rect 13537 134330 13603 134333
rect 38653 134330 38719 134333
rect 13537 134328 16100 134330
rect 13537 134272 13542 134328
rect 13598 134272 16100 134328
rect 13537 134270 16100 134272
rect 36892 134328 38719 134330
rect 36892 134272 38658 134328
rect 38714 134272 38719 134328
rect 36892 134270 38719 134272
rect 13537 134267 13603 134270
rect 38653 134267 38719 134270
rect 42701 134330 42767 134333
rect 66253 134330 66319 134333
rect 42701 134328 44068 134330
rect 42701 134272 42706 134328
rect 42762 134272 44068 134328
rect 42701 134270 44068 134272
rect 64860 134328 66319 134330
rect 64860 134272 66258 134328
rect 66314 134272 66319 134328
rect 64860 134270 66319 134272
rect 42701 134267 42767 134270
rect 66253 134267 66319 134270
rect 70301 134330 70367 134333
rect 95233 134330 95299 134333
rect 70301 134328 72036 134330
rect 70301 134272 70306 134328
rect 70362 134272 72036 134328
rect 70301 134270 72036 134272
rect 92828 134328 95299 134330
rect 92828 134272 95238 134328
rect 95294 134272 95299 134328
rect 92828 134270 95299 134272
rect 70301 134267 70367 134270
rect 95233 134267 95299 134270
rect 97901 134330 97967 134333
rect 122833 134330 122899 134333
rect 97901 134328 100188 134330
rect 97901 134272 97906 134328
rect 97962 134272 100188 134328
rect 97901 134270 100188 134272
rect 120796 134328 122899 134330
rect 120796 134272 122838 134328
rect 122894 134272 122899 134328
rect 120796 134270 122899 134272
rect 97901 134267 97967 134270
rect 122833 134267 122899 134270
rect 126881 134330 126947 134333
rect 150433 134330 150499 134333
rect 126881 134328 128156 134330
rect 126881 134272 126886 134328
rect 126942 134272 128156 134328
rect 126881 134270 128156 134272
rect 148948 134328 150499 134330
rect 148948 134272 150438 134328
rect 150494 134272 150499 134328
rect 148948 134270 150499 134272
rect 126881 134267 126947 134270
rect 150433 134267 150499 134270
rect 154481 134330 154547 134333
rect 178033 134330 178099 134333
rect 154481 134328 156124 134330
rect 154481 134272 154486 134328
rect 154542 134272 156124 134328
rect 154481 134270 156124 134272
rect 176916 134328 178099 134330
rect 176916 134272 178038 134328
rect 178094 134272 178099 134328
rect 176916 134270 178099 134272
rect 154481 134267 154547 134270
rect 178033 134267 178099 134270
rect 182081 134330 182147 134333
rect 207013 134330 207079 134333
rect 182081 134328 184092 134330
rect 182081 134272 182086 134328
rect 182142 134272 184092 134328
rect 182081 134270 184092 134272
rect 204884 134328 207079 134330
rect 204884 134272 207018 134328
rect 207074 134272 207079 134328
rect 204884 134270 207079 134272
rect 182081 134267 182147 134270
rect 207013 134267 207079 134270
rect 209681 134330 209747 134333
rect 234705 134330 234771 134333
rect 209681 134328 212060 134330
rect 209681 134272 209686 134328
rect 209742 134272 212060 134328
rect 209681 134270 212060 134272
rect 232852 134328 234771 134330
rect 232852 134272 234710 134328
rect 234766 134272 234771 134328
rect 232852 134270 234771 134272
rect 209681 134267 209747 134270
rect 234705 134267 234771 134270
rect 238661 134330 238727 134333
rect 262213 134330 262279 134333
rect 238661 134328 240212 134330
rect 238661 134272 238666 134328
rect 238722 134272 240212 134328
rect 238661 134270 240212 134272
rect 260820 134328 262279 134330
rect 260820 134272 262218 134328
rect 262274 134272 262279 134328
rect 260820 134270 262279 134272
rect 238661 134267 238727 134270
rect 262213 134267 262279 134270
rect 266261 134330 266327 134333
rect 291193 134330 291259 134333
rect 266261 134328 268180 134330
rect 266261 134272 266266 134328
rect 266322 134272 268180 134328
rect 266261 134270 268180 134272
rect 288788 134328 291259 134330
rect 288788 134272 291198 134328
rect 291254 134272 291259 134328
rect 288788 134270 291259 134272
rect 266261 134267 266327 134270
rect 291193 134267 291259 134270
rect 293861 134330 293927 134333
rect 318793 134330 318859 134333
rect 293861 134328 296148 134330
rect 293861 134272 293866 134328
rect 293922 134272 296148 134328
rect 293861 134270 296148 134272
rect 316940 134328 318859 134330
rect 316940 134272 318798 134328
rect 318854 134272 318859 134328
rect 316940 134270 318859 134272
rect 293861 134267 293927 134270
rect 318793 134267 318859 134270
rect 322841 134330 322907 134333
rect 346393 134330 346459 134333
rect 322841 134328 324116 134330
rect 322841 134272 322846 134328
rect 322902 134272 324116 134328
rect 322841 134270 324116 134272
rect 344908 134328 346459 134330
rect 344908 134272 346398 134328
rect 346454 134272 346459 134328
rect 344908 134270 346459 134272
rect 322841 134267 322907 134270
rect 346393 134267 346459 134270
rect 350441 134330 350507 134333
rect 375373 134330 375439 134333
rect 350441 134328 352084 134330
rect 350441 134272 350446 134328
rect 350502 134272 352084 134328
rect 350441 134270 352084 134272
rect 372876 134328 375439 134330
rect 372876 134272 375378 134328
rect 375434 134272 375439 134328
rect 372876 134270 375439 134272
rect 350441 134267 350507 134270
rect 375373 134267 375439 134270
rect 378041 134330 378107 134333
rect 402973 134330 403039 134333
rect 378041 134328 380052 134330
rect 378041 134272 378046 134328
rect 378102 134272 380052 134328
rect 378041 134270 380052 134272
rect 400844 134328 403039 134330
rect 400844 134272 402978 134328
rect 403034 134272 403039 134328
rect 400844 134270 403039 134272
rect 378041 134267 378107 134270
rect 402973 134267 403039 134270
rect 405641 134330 405707 134333
rect 430573 134330 430639 134333
rect 405641 134328 408204 134330
rect 405641 134272 405646 134328
rect 405702 134272 408204 134328
rect 405641 134270 408204 134272
rect 428812 134328 430639 134330
rect 428812 134272 430578 134328
rect 430634 134272 430639 134328
rect 428812 134270 430639 134272
rect 405641 134267 405707 134270
rect 430573 134267 430639 134270
rect 434621 134330 434687 134333
rect 458173 134330 458239 134333
rect 434621 134328 436172 134330
rect 434621 134272 434626 134328
rect 434682 134272 436172 134328
rect 434621 134270 436172 134272
rect 456964 134328 458239 134330
rect 456964 134272 458178 134328
rect 458234 134272 458239 134328
rect 456964 134270 458239 134272
rect 434621 134267 434687 134270
rect 458173 134267 458239 134270
rect 462221 134330 462287 134333
rect 487153 134330 487219 134333
rect 462221 134328 464140 134330
rect 462221 134272 462226 134328
rect 462282 134272 464140 134328
rect 462221 134270 464140 134272
rect 484932 134328 487219 134330
rect 484932 134272 487158 134328
rect 487214 134272 487219 134328
rect 484932 134270 487219 134272
rect 462221 134267 462287 134270
rect 487153 134267 487219 134270
rect 489821 134330 489887 134333
rect 514753 134330 514819 134333
rect 489821 134328 492108 134330
rect 489821 134272 489826 134328
rect 489882 134272 492108 134328
rect 489821 134270 492108 134272
rect 512900 134328 514819 134330
rect 512900 134272 514758 134328
rect 514814 134272 514819 134328
rect 512900 134270 514819 134272
rect 489821 134267 489887 134270
rect 514753 134267 514819 134270
rect 518801 134330 518867 134333
rect 542353 134330 542419 134333
rect 518801 134328 520076 134330
rect 518801 134272 518806 134328
rect 518862 134272 520076 134328
rect 518801 134270 520076 134272
rect 540868 134328 542419 134330
rect 540868 134272 542358 134328
rect 542414 134272 542419 134328
rect 540868 134270 542419 134272
rect 518801 134267 518867 134270
rect 542353 134267 542419 134270
rect 546401 134330 546467 134333
rect 571333 134330 571399 134333
rect 546401 134328 548044 134330
rect 546401 134272 546406 134328
rect 546462 134272 548044 134328
rect 546401 134270 548044 134272
rect 568836 134328 571399 134330
rect 568836 134272 571338 134328
rect 571394 134272 571399 134328
rect 568836 134270 571399 134272
rect 546401 134267 546467 134270
rect 571333 134267 571399 134270
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 344645 122770 344711 122773
rect 361614 122770 361620 122772
rect 344645 122768 361620 122770
rect 344645 122712 344650 122768
rect 344706 122712 361620 122768
rect 344645 122710 361620 122712
rect 344645 122707 344711 122710
rect 361614 122708 361620 122710
rect 361684 122708 361690 122772
rect 428641 122770 428707 122773
rect 445702 122770 445708 122772
rect 428641 122768 445708 122770
rect 428641 122712 428646 122768
rect 428702 122712 445708 122768
rect 428641 122710 445708 122712
rect 428641 122707 428707 122710
rect 445702 122708 445708 122710
rect 445772 122708 445778 122772
rect 194777 117332 194843 117333
rect 194726 117330 194732 117332
rect 194686 117270 194732 117330
rect 194796 117328 194843 117332
rect 194838 117272 194843 117328
rect 194726 117268 194732 117270
rect 194796 117268 194843 117272
rect 194777 117267 194843 117268
rect 324221 117332 324287 117333
rect 324221 117328 324268 117332
rect 324332 117330 324338 117332
rect 324221 117272 324226 117328
rect 324221 117268 324268 117272
rect 324332 117270 324378 117330
rect 324332 117268 324338 117270
rect 324221 117267 324287 117268
rect 209681 116514 209747 116517
rect 260414 116514 260420 116516
rect 209681 116512 260420 116514
rect 209681 116456 209686 116512
rect 209742 116456 260420 116512
rect 209681 116454 260420 116456
rect 209681 116451 209747 116454
rect 260414 116452 260420 116454
rect 260484 116452 260490 116516
rect 126881 116378 126947 116381
rect 176326 116378 176332 116380
rect 126881 116376 176332 116378
rect 126881 116320 126886 116376
rect 126942 116320 176332 116376
rect 126881 116318 176332 116320
rect 126881 116315 126947 116318
rect 176326 116316 176332 116318
rect 176396 116316 176402 116380
rect 182081 116378 182147 116381
rect 234705 116378 234771 116381
rect 182081 116376 234771 116378
rect 182081 116320 182086 116376
rect 182142 116320 234710 116376
rect 234766 116320 234771 116376
rect 182081 116318 234771 116320
rect 182081 116315 182147 116318
rect 234705 116315 234771 116318
rect 42701 116242 42767 116245
rect 92422 116242 92428 116244
rect 42701 116240 92428 116242
rect 42701 116184 42706 116240
rect 42762 116184 92428 116240
rect 42701 116182 92428 116184
rect 42701 116179 42767 116182
rect 92422 116180 92428 116182
rect 92492 116180 92498 116244
rect 97901 116242 97967 116245
rect 148358 116242 148364 116244
rect 97901 116240 148364 116242
rect 97901 116184 97906 116240
rect 97962 116184 148364 116240
rect 97901 116182 148364 116184
rect 97901 116179 97967 116182
rect 148358 116180 148364 116182
rect 148428 116180 148434 116244
rect 378041 116242 378107 116245
rect 430573 116242 430639 116245
rect 378041 116240 430639 116242
rect 378041 116184 378046 116240
rect 378102 116184 430578 116240
rect 430634 116184 430639 116240
rect 378041 116182 430639 116184
rect 378041 116179 378107 116182
rect 430573 116179 430639 116182
rect 489821 116242 489887 116245
rect 540462 116242 540468 116244
rect 489821 116240 540468 116242
rect 489821 116184 489826 116240
rect 489882 116184 540468 116240
rect 489821 116182 540468 116184
rect 489821 116179 489887 116182
rect 540462 116180 540468 116182
rect 540532 116180 540538 116244
rect 13537 116106 13603 116109
rect 64454 116106 64460 116108
rect 13537 116104 64460 116106
rect 13537 116048 13542 116104
rect 13598 116048 64460 116104
rect 13537 116046 64460 116048
rect 13537 116043 13603 116046
rect 64454 116044 64460 116046
rect 64524 116044 64530 116108
rect 70301 116106 70367 116109
rect 122833 116106 122899 116109
rect 70301 116104 122899 116106
rect 70301 116048 70306 116104
rect 70362 116048 122838 116104
rect 122894 116048 122899 116104
rect 70301 116046 122899 116048
rect 70301 116043 70367 116046
rect 122833 116043 122899 116046
rect 154481 116106 154547 116109
rect 207013 116106 207079 116109
rect 154481 116104 207079 116106
rect 154481 116048 154486 116104
rect 154542 116048 207018 116104
rect 207074 116048 207079 116104
rect 154481 116046 207079 116048
rect 154481 116043 154547 116046
rect 207013 116043 207079 116046
rect 266261 116106 266327 116109
rect 318793 116106 318859 116109
rect 266261 116104 318859 116106
rect 266261 116048 266266 116104
rect 266322 116048 318798 116104
rect 318854 116048 318859 116104
rect 266261 116046 318859 116048
rect 266261 116043 266327 116046
rect 318793 116043 318859 116046
rect 350441 116106 350507 116109
rect 402973 116106 403039 116109
rect 350441 116104 403039 116106
rect 350441 116048 350446 116104
rect 350502 116048 402978 116104
rect 403034 116048 403039 116104
rect 350441 116046 403039 116048
rect 350441 116043 350507 116046
rect 402973 116043 403039 116046
rect 408534 116044 408540 116108
rect 408604 116106 408610 116108
rect 458173 116106 458239 116109
rect 408604 116104 458239 116106
rect 408604 116048 458178 116104
rect 458234 116048 458239 116104
rect 408604 116046 458239 116048
rect 408604 116044 408610 116046
rect 458173 116043 458239 116046
rect 462221 116106 462287 116109
rect 514753 116106 514819 116109
rect 462221 116104 514819 116106
rect 462221 116048 462226 116104
rect 462282 116048 514758 116104
rect 514814 116048 514819 116104
rect 462221 116046 514819 116048
rect 462221 116043 462287 116046
rect 514753 116043 514819 116046
rect 520590 116044 520596 116108
rect 520660 116106 520666 116108
rect 571333 116106 571399 116109
rect 520660 116104 571399 116106
rect 520660 116048 571338 116104
rect 571394 116048 571399 116104
rect 520660 116046 571399 116048
rect 520660 116044 520666 116046
rect 571333 116043 571399 116046
rect 580073 112842 580139 112845
rect 583520 112842 584960 112932
rect 580073 112840 584960 112842
rect 580073 112784 580078 112840
rect 580134 112784 584960 112840
rect 580073 112782 584960 112784
rect 580073 112779 580139 112782
rect 583520 112692 584960 112782
rect -960 110516 480 110756
rect 64454 108292 64460 108356
rect 64524 108292 64530 108356
rect 70301 108354 70367 108357
rect 70301 108352 72066 108354
rect 70301 108296 70306 108352
rect 70362 108296 72066 108352
rect 70301 108294 72066 108296
rect 13537 107810 13603 107813
rect 38653 107810 38719 107813
rect 13537 107808 16100 107810
rect 13537 107752 13542 107808
rect 13598 107752 16100 107808
rect 13537 107750 16100 107752
rect 36892 107808 38719 107810
rect 36892 107752 38658 107808
rect 38714 107752 38719 107808
rect 36892 107750 38719 107752
rect 13537 107747 13603 107750
rect 38653 107747 38719 107750
rect 42701 107810 42767 107813
rect 42701 107808 44068 107810
rect 42701 107752 42706 107808
rect 42762 107752 44068 107808
rect 64462 107780 64522 108292
rect 70301 108291 70367 108294
rect 72006 107780 72066 108294
rect 92422 108292 92428 108356
rect 92492 108292 92498 108356
rect 148358 108292 148364 108356
rect 148428 108292 148434 108356
rect 176326 108292 176332 108356
rect 176396 108292 176402 108356
rect 260414 108292 260420 108356
rect 260484 108292 260490 108356
rect 408534 108292 408540 108356
rect 408604 108292 408610 108356
rect 458173 108354 458239 108357
rect 456934 108352 458239 108354
rect 456934 108296 458178 108352
rect 458234 108296 458239 108352
rect 456934 108294 458239 108296
rect 92430 107780 92490 108292
rect 97901 107810 97967 107813
rect 122833 107810 122899 107813
rect 97901 107808 100188 107810
rect 42701 107750 44068 107752
rect 97901 107752 97906 107808
rect 97962 107752 100188 107808
rect 97901 107750 100188 107752
rect 120796 107808 122899 107810
rect 120796 107752 122838 107808
rect 122894 107752 122899 107808
rect 120796 107750 122899 107752
rect 42701 107747 42767 107750
rect 97901 107747 97967 107750
rect 122833 107747 122899 107750
rect 126881 107810 126947 107813
rect 126881 107808 128156 107810
rect 126881 107752 126886 107808
rect 126942 107752 128156 107808
rect 148366 107780 148426 108292
rect 154481 107810 154547 107813
rect 154481 107808 156124 107810
rect 126881 107750 128156 107752
rect 154481 107752 154486 107808
rect 154542 107752 156124 107808
rect 176334 107780 176394 108292
rect 182081 107810 182147 107813
rect 207013 107810 207079 107813
rect 182081 107808 184092 107810
rect 154481 107750 156124 107752
rect 182081 107752 182086 107808
rect 182142 107752 184092 107808
rect 182081 107750 184092 107752
rect 204884 107808 207079 107810
rect 204884 107752 207018 107808
rect 207074 107752 207079 107808
rect 204884 107750 207079 107752
rect 126881 107747 126947 107750
rect 154481 107747 154547 107750
rect 182081 107747 182147 107750
rect 207013 107747 207079 107750
rect 209681 107810 209747 107813
rect 234705 107810 234771 107813
rect 209681 107808 212060 107810
rect 209681 107752 209686 107808
rect 209742 107752 212060 107808
rect 209681 107750 212060 107752
rect 232852 107808 234771 107810
rect 232852 107752 234710 107808
rect 234766 107752 234771 107808
rect 232852 107750 234771 107752
rect 209681 107747 209747 107750
rect 234705 107747 234771 107750
rect 238661 107810 238727 107813
rect 238661 107808 240212 107810
rect 238661 107752 238666 107808
rect 238722 107752 240212 107808
rect 260422 107780 260482 108292
rect 266261 107810 266327 107813
rect 291193 107810 291259 107813
rect 266261 107808 268180 107810
rect 238661 107750 240212 107752
rect 266261 107752 266266 107808
rect 266322 107752 268180 107808
rect 266261 107750 268180 107752
rect 288788 107808 291259 107810
rect 288788 107752 291198 107808
rect 291254 107752 291259 107808
rect 288788 107750 291259 107752
rect 238661 107747 238727 107750
rect 266261 107747 266327 107750
rect 291193 107747 291259 107750
rect 293861 107810 293927 107813
rect 318793 107810 318859 107813
rect 293861 107808 296148 107810
rect 293861 107752 293866 107808
rect 293922 107752 296148 107808
rect 293861 107750 296148 107752
rect 316940 107808 318859 107810
rect 316940 107752 318798 107808
rect 318854 107752 318859 107808
rect 316940 107750 318859 107752
rect 293861 107747 293927 107750
rect 318793 107747 318859 107750
rect 322841 107810 322907 107813
rect 346393 107810 346459 107813
rect 322841 107808 324116 107810
rect 322841 107752 322846 107808
rect 322902 107752 324116 107808
rect 322841 107750 324116 107752
rect 344908 107808 346459 107810
rect 344908 107752 346398 107808
rect 346454 107752 346459 107808
rect 344908 107750 346459 107752
rect 322841 107747 322907 107750
rect 346393 107747 346459 107750
rect 350441 107810 350507 107813
rect 375373 107810 375439 107813
rect 350441 107808 352084 107810
rect 350441 107752 350446 107808
rect 350502 107752 352084 107808
rect 350441 107750 352084 107752
rect 372876 107808 375439 107810
rect 372876 107752 375378 107808
rect 375434 107752 375439 107808
rect 372876 107750 375439 107752
rect 350441 107747 350507 107750
rect 375373 107747 375439 107750
rect 378041 107810 378107 107813
rect 402973 107810 403039 107813
rect 378041 107808 380052 107810
rect 378041 107752 378046 107808
rect 378102 107752 380052 107808
rect 378041 107750 380052 107752
rect 400844 107808 403039 107810
rect 400844 107752 402978 107808
rect 403034 107752 403039 107808
rect 408542 107780 408602 108292
rect 430573 107810 430639 107813
rect 428812 107808 430639 107810
rect 400844 107750 403039 107752
rect 428812 107752 430578 107808
rect 430634 107752 430639 107808
rect 428812 107750 430639 107752
rect 378041 107747 378107 107750
rect 402973 107747 403039 107750
rect 430573 107747 430639 107750
rect 434621 107810 434687 107813
rect 434621 107808 436172 107810
rect 434621 107752 434626 107808
rect 434682 107752 436172 107808
rect 456934 107780 456994 108294
rect 458173 108291 458239 108294
rect 520590 108292 520596 108356
rect 520660 108292 520666 108356
rect 540462 108292 540468 108356
rect 540532 108292 540538 108356
rect 462221 107810 462287 107813
rect 487153 107810 487219 107813
rect 462221 107808 464140 107810
rect 434621 107750 436172 107752
rect 462221 107752 462226 107808
rect 462282 107752 464140 107808
rect 462221 107750 464140 107752
rect 484932 107808 487219 107810
rect 484932 107752 487158 107808
rect 487214 107752 487219 107808
rect 484932 107750 487219 107752
rect 434621 107747 434687 107750
rect 462221 107747 462287 107750
rect 487153 107747 487219 107750
rect 489821 107810 489887 107813
rect 514753 107810 514819 107813
rect 489821 107808 492108 107810
rect 489821 107752 489826 107808
rect 489882 107752 492108 107808
rect 489821 107750 492108 107752
rect 512900 107808 514819 107810
rect 512900 107752 514758 107808
rect 514814 107752 514819 107808
rect 520598 107780 520658 108292
rect 540470 107780 540530 108292
rect 546401 107810 546467 107813
rect 571333 107810 571399 107813
rect 546401 107808 548044 107810
rect 512900 107750 514819 107752
rect 489821 107747 489887 107750
rect 514753 107747 514819 107750
rect 546401 107752 546406 107808
rect 546462 107752 548044 107808
rect 546401 107750 548044 107752
rect 568836 107808 571399 107810
rect 568836 107752 571338 107808
rect 571394 107752 571399 107808
rect 568836 107750 571399 107752
rect 546401 107747 546467 107750
rect 571333 107747 571399 107750
rect 583520 99364 584960 99604
rect -960 97610 480 97700
rect 4061 97610 4127 97613
rect -960 97608 4127 97610
rect -960 97552 4066 97608
rect 4122 97552 4127 97608
rect -960 97550 4127 97552
rect -960 97460 480 97550
rect 4061 97547 4127 97550
rect 156321 95162 156387 95165
rect 194726 95162 194732 95164
rect 156321 95160 194732 95162
rect 156321 95104 156326 95160
rect 156382 95104 194732 95160
rect 156321 95102 194732 95104
rect 156321 95099 156387 95102
rect 194726 95100 194732 95102
rect 194796 95100 194802 95164
rect 306925 95162 306991 95165
rect 324262 95162 324268 95164
rect 306925 95160 324268 95162
rect 306925 95104 306930 95160
rect 306986 95104 324268 95160
rect 306925 95102 324268 95104
rect 306925 95099 306991 95102
rect 324262 95100 324268 95102
rect 324332 95100 324338 95164
rect 322841 89042 322907 89045
rect 372286 89042 372292 89044
rect 322841 89040 372292 89042
rect 322841 88984 322846 89040
rect 322902 88984 372292 89040
rect 322841 88982 372292 88984
rect 322841 88979 322907 88982
rect 372286 88980 372292 88982
rect 372356 88980 372362 89044
rect 44582 88844 44588 88908
rect 44652 88906 44658 88908
rect 95233 88906 95299 88909
rect 44652 88904 95299 88906
rect 44652 88848 95238 88904
rect 95294 88848 95299 88904
rect 44652 88846 95299 88848
rect 44652 88844 44658 88846
rect 95233 88843 95299 88846
rect 97901 88906 97967 88909
rect 150433 88906 150499 88909
rect 97901 88904 150499 88906
rect 97901 88848 97906 88904
rect 97962 88848 150438 88904
rect 150494 88848 150499 88904
rect 97901 88846 150499 88848
rect 97901 88843 97967 88846
rect 150433 88843 150499 88846
rect 154481 88906 154547 88909
rect 207013 88906 207079 88909
rect 154481 88904 207079 88906
rect 154481 88848 154486 88904
rect 154542 88848 207018 88904
rect 207074 88848 207079 88904
rect 154481 88846 207079 88848
rect 154481 88843 154547 88846
rect 207013 88843 207079 88846
rect 238661 88906 238727 88909
rect 288382 88906 288388 88908
rect 238661 88904 288388 88906
rect 238661 88848 238666 88904
rect 238722 88848 288388 88904
rect 238661 88846 288388 88848
rect 238661 88843 238727 88846
rect 288382 88844 288388 88846
rect 288452 88844 288458 88908
rect 296846 88844 296852 88908
rect 296916 88906 296922 88908
rect 346393 88906 346459 88909
rect 296916 88904 346459 88906
rect 296916 88848 346398 88904
rect 346454 88848 346459 88904
rect 296916 88846 346459 88848
rect 296916 88844 296922 88846
rect 346393 88843 346459 88846
rect 378041 88906 378107 88909
rect 430573 88906 430639 88909
rect 378041 88904 430639 88906
rect 378041 88848 378046 88904
rect 378102 88848 430578 88904
rect 430634 88848 430639 88904
rect 378041 88846 430639 88848
rect 378041 88843 378107 88846
rect 430573 88843 430639 88846
rect 434621 88906 434687 88909
rect 484342 88906 484348 88908
rect 434621 88904 484348 88906
rect 434621 88848 434626 88904
rect 434682 88848 484348 88904
rect 434621 88846 484348 88848
rect 434621 88843 434687 88846
rect 484342 88844 484348 88846
rect 484412 88844 484418 88908
rect 13537 88770 13603 88773
rect 66253 88770 66319 88773
rect 13537 88768 66319 88770
rect 13537 88712 13542 88768
rect 13598 88712 66258 88768
rect 66314 88712 66319 88768
rect 13537 88710 66319 88712
rect 13537 88707 13603 88710
rect 66253 88707 66319 88710
rect 70301 88770 70367 88773
rect 122833 88770 122899 88773
rect 70301 88768 122899 88770
rect 70301 88712 70306 88768
rect 70362 88712 122838 88768
rect 122894 88712 122899 88768
rect 70301 88710 122899 88712
rect 70301 88707 70367 88710
rect 122833 88707 122899 88710
rect 126881 88770 126947 88773
rect 176326 88770 176332 88772
rect 126881 88768 176332 88770
rect 126881 88712 126886 88768
rect 126942 88712 176332 88768
rect 126881 88710 176332 88712
rect 126881 88707 126947 88710
rect 176326 88708 176332 88710
rect 176396 88708 176402 88772
rect 182081 88770 182147 88773
rect 234705 88770 234771 88773
rect 182081 88768 234771 88770
rect 182081 88712 182086 88768
rect 182142 88712 234710 88768
rect 234766 88712 234771 88768
rect 182081 88710 234771 88712
rect 182081 88707 182147 88710
rect 234705 88707 234771 88710
rect 266261 88770 266327 88773
rect 318793 88770 318859 88773
rect 266261 88768 318859 88770
rect 266261 88712 266266 88768
rect 266322 88712 318798 88768
rect 318854 88712 318859 88768
rect 266261 88710 318859 88712
rect 266261 88707 266327 88710
rect 318793 88707 318859 88710
rect 350441 88770 350507 88773
rect 402973 88770 403039 88773
rect 350441 88768 403039 88770
rect 350441 88712 350446 88768
rect 350502 88712 402978 88768
rect 403034 88712 403039 88768
rect 350441 88710 403039 88712
rect 350441 88707 350507 88710
rect 402973 88707 403039 88710
rect 462221 88770 462287 88773
rect 514753 88770 514819 88773
rect 462221 88768 514819 88770
rect 462221 88712 462226 88768
rect 462282 88712 514758 88768
rect 514814 88712 514819 88768
rect 462221 88710 514819 88712
rect 462221 88707 462287 88710
rect 514753 88707 514819 88710
rect 520590 88708 520596 88772
rect 520660 88770 520666 88772
rect 571333 88770 571399 88773
rect 520660 88768 571399 88770
rect 520660 88712 571338 88768
rect 571394 88712 571399 88768
rect 520660 88710 571399 88712
rect 520660 88708 520666 88710
rect 571333 88707 571399 88710
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 44582 80820 44588 80884
rect 44652 80820 44658 80884
rect 176326 80820 176332 80884
rect 176396 80820 176402 80884
rect 288382 80820 288388 80884
rect 288452 80820 288458 80884
rect 296478 80820 296484 80884
rect 296548 80820 296554 80884
rect 372286 80820 372292 80884
rect 372356 80820 372362 80884
rect 484342 80820 484348 80884
rect 484412 80820 484418 80884
rect 520590 80820 520596 80884
rect 520660 80820 520666 80884
rect 13537 80338 13603 80341
rect 38653 80338 38719 80341
rect 13537 80336 16100 80338
rect 13537 80280 13542 80336
rect 13598 80280 16100 80336
rect 13537 80278 16100 80280
rect 36892 80336 38719 80338
rect 36892 80280 38658 80336
rect 38714 80280 38719 80336
rect 44590 80308 44650 80820
rect 66253 80338 66319 80341
rect 64860 80336 66319 80338
rect 36892 80278 38719 80280
rect 64860 80280 66258 80336
rect 66314 80280 66319 80336
rect 64860 80278 66319 80280
rect 13537 80275 13603 80278
rect 38653 80275 38719 80278
rect 66253 80275 66319 80278
rect 70301 80338 70367 80341
rect 95233 80338 95299 80341
rect 70301 80336 72036 80338
rect 70301 80280 70306 80336
rect 70362 80280 72036 80336
rect 70301 80278 72036 80280
rect 92828 80336 95299 80338
rect 92828 80280 95238 80336
rect 95294 80280 95299 80336
rect 92828 80278 95299 80280
rect 70301 80275 70367 80278
rect 95233 80275 95299 80278
rect 97901 80338 97967 80341
rect 122833 80338 122899 80341
rect 97901 80336 100188 80338
rect 97901 80280 97906 80336
rect 97962 80280 100188 80336
rect 97901 80278 100188 80280
rect 120796 80336 122899 80338
rect 120796 80280 122838 80336
rect 122894 80280 122899 80336
rect 120796 80278 122899 80280
rect 97901 80275 97967 80278
rect 122833 80275 122899 80278
rect 126881 80338 126947 80341
rect 150433 80338 150499 80341
rect 126881 80336 128156 80338
rect 126881 80280 126886 80336
rect 126942 80280 128156 80336
rect 126881 80278 128156 80280
rect 148948 80336 150499 80338
rect 148948 80280 150438 80336
rect 150494 80280 150499 80336
rect 148948 80278 150499 80280
rect 126881 80275 126947 80278
rect 150433 80275 150499 80278
rect 154481 80338 154547 80341
rect 154481 80336 156124 80338
rect 154481 80280 154486 80336
rect 154542 80280 156124 80336
rect 176334 80308 176394 80820
rect 182081 80338 182147 80341
rect 207013 80338 207079 80341
rect 182081 80336 184092 80338
rect 154481 80278 156124 80280
rect 182081 80280 182086 80336
rect 182142 80280 184092 80336
rect 182081 80278 184092 80280
rect 204884 80336 207079 80338
rect 204884 80280 207018 80336
rect 207074 80280 207079 80336
rect 204884 80278 207079 80280
rect 154481 80275 154547 80278
rect 182081 80275 182147 80278
rect 207013 80275 207079 80278
rect 209681 80338 209747 80341
rect 234705 80338 234771 80341
rect 209681 80336 212060 80338
rect 209681 80280 209686 80336
rect 209742 80280 212060 80336
rect 209681 80278 212060 80280
rect 232852 80336 234771 80338
rect 232852 80280 234710 80336
rect 234766 80280 234771 80336
rect 232852 80278 234771 80280
rect 209681 80275 209747 80278
rect 234705 80275 234771 80278
rect 238661 80338 238727 80341
rect 262213 80338 262279 80341
rect 238661 80336 239690 80338
rect 238661 80280 238666 80336
rect 238722 80280 239690 80336
rect 238661 80278 239690 80280
rect 260820 80336 262279 80338
rect 260820 80280 262218 80336
rect 262274 80280 262279 80336
rect 260820 80278 262279 80280
rect 238661 80275 238727 80278
rect 239630 80270 239690 80278
rect 262213 80275 262279 80278
rect 266261 80338 266327 80341
rect 266261 80336 268180 80338
rect 266261 80280 266266 80336
rect 266322 80280 268180 80336
rect 288390 80308 288450 80820
rect 296486 80308 296546 80820
rect 318793 80338 318859 80341
rect 316940 80336 318859 80338
rect 266261 80278 268180 80280
rect 316940 80280 318798 80336
rect 318854 80280 318859 80336
rect 316940 80278 318859 80280
rect 266261 80275 266327 80278
rect 318793 80275 318859 80278
rect 322841 80338 322907 80341
rect 346393 80338 346459 80341
rect 322841 80336 324116 80338
rect 322841 80280 322846 80336
rect 322902 80280 324116 80336
rect 322841 80278 324116 80280
rect 344908 80336 346459 80338
rect 344908 80280 346398 80336
rect 346454 80280 346459 80336
rect 344908 80278 346459 80280
rect 322841 80275 322907 80278
rect 346393 80275 346459 80278
rect 350441 80338 350507 80341
rect 350441 80336 352084 80338
rect 350441 80280 350446 80336
rect 350502 80280 352084 80336
rect 372294 80308 372354 80820
rect 378041 80338 378107 80341
rect 402973 80338 403039 80341
rect 378041 80336 380052 80338
rect 350441 80278 352084 80280
rect 378041 80280 378046 80336
rect 378102 80280 380052 80336
rect 378041 80278 380052 80280
rect 400844 80336 403039 80338
rect 400844 80280 402978 80336
rect 403034 80280 403039 80336
rect 400844 80278 403039 80280
rect 350441 80275 350507 80278
rect 378041 80275 378107 80278
rect 402973 80275 403039 80278
rect 405641 80338 405707 80341
rect 430573 80338 430639 80341
rect 405641 80336 408204 80338
rect 405641 80280 405646 80336
rect 405702 80280 408204 80336
rect 405641 80278 408204 80280
rect 428812 80336 430639 80338
rect 428812 80280 430578 80336
rect 430634 80280 430639 80336
rect 428812 80278 430639 80280
rect 405641 80275 405707 80278
rect 430573 80275 430639 80278
rect 434621 80338 434687 80341
rect 458173 80338 458239 80341
rect 434621 80336 436172 80338
rect 434621 80280 434626 80336
rect 434682 80280 436172 80336
rect 434621 80278 436172 80280
rect 456964 80336 458239 80338
rect 456964 80280 458178 80336
rect 458234 80280 458239 80336
rect 456964 80278 458239 80280
rect 434621 80275 434687 80278
rect 458173 80275 458239 80278
rect 462221 80338 462287 80341
rect 462221 80336 464140 80338
rect 462221 80280 462226 80336
rect 462282 80280 464140 80336
rect 484350 80308 484410 80820
rect 489821 80338 489887 80341
rect 514753 80338 514819 80341
rect 489821 80336 492108 80338
rect 462221 80278 464140 80280
rect 489821 80280 489826 80336
rect 489882 80280 492108 80336
rect 489821 80278 492108 80280
rect 512900 80336 514819 80338
rect 512900 80280 514758 80336
rect 514814 80280 514819 80336
rect 520598 80308 520658 80820
rect 542353 80338 542419 80341
rect 540868 80336 542419 80338
rect 512900 80278 514819 80280
rect 540868 80280 542358 80336
rect 542414 80280 542419 80336
rect 540868 80278 542419 80280
rect 462221 80275 462287 80278
rect 489821 80275 489887 80278
rect 514753 80275 514819 80278
rect 542353 80275 542419 80278
rect 546401 80338 546467 80341
rect 571333 80338 571399 80341
rect 546401 80336 548044 80338
rect 546401 80280 546406 80336
rect 546462 80280 548044 80336
rect 546401 80278 548044 80280
rect 568836 80336 571399 80338
rect 568836 80280 571338 80336
rect 571394 80280 571399 80336
rect 568836 80278 571399 80280
rect 546401 80275 546467 80278
rect 571333 80275 571399 80278
rect 239630 80210 240212 80270
rect 580073 72994 580139 72997
rect 583520 72994 584960 73084
rect 580073 72992 584960 72994
rect 580073 72936 580078 72992
rect 580134 72936 584960 72992
rect 580073 72934 584960 72936
rect 580073 72931 580139 72934
rect 583520 72844 584960 72934
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58578 480 58668
rect 3325 58578 3391 58581
rect -960 58576 3391 58578
rect -960 58520 3330 58576
rect 3386 58520 3391 58576
rect -960 58518 3391 58520
rect -960 58428 480 58518
rect 3325 58515 3391 58518
rect 13537 53818 13603 53821
rect 38653 53818 38719 53821
rect 13537 53816 16100 53818
rect 13537 53760 13542 53816
rect 13598 53760 16100 53816
rect 13537 53758 16100 53760
rect 36892 53816 38719 53818
rect 36892 53760 38658 53816
rect 38714 53760 38719 53816
rect 36892 53758 38719 53760
rect 13537 53755 13603 53758
rect 38653 53755 38719 53758
rect 42701 53818 42767 53821
rect 97901 53818 97967 53821
rect 122833 53818 122899 53821
rect 42701 53816 44068 53818
rect 42701 53760 42706 53816
rect 42762 53760 44068 53816
rect 97901 53816 100188 53818
rect 42701 53758 44068 53760
rect 42701 53755 42767 53758
rect 64462 53412 64522 53788
rect 64454 53348 64460 53412
rect 64524 53348 64530 53412
rect 70301 53274 70367 53277
rect 72006 53274 72066 53788
rect 92430 53276 92490 53788
rect 97901 53760 97906 53816
rect 97962 53760 100188 53816
rect 97901 53758 100188 53760
rect 120796 53816 122899 53818
rect 120796 53760 122838 53816
rect 122894 53760 122899 53816
rect 120796 53758 122899 53760
rect 97901 53755 97967 53758
rect 122833 53755 122899 53758
rect 126881 53818 126947 53821
rect 154481 53818 154547 53821
rect 182081 53818 182147 53821
rect 207013 53818 207079 53821
rect 126881 53816 128156 53818
rect 126881 53760 126886 53816
rect 126942 53760 128156 53816
rect 154481 53816 156124 53818
rect 126881 53758 128156 53760
rect 126881 53755 126947 53758
rect 148366 53276 148426 53788
rect 154481 53760 154486 53816
rect 154542 53760 156124 53816
rect 182081 53816 184092 53818
rect 154481 53758 156124 53760
rect 154481 53755 154547 53758
rect 176334 53276 176394 53788
rect 182081 53760 182086 53816
rect 182142 53760 184092 53816
rect 182081 53758 184092 53760
rect 204884 53816 207079 53818
rect 204884 53760 207018 53816
rect 207074 53760 207079 53816
rect 204884 53758 207079 53760
rect 182081 53755 182147 53758
rect 207013 53755 207079 53758
rect 209681 53818 209747 53821
rect 234705 53818 234771 53821
rect 209681 53816 212060 53818
rect 209681 53760 209686 53816
rect 209742 53760 212060 53816
rect 209681 53758 212060 53760
rect 232852 53816 234771 53818
rect 232852 53760 234710 53816
rect 234766 53760 234771 53816
rect 232852 53758 234771 53760
rect 209681 53755 209747 53758
rect 234705 53755 234771 53758
rect 238661 53818 238727 53821
rect 266261 53818 266327 53821
rect 293861 53818 293927 53821
rect 318793 53818 318859 53821
rect 238661 53816 240212 53818
rect 238661 53760 238666 53816
rect 238722 53760 240212 53816
rect 266261 53816 268180 53818
rect 238661 53758 240212 53760
rect 238661 53755 238727 53758
rect 260422 53276 260482 53788
rect 266261 53760 266266 53816
rect 266322 53760 268180 53816
rect 293861 53816 296148 53818
rect 266261 53758 268180 53760
rect 266261 53755 266327 53758
rect 288390 53276 288450 53788
rect 293861 53760 293866 53816
rect 293922 53760 296148 53816
rect 293861 53758 296148 53760
rect 316940 53816 318859 53818
rect 316940 53760 318798 53816
rect 318854 53760 318859 53816
rect 316940 53758 318859 53760
rect 293861 53755 293927 53758
rect 318793 53755 318859 53758
rect 322841 53818 322907 53821
rect 350441 53818 350507 53821
rect 378041 53818 378107 53821
rect 402973 53818 403039 53821
rect 322841 53816 324116 53818
rect 322841 53760 322846 53816
rect 322902 53760 324116 53816
rect 350441 53816 352084 53818
rect 322841 53758 324116 53760
rect 322841 53755 322907 53758
rect 344326 53276 344386 53788
rect 350441 53760 350446 53816
rect 350502 53760 352084 53816
rect 378041 53816 380052 53818
rect 350441 53758 352084 53760
rect 350441 53755 350507 53758
rect 372294 53276 372354 53788
rect 378041 53760 378046 53816
rect 378102 53760 380052 53816
rect 378041 53758 380052 53760
rect 400844 53816 403039 53818
rect 400844 53760 402978 53816
rect 403034 53760 403039 53816
rect 400844 53758 403039 53760
rect 378041 53755 378107 53758
rect 402973 53755 403039 53758
rect 405641 53818 405707 53821
rect 430573 53818 430639 53821
rect 405641 53816 408204 53818
rect 405641 53760 405646 53816
rect 405702 53760 408204 53816
rect 405641 53758 408204 53760
rect 428812 53816 430639 53818
rect 428812 53760 430578 53816
rect 430634 53760 430639 53816
rect 428812 53758 430639 53760
rect 405641 53755 405707 53758
rect 430573 53755 430639 53758
rect 434621 53818 434687 53821
rect 462221 53818 462287 53821
rect 489821 53818 489887 53821
rect 514753 53818 514819 53821
rect 542353 53818 542419 53821
rect 571333 53818 571399 53821
rect 434621 53816 436172 53818
rect 434621 53760 434626 53816
rect 434682 53760 436172 53816
rect 462221 53816 464140 53818
rect 434621 53758 436172 53760
rect 434621 53755 434687 53758
rect 456382 53276 456442 53788
rect 462221 53760 462226 53816
rect 462282 53760 464140 53816
rect 489821 53816 492108 53818
rect 462221 53758 464140 53760
rect 462221 53755 462287 53758
rect 484350 53276 484410 53788
rect 489821 53760 489826 53816
rect 489882 53760 492108 53816
rect 489821 53758 492108 53760
rect 512900 53816 514819 53818
rect 512900 53760 514758 53816
rect 514814 53760 514819 53816
rect 540868 53816 542419 53818
rect 512900 53758 514819 53760
rect 489821 53755 489887 53758
rect 514753 53755 514819 53758
rect 520598 53276 520658 53788
rect 540868 53760 542358 53816
rect 542414 53760 542419 53816
rect 568836 53816 571399 53818
rect 540868 53758 542419 53760
rect 542353 53755 542419 53758
rect 70301 53272 72066 53274
rect 70301 53216 70306 53272
rect 70362 53216 72066 53272
rect 70301 53214 72066 53216
rect 70301 53211 70367 53214
rect 92422 53212 92428 53276
rect 92492 53212 92498 53276
rect 148358 53212 148364 53276
rect 148428 53212 148434 53276
rect 176326 53212 176332 53276
rect 176396 53212 176402 53276
rect 260414 53212 260420 53276
rect 260484 53212 260490 53276
rect 288382 53212 288388 53276
rect 288452 53212 288458 53276
rect 344318 53212 344324 53276
rect 344388 53212 344394 53276
rect 372286 53212 372292 53276
rect 372356 53212 372362 53276
rect 456374 53212 456380 53276
rect 456444 53212 456450 53276
rect 484342 53212 484348 53276
rect 484412 53212 484418 53276
rect 520590 53212 520596 53276
rect 520660 53212 520666 53276
rect 546401 53274 546467 53277
rect 548014 53274 548074 53788
rect 568836 53760 571338 53816
rect 571394 53760 571399 53816
rect 568836 53758 571399 53760
rect 571333 53755 571399 53758
rect 546401 53272 548074 53274
rect 546401 53216 546406 53272
rect 546462 53216 548074 53272
rect 546401 53214 548074 53216
rect 546401 53211 546467 53214
rect 583520 46188 584960 46428
rect -960 45522 480 45612
rect 2957 45522 3023 45525
rect -960 45520 3023 45522
rect -960 45464 2962 45520
rect 3018 45464 3023 45520
rect -960 45462 3023 45464
rect -960 45372 480 45462
rect 2957 45459 3023 45462
rect 13537 45386 13603 45389
rect 63902 45386 63908 45388
rect 13537 45384 63908 45386
rect 13537 45328 13542 45384
rect 13598 45328 63908 45384
rect 13537 45326 63908 45328
rect 13537 45323 13603 45326
rect 63902 45324 63908 45326
rect 63972 45324 63978 45388
rect 70301 45386 70367 45389
rect 122833 45386 122899 45389
rect 70301 45384 122899 45386
rect 70301 45328 70306 45384
rect 70362 45328 122838 45384
rect 122894 45328 122899 45384
rect 70301 45326 122899 45328
rect 70301 45323 70367 45326
rect 122833 45323 122899 45326
rect 126881 45386 126947 45389
rect 175222 45386 175228 45388
rect 126881 45384 175228 45386
rect 126881 45328 126886 45384
rect 126942 45328 175228 45384
rect 126881 45326 175228 45328
rect 126881 45323 126947 45326
rect 175222 45324 175228 45326
rect 175292 45324 175298 45388
rect 182081 45386 182147 45389
rect 234705 45386 234771 45389
rect 182081 45384 234771 45386
rect 182081 45328 182086 45384
rect 182142 45328 234710 45384
rect 234766 45328 234771 45384
rect 182081 45326 234771 45328
rect 182081 45323 182147 45326
rect 234705 45323 234771 45326
rect 266261 45386 266327 45389
rect 318793 45386 318859 45389
rect 266261 45384 318859 45386
rect 266261 45328 266266 45384
rect 266322 45328 318798 45384
rect 318854 45328 318859 45384
rect 266261 45326 318859 45328
rect 266261 45323 266327 45326
rect 318793 45323 318859 45326
rect 350441 45386 350507 45389
rect 402973 45386 403039 45389
rect 350441 45384 403039 45386
rect 350441 45328 350446 45384
rect 350502 45328 402978 45384
rect 403034 45328 403039 45384
rect 350441 45326 403039 45328
rect 350441 45323 350507 45326
rect 402973 45323 403039 45326
rect 405641 45386 405707 45389
rect 455454 45386 455460 45388
rect 405641 45384 455460 45386
rect 405641 45328 405646 45384
rect 405702 45328 455460 45384
rect 405641 45326 455460 45328
rect 405641 45323 405707 45326
rect 455454 45324 455460 45326
rect 455524 45324 455530 45388
rect 462221 45386 462287 45389
rect 514753 45386 514819 45389
rect 462221 45384 514819 45386
rect 462221 45328 462226 45384
rect 462282 45328 514758 45384
rect 514814 45328 514819 45384
rect 462221 45326 514819 45328
rect 462221 45323 462287 45326
rect 514753 45323 514819 45326
rect 520774 45324 520780 45388
rect 520844 45386 520850 45388
rect 571333 45386 571399 45389
rect 520844 45384 571399 45386
rect 520844 45328 571338 45384
rect 571394 45328 571399 45384
rect 520844 45326 571399 45328
rect 520844 45324 520850 45326
rect 571333 45323 571399 45326
rect 42701 45250 42767 45253
rect 91134 45250 91140 45252
rect 42701 45248 91140 45250
rect 42701 45192 42706 45248
rect 42762 45192 91140 45248
rect 42701 45190 91140 45192
rect 42701 45187 42767 45190
rect 91134 45188 91140 45190
rect 91204 45188 91210 45252
rect 97901 45250 97967 45253
rect 147622 45250 147628 45252
rect 97901 45248 147628 45250
rect 97901 45192 97906 45248
rect 97962 45192 147628 45248
rect 97901 45190 147628 45192
rect 97901 45187 97967 45190
rect 147622 45188 147628 45190
rect 147692 45188 147698 45252
rect 154481 45250 154547 45253
rect 207013 45250 207079 45253
rect 154481 45248 207079 45250
rect 154481 45192 154486 45248
rect 154542 45192 207018 45248
rect 207074 45192 207079 45248
rect 154481 45190 207079 45192
rect 154481 45187 154547 45190
rect 207013 45187 207079 45190
rect 209681 45250 209747 45253
rect 259494 45250 259500 45252
rect 209681 45248 259500 45250
rect 209681 45192 209686 45248
rect 209742 45192 259500 45248
rect 209681 45190 259500 45192
rect 209681 45187 209747 45190
rect 259494 45188 259500 45190
rect 259564 45188 259570 45252
rect 293861 45250 293927 45253
rect 343582 45250 343588 45252
rect 293861 45248 343588 45250
rect 293861 45192 293866 45248
rect 293922 45192 343588 45248
rect 293861 45190 343588 45192
rect 293861 45187 293927 45190
rect 343582 45188 343588 45190
rect 343652 45188 343658 45252
rect 378041 45250 378107 45253
rect 430573 45250 430639 45253
rect 378041 45248 430639 45250
rect 378041 45192 378046 45248
rect 378102 45192 430578 45248
rect 430634 45192 430639 45248
rect 378041 45190 430639 45192
rect 378041 45187 378107 45190
rect 430573 45187 430639 45190
rect 434621 45250 434687 45253
rect 483054 45250 483060 45252
rect 434621 45248 483060 45250
rect 434621 45192 434626 45248
rect 434682 45192 483060 45248
rect 434621 45190 483060 45192
rect 434621 45187 434687 45190
rect 483054 45188 483060 45190
rect 483124 45188 483130 45252
rect 238661 45114 238727 45117
rect 287094 45114 287100 45116
rect 238661 45112 287100 45114
rect 238661 45056 238666 45112
rect 238722 45056 287100 45112
rect 238661 45054 287100 45056
rect 238661 45051 238727 45054
rect 287094 45052 287100 45054
rect 287164 45052 287170 45116
rect 322841 45114 322907 45117
rect 371182 45114 371188 45116
rect 322841 45112 371188 45114
rect 322841 45056 322846 45112
rect 322902 45056 371188 45112
rect 322841 45054 371188 45056
rect 322841 45051 322907 45054
rect 371182 45052 371188 45054
rect 371252 45052 371258 45116
rect 53373 37906 53439 37909
rect 580206 37906 580212 37908
rect 53373 37904 580212 37906
rect 53373 37848 53378 37904
rect 53434 37848 580212 37904
rect 53373 37846 580212 37848
rect 53373 37843 53439 37846
rect 580206 37844 580212 37846
rect 580276 37844 580282 37908
rect 249742 36484 249748 36548
rect 249812 36546 249818 36548
rect 250069 36546 250135 36549
rect 249812 36544 250135 36546
rect 249812 36488 250074 36544
rect 250130 36488 250135 36544
rect 249812 36486 250135 36488
rect 249812 36484 249818 36486
rect 250069 36483 250135 36486
rect 455454 36484 455460 36548
rect 455524 36546 455530 36548
rect 456333 36546 456399 36549
rect 455524 36544 456399 36546
rect 455524 36488 456338 36544
rect 456394 36488 456399 36544
rect 455524 36486 456399 36488
rect 455524 36484 455530 36486
rect 456333 36483 456399 36486
rect 557574 36484 557580 36548
rect 557644 36546 557650 36548
rect 557993 36546 558059 36549
rect 557644 36544 558059 36546
rect 557644 36488 557998 36544
rect 558054 36488 558059 36544
rect 557644 36486 558059 36488
rect 557644 36484 557650 36486
rect 557993 36483 558059 36486
rect 64229 35186 64295 35189
rect 61916 35184 64295 35186
rect 61916 35128 64234 35184
rect 64290 35128 64295 35184
rect 61916 35126 64295 35128
rect 64229 35123 64295 35126
rect 296846 34988 296852 35052
rect 296916 35050 296922 35052
rect 346393 35050 346459 35053
rect 296916 35048 346459 35050
rect 296916 34992 346398 35048
rect 346454 34992 346459 35048
rect 296916 34990 346459 34992
rect 296916 34988 296922 34990
rect 346393 34987 346459 34990
rect 70301 34914 70367 34917
rect 122833 34914 122899 34917
rect 70301 34912 122899 34914
rect 70301 34856 70306 34912
rect 70362 34856 122838 34912
rect 122894 34856 122899 34912
rect 70301 34854 122899 34856
rect 70301 34851 70367 34854
rect 122833 34851 122899 34854
rect 128486 34852 128492 34916
rect 128556 34914 128562 34916
rect 178033 34914 178099 34917
rect 128556 34912 178099 34914
rect 128556 34856 178038 34912
rect 178094 34856 178099 34912
rect 128556 34854 178099 34856
rect 128556 34852 128562 34854
rect 178033 34851 178099 34854
rect 182081 34914 182147 34917
rect 234613 34914 234679 34917
rect 182081 34912 234679 34914
rect 182081 34856 182086 34912
rect 182142 34856 234618 34912
rect 234674 34856 234679 34912
rect 182081 34854 234679 34856
rect 182081 34851 182147 34854
rect 234613 34851 234679 34854
rect 240542 34852 240548 34916
rect 240612 34914 240618 34916
rect 291193 34914 291259 34917
rect 240612 34912 291259 34914
rect 240612 34856 291198 34912
rect 291254 34856 291259 34912
rect 240612 34854 291259 34856
rect 240612 34852 240618 34854
rect 291193 34851 291259 34854
rect 324630 34852 324636 34916
rect 324700 34914 324706 34916
rect 375373 34914 375439 34917
rect 324700 34912 375439 34914
rect 324700 34856 375378 34912
rect 375434 34856 375439 34912
rect 324700 34854 375439 34856
rect 324700 34852 324706 34854
rect 375373 34851 375439 34854
rect 378041 34914 378107 34917
rect 430573 34914 430639 34917
rect 378041 34912 430639 34914
rect 378041 34856 378046 34912
rect 378102 34856 430578 34912
rect 430634 34856 430639 34912
rect 378041 34854 430639 34856
rect 378041 34851 378107 34854
rect 430573 34851 430639 34854
rect 436502 34852 436508 34916
rect 436572 34914 436578 34916
rect 487153 34914 487219 34917
rect 436572 34912 487219 34914
rect 436572 34856 487158 34912
rect 487214 34856 487219 34912
rect 436572 34854 487219 34856
rect 436572 34852 436578 34854
rect 487153 34851 487219 34854
rect 492622 34852 492628 34916
rect 492692 34914 492698 34916
rect 542353 34914 542419 34917
rect 492692 34912 542419 34914
rect 492692 34856 542358 34912
rect 542414 34856 542419 34912
rect 492692 34854 542419 34856
rect 492692 34852 492698 34854
rect 542353 34851 542419 34854
rect 97901 34778 97967 34781
rect 150433 34778 150499 34781
rect 97901 34776 150499 34778
rect 97901 34720 97906 34776
rect 97962 34720 150438 34776
rect 150494 34720 150499 34776
rect 97901 34718 150499 34720
rect 97901 34715 97967 34718
rect 150433 34715 150499 34718
rect 154481 34778 154547 34781
rect 207013 34778 207079 34781
rect 154481 34776 207079 34778
rect 154481 34720 154486 34776
rect 154542 34720 207018 34776
rect 207074 34720 207079 34776
rect 154481 34718 207079 34720
rect 154481 34715 154547 34718
rect 207013 34715 207079 34718
rect 212574 34716 212580 34780
rect 212644 34778 212650 34780
rect 262213 34778 262279 34781
rect 212644 34776 262279 34778
rect 212644 34720 262218 34776
rect 262274 34720 262279 34776
rect 212644 34718 262279 34720
rect 212644 34716 212650 34718
rect 262213 34715 262279 34718
rect 266261 34778 266327 34781
rect 318793 34778 318859 34781
rect 266261 34776 318859 34778
rect 266261 34720 266266 34776
rect 266322 34720 318798 34776
rect 318854 34720 318859 34776
rect 266261 34718 318859 34720
rect 266261 34715 266327 34718
rect 318793 34715 318859 34718
rect 350441 34778 350507 34781
rect 402973 34778 403039 34781
rect 350441 34776 403039 34778
rect 350441 34720 350446 34776
rect 350502 34720 402978 34776
rect 403034 34720 403039 34776
rect 350441 34718 403039 34720
rect 350441 34715 350507 34718
rect 402973 34715 403039 34718
rect 408534 34716 408540 34780
rect 408604 34778 408610 34780
rect 458173 34778 458239 34781
rect 408604 34776 458239 34778
rect 408604 34720 458178 34776
rect 458234 34720 458239 34776
rect 408604 34718 458239 34720
rect 408604 34716 408610 34718
rect 458173 34715 458239 34718
rect 462221 34778 462287 34781
rect 514753 34778 514819 34781
rect 462221 34776 514819 34778
rect 462221 34720 462226 34776
rect 462282 34720 514758 34776
rect 514814 34720 514819 34776
rect 462221 34718 514819 34720
rect 462221 34715 462287 34718
rect 514753 34715 514819 34718
rect 520590 34716 520596 34780
rect 520660 34778 520666 34780
rect 571333 34778 571399 34781
rect 520660 34776 571399 34778
rect 520660 34720 571338 34776
rect 571394 34720 571399 34776
rect 520660 34718 571399 34720
rect 520660 34716 520666 34718
rect 571333 34715 571399 34718
rect 11881 34506 11947 34509
rect 11881 34504 16100 34506
rect 11881 34448 11886 34504
rect 11942 34448 16100 34504
rect 11881 34446 16100 34448
rect 11881 34443 11947 34446
rect 61285 34370 61351 34373
rect 61285 34368 61394 34370
rect 61285 34312 61290 34368
rect 61346 34312 61394 34368
rect 61285 34307 61394 34312
rect 61334 33796 61394 34307
rect 13445 33146 13511 33149
rect 580901 33146 580967 33149
rect 583520 33146 584960 33236
rect 13445 33144 16100 33146
rect 13445 33088 13450 33144
rect 13506 33088 16100 33144
rect 13445 33086 16100 33088
rect 580901 33144 584960 33146
rect 580901 33088 580906 33144
rect 580962 33088 584960 33144
rect 580901 33086 584960 33088
rect 13445 33083 13511 33086
rect 580901 33083 580967 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 64413 31650 64479 31653
rect 61916 31648 64479 31650
rect 61916 31592 64418 31648
rect 64474 31592 64479 31648
rect 61916 31590 64479 31592
rect 64413 31587 64479 31590
rect 12433 31106 12499 31109
rect 12433 31104 16100 31106
rect 12433 31048 12438 31104
rect 12494 31048 16100 31104
rect 12433 31046 16100 31048
rect 12433 31043 12499 31046
rect 64137 30290 64203 30293
rect 61916 30288 64203 30290
rect 61916 30232 64142 30288
rect 64198 30232 64203 30288
rect 61916 30230 64203 30232
rect 64137 30227 64203 30230
rect 13537 29746 13603 29749
rect 13537 29744 16100 29746
rect 13537 29688 13542 29744
rect 13598 29688 16100 29744
rect 13537 29686 16100 29688
rect 13537 29683 13603 29686
rect 64229 28386 64295 28389
rect 61916 28384 64295 28386
rect 61916 28328 64234 28384
rect 64290 28328 64295 28384
rect 61916 28326 64295 28328
rect 64229 28323 64295 28326
rect 13629 27706 13695 27709
rect 13629 27704 16100 27706
rect 13629 27648 13634 27704
rect 13690 27648 16100 27704
rect 13629 27646 16100 27648
rect 13629 27643 13695 27646
rect 63493 27026 63559 27029
rect 61916 27024 63559 27026
rect 61916 26968 63498 27024
rect 63554 26968 63559 27024
rect 61916 26966 63559 26968
rect 63493 26963 63559 26966
rect 70301 26890 70367 26893
rect 70301 26888 72066 26890
rect 70301 26832 70306 26888
rect 70362 26832 72066 26888
rect 70301 26830 72066 26832
rect 70301 26827 70367 26830
rect 13721 26346 13787 26349
rect 13721 26344 16100 26346
rect 13721 26288 13726 26344
rect 13782 26288 16100 26344
rect 72006 26316 72066 26830
rect 128486 26828 128492 26892
rect 128556 26828 128562 26892
rect 212574 26828 212580 26892
rect 212644 26828 212650 26892
rect 240542 26828 240548 26892
rect 240612 26828 240618 26892
rect 296478 26828 296484 26892
rect 296548 26828 296554 26892
rect 324630 26828 324636 26892
rect 324700 26828 324706 26892
rect 408534 26828 408540 26892
rect 408604 26828 408610 26892
rect 436502 26828 436508 26892
rect 436572 26828 436578 26892
rect 458173 26890 458239 26893
rect 456934 26888 458239 26890
rect 456934 26832 458178 26888
rect 458234 26832 458239 26888
rect 456934 26830 458239 26832
rect 95233 26346 95299 26349
rect 92828 26344 95299 26346
rect 13721 26286 16100 26288
rect 92828 26288 95238 26344
rect 95294 26288 95299 26344
rect 92828 26286 95299 26288
rect 13721 26283 13787 26286
rect 95233 26283 95299 26286
rect 97901 26346 97967 26349
rect 122833 26346 122899 26349
rect 97901 26344 100188 26346
rect 97901 26288 97906 26344
rect 97962 26288 100188 26344
rect 97901 26286 100188 26288
rect 120796 26344 122899 26346
rect 120796 26288 122838 26344
rect 122894 26288 122899 26344
rect 128494 26316 128554 26828
rect 150433 26346 150499 26349
rect 148948 26344 150499 26346
rect 120796 26286 122899 26288
rect 148948 26288 150438 26344
rect 150494 26288 150499 26344
rect 148948 26286 150499 26288
rect 97901 26283 97967 26286
rect 122833 26283 122899 26286
rect 150433 26283 150499 26286
rect 154481 26346 154547 26349
rect 178033 26346 178099 26349
rect 154481 26344 156124 26346
rect 154481 26288 154486 26344
rect 154542 26288 156124 26344
rect 154481 26286 156124 26288
rect 176916 26344 178099 26346
rect 176916 26288 178038 26344
rect 178094 26288 178099 26344
rect 176916 26286 178099 26288
rect 154481 26283 154547 26286
rect 178033 26283 178099 26286
rect 182081 26346 182147 26349
rect 207013 26346 207079 26349
rect 182081 26344 184092 26346
rect 182081 26288 182086 26344
rect 182142 26288 184092 26344
rect 182081 26286 184092 26288
rect 204884 26344 207079 26346
rect 204884 26288 207018 26344
rect 207074 26288 207079 26344
rect 212582 26316 212642 26828
rect 234613 26346 234679 26349
rect 232852 26344 234679 26346
rect 204884 26286 207079 26288
rect 232852 26288 234618 26344
rect 234674 26288 234679 26344
rect 240550 26316 240610 26828
rect 262213 26346 262279 26349
rect 260820 26344 262279 26346
rect 232852 26286 234679 26288
rect 260820 26288 262218 26344
rect 262274 26288 262279 26344
rect 260820 26286 262279 26288
rect 182081 26283 182147 26286
rect 207013 26283 207079 26286
rect 234613 26283 234679 26286
rect 262213 26283 262279 26286
rect 266261 26346 266327 26349
rect 291193 26346 291259 26349
rect 266261 26344 268180 26346
rect 266261 26288 266266 26344
rect 266322 26288 268180 26344
rect 266261 26286 268180 26288
rect 288788 26344 291259 26346
rect 288788 26288 291198 26344
rect 291254 26288 291259 26344
rect 296486 26316 296546 26828
rect 318793 26346 318859 26349
rect 316940 26344 318859 26346
rect 288788 26286 291259 26288
rect 316940 26288 318798 26344
rect 318854 26288 318859 26344
rect 324638 26316 324698 26828
rect 346393 26346 346459 26349
rect 344908 26344 346459 26346
rect 316940 26286 318859 26288
rect 344908 26288 346398 26344
rect 346454 26288 346459 26344
rect 344908 26286 346459 26288
rect 266261 26283 266327 26286
rect 291193 26283 291259 26286
rect 318793 26283 318859 26286
rect 346393 26283 346459 26286
rect 350441 26346 350507 26349
rect 375373 26346 375439 26349
rect 350441 26344 352084 26346
rect 350441 26288 350446 26344
rect 350502 26288 352084 26344
rect 350441 26286 352084 26288
rect 372876 26344 375439 26346
rect 372876 26288 375378 26344
rect 375434 26288 375439 26344
rect 372876 26286 375439 26288
rect 350441 26283 350507 26286
rect 375373 26283 375439 26286
rect 378041 26346 378107 26349
rect 402973 26346 403039 26349
rect 378041 26344 380052 26346
rect 378041 26288 378046 26344
rect 378102 26288 380052 26344
rect 378041 26286 380052 26288
rect 400844 26344 403039 26346
rect 400844 26288 402978 26344
rect 403034 26288 403039 26344
rect 408542 26316 408602 26828
rect 430573 26346 430639 26349
rect 428812 26344 430639 26346
rect 400844 26286 403039 26288
rect 428812 26288 430578 26344
rect 430634 26288 430639 26344
rect 436510 26316 436570 26828
rect 456934 26316 456994 26830
rect 458173 26827 458239 26830
rect 492622 26828 492628 26892
rect 492692 26828 492698 26892
rect 520590 26828 520596 26892
rect 520660 26828 520666 26892
rect 462221 26346 462287 26349
rect 487153 26346 487219 26349
rect 462221 26344 464140 26346
rect 428812 26286 430639 26288
rect 378041 26283 378107 26286
rect 402973 26283 403039 26286
rect 430573 26283 430639 26286
rect 462221 26288 462226 26344
rect 462282 26288 464140 26344
rect 462221 26286 464140 26288
rect 484932 26344 487219 26346
rect 484932 26288 487158 26344
rect 487214 26288 487219 26344
rect 492630 26316 492690 26828
rect 514753 26346 514819 26349
rect 512900 26344 514819 26346
rect 484932 26286 487219 26288
rect 512900 26288 514758 26344
rect 514814 26288 514819 26344
rect 520598 26316 520658 26828
rect 542353 26346 542419 26349
rect 540868 26344 542419 26346
rect 512900 26286 514819 26288
rect 540868 26288 542358 26344
rect 542414 26288 542419 26344
rect 540868 26286 542419 26288
rect 462221 26283 462287 26286
rect 487153 26283 487219 26286
rect 514753 26283 514819 26286
rect 542353 26283 542419 26286
rect 546401 26346 546467 26349
rect 571333 26346 571399 26349
rect 546401 26344 548044 26346
rect 546401 26288 546406 26344
rect 546462 26288 548044 26344
rect 546401 26286 548044 26288
rect 568836 26344 571399 26346
rect 568836 26288 571338 26344
rect 571394 26288 571399 26344
rect 568836 26286 571399 26288
rect 546401 26283 546467 26286
rect 571333 26283 571399 26286
rect 64229 24986 64295 24989
rect 61916 24984 64295 24986
rect 61916 24928 64234 24984
rect 64290 24928 64295 24984
rect 61916 24926 64295 24928
rect 64229 24923 64295 24926
rect 13721 24170 13787 24173
rect 13721 24168 16100 24170
rect 13721 24112 13726 24168
rect 13782 24112 16100 24168
rect 13721 24110 16100 24112
rect 13721 24107 13787 24110
rect 64413 23626 64479 23629
rect 61916 23624 64479 23626
rect 61916 23568 64418 23624
rect 64474 23568 64479 23624
rect 61916 23566 64479 23568
rect 64413 23563 64479 23566
rect 12433 22946 12499 22949
rect 12433 22944 16100 22946
rect 12433 22888 12438 22944
rect 12494 22888 16100 22944
rect 12433 22886 16100 22888
rect 12433 22883 12499 22886
rect 63585 21450 63651 21453
rect 61916 21448 63651 21450
rect 61916 21392 63590 21448
rect 63646 21392 63651 21448
rect 61916 21390 63651 21392
rect 63585 21387 63651 21390
rect 12433 20906 12499 20909
rect 12433 20904 16100 20906
rect 12433 20848 12438 20904
rect 12494 20848 16100 20904
rect 12433 20846 16100 20848
rect 12433 20843 12499 20846
rect 63718 20226 63724 20228
rect 61916 20166 63724 20226
rect 63718 20164 63724 20166
rect 63788 20164 63794 20228
rect 583520 19668 584960 19908
rect 12433 19546 12499 19549
rect 12433 19544 16100 19546
rect -960 19410 480 19500
rect 12433 19488 12438 19544
rect 12494 19488 16100 19544
rect 12433 19486 16100 19488
rect 12433 19483 12499 19486
rect 3785 19410 3851 19413
rect -960 19408 3851 19410
rect -960 19352 3790 19408
rect 3846 19352 3851 19408
rect -960 19350 3851 19352
rect -960 19260 480 19350
rect 3785 19347 3851 19350
rect 63493 18186 63559 18189
rect 61916 18184 63559 18186
rect 61916 18128 63498 18184
rect 63554 18128 63559 18184
rect 61916 18126 63559 18128
rect 63493 18123 63559 18126
rect 12433 17506 12499 17509
rect 12433 17504 16100 17506
rect 12433 17448 12438 17504
rect 12494 17448 16100 17504
rect 12433 17446 16100 17448
rect 12433 17443 12499 17446
rect 64321 16826 64387 16829
rect 61916 16824 64387 16826
rect 61916 16768 64326 16824
rect 64382 16768 64387 16824
rect 61916 16766 64387 16768
rect 64321 16763 64387 16766
rect 45001 13698 45067 13701
rect 580574 13698 580580 13700
rect 45001 13696 580580 13698
rect 45001 13640 45006 13696
rect 45062 13640 580580 13696
rect 45001 13638 580580 13640
rect 45001 13635 45067 13638
rect 580574 13636 580580 13638
rect 580644 13636 580650 13700
rect 61101 13562 61167 13565
rect 580390 13562 580396 13564
rect 61101 13560 580396 13562
rect 61101 13504 61106 13560
rect 61162 13504 580396 13560
rect 61101 13502 580396 13504
rect 61101 13499 61167 13502
rect 580390 13500 580396 13502
rect 580460 13500 580466 13564
rect 232589 13426 232655 13429
rect 249742 13426 249748 13428
rect 232589 13424 249748 13426
rect 232589 13368 232594 13424
rect 232650 13368 249748 13424
rect 232589 13366 249748 13368
rect 232589 13363 232655 13366
rect 249742 13364 249748 13366
rect 249812 13364 249818 13428
rect 418337 13426 418403 13429
rect 455454 13426 455460 13428
rect 418337 13424 455460 13426
rect 418337 13368 418342 13424
rect 418398 13368 455460 13424
rect 418337 13366 455460 13368
rect 418337 13363 418403 13366
rect 455454 13364 455460 13366
rect 455524 13364 455530 13428
rect 540605 13426 540671 13429
rect 557574 13426 557580 13428
rect 540605 13424 557580 13426
rect 540605 13368 540610 13424
rect 540666 13368 557580 13424
rect 540605 13366 557580 13368
rect 540605 13363 540671 13366
rect 557574 13364 557580 13366
rect 557644 13364 557650 13428
rect -960 6490 480 6580
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6716
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 580212 697172 580276 697236
rect 165660 684524 165724 684588
rect 259500 684524 259564 684588
rect 361620 684524 361684 684588
rect 445708 684524 445772 684588
rect 557580 684524 557644 684588
rect 580396 670652 580460 670716
rect 165660 662356 165724 662420
rect 259500 662356 259564 662420
rect 361620 662356 361684 662420
rect 445708 662356 445772 662420
rect 557580 662356 557644 662420
rect 81388 657324 81452 657388
rect 128308 657324 128372 657388
rect 194732 657384 194796 657388
rect 194732 657328 194782 657384
rect 194782 657328 194796 657384
rect 194732 657324 194796 657328
rect 277532 657324 277596 657388
rect 390876 657384 390940 657388
rect 390876 657328 390890 657384
rect 390890 657328 390940 657384
rect 390876 657324 390940 657328
rect 473492 657324 473556 657388
rect 520228 657248 520292 657252
rect 520228 657192 520242 657248
rect 520242 657192 520292 657248
rect 520228 657188 520292 657192
rect 176332 655964 176396 656028
rect 456380 655964 456444 656028
rect 568436 655964 568500 656028
rect 176332 648212 176396 648276
rect 456380 648212 456444 648276
rect 568436 648212 568500 648276
rect 580580 643996 580644 644060
rect 81388 634748 81452 634812
rect 128308 634748 128372 634812
rect 194732 634748 194796 634812
rect 277164 634748 277228 634812
rect 390876 634748 390940 634812
rect 473492 634748 473556 634812
rect 520228 634748 520292 634812
rect 165660 630396 165724 630460
rect 259500 630396 259564 630460
rect 361620 630396 361684 630460
rect 445708 630396 445772 630460
rect 557580 630396 557644 630460
rect 165660 608500 165724 608564
rect 259500 608500 259564 608564
rect 361620 608500 361684 608564
rect 445708 608500 445772 608564
rect 557580 608500 557644 608564
rect 128308 603332 128372 603396
rect 194732 603392 194796 603396
rect 194732 603336 194782 603392
rect 194782 603336 194796 603392
rect 194732 603332 194796 603336
rect 390876 603392 390940 603396
rect 390876 603336 390890 603392
rect 390890 603336 390940 603392
rect 390876 603332 390940 603336
rect 288388 602244 288452 602308
rect 484348 602244 484412 602308
rect 92428 602108 92492 602172
rect 148364 602108 148428 602172
rect 260420 602108 260484 602172
rect 344324 602108 344388 602172
rect 456380 602108 456444 602172
rect 492812 602108 492876 602172
rect 64460 601972 64524 602036
rect 176332 601972 176396 602036
rect 372292 601972 372356 602036
rect 520596 601972 520660 602036
rect 64460 594220 64524 594284
rect 92428 594220 92492 594284
rect 148364 594220 148428 594284
rect 176332 594220 176396 594284
rect 260420 594220 260484 594284
rect 288388 594220 288452 594284
rect 344324 594220 344388 594284
rect 372292 594220 372356 594284
rect 456380 594220 456444 594284
rect 484348 594220 484412 594284
rect 492628 594220 492692 594284
rect 520596 594220 520660 594284
rect 128124 580892 128188 580956
rect 194732 580892 194796 580956
rect 390876 580892 390940 580956
rect 165660 576404 165724 576468
rect 259500 576404 259564 576468
rect 361620 576404 361684 576468
rect 445708 576404 445772 576468
rect 557580 576404 557644 576468
rect 165660 554644 165724 554708
rect 259500 554644 259564 554708
rect 361620 554644 361684 554708
rect 445708 554644 445772 554708
rect 557580 554644 557644 554708
rect 128308 549340 128372 549404
rect 194732 549400 194796 549404
rect 194732 549344 194782 549400
rect 194782 549344 194796 549400
rect 194732 549340 194796 549344
rect 390876 549400 390940 549404
rect 390876 549344 390890 549400
rect 390890 549344 390940 549400
rect 390876 549340 390940 549344
rect 288388 548252 288452 548316
rect 372292 548252 372356 548316
rect 92428 548116 92492 548180
rect 148364 548116 148428 548180
rect 212580 548116 212644 548180
rect 296852 548116 296916 548180
rect 484348 548116 484412 548180
rect 540468 548116 540532 548180
rect 64460 547980 64524 548044
rect 176332 547980 176396 548044
rect 408540 547980 408604 548044
rect 520596 547980 520660 548044
rect 64460 540228 64524 540292
rect 92428 540228 92492 540292
rect 148364 540228 148428 540292
rect 176332 540228 176396 540292
rect 212580 540228 212644 540292
rect 288388 540228 288452 540292
rect 296484 540228 296548 540292
rect 372292 540228 372356 540292
rect 408540 540228 408604 540292
rect 484348 540228 484412 540292
rect 520596 540228 520660 540292
rect 540468 540228 540532 540292
rect 128308 527036 128372 527100
rect 194732 527036 194796 527100
rect 390876 527036 390940 527100
rect 165660 522412 165724 522476
rect 259500 522412 259564 522476
rect 361620 522412 361684 522476
rect 445708 522412 445772 522476
rect 557580 522412 557644 522476
rect 44588 520916 44652 520980
rect 176332 520916 176396 520980
rect 288388 520916 288452 520980
rect 484348 520916 484412 520980
rect 212580 520780 212644 520844
rect 296852 520780 296916 520844
rect 408540 520780 408604 520844
rect 492812 520780 492876 520844
rect 372292 520644 372356 520708
rect 520596 520644 520660 520708
rect 44588 512756 44652 512820
rect 176332 512756 176396 512820
rect 212580 512756 212644 512820
rect 288388 512756 288452 512820
rect 296484 512756 296548 512820
rect 372292 512756 372356 512820
rect 408540 512756 408604 512820
rect 484348 512756 484412 512820
rect 492628 512756 492692 512820
rect 520596 512756 520660 512820
rect 165660 500788 165724 500852
rect 259500 500788 259564 500852
rect 361620 500788 361684 500852
rect 445708 500788 445772 500852
rect 557580 500788 557644 500852
rect 194732 495544 194796 495548
rect 194732 495488 194782 495544
rect 194782 495488 194796 495544
rect 194732 495484 194796 495488
rect 390876 495544 390940 495548
rect 390876 495488 390890 495544
rect 390890 495488 390940 495544
rect 390876 495484 390940 495488
rect 128308 495212 128372 495276
rect 64460 485148 64524 485212
rect 92428 485148 92492 485212
rect 148364 485148 148428 485212
rect 176332 485148 176396 485212
rect 212580 485148 212644 485212
rect 288388 485148 288452 485212
rect 296484 485148 296548 485212
rect 372292 485148 372356 485212
rect 408540 485148 408604 485212
rect 484348 485148 484412 485212
rect 520596 485148 520660 485212
rect 540468 485148 540532 485212
rect 64460 477260 64524 477324
rect 176332 477260 176396 477324
rect 408540 477260 408604 477324
rect 520596 477260 520660 477324
rect 92428 477124 92492 477188
rect 148364 477124 148428 477188
rect 212580 477124 212644 477188
rect 296852 477124 296916 477188
rect 484348 477124 484412 477188
rect 540468 477124 540532 477188
rect 288388 476988 288452 477052
rect 372292 476988 372356 477052
rect 128308 473180 128372 473244
rect 194732 473180 194796 473244
rect 390876 473180 390940 473244
rect 81388 468420 81452 468484
rect 165660 468420 165724 468484
rect 259500 468420 259564 468484
rect 361620 468420 361684 468484
rect 445708 468420 445772 468484
rect 455460 468420 455524 468484
rect 557580 468420 557644 468484
rect 212580 466924 212644 466988
rect 408540 466924 408604 466988
rect 44588 466788 44652 466852
rect 240548 466788 240612 466852
rect 296852 466788 296916 466852
rect 436508 466788 436572 466852
rect 492812 466788 492876 466852
rect 128492 466652 128556 466716
rect 324636 466652 324700 466716
rect 520596 466652 520660 466716
rect 44588 458764 44652 458828
rect 128492 458764 128556 458828
rect 212580 458764 212644 458828
rect 240548 458764 240612 458828
rect 296484 458764 296548 458828
rect 324636 458764 324700 458828
rect 408540 458764 408604 458828
rect 436508 458764 436572 458828
rect 492628 458764 492692 458828
rect 520596 458764 520660 458828
rect 81388 445572 81452 445636
rect 165660 445572 165724 445636
rect 259500 445572 259564 445636
rect 361620 445572 361684 445636
rect 455460 445572 455524 445636
rect 557580 445572 557644 445636
rect 445708 445436 445772 445500
rect 128308 441628 128372 441692
rect 194732 441688 194796 441692
rect 194732 441632 194782 441688
rect 194782 441632 194796 441688
rect 194732 441628 194796 441632
rect 390876 441688 390940 441692
rect 390876 441632 390890 441688
rect 390890 441632 390940 441688
rect 390876 441628 390940 441632
rect 64460 431156 64524 431220
rect 92428 431156 92492 431220
rect 148364 431156 148428 431220
rect 176332 431156 176396 431220
rect 260420 431156 260484 431220
rect 288388 431156 288452 431220
rect 344324 431156 344388 431220
rect 372292 431156 372356 431220
rect 456380 431156 456444 431220
rect 484348 431156 484412 431220
rect 492628 431156 492692 431220
rect 520596 431156 520660 431220
rect 64460 423268 64524 423332
rect 176332 423268 176396 423332
rect 372292 423268 372356 423332
rect 520596 423268 520660 423332
rect 92428 423132 92492 423196
rect 148364 423132 148428 423196
rect 260420 423132 260484 423196
rect 344324 423132 344388 423196
rect 456380 423132 456444 423196
rect 492628 423132 492692 423196
rect 288388 422996 288452 423060
rect 484348 422996 484412 423060
rect 128308 419460 128372 419524
rect 194732 419460 194796 419524
rect 390876 419460 390940 419524
rect 81388 414428 81452 414492
rect 165660 414428 165724 414492
rect 259500 414428 259564 414492
rect 361620 414428 361684 414492
rect 445708 414428 445772 414492
rect 455460 414428 455524 414492
rect 557580 414428 557644 414492
rect 44588 403684 44652 403748
rect 128492 403684 128556 403748
rect 212580 403684 212644 403748
rect 240548 403684 240612 403748
rect 296484 403684 296548 403748
rect 324636 403684 324700 403748
rect 408540 403684 408604 403748
rect 436508 403684 436572 403748
rect 492628 403684 492692 403748
rect 520596 403684 520660 403748
rect 128492 395932 128556 395996
rect 408540 395932 408604 395996
rect 520596 395932 520660 395996
rect 44588 395796 44652 395860
rect 240548 395796 240612 395860
rect 324636 395796 324700 395860
rect 436508 395796 436572 395860
rect 492628 395796 492692 395860
rect 212580 395660 212644 395724
rect 296852 395660 296916 395724
rect 81388 391852 81452 391916
rect 165660 391852 165724 391916
rect 259500 391852 259564 391916
rect 361620 391852 361684 391916
rect 455460 391852 455524 391916
rect 557580 391852 557644 391916
rect 445708 391716 445772 391780
rect 128308 387364 128372 387428
rect 194732 387424 194796 387428
rect 194732 387368 194782 387424
rect 194782 387368 194796 387424
rect 194732 387364 194796 387368
rect 390876 387424 390940 387428
rect 390876 387368 390890 387424
rect 390890 387368 390940 387424
rect 390876 387364 390940 387368
rect 176332 377164 176396 377228
rect 456380 377164 456444 377228
rect 568436 377164 568500 377228
rect 175228 369276 175292 369340
rect 455460 369276 455524 369340
rect 566964 369276 567028 369340
rect 128308 365604 128372 365668
rect 194732 365604 194796 365668
rect 390876 365604 390940 365668
rect 165660 360436 165724 360500
rect 259500 360436 259564 360500
rect 361620 360436 361684 360500
rect 445708 360436 445772 360500
rect 557580 360436 557644 360500
rect 44588 349692 44652 349756
rect 128492 349692 128556 349756
rect 212580 349692 212644 349756
rect 240548 349692 240612 349756
rect 296484 349692 296548 349756
rect 324636 349692 324700 349756
rect 408540 349692 408604 349756
rect 436508 349692 436572 349756
rect 492628 349692 492692 349756
rect 520596 349692 520660 349756
rect 408540 341940 408604 342004
rect 520596 341940 520660 342004
rect 240548 341804 240612 341868
rect 324636 341804 324700 341868
rect 436508 341804 436572 341868
rect 492628 341804 492692 341868
rect 44588 341668 44652 341732
rect 128492 341668 128556 341732
rect 212580 341668 212644 341732
rect 296852 341668 296916 341732
rect 165660 337996 165724 338060
rect 259500 337996 259564 338060
rect 361620 337996 361684 338060
rect 445708 337996 445772 338060
rect 557580 337996 557644 338060
rect 128308 333236 128372 333300
rect 194732 333296 194796 333300
rect 194732 333240 194782 333296
rect 194782 333240 194796 333296
rect 194732 333236 194796 333240
rect 390876 333296 390940 333300
rect 390876 333240 390890 333296
rect 390890 333240 390940 333296
rect 390876 333236 390940 333240
rect 568436 323308 568500 323372
rect 176332 323172 176396 323236
rect 456380 323172 456444 323236
rect 175228 315284 175292 315348
rect 455460 315284 455524 315348
rect 566964 315284 567028 315348
rect 128308 311748 128372 311812
rect 194732 311748 194796 311812
rect 390876 311748 390940 311812
rect 165660 306444 165724 306508
rect 259500 306444 259564 306508
rect 361620 306444 361684 306508
rect 445708 306444 445772 306508
rect 557580 306444 557644 306508
rect 44588 295700 44652 295764
rect 176332 295700 176396 295764
rect 212580 295700 212644 295764
rect 288388 295700 288452 295764
rect 296484 295700 296548 295764
rect 372292 295700 372356 295764
rect 408540 295700 408604 295764
rect 484348 295700 484412 295764
rect 492628 295700 492692 295764
rect 520596 295700 520660 295764
rect 176332 287948 176396 288012
rect 372292 287948 372356 288012
rect 520596 287948 520660 288012
rect 44588 287812 44652 287876
rect 212580 287812 212644 287876
rect 296852 287812 296916 287876
rect 408540 287812 408604 287876
rect 492628 287812 492692 287876
rect 288388 287676 288452 287740
rect 484348 287676 484412 287740
rect 165660 284140 165724 284204
rect 259500 284140 259564 284204
rect 361620 284140 361684 284204
rect 445708 284140 445772 284204
rect 557580 284140 557644 284204
rect 277348 279788 277412 279852
rect 81388 279244 81452 279308
rect 128308 279244 128372 279308
rect 194732 279304 194796 279308
rect 194732 279248 194782 279304
rect 194782 279248 194796 279304
rect 194732 279244 194796 279248
rect 390876 279304 390940 279308
rect 390876 279248 390890 279304
rect 390890 279248 390940 279304
rect 390876 279244 390940 279248
rect 473492 279244 473556 279308
rect 520228 279304 520292 279308
rect 520228 279248 520242 279304
rect 520242 279248 520292 279304
rect 520228 279244 520292 279248
rect 176332 278020 176396 278084
rect 456380 278020 456444 278084
rect 566964 278020 567028 278084
rect 176332 270268 176396 270332
rect 456380 270268 456444 270332
rect 568436 270132 568500 270196
rect 81388 256532 81452 256596
rect 128308 256532 128372 256596
rect 194732 256532 194796 256596
rect 277164 256532 277228 256596
rect 390876 256532 390940 256596
rect 473492 256532 473556 256596
rect 520228 256532 520292 256596
rect 165660 252588 165724 252652
rect 259500 252588 259564 252652
rect 361620 252588 361684 252652
rect 445708 252588 445772 252652
rect 557580 252588 557644 252652
rect 165660 230420 165724 230484
rect 259500 230420 259564 230484
rect 361620 230420 361684 230484
rect 445708 230420 445772 230484
rect 557580 230420 557644 230484
rect 128308 225252 128372 225316
rect 194732 225312 194796 225316
rect 194732 225256 194782 225312
rect 194782 225256 194796 225312
rect 194732 225252 194796 225256
rect 288388 224300 288452 224364
rect 92428 224164 92492 224228
rect 148364 224164 148428 224228
rect 260420 224164 260484 224228
rect 492628 224164 492692 224228
rect 64460 224028 64524 224092
rect 176332 224028 176396 224092
rect 520596 224028 520660 224092
rect 64460 216276 64524 216340
rect 92428 216276 92492 216340
rect 148364 216276 148428 216340
rect 176332 216276 176396 216340
rect 260420 216276 260484 216340
rect 288388 216276 288452 216340
rect 492628 216276 492692 216340
rect 520596 216276 520660 216340
rect 128308 202812 128372 202876
rect 194732 202812 194796 202876
rect 63724 201452 63788 201516
rect 259500 198460 259564 198524
rect 361620 198460 361684 198524
rect 445708 198460 445772 198524
rect 259500 176564 259564 176628
rect 361620 176564 361684 176628
rect 445708 176564 445772 176628
rect 148364 170580 148428 170644
rect 128492 170308 128556 170372
rect 372292 170308 372356 170372
rect 344324 170172 344388 170236
rect 540468 170172 540532 170236
rect 408540 170036 408604 170100
rect 520596 170036 520660 170100
rect 128492 162284 128556 162348
rect 148364 162284 148428 162348
rect 344324 162284 344388 162348
rect 372292 162284 372356 162348
rect 408540 162284 408604 162348
rect 520596 162284 520660 162348
rect 540468 162284 540532 162348
rect 361620 144468 361684 144532
rect 445708 144468 445772 144532
rect 361620 122708 361684 122772
rect 445708 122708 445772 122772
rect 194732 117328 194796 117332
rect 194732 117272 194782 117328
rect 194782 117272 194796 117328
rect 194732 117268 194796 117272
rect 324268 117328 324332 117332
rect 324268 117272 324282 117328
rect 324282 117272 324332 117328
rect 324268 117268 324332 117272
rect 260420 116452 260484 116516
rect 176332 116316 176396 116380
rect 92428 116180 92492 116244
rect 148364 116180 148428 116244
rect 540468 116180 540532 116244
rect 64460 116044 64524 116108
rect 408540 116044 408604 116108
rect 520596 116044 520660 116108
rect 64460 108292 64524 108356
rect 92428 108292 92492 108356
rect 148364 108292 148428 108356
rect 176332 108292 176396 108356
rect 260420 108292 260484 108356
rect 408540 108292 408604 108356
rect 520596 108292 520660 108356
rect 540468 108292 540532 108356
rect 194732 95100 194796 95164
rect 324268 95100 324332 95164
rect 372292 88980 372356 89044
rect 44588 88844 44652 88908
rect 288388 88844 288452 88908
rect 296852 88844 296916 88908
rect 484348 88844 484412 88908
rect 176332 88708 176396 88772
rect 520596 88708 520660 88772
rect 44588 80820 44652 80884
rect 176332 80820 176396 80884
rect 288388 80820 288452 80884
rect 296484 80820 296548 80884
rect 372292 80820 372356 80884
rect 484348 80820 484412 80884
rect 520596 80820 520660 80884
rect 64460 53348 64524 53412
rect 92428 53212 92492 53276
rect 148364 53212 148428 53276
rect 176332 53212 176396 53276
rect 260420 53212 260484 53276
rect 288388 53212 288452 53276
rect 344324 53212 344388 53276
rect 372292 53212 372356 53276
rect 456380 53212 456444 53276
rect 484348 53212 484412 53276
rect 520596 53212 520660 53276
rect 63908 45324 63972 45388
rect 175228 45324 175292 45388
rect 455460 45324 455524 45388
rect 520780 45324 520844 45388
rect 91140 45188 91204 45252
rect 147628 45188 147692 45252
rect 259500 45188 259564 45252
rect 343588 45188 343652 45252
rect 483060 45188 483124 45252
rect 287100 45052 287164 45116
rect 371188 45052 371252 45116
rect 580212 37844 580276 37908
rect 249748 36484 249812 36548
rect 455460 36484 455524 36548
rect 557580 36484 557644 36548
rect 296852 34988 296916 35052
rect 128492 34852 128556 34916
rect 240548 34852 240612 34916
rect 324636 34852 324700 34916
rect 436508 34852 436572 34916
rect 492628 34852 492692 34916
rect 212580 34716 212644 34780
rect 408540 34716 408604 34780
rect 520596 34716 520660 34780
rect 128492 26828 128556 26892
rect 212580 26828 212644 26892
rect 240548 26828 240612 26892
rect 296484 26828 296548 26892
rect 324636 26828 324700 26892
rect 408540 26828 408604 26892
rect 436508 26828 436572 26892
rect 492628 26828 492692 26892
rect 520596 26828 520660 26892
rect 63724 20164 63788 20228
rect 580580 13636 580644 13700
rect 580396 13500 580460 13564
rect 249748 13364 249812 13428
rect 455460 13364 455524 13428
rect 557580 13364 557644 13428
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 -7066 -8106 711002
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 -6106 -7146 710042
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 -5146 -6186 709082
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 -4186 -5226 708122
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 -3226 -4266 707162
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 -2266 -3306 706202
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 698454 -2346 705242
rect 37994 705798 38614 711590
rect 37994 705562 38026 705798
rect 38262 705562 38346 705798
rect 38582 705562 38614 705798
rect 37994 705478 38614 705562
rect 37994 705242 38026 705478
rect 38262 705242 38346 705478
rect 38582 705242 38614 705478
rect -2966 698218 -2934 698454
rect -2698 698218 -2614 698454
rect -2378 698218 -2346 698454
rect -2966 698134 -2346 698218
rect -2966 697898 -2934 698134
rect -2698 697898 -2614 698134
rect -2378 697898 -2346 698134
rect -2966 671454 -2346 697898
rect -2966 671218 -2934 671454
rect -2698 671218 -2614 671454
rect -2378 671218 -2346 671454
rect -2966 671134 -2346 671218
rect -2966 670898 -2934 671134
rect -2698 670898 -2614 671134
rect -2378 670898 -2346 671134
rect -2966 644454 -2346 670898
rect -2966 644218 -2934 644454
rect -2698 644218 -2614 644454
rect -2378 644218 -2346 644454
rect -2966 644134 -2346 644218
rect -2966 643898 -2934 644134
rect -2698 643898 -2614 644134
rect -2378 643898 -2346 644134
rect -2966 617454 -2346 643898
rect -2966 617218 -2934 617454
rect -2698 617218 -2614 617454
rect -2378 617218 -2346 617454
rect -2966 617134 -2346 617218
rect -2966 616898 -2934 617134
rect -2698 616898 -2614 617134
rect -2378 616898 -2346 617134
rect -2966 590454 -2346 616898
rect -2966 590218 -2934 590454
rect -2698 590218 -2614 590454
rect -2378 590218 -2346 590454
rect -2966 590134 -2346 590218
rect -2966 589898 -2934 590134
rect -2698 589898 -2614 590134
rect -2378 589898 -2346 590134
rect -2966 563454 -2346 589898
rect -2966 563218 -2934 563454
rect -2698 563218 -2614 563454
rect -2378 563218 -2346 563454
rect -2966 563134 -2346 563218
rect -2966 562898 -2934 563134
rect -2698 562898 -2614 563134
rect -2378 562898 -2346 563134
rect -2966 536454 -2346 562898
rect -2966 536218 -2934 536454
rect -2698 536218 -2614 536454
rect -2378 536218 -2346 536454
rect -2966 536134 -2346 536218
rect -2966 535898 -2934 536134
rect -2698 535898 -2614 536134
rect -2378 535898 -2346 536134
rect -2966 509454 -2346 535898
rect -2966 509218 -2934 509454
rect -2698 509218 -2614 509454
rect -2378 509218 -2346 509454
rect -2966 509134 -2346 509218
rect -2966 508898 -2934 509134
rect -2698 508898 -2614 509134
rect -2378 508898 -2346 509134
rect -2966 482454 -2346 508898
rect -2966 482218 -2934 482454
rect -2698 482218 -2614 482454
rect -2378 482218 -2346 482454
rect -2966 482134 -2346 482218
rect -2966 481898 -2934 482134
rect -2698 481898 -2614 482134
rect -2378 481898 -2346 482134
rect -2966 455454 -2346 481898
rect -2966 455218 -2934 455454
rect -2698 455218 -2614 455454
rect -2378 455218 -2346 455454
rect -2966 455134 -2346 455218
rect -2966 454898 -2934 455134
rect -2698 454898 -2614 455134
rect -2378 454898 -2346 455134
rect -2966 428454 -2346 454898
rect -2966 428218 -2934 428454
rect -2698 428218 -2614 428454
rect -2378 428218 -2346 428454
rect -2966 428134 -2346 428218
rect -2966 427898 -2934 428134
rect -2698 427898 -2614 428134
rect -2378 427898 -2346 428134
rect -2966 401454 -2346 427898
rect -2966 401218 -2934 401454
rect -2698 401218 -2614 401454
rect -2378 401218 -2346 401454
rect -2966 401134 -2346 401218
rect -2966 400898 -2934 401134
rect -2698 400898 -2614 401134
rect -2378 400898 -2346 401134
rect -2966 374454 -2346 400898
rect -2966 374218 -2934 374454
rect -2698 374218 -2614 374454
rect -2378 374218 -2346 374454
rect -2966 374134 -2346 374218
rect -2966 373898 -2934 374134
rect -2698 373898 -2614 374134
rect -2378 373898 -2346 374134
rect -2966 347454 -2346 373898
rect -2966 347218 -2934 347454
rect -2698 347218 -2614 347454
rect -2378 347218 -2346 347454
rect -2966 347134 -2346 347218
rect -2966 346898 -2934 347134
rect -2698 346898 -2614 347134
rect -2378 346898 -2346 347134
rect -2966 320454 -2346 346898
rect -2966 320218 -2934 320454
rect -2698 320218 -2614 320454
rect -2378 320218 -2346 320454
rect -2966 320134 -2346 320218
rect -2966 319898 -2934 320134
rect -2698 319898 -2614 320134
rect -2378 319898 -2346 320134
rect -2966 293454 -2346 319898
rect -2966 293218 -2934 293454
rect -2698 293218 -2614 293454
rect -2378 293218 -2346 293454
rect -2966 293134 -2346 293218
rect -2966 292898 -2934 293134
rect -2698 292898 -2614 293134
rect -2378 292898 -2346 293134
rect -2966 266454 -2346 292898
rect -2966 266218 -2934 266454
rect -2698 266218 -2614 266454
rect -2378 266218 -2346 266454
rect -2966 266134 -2346 266218
rect -2966 265898 -2934 266134
rect -2698 265898 -2614 266134
rect -2378 265898 -2346 266134
rect -2966 239454 -2346 265898
rect -2966 239218 -2934 239454
rect -2698 239218 -2614 239454
rect -2378 239218 -2346 239454
rect -2966 239134 -2346 239218
rect -2966 238898 -2934 239134
rect -2698 238898 -2614 239134
rect -2378 238898 -2346 239134
rect -2966 212454 -2346 238898
rect -2966 212218 -2934 212454
rect -2698 212218 -2614 212454
rect -2378 212218 -2346 212454
rect -2966 212134 -2346 212218
rect -2966 211898 -2934 212134
rect -2698 211898 -2614 212134
rect -2378 211898 -2346 212134
rect -2966 185454 -2346 211898
rect -2966 185218 -2934 185454
rect -2698 185218 -2614 185454
rect -2378 185218 -2346 185454
rect -2966 185134 -2346 185218
rect -2966 184898 -2934 185134
rect -2698 184898 -2614 185134
rect -2378 184898 -2346 185134
rect -2966 158454 -2346 184898
rect -2966 158218 -2934 158454
rect -2698 158218 -2614 158454
rect -2378 158218 -2346 158454
rect -2966 158134 -2346 158218
rect -2966 157898 -2934 158134
rect -2698 157898 -2614 158134
rect -2378 157898 -2346 158134
rect -2966 131454 -2346 157898
rect -2966 131218 -2934 131454
rect -2698 131218 -2614 131454
rect -2378 131218 -2346 131454
rect -2966 131134 -2346 131218
rect -2966 130898 -2934 131134
rect -2698 130898 -2614 131134
rect -2378 130898 -2346 131134
rect -2966 104454 -2346 130898
rect -2966 104218 -2934 104454
rect -2698 104218 -2614 104454
rect -2378 104218 -2346 104454
rect -2966 104134 -2346 104218
rect -2966 103898 -2934 104134
rect -2698 103898 -2614 104134
rect -2378 103898 -2346 104134
rect -2966 77454 -2346 103898
rect -2966 77218 -2934 77454
rect -2698 77218 -2614 77454
rect -2378 77218 -2346 77454
rect -2966 77134 -2346 77218
rect -2966 76898 -2934 77134
rect -2698 76898 -2614 77134
rect -2378 76898 -2346 77134
rect -2966 50454 -2346 76898
rect -2966 50218 -2934 50454
rect -2698 50218 -2614 50454
rect -2378 50218 -2346 50454
rect -2966 50134 -2346 50218
rect -2966 49898 -2934 50134
rect -2698 49898 -2614 50134
rect -2378 49898 -2346 50134
rect -2966 23454 -2346 49898
rect -2966 23218 -2934 23454
rect -2698 23218 -2614 23454
rect -2378 23218 -2346 23454
rect -2966 23134 -2346 23218
rect -2966 22898 -2934 23134
rect -2698 22898 -2614 23134
rect -2378 22898 -2346 23134
rect -2966 -1306 -2346 22898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 701829 -1386 704282
rect -2006 701593 -1974 701829
rect -1738 701593 -1654 701829
rect -1418 701593 -1386 701829
rect -2006 701509 -1386 701593
rect -2006 701273 -1974 701509
rect -1738 701273 -1654 701509
rect -1418 701273 -1386 701509
rect -2006 674829 -1386 701273
rect 37994 698454 38614 705242
rect 37994 698218 38026 698454
rect 38262 698218 38346 698454
rect 38582 698218 38614 698454
rect 37994 698134 38614 698218
rect 37994 697898 38026 698134
rect 38262 697898 38346 698134
rect 38582 697898 38614 698134
rect 37994 687000 38614 697898
rect 41494 704838 42114 711590
rect 41494 704602 41526 704838
rect 41762 704602 41846 704838
rect 42082 704602 42114 704838
rect 41494 704518 42114 704602
rect 41494 704282 41526 704518
rect 41762 704282 41846 704518
rect 42082 704282 42114 704518
rect 41494 701829 42114 704282
rect 41494 701593 41526 701829
rect 41762 701593 41846 701829
rect 42082 701593 42114 701829
rect 41494 701509 42114 701593
rect 41494 701273 41526 701509
rect 41762 701273 41846 701509
rect 42082 701273 42114 701509
rect 41494 687000 42114 701273
rect 65994 705798 66614 711590
rect 65994 705562 66026 705798
rect 66262 705562 66346 705798
rect 66582 705562 66614 705798
rect 65994 705478 66614 705562
rect 65994 705242 66026 705478
rect 66262 705242 66346 705478
rect 66582 705242 66614 705478
rect 65994 698454 66614 705242
rect 65994 698218 66026 698454
rect 66262 698218 66346 698454
rect 66582 698218 66614 698454
rect 65994 698134 66614 698218
rect 65994 697898 66026 698134
rect 66262 697898 66346 698134
rect 66582 697898 66614 698134
rect 65994 687000 66614 697898
rect 69494 704838 70114 711590
rect 69494 704602 69526 704838
rect 69762 704602 69846 704838
rect 70082 704602 70114 704838
rect 69494 704518 70114 704602
rect 69494 704282 69526 704518
rect 69762 704282 69846 704518
rect 70082 704282 70114 704518
rect 69494 701829 70114 704282
rect 69494 701593 69526 701829
rect 69762 701593 69846 701829
rect 70082 701593 70114 701829
rect 69494 701509 70114 701593
rect 69494 701273 69526 701509
rect 69762 701273 69846 701509
rect 70082 701273 70114 701509
rect 69494 687000 70114 701273
rect 93994 705798 94614 711590
rect 93994 705562 94026 705798
rect 94262 705562 94346 705798
rect 94582 705562 94614 705798
rect 93994 705478 94614 705562
rect 93994 705242 94026 705478
rect 94262 705242 94346 705478
rect 94582 705242 94614 705478
rect 93994 698454 94614 705242
rect 93994 698218 94026 698454
rect 94262 698218 94346 698454
rect 94582 698218 94614 698454
rect 93994 698134 94614 698218
rect 93994 697898 94026 698134
rect 94262 697898 94346 698134
rect 94582 697898 94614 698134
rect 93994 687000 94614 697898
rect 97494 704838 98114 711590
rect 97494 704602 97526 704838
rect 97762 704602 97846 704838
rect 98082 704602 98114 704838
rect 97494 704518 98114 704602
rect 97494 704282 97526 704518
rect 97762 704282 97846 704518
rect 98082 704282 98114 704518
rect 97494 701829 98114 704282
rect 97494 701593 97526 701829
rect 97762 701593 97846 701829
rect 98082 701593 98114 701829
rect 97494 701509 98114 701593
rect 97494 701273 97526 701509
rect 97762 701273 97846 701509
rect 98082 701273 98114 701509
rect 97494 687000 98114 701273
rect 121994 705798 122614 711590
rect 121994 705562 122026 705798
rect 122262 705562 122346 705798
rect 122582 705562 122614 705798
rect 121994 705478 122614 705562
rect 121994 705242 122026 705478
rect 122262 705242 122346 705478
rect 122582 705242 122614 705478
rect 121994 698454 122614 705242
rect 121994 698218 122026 698454
rect 122262 698218 122346 698454
rect 122582 698218 122614 698454
rect 121994 698134 122614 698218
rect 121994 697898 122026 698134
rect 122262 697898 122346 698134
rect 122582 697898 122614 698134
rect 121994 687000 122614 697898
rect 125494 704838 126114 711590
rect 125494 704602 125526 704838
rect 125762 704602 125846 704838
rect 126082 704602 126114 704838
rect 125494 704518 126114 704602
rect 125494 704282 125526 704518
rect 125762 704282 125846 704518
rect 126082 704282 126114 704518
rect 125494 701829 126114 704282
rect 125494 701593 125526 701829
rect 125762 701593 125846 701829
rect 126082 701593 126114 701829
rect 125494 701509 126114 701593
rect 125494 701273 125526 701509
rect 125762 701273 125846 701509
rect 126082 701273 126114 701509
rect 125494 687000 126114 701273
rect 149994 705798 150614 711590
rect 149994 705562 150026 705798
rect 150262 705562 150346 705798
rect 150582 705562 150614 705798
rect 149994 705478 150614 705562
rect 149994 705242 150026 705478
rect 150262 705242 150346 705478
rect 150582 705242 150614 705478
rect 149994 698454 150614 705242
rect 149994 698218 150026 698454
rect 150262 698218 150346 698454
rect 150582 698218 150614 698454
rect 149994 698134 150614 698218
rect 149994 697898 150026 698134
rect 150262 697898 150346 698134
rect 150582 697898 150614 698134
rect 149994 687000 150614 697898
rect 153494 704838 154114 711590
rect 153494 704602 153526 704838
rect 153762 704602 153846 704838
rect 154082 704602 154114 704838
rect 153494 704518 154114 704602
rect 153494 704282 153526 704518
rect 153762 704282 153846 704518
rect 154082 704282 154114 704518
rect 153494 701829 154114 704282
rect 153494 701593 153526 701829
rect 153762 701593 153846 701829
rect 154082 701593 154114 701829
rect 153494 701509 154114 701593
rect 153494 701273 153526 701509
rect 153762 701273 153846 701509
rect 154082 701273 154114 701509
rect 153494 687000 154114 701273
rect 177994 705798 178614 711590
rect 177994 705562 178026 705798
rect 178262 705562 178346 705798
rect 178582 705562 178614 705798
rect 177994 705478 178614 705562
rect 177994 705242 178026 705478
rect 178262 705242 178346 705478
rect 178582 705242 178614 705478
rect 177994 698454 178614 705242
rect 177994 698218 178026 698454
rect 178262 698218 178346 698454
rect 178582 698218 178614 698454
rect 177994 698134 178614 698218
rect 177994 697898 178026 698134
rect 178262 697898 178346 698134
rect 178582 697898 178614 698134
rect 177994 687000 178614 697898
rect 181494 704838 182114 711590
rect 181494 704602 181526 704838
rect 181762 704602 181846 704838
rect 182082 704602 182114 704838
rect 181494 704518 182114 704602
rect 181494 704282 181526 704518
rect 181762 704282 181846 704518
rect 182082 704282 182114 704518
rect 181494 701829 182114 704282
rect 181494 701593 181526 701829
rect 181762 701593 181846 701829
rect 182082 701593 182114 701829
rect 181494 701509 182114 701593
rect 181494 701273 181526 701509
rect 181762 701273 181846 701509
rect 182082 701273 182114 701509
rect 181494 687000 182114 701273
rect 205994 705798 206614 711590
rect 205994 705562 206026 705798
rect 206262 705562 206346 705798
rect 206582 705562 206614 705798
rect 205994 705478 206614 705562
rect 205994 705242 206026 705478
rect 206262 705242 206346 705478
rect 206582 705242 206614 705478
rect 205994 698454 206614 705242
rect 205994 698218 206026 698454
rect 206262 698218 206346 698454
rect 206582 698218 206614 698454
rect 205994 698134 206614 698218
rect 205994 697898 206026 698134
rect 206262 697898 206346 698134
rect 206582 697898 206614 698134
rect 205994 687000 206614 697898
rect 209494 704838 210114 711590
rect 209494 704602 209526 704838
rect 209762 704602 209846 704838
rect 210082 704602 210114 704838
rect 209494 704518 210114 704602
rect 209494 704282 209526 704518
rect 209762 704282 209846 704518
rect 210082 704282 210114 704518
rect 209494 701829 210114 704282
rect 209494 701593 209526 701829
rect 209762 701593 209846 701829
rect 210082 701593 210114 701829
rect 209494 701509 210114 701593
rect 209494 701273 209526 701509
rect 209762 701273 209846 701509
rect 210082 701273 210114 701509
rect 209494 687000 210114 701273
rect 233994 705798 234614 711590
rect 233994 705562 234026 705798
rect 234262 705562 234346 705798
rect 234582 705562 234614 705798
rect 233994 705478 234614 705562
rect 233994 705242 234026 705478
rect 234262 705242 234346 705478
rect 234582 705242 234614 705478
rect 233994 698454 234614 705242
rect 233994 698218 234026 698454
rect 234262 698218 234346 698454
rect 234582 698218 234614 698454
rect 233994 698134 234614 698218
rect 233994 697898 234026 698134
rect 234262 697898 234346 698134
rect 234582 697898 234614 698134
rect 233994 687000 234614 697898
rect 237494 704838 238114 711590
rect 237494 704602 237526 704838
rect 237762 704602 237846 704838
rect 238082 704602 238114 704838
rect 237494 704518 238114 704602
rect 237494 704282 237526 704518
rect 237762 704282 237846 704518
rect 238082 704282 238114 704518
rect 237494 701829 238114 704282
rect 237494 701593 237526 701829
rect 237762 701593 237846 701829
rect 238082 701593 238114 701829
rect 237494 701509 238114 701593
rect 237494 701273 237526 701509
rect 237762 701273 237846 701509
rect 238082 701273 238114 701509
rect 237494 687000 238114 701273
rect 261994 705798 262614 711590
rect 261994 705562 262026 705798
rect 262262 705562 262346 705798
rect 262582 705562 262614 705798
rect 261994 705478 262614 705562
rect 261994 705242 262026 705478
rect 262262 705242 262346 705478
rect 262582 705242 262614 705478
rect 261994 698454 262614 705242
rect 261994 698218 262026 698454
rect 262262 698218 262346 698454
rect 262582 698218 262614 698454
rect 261994 698134 262614 698218
rect 261994 697898 262026 698134
rect 262262 697898 262346 698134
rect 262582 697898 262614 698134
rect 261994 687000 262614 697898
rect 265494 704838 266114 711590
rect 265494 704602 265526 704838
rect 265762 704602 265846 704838
rect 266082 704602 266114 704838
rect 265494 704518 266114 704602
rect 265494 704282 265526 704518
rect 265762 704282 265846 704518
rect 266082 704282 266114 704518
rect 265494 701829 266114 704282
rect 265494 701593 265526 701829
rect 265762 701593 265846 701829
rect 266082 701593 266114 701829
rect 265494 701509 266114 701593
rect 265494 701273 265526 701509
rect 265762 701273 265846 701509
rect 266082 701273 266114 701509
rect 265494 687000 266114 701273
rect 289994 705798 290614 711590
rect 289994 705562 290026 705798
rect 290262 705562 290346 705798
rect 290582 705562 290614 705798
rect 289994 705478 290614 705562
rect 289994 705242 290026 705478
rect 290262 705242 290346 705478
rect 290582 705242 290614 705478
rect 289994 698454 290614 705242
rect 289994 698218 290026 698454
rect 290262 698218 290346 698454
rect 290582 698218 290614 698454
rect 289994 698134 290614 698218
rect 289994 697898 290026 698134
rect 290262 697898 290346 698134
rect 290582 697898 290614 698134
rect 289994 687000 290614 697898
rect 293494 704838 294114 711590
rect 293494 704602 293526 704838
rect 293762 704602 293846 704838
rect 294082 704602 294114 704838
rect 293494 704518 294114 704602
rect 293494 704282 293526 704518
rect 293762 704282 293846 704518
rect 294082 704282 294114 704518
rect 293494 701829 294114 704282
rect 293494 701593 293526 701829
rect 293762 701593 293846 701829
rect 294082 701593 294114 701829
rect 293494 701509 294114 701593
rect 293494 701273 293526 701509
rect 293762 701273 293846 701509
rect 294082 701273 294114 701509
rect 293494 687000 294114 701273
rect 317994 705798 318614 711590
rect 317994 705562 318026 705798
rect 318262 705562 318346 705798
rect 318582 705562 318614 705798
rect 317994 705478 318614 705562
rect 317994 705242 318026 705478
rect 318262 705242 318346 705478
rect 318582 705242 318614 705478
rect 317994 698454 318614 705242
rect 317994 698218 318026 698454
rect 318262 698218 318346 698454
rect 318582 698218 318614 698454
rect 317994 698134 318614 698218
rect 317994 697898 318026 698134
rect 318262 697898 318346 698134
rect 318582 697898 318614 698134
rect 317994 687000 318614 697898
rect 321494 704838 322114 711590
rect 321494 704602 321526 704838
rect 321762 704602 321846 704838
rect 322082 704602 322114 704838
rect 321494 704518 322114 704602
rect 321494 704282 321526 704518
rect 321762 704282 321846 704518
rect 322082 704282 322114 704518
rect 321494 701829 322114 704282
rect 321494 701593 321526 701829
rect 321762 701593 321846 701829
rect 322082 701593 322114 701829
rect 321494 701509 322114 701593
rect 321494 701273 321526 701509
rect 321762 701273 321846 701509
rect 322082 701273 322114 701509
rect 321494 687000 322114 701273
rect 345994 705798 346614 711590
rect 345994 705562 346026 705798
rect 346262 705562 346346 705798
rect 346582 705562 346614 705798
rect 345994 705478 346614 705562
rect 345994 705242 346026 705478
rect 346262 705242 346346 705478
rect 346582 705242 346614 705478
rect 345994 698454 346614 705242
rect 345994 698218 346026 698454
rect 346262 698218 346346 698454
rect 346582 698218 346614 698454
rect 345994 698134 346614 698218
rect 345994 697898 346026 698134
rect 346262 697898 346346 698134
rect 346582 697898 346614 698134
rect 345994 687000 346614 697898
rect 349494 704838 350114 711590
rect 349494 704602 349526 704838
rect 349762 704602 349846 704838
rect 350082 704602 350114 704838
rect 349494 704518 350114 704602
rect 349494 704282 349526 704518
rect 349762 704282 349846 704518
rect 350082 704282 350114 704518
rect 349494 701829 350114 704282
rect 349494 701593 349526 701829
rect 349762 701593 349846 701829
rect 350082 701593 350114 701829
rect 349494 701509 350114 701593
rect 349494 701273 349526 701509
rect 349762 701273 349846 701509
rect 350082 701273 350114 701509
rect 349494 687000 350114 701273
rect 373994 705798 374614 711590
rect 373994 705562 374026 705798
rect 374262 705562 374346 705798
rect 374582 705562 374614 705798
rect 373994 705478 374614 705562
rect 373994 705242 374026 705478
rect 374262 705242 374346 705478
rect 374582 705242 374614 705478
rect 373994 698454 374614 705242
rect 373994 698218 374026 698454
rect 374262 698218 374346 698454
rect 374582 698218 374614 698454
rect 373994 698134 374614 698218
rect 373994 697898 374026 698134
rect 374262 697898 374346 698134
rect 374582 697898 374614 698134
rect 373994 687000 374614 697898
rect 377494 704838 378114 711590
rect 377494 704602 377526 704838
rect 377762 704602 377846 704838
rect 378082 704602 378114 704838
rect 377494 704518 378114 704602
rect 377494 704282 377526 704518
rect 377762 704282 377846 704518
rect 378082 704282 378114 704518
rect 377494 701829 378114 704282
rect 377494 701593 377526 701829
rect 377762 701593 377846 701829
rect 378082 701593 378114 701829
rect 377494 701509 378114 701593
rect 377494 701273 377526 701509
rect 377762 701273 377846 701509
rect 378082 701273 378114 701509
rect 377494 687000 378114 701273
rect 401994 705798 402614 711590
rect 401994 705562 402026 705798
rect 402262 705562 402346 705798
rect 402582 705562 402614 705798
rect 401994 705478 402614 705562
rect 401994 705242 402026 705478
rect 402262 705242 402346 705478
rect 402582 705242 402614 705478
rect 401994 698454 402614 705242
rect 401994 698218 402026 698454
rect 402262 698218 402346 698454
rect 402582 698218 402614 698454
rect 401994 698134 402614 698218
rect 401994 697898 402026 698134
rect 402262 697898 402346 698134
rect 402582 697898 402614 698134
rect 401994 687000 402614 697898
rect 405494 704838 406114 711590
rect 405494 704602 405526 704838
rect 405762 704602 405846 704838
rect 406082 704602 406114 704838
rect 405494 704518 406114 704602
rect 405494 704282 405526 704518
rect 405762 704282 405846 704518
rect 406082 704282 406114 704518
rect 405494 701829 406114 704282
rect 405494 701593 405526 701829
rect 405762 701593 405846 701829
rect 406082 701593 406114 701829
rect 405494 701509 406114 701593
rect 405494 701273 405526 701509
rect 405762 701273 405846 701509
rect 406082 701273 406114 701509
rect 405494 687000 406114 701273
rect 429994 705798 430614 711590
rect 429994 705562 430026 705798
rect 430262 705562 430346 705798
rect 430582 705562 430614 705798
rect 429994 705478 430614 705562
rect 429994 705242 430026 705478
rect 430262 705242 430346 705478
rect 430582 705242 430614 705478
rect 429994 698454 430614 705242
rect 429994 698218 430026 698454
rect 430262 698218 430346 698454
rect 430582 698218 430614 698454
rect 429994 698134 430614 698218
rect 429994 697898 430026 698134
rect 430262 697898 430346 698134
rect 430582 697898 430614 698134
rect 429994 687000 430614 697898
rect 433494 704838 434114 711590
rect 433494 704602 433526 704838
rect 433762 704602 433846 704838
rect 434082 704602 434114 704838
rect 433494 704518 434114 704602
rect 433494 704282 433526 704518
rect 433762 704282 433846 704518
rect 434082 704282 434114 704518
rect 433494 701829 434114 704282
rect 433494 701593 433526 701829
rect 433762 701593 433846 701829
rect 434082 701593 434114 701829
rect 433494 701509 434114 701593
rect 433494 701273 433526 701509
rect 433762 701273 433846 701509
rect 434082 701273 434114 701509
rect 433494 687000 434114 701273
rect 457994 705798 458614 711590
rect 457994 705562 458026 705798
rect 458262 705562 458346 705798
rect 458582 705562 458614 705798
rect 457994 705478 458614 705562
rect 457994 705242 458026 705478
rect 458262 705242 458346 705478
rect 458582 705242 458614 705478
rect 457994 698454 458614 705242
rect 457994 698218 458026 698454
rect 458262 698218 458346 698454
rect 458582 698218 458614 698454
rect 457994 698134 458614 698218
rect 457994 697898 458026 698134
rect 458262 697898 458346 698134
rect 458582 697898 458614 698134
rect 457994 687000 458614 697898
rect 461494 704838 462114 711590
rect 461494 704602 461526 704838
rect 461762 704602 461846 704838
rect 462082 704602 462114 704838
rect 461494 704518 462114 704602
rect 461494 704282 461526 704518
rect 461762 704282 461846 704518
rect 462082 704282 462114 704518
rect 461494 701829 462114 704282
rect 461494 701593 461526 701829
rect 461762 701593 461846 701829
rect 462082 701593 462114 701829
rect 461494 701509 462114 701593
rect 461494 701273 461526 701509
rect 461762 701273 461846 701509
rect 462082 701273 462114 701509
rect 461494 687000 462114 701273
rect 485994 705798 486614 711590
rect 485994 705562 486026 705798
rect 486262 705562 486346 705798
rect 486582 705562 486614 705798
rect 485994 705478 486614 705562
rect 485994 705242 486026 705478
rect 486262 705242 486346 705478
rect 486582 705242 486614 705478
rect 485994 698454 486614 705242
rect 485994 698218 486026 698454
rect 486262 698218 486346 698454
rect 486582 698218 486614 698454
rect 485994 698134 486614 698218
rect 485994 697898 486026 698134
rect 486262 697898 486346 698134
rect 486582 697898 486614 698134
rect 485994 687000 486614 697898
rect 489494 704838 490114 711590
rect 489494 704602 489526 704838
rect 489762 704602 489846 704838
rect 490082 704602 490114 704838
rect 489494 704518 490114 704602
rect 489494 704282 489526 704518
rect 489762 704282 489846 704518
rect 490082 704282 490114 704518
rect 489494 701829 490114 704282
rect 489494 701593 489526 701829
rect 489762 701593 489846 701829
rect 490082 701593 490114 701829
rect 489494 701509 490114 701593
rect 489494 701273 489526 701509
rect 489762 701273 489846 701509
rect 490082 701273 490114 701509
rect 489494 687000 490114 701273
rect 513994 705798 514614 711590
rect 513994 705562 514026 705798
rect 514262 705562 514346 705798
rect 514582 705562 514614 705798
rect 513994 705478 514614 705562
rect 513994 705242 514026 705478
rect 514262 705242 514346 705478
rect 514582 705242 514614 705478
rect 513994 698454 514614 705242
rect 513994 698218 514026 698454
rect 514262 698218 514346 698454
rect 514582 698218 514614 698454
rect 513994 698134 514614 698218
rect 513994 697898 514026 698134
rect 514262 697898 514346 698134
rect 514582 697898 514614 698134
rect 513994 687000 514614 697898
rect 517494 704838 518114 711590
rect 517494 704602 517526 704838
rect 517762 704602 517846 704838
rect 518082 704602 518114 704838
rect 517494 704518 518114 704602
rect 517494 704282 517526 704518
rect 517762 704282 517846 704518
rect 518082 704282 518114 704518
rect 517494 701829 518114 704282
rect 517494 701593 517526 701829
rect 517762 701593 517846 701829
rect 518082 701593 518114 701829
rect 517494 701509 518114 701593
rect 517494 701273 517526 701509
rect 517762 701273 517846 701509
rect 518082 701273 518114 701509
rect 517494 687000 518114 701273
rect 541994 705798 542614 711590
rect 541994 705562 542026 705798
rect 542262 705562 542346 705798
rect 542582 705562 542614 705798
rect 541994 705478 542614 705562
rect 541994 705242 542026 705478
rect 542262 705242 542346 705478
rect 542582 705242 542614 705478
rect 541994 698454 542614 705242
rect 541994 698218 542026 698454
rect 542262 698218 542346 698454
rect 542582 698218 542614 698454
rect 541994 698134 542614 698218
rect 541994 697898 542026 698134
rect 542262 697898 542346 698134
rect 542582 697898 542614 698134
rect 541994 687000 542614 697898
rect 545494 704838 546114 711590
rect 545494 704602 545526 704838
rect 545762 704602 545846 704838
rect 546082 704602 546114 704838
rect 545494 704518 546114 704602
rect 545494 704282 545526 704518
rect 545762 704282 545846 704518
rect 546082 704282 546114 704518
rect 545494 701829 546114 704282
rect 545494 701593 545526 701829
rect 545762 701593 545846 701829
rect 546082 701593 546114 701829
rect 545494 701509 546114 701593
rect 545494 701273 545526 701509
rect 545762 701273 545846 701509
rect 546082 701273 546114 701509
rect 545494 687000 546114 701273
rect 569994 705798 570614 711590
rect 569994 705562 570026 705798
rect 570262 705562 570346 705798
rect 570582 705562 570614 705798
rect 569994 705478 570614 705562
rect 569994 705242 570026 705478
rect 570262 705242 570346 705478
rect 570582 705242 570614 705478
rect 569994 698454 570614 705242
rect 569994 698218 570026 698454
rect 570262 698218 570346 698454
rect 570582 698218 570614 698454
rect 569994 698134 570614 698218
rect 569994 697898 570026 698134
rect 570262 697898 570346 698134
rect 570582 697898 570614 698134
rect 569994 687000 570614 697898
rect 573494 704838 574114 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 573494 704602 573526 704838
rect 573762 704602 573846 704838
rect 574082 704602 574114 704838
rect 573494 704518 574114 704602
rect 573494 704282 573526 704518
rect 573762 704282 573846 704518
rect 574082 704282 574114 704518
rect 573494 701829 574114 704282
rect 573494 701593 573526 701829
rect 573762 701593 573846 701829
rect 574082 701593 574114 701829
rect 573494 701509 574114 701593
rect 573494 701273 573526 701509
rect 573762 701273 573846 701509
rect 574082 701273 574114 701509
rect 165659 684588 165725 684589
rect 165659 684524 165660 684588
rect 165724 684524 165725 684588
rect 165659 684523 165725 684524
rect 259499 684588 259565 684589
rect 259499 684524 259500 684588
rect 259564 684524 259565 684588
rect 259499 684523 259565 684524
rect 361619 684588 361685 684589
rect 361619 684524 361620 684588
rect 361684 684524 361685 684588
rect 361619 684523 361685 684524
rect 445707 684588 445773 684589
rect 445707 684524 445708 684588
rect 445772 684524 445773 684588
rect 445707 684523 445773 684524
rect 557579 684588 557645 684589
rect 557579 684524 557580 684588
rect 557644 684524 557645 684588
rect 557579 684523 557645 684524
rect -2006 674593 -1974 674829
rect -1738 674593 -1654 674829
rect -1418 674593 -1386 674829
rect -2006 674509 -1386 674593
rect -2006 674273 -1974 674509
rect -1738 674273 -1654 674509
rect -1418 674273 -1386 674509
rect -2006 647829 -1386 674273
rect 20076 674829 20396 674861
rect 20076 674593 20118 674829
rect 20354 674593 20396 674829
rect 20076 674509 20396 674593
rect 20076 674273 20118 674509
rect 20354 674273 20396 674509
rect 20076 674241 20396 674273
rect 26340 674829 26660 674861
rect 26340 674593 26382 674829
rect 26618 674593 26660 674829
rect 26340 674509 26660 674593
rect 26340 674273 26382 674509
rect 26618 674273 26660 674509
rect 26340 674241 26660 674273
rect 32604 674829 32924 674861
rect 32604 674593 32646 674829
rect 32882 674593 32924 674829
rect 32604 674509 32924 674593
rect 32604 674273 32646 674509
rect 32882 674273 32924 674509
rect 32604 674241 32924 674273
rect 48076 674829 48396 674861
rect 48076 674593 48118 674829
rect 48354 674593 48396 674829
rect 48076 674509 48396 674593
rect 48076 674273 48118 674509
rect 48354 674273 48396 674509
rect 48076 674241 48396 674273
rect 54340 674829 54660 674861
rect 54340 674593 54382 674829
rect 54618 674593 54660 674829
rect 54340 674509 54660 674593
rect 54340 674273 54382 674509
rect 54618 674273 54660 674509
rect 54340 674241 54660 674273
rect 60604 674829 60924 674861
rect 60604 674593 60646 674829
rect 60882 674593 60924 674829
rect 60604 674509 60924 674593
rect 60604 674273 60646 674509
rect 60882 674273 60924 674509
rect 60604 674241 60924 674273
rect 76076 674829 76396 674861
rect 76076 674593 76118 674829
rect 76354 674593 76396 674829
rect 76076 674509 76396 674593
rect 76076 674273 76118 674509
rect 76354 674273 76396 674509
rect 76076 674241 76396 674273
rect 82340 674829 82660 674861
rect 82340 674593 82382 674829
rect 82618 674593 82660 674829
rect 82340 674509 82660 674593
rect 82340 674273 82382 674509
rect 82618 674273 82660 674509
rect 82340 674241 82660 674273
rect 88604 674829 88924 674861
rect 88604 674593 88646 674829
rect 88882 674593 88924 674829
rect 88604 674509 88924 674593
rect 88604 674273 88646 674509
rect 88882 674273 88924 674509
rect 88604 674241 88924 674273
rect 104076 674829 104396 674861
rect 104076 674593 104118 674829
rect 104354 674593 104396 674829
rect 104076 674509 104396 674593
rect 104076 674273 104118 674509
rect 104354 674273 104396 674509
rect 104076 674241 104396 674273
rect 110340 674829 110660 674861
rect 110340 674593 110382 674829
rect 110618 674593 110660 674829
rect 110340 674509 110660 674593
rect 110340 674273 110382 674509
rect 110618 674273 110660 674509
rect 110340 674241 110660 674273
rect 116604 674829 116924 674861
rect 116604 674593 116646 674829
rect 116882 674593 116924 674829
rect 116604 674509 116924 674593
rect 116604 674273 116646 674509
rect 116882 674273 116924 674509
rect 116604 674241 116924 674273
rect 132076 674829 132396 674861
rect 132076 674593 132118 674829
rect 132354 674593 132396 674829
rect 132076 674509 132396 674593
rect 132076 674273 132118 674509
rect 132354 674273 132396 674509
rect 132076 674241 132396 674273
rect 138340 674829 138660 674861
rect 138340 674593 138382 674829
rect 138618 674593 138660 674829
rect 138340 674509 138660 674593
rect 138340 674273 138382 674509
rect 138618 674273 138660 674509
rect 138340 674241 138660 674273
rect 144604 674829 144924 674861
rect 144604 674593 144646 674829
rect 144882 674593 144924 674829
rect 144604 674509 144924 674593
rect 144604 674273 144646 674509
rect 144882 674273 144924 674509
rect 144604 674241 144924 674273
rect 160076 674829 160396 674861
rect 160076 674593 160118 674829
rect 160354 674593 160396 674829
rect 160076 674509 160396 674593
rect 160076 674273 160118 674509
rect 160354 674273 160396 674509
rect 160076 674241 160396 674273
rect 23208 671454 23528 671486
rect 23208 671218 23250 671454
rect 23486 671218 23528 671454
rect 23208 671134 23528 671218
rect 23208 670898 23250 671134
rect 23486 670898 23528 671134
rect 23208 670866 23528 670898
rect 29472 671454 29792 671486
rect 29472 671218 29514 671454
rect 29750 671218 29792 671454
rect 29472 671134 29792 671218
rect 29472 670898 29514 671134
rect 29750 670898 29792 671134
rect 29472 670866 29792 670898
rect 51208 671454 51528 671486
rect 51208 671218 51250 671454
rect 51486 671218 51528 671454
rect 51208 671134 51528 671218
rect 51208 670898 51250 671134
rect 51486 670898 51528 671134
rect 51208 670866 51528 670898
rect 57472 671454 57792 671486
rect 57472 671218 57514 671454
rect 57750 671218 57792 671454
rect 57472 671134 57792 671218
rect 57472 670898 57514 671134
rect 57750 670898 57792 671134
rect 57472 670866 57792 670898
rect 79208 671454 79528 671486
rect 79208 671218 79250 671454
rect 79486 671218 79528 671454
rect 79208 671134 79528 671218
rect 79208 670898 79250 671134
rect 79486 670898 79528 671134
rect 79208 670866 79528 670898
rect 85472 671454 85792 671486
rect 85472 671218 85514 671454
rect 85750 671218 85792 671454
rect 85472 671134 85792 671218
rect 85472 670898 85514 671134
rect 85750 670898 85792 671134
rect 85472 670866 85792 670898
rect 107208 671454 107528 671486
rect 107208 671218 107250 671454
rect 107486 671218 107528 671454
rect 107208 671134 107528 671218
rect 107208 670898 107250 671134
rect 107486 670898 107528 671134
rect 107208 670866 107528 670898
rect 113472 671454 113792 671486
rect 113472 671218 113514 671454
rect 113750 671218 113792 671454
rect 113472 671134 113792 671218
rect 113472 670898 113514 671134
rect 113750 670898 113792 671134
rect 113472 670866 113792 670898
rect 135208 671454 135528 671486
rect 135208 671218 135250 671454
rect 135486 671218 135528 671454
rect 135208 671134 135528 671218
rect 135208 670898 135250 671134
rect 135486 670898 135528 671134
rect 135208 670866 135528 670898
rect 141472 671454 141792 671486
rect 141472 671218 141514 671454
rect 141750 671218 141792 671454
rect 141472 671134 141792 671218
rect 141472 670898 141514 671134
rect 141750 670898 141792 671134
rect 141472 670866 141792 670898
rect 163208 671454 163528 671486
rect 163208 671218 163250 671454
rect 163486 671218 163528 671454
rect 163208 671134 163528 671218
rect 163208 670898 163250 671134
rect 163486 670898 163528 671134
rect 163208 670866 163528 670898
rect 165662 662421 165722 684523
rect 166340 674829 166660 674861
rect 166340 674593 166382 674829
rect 166618 674593 166660 674829
rect 166340 674509 166660 674593
rect 166340 674273 166382 674509
rect 166618 674273 166660 674509
rect 166340 674241 166660 674273
rect 172604 674829 172924 674861
rect 172604 674593 172646 674829
rect 172882 674593 172924 674829
rect 172604 674509 172924 674593
rect 172604 674273 172646 674509
rect 172882 674273 172924 674509
rect 172604 674241 172924 674273
rect 188076 674829 188396 674861
rect 188076 674593 188118 674829
rect 188354 674593 188396 674829
rect 188076 674509 188396 674593
rect 188076 674273 188118 674509
rect 188354 674273 188396 674509
rect 188076 674241 188396 674273
rect 194340 674829 194660 674861
rect 194340 674593 194382 674829
rect 194618 674593 194660 674829
rect 194340 674509 194660 674593
rect 194340 674273 194382 674509
rect 194618 674273 194660 674509
rect 194340 674241 194660 674273
rect 200604 674829 200924 674861
rect 200604 674593 200646 674829
rect 200882 674593 200924 674829
rect 200604 674509 200924 674593
rect 200604 674273 200646 674509
rect 200882 674273 200924 674509
rect 200604 674241 200924 674273
rect 216076 674829 216396 674861
rect 216076 674593 216118 674829
rect 216354 674593 216396 674829
rect 216076 674509 216396 674593
rect 216076 674273 216118 674509
rect 216354 674273 216396 674509
rect 216076 674241 216396 674273
rect 222340 674829 222660 674861
rect 222340 674593 222382 674829
rect 222618 674593 222660 674829
rect 222340 674509 222660 674593
rect 222340 674273 222382 674509
rect 222618 674273 222660 674509
rect 222340 674241 222660 674273
rect 228604 674829 228924 674861
rect 228604 674593 228646 674829
rect 228882 674593 228924 674829
rect 228604 674509 228924 674593
rect 228604 674273 228646 674509
rect 228882 674273 228924 674509
rect 228604 674241 228924 674273
rect 244076 674829 244396 674861
rect 244076 674593 244118 674829
rect 244354 674593 244396 674829
rect 244076 674509 244396 674593
rect 244076 674273 244118 674509
rect 244354 674273 244396 674509
rect 244076 674241 244396 674273
rect 250340 674829 250660 674861
rect 250340 674593 250382 674829
rect 250618 674593 250660 674829
rect 250340 674509 250660 674593
rect 250340 674273 250382 674509
rect 250618 674273 250660 674509
rect 250340 674241 250660 674273
rect 256604 674829 256924 674861
rect 256604 674593 256646 674829
rect 256882 674593 256924 674829
rect 256604 674509 256924 674593
rect 256604 674273 256646 674509
rect 256882 674273 256924 674509
rect 256604 674241 256924 674273
rect 169472 671454 169792 671486
rect 169472 671218 169514 671454
rect 169750 671218 169792 671454
rect 169472 671134 169792 671218
rect 169472 670898 169514 671134
rect 169750 670898 169792 671134
rect 169472 670866 169792 670898
rect 191208 671454 191528 671486
rect 191208 671218 191250 671454
rect 191486 671218 191528 671454
rect 191208 671134 191528 671218
rect 191208 670898 191250 671134
rect 191486 670898 191528 671134
rect 191208 670866 191528 670898
rect 197472 671454 197792 671486
rect 197472 671218 197514 671454
rect 197750 671218 197792 671454
rect 197472 671134 197792 671218
rect 197472 670898 197514 671134
rect 197750 670898 197792 671134
rect 197472 670866 197792 670898
rect 219208 671454 219528 671486
rect 219208 671218 219250 671454
rect 219486 671218 219528 671454
rect 219208 671134 219528 671218
rect 219208 670898 219250 671134
rect 219486 670898 219528 671134
rect 219208 670866 219528 670898
rect 225472 671454 225792 671486
rect 225472 671218 225514 671454
rect 225750 671218 225792 671454
rect 225472 671134 225792 671218
rect 225472 670898 225514 671134
rect 225750 670898 225792 671134
rect 225472 670866 225792 670898
rect 247208 671454 247528 671486
rect 247208 671218 247250 671454
rect 247486 671218 247528 671454
rect 247208 671134 247528 671218
rect 247208 670898 247250 671134
rect 247486 670898 247528 671134
rect 247208 670866 247528 670898
rect 253472 671454 253792 671486
rect 253472 671218 253514 671454
rect 253750 671218 253792 671454
rect 253472 671134 253792 671218
rect 253472 670898 253514 671134
rect 253750 670898 253792 671134
rect 253472 670866 253792 670898
rect 259502 662421 259562 684523
rect 272076 674829 272396 674861
rect 272076 674593 272118 674829
rect 272354 674593 272396 674829
rect 272076 674509 272396 674593
rect 272076 674273 272118 674509
rect 272354 674273 272396 674509
rect 272076 674241 272396 674273
rect 278340 674829 278660 674861
rect 278340 674593 278382 674829
rect 278618 674593 278660 674829
rect 278340 674509 278660 674593
rect 278340 674273 278382 674509
rect 278618 674273 278660 674509
rect 278340 674241 278660 674273
rect 284604 674829 284924 674861
rect 284604 674593 284646 674829
rect 284882 674593 284924 674829
rect 284604 674509 284924 674593
rect 284604 674273 284646 674509
rect 284882 674273 284924 674509
rect 284604 674241 284924 674273
rect 300076 674829 300396 674861
rect 300076 674593 300118 674829
rect 300354 674593 300396 674829
rect 300076 674509 300396 674593
rect 300076 674273 300118 674509
rect 300354 674273 300396 674509
rect 300076 674241 300396 674273
rect 306340 674829 306660 674861
rect 306340 674593 306382 674829
rect 306618 674593 306660 674829
rect 306340 674509 306660 674593
rect 306340 674273 306382 674509
rect 306618 674273 306660 674509
rect 306340 674241 306660 674273
rect 312604 674829 312924 674861
rect 312604 674593 312646 674829
rect 312882 674593 312924 674829
rect 312604 674509 312924 674593
rect 312604 674273 312646 674509
rect 312882 674273 312924 674509
rect 312604 674241 312924 674273
rect 328076 674829 328396 674861
rect 328076 674593 328118 674829
rect 328354 674593 328396 674829
rect 328076 674509 328396 674593
rect 328076 674273 328118 674509
rect 328354 674273 328396 674509
rect 328076 674241 328396 674273
rect 334340 674829 334660 674861
rect 334340 674593 334382 674829
rect 334618 674593 334660 674829
rect 334340 674509 334660 674593
rect 334340 674273 334382 674509
rect 334618 674273 334660 674509
rect 334340 674241 334660 674273
rect 340604 674829 340924 674861
rect 340604 674593 340646 674829
rect 340882 674593 340924 674829
rect 340604 674509 340924 674593
rect 340604 674273 340646 674509
rect 340882 674273 340924 674509
rect 340604 674241 340924 674273
rect 356076 674829 356396 674861
rect 356076 674593 356118 674829
rect 356354 674593 356396 674829
rect 356076 674509 356396 674593
rect 356076 674273 356118 674509
rect 356354 674273 356396 674509
rect 356076 674241 356396 674273
rect 275208 671454 275528 671486
rect 275208 671218 275250 671454
rect 275486 671218 275528 671454
rect 275208 671134 275528 671218
rect 275208 670898 275250 671134
rect 275486 670898 275528 671134
rect 275208 670866 275528 670898
rect 281472 671454 281792 671486
rect 281472 671218 281514 671454
rect 281750 671218 281792 671454
rect 281472 671134 281792 671218
rect 281472 670898 281514 671134
rect 281750 670898 281792 671134
rect 281472 670866 281792 670898
rect 303208 671454 303528 671486
rect 303208 671218 303250 671454
rect 303486 671218 303528 671454
rect 303208 671134 303528 671218
rect 303208 670898 303250 671134
rect 303486 670898 303528 671134
rect 303208 670866 303528 670898
rect 309472 671454 309792 671486
rect 309472 671218 309514 671454
rect 309750 671218 309792 671454
rect 309472 671134 309792 671218
rect 309472 670898 309514 671134
rect 309750 670898 309792 671134
rect 309472 670866 309792 670898
rect 331208 671454 331528 671486
rect 331208 671218 331250 671454
rect 331486 671218 331528 671454
rect 331208 671134 331528 671218
rect 331208 670898 331250 671134
rect 331486 670898 331528 671134
rect 331208 670866 331528 670898
rect 337472 671454 337792 671486
rect 337472 671218 337514 671454
rect 337750 671218 337792 671454
rect 337472 671134 337792 671218
rect 337472 670898 337514 671134
rect 337750 670898 337792 671134
rect 337472 670866 337792 670898
rect 359208 671454 359528 671486
rect 359208 671218 359250 671454
rect 359486 671218 359528 671454
rect 359208 671134 359528 671218
rect 359208 670898 359250 671134
rect 359486 670898 359528 671134
rect 359208 670866 359528 670898
rect 361622 662421 361682 684523
rect 362340 674829 362660 674861
rect 362340 674593 362382 674829
rect 362618 674593 362660 674829
rect 362340 674509 362660 674593
rect 362340 674273 362382 674509
rect 362618 674273 362660 674509
rect 362340 674241 362660 674273
rect 368604 674829 368924 674861
rect 368604 674593 368646 674829
rect 368882 674593 368924 674829
rect 368604 674509 368924 674593
rect 368604 674273 368646 674509
rect 368882 674273 368924 674509
rect 368604 674241 368924 674273
rect 384076 674829 384396 674861
rect 384076 674593 384118 674829
rect 384354 674593 384396 674829
rect 384076 674509 384396 674593
rect 384076 674273 384118 674509
rect 384354 674273 384396 674509
rect 384076 674241 384396 674273
rect 390340 674829 390660 674861
rect 390340 674593 390382 674829
rect 390618 674593 390660 674829
rect 390340 674509 390660 674593
rect 390340 674273 390382 674509
rect 390618 674273 390660 674509
rect 390340 674241 390660 674273
rect 396604 674829 396924 674861
rect 396604 674593 396646 674829
rect 396882 674593 396924 674829
rect 396604 674509 396924 674593
rect 396604 674273 396646 674509
rect 396882 674273 396924 674509
rect 396604 674241 396924 674273
rect 412076 674829 412396 674861
rect 412076 674593 412118 674829
rect 412354 674593 412396 674829
rect 412076 674509 412396 674593
rect 412076 674273 412118 674509
rect 412354 674273 412396 674509
rect 412076 674241 412396 674273
rect 418340 674829 418660 674861
rect 418340 674593 418382 674829
rect 418618 674593 418660 674829
rect 418340 674509 418660 674593
rect 418340 674273 418382 674509
rect 418618 674273 418660 674509
rect 418340 674241 418660 674273
rect 424604 674829 424924 674861
rect 424604 674593 424646 674829
rect 424882 674593 424924 674829
rect 424604 674509 424924 674593
rect 424604 674273 424646 674509
rect 424882 674273 424924 674509
rect 424604 674241 424924 674273
rect 440076 674829 440396 674861
rect 440076 674593 440118 674829
rect 440354 674593 440396 674829
rect 440076 674509 440396 674593
rect 440076 674273 440118 674509
rect 440354 674273 440396 674509
rect 440076 674241 440396 674273
rect 365472 671454 365792 671486
rect 365472 671218 365514 671454
rect 365750 671218 365792 671454
rect 365472 671134 365792 671218
rect 365472 670898 365514 671134
rect 365750 670898 365792 671134
rect 365472 670866 365792 670898
rect 387208 671454 387528 671486
rect 387208 671218 387250 671454
rect 387486 671218 387528 671454
rect 387208 671134 387528 671218
rect 387208 670898 387250 671134
rect 387486 670898 387528 671134
rect 387208 670866 387528 670898
rect 393472 671454 393792 671486
rect 393472 671218 393514 671454
rect 393750 671218 393792 671454
rect 393472 671134 393792 671218
rect 393472 670898 393514 671134
rect 393750 670898 393792 671134
rect 393472 670866 393792 670898
rect 415208 671454 415528 671486
rect 415208 671218 415250 671454
rect 415486 671218 415528 671454
rect 415208 671134 415528 671218
rect 415208 670898 415250 671134
rect 415486 670898 415528 671134
rect 415208 670866 415528 670898
rect 421472 671454 421792 671486
rect 421472 671218 421514 671454
rect 421750 671218 421792 671454
rect 421472 671134 421792 671218
rect 421472 670898 421514 671134
rect 421750 670898 421792 671134
rect 421472 670866 421792 670898
rect 443208 671454 443528 671486
rect 443208 671218 443250 671454
rect 443486 671218 443528 671454
rect 443208 671134 443528 671218
rect 443208 670898 443250 671134
rect 443486 670898 443528 671134
rect 443208 670866 443528 670898
rect 445710 662421 445770 684523
rect 446340 674829 446660 674861
rect 446340 674593 446382 674829
rect 446618 674593 446660 674829
rect 446340 674509 446660 674593
rect 446340 674273 446382 674509
rect 446618 674273 446660 674509
rect 446340 674241 446660 674273
rect 452604 674829 452924 674861
rect 452604 674593 452646 674829
rect 452882 674593 452924 674829
rect 452604 674509 452924 674593
rect 452604 674273 452646 674509
rect 452882 674273 452924 674509
rect 452604 674241 452924 674273
rect 468076 674829 468396 674861
rect 468076 674593 468118 674829
rect 468354 674593 468396 674829
rect 468076 674509 468396 674593
rect 468076 674273 468118 674509
rect 468354 674273 468396 674509
rect 468076 674241 468396 674273
rect 474340 674829 474660 674861
rect 474340 674593 474382 674829
rect 474618 674593 474660 674829
rect 474340 674509 474660 674593
rect 474340 674273 474382 674509
rect 474618 674273 474660 674509
rect 474340 674241 474660 674273
rect 480604 674829 480924 674861
rect 480604 674593 480646 674829
rect 480882 674593 480924 674829
rect 480604 674509 480924 674593
rect 480604 674273 480646 674509
rect 480882 674273 480924 674509
rect 480604 674241 480924 674273
rect 496076 674829 496396 674861
rect 496076 674593 496118 674829
rect 496354 674593 496396 674829
rect 496076 674509 496396 674593
rect 496076 674273 496118 674509
rect 496354 674273 496396 674509
rect 496076 674241 496396 674273
rect 502340 674829 502660 674861
rect 502340 674593 502382 674829
rect 502618 674593 502660 674829
rect 502340 674509 502660 674593
rect 502340 674273 502382 674509
rect 502618 674273 502660 674509
rect 502340 674241 502660 674273
rect 508604 674829 508924 674861
rect 508604 674593 508646 674829
rect 508882 674593 508924 674829
rect 508604 674509 508924 674593
rect 508604 674273 508646 674509
rect 508882 674273 508924 674509
rect 508604 674241 508924 674273
rect 524076 674829 524396 674861
rect 524076 674593 524118 674829
rect 524354 674593 524396 674829
rect 524076 674509 524396 674593
rect 524076 674273 524118 674509
rect 524354 674273 524396 674509
rect 524076 674241 524396 674273
rect 530340 674829 530660 674861
rect 530340 674593 530382 674829
rect 530618 674593 530660 674829
rect 530340 674509 530660 674593
rect 530340 674273 530382 674509
rect 530618 674273 530660 674509
rect 530340 674241 530660 674273
rect 536604 674829 536924 674861
rect 536604 674593 536646 674829
rect 536882 674593 536924 674829
rect 536604 674509 536924 674593
rect 536604 674273 536646 674509
rect 536882 674273 536924 674509
rect 536604 674241 536924 674273
rect 552076 674829 552396 674861
rect 552076 674593 552118 674829
rect 552354 674593 552396 674829
rect 552076 674509 552396 674593
rect 552076 674273 552118 674509
rect 552354 674273 552396 674509
rect 552076 674241 552396 674273
rect 449472 671454 449792 671486
rect 449472 671218 449514 671454
rect 449750 671218 449792 671454
rect 449472 671134 449792 671218
rect 449472 670898 449514 671134
rect 449750 670898 449792 671134
rect 449472 670866 449792 670898
rect 471208 671454 471528 671486
rect 471208 671218 471250 671454
rect 471486 671218 471528 671454
rect 471208 671134 471528 671218
rect 471208 670898 471250 671134
rect 471486 670898 471528 671134
rect 471208 670866 471528 670898
rect 477472 671454 477792 671486
rect 477472 671218 477514 671454
rect 477750 671218 477792 671454
rect 477472 671134 477792 671218
rect 477472 670898 477514 671134
rect 477750 670898 477792 671134
rect 477472 670866 477792 670898
rect 499208 671454 499528 671486
rect 499208 671218 499250 671454
rect 499486 671218 499528 671454
rect 499208 671134 499528 671218
rect 499208 670898 499250 671134
rect 499486 670898 499528 671134
rect 499208 670866 499528 670898
rect 505472 671454 505792 671486
rect 505472 671218 505514 671454
rect 505750 671218 505792 671454
rect 505472 671134 505792 671218
rect 505472 670898 505514 671134
rect 505750 670898 505792 671134
rect 505472 670866 505792 670898
rect 527208 671454 527528 671486
rect 527208 671218 527250 671454
rect 527486 671218 527528 671454
rect 527208 671134 527528 671218
rect 527208 670898 527250 671134
rect 527486 670898 527528 671134
rect 527208 670866 527528 670898
rect 533472 671454 533792 671486
rect 533472 671218 533514 671454
rect 533750 671218 533792 671454
rect 533472 671134 533792 671218
rect 533472 670898 533514 671134
rect 533750 670898 533792 671134
rect 533472 670866 533792 670898
rect 555208 671454 555528 671486
rect 555208 671218 555250 671454
rect 555486 671218 555528 671454
rect 555208 671134 555528 671218
rect 555208 670898 555250 671134
rect 555486 670898 555528 671134
rect 555208 670866 555528 670898
rect 557582 662421 557642 684523
rect 558340 674829 558660 674861
rect 558340 674593 558382 674829
rect 558618 674593 558660 674829
rect 558340 674509 558660 674593
rect 558340 674273 558382 674509
rect 558618 674273 558660 674509
rect 558340 674241 558660 674273
rect 564604 674829 564924 674861
rect 564604 674593 564646 674829
rect 564882 674593 564924 674829
rect 564604 674509 564924 674593
rect 564604 674273 564646 674509
rect 564882 674273 564924 674509
rect 564604 674241 564924 674273
rect 573494 674829 574114 701273
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 701829 585930 704282
rect 585310 701593 585342 701829
rect 585578 701593 585662 701829
rect 585898 701593 585930 701829
rect 585310 701509 585930 701593
rect 585310 701273 585342 701509
rect 585578 701273 585662 701509
rect 585898 701273 585930 701509
rect 580211 697236 580277 697237
rect 580211 697172 580212 697236
rect 580276 697172 580277 697236
rect 580211 697171 580277 697172
rect 573494 674593 573526 674829
rect 573762 674593 573846 674829
rect 574082 674593 574114 674829
rect 573494 674509 574114 674593
rect 573494 674273 573526 674509
rect 573762 674273 573846 674509
rect 574082 674273 574114 674509
rect 561472 671454 561792 671486
rect 561472 671218 561514 671454
rect 561750 671218 561792 671454
rect 561472 671134 561792 671218
rect 561472 670898 561514 671134
rect 561750 670898 561792 671134
rect 561472 670866 561792 670898
rect 165659 662420 165725 662421
rect 165659 662356 165660 662420
rect 165724 662356 165725 662420
rect 165659 662355 165725 662356
rect 259499 662420 259565 662421
rect 259499 662356 259500 662420
rect 259564 662356 259565 662420
rect 259499 662355 259565 662356
rect 361619 662420 361685 662421
rect 361619 662356 361620 662420
rect 361684 662356 361685 662420
rect 361619 662355 361685 662356
rect 445707 662420 445773 662421
rect 445707 662356 445708 662420
rect 445772 662356 445773 662420
rect 445707 662355 445773 662356
rect 557579 662420 557645 662421
rect 557579 662356 557580 662420
rect 557644 662356 557645 662420
rect 557579 662355 557645 662356
rect 81387 657388 81453 657389
rect 81387 657324 81388 657388
rect 81452 657324 81453 657388
rect 81387 657323 81453 657324
rect 128307 657388 128373 657389
rect 128307 657324 128308 657388
rect 128372 657324 128373 657388
rect 128307 657323 128373 657324
rect 194731 657388 194797 657389
rect 194731 657324 194732 657388
rect 194796 657324 194797 657388
rect 194731 657323 194797 657324
rect 277531 657388 277597 657389
rect 277531 657324 277532 657388
rect 277596 657324 277597 657388
rect 277531 657323 277597 657324
rect 390875 657388 390941 657389
rect 390875 657324 390876 657388
rect 390940 657324 390941 657388
rect 390875 657323 390941 657324
rect 473491 657388 473557 657389
rect 473491 657324 473492 657388
rect 473556 657324 473557 657388
rect 473491 657323 473557 657324
rect -2006 647593 -1974 647829
rect -1738 647593 -1654 647829
rect -1418 647593 -1386 647829
rect -2006 647509 -1386 647593
rect -2006 647273 -1974 647509
rect -1738 647273 -1654 647509
rect -1418 647273 -1386 647509
rect -2006 620829 -1386 647273
rect 20076 647829 20396 647861
rect 20076 647593 20118 647829
rect 20354 647593 20396 647829
rect 20076 647509 20396 647593
rect 20076 647273 20118 647509
rect 20354 647273 20396 647509
rect 20076 647241 20396 647273
rect 26340 647829 26660 647861
rect 26340 647593 26382 647829
rect 26618 647593 26660 647829
rect 26340 647509 26660 647593
rect 26340 647273 26382 647509
rect 26618 647273 26660 647509
rect 26340 647241 26660 647273
rect 32604 647829 32924 647861
rect 32604 647593 32646 647829
rect 32882 647593 32924 647829
rect 32604 647509 32924 647593
rect 32604 647273 32646 647509
rect 32882 647273 32924 647509
rect 32604 647241 32924 647273
rect 48076 647829 48396 647861
rect 48076 647593 48118 647829
rect 48354 647593 48396 647829
rect 48076 647509 48396 647593
rect 48076 647273 48118 647509
rect 48354 647273 48396 647509
rect 48076 647241 48396 647273
rect 54340 647829 54660 647861
rect 54340 647593 54382 647829
rect 54618 647593 54660 647829
rect 54340 647509 54660 647593
rect 54340 647273 54382 647509
rect 54618 647273 54660 647509
rect 54340 647241 54660 647273
rect 60604 647829 60924 647861
rect 60604 647593 60646 647829
rect 60882 647593 60924 647829
rect 60604 647509 60924 647593
rect 60604 647273 60646 647509
rect 60882 647273 60924 647509
rect 60604 647241 60924 647273
rect 76076 647829 76396 647861
rect 76076 647593 76118 647829
rect 76354 647593 76396 647829
rect 76076 647509 76396 647593
rect 76076 647273 76118 647509
rect 76354 647273 76396 647509
rect 76076 647241 76396 647273
rect 23208 644454 23528 644486
rect 23208 644218 23250 644454
rect 23486 644218 23528 644454
rect 23208 644134 23528 644218
rect 23208 643898 23250 644134
rect 23486 643898 23528 644134
rect 23208 643866 23528 643898
rect 29472 644454 29792 644486
rect 29472 644218 29514 644454
rect 29750 644218 29792 644454
rect 29472 644134 29792 644218
rect 29472 643898 29514 644134
rect 29750 643898 29792 644134
rect 29472 643866 29792 643898
rect 51208 644454 51528 644486
rect 51208 644218 51250 644454
rect 51486 644218 51528 644454
rect 51208 644134 51528 644218
rect 51208 643898 51250 644134
rect 51486 643898 51528 644134
rect 51208 643866 51528 643898
rect 57472 644454 57792 644486
rect 57472 644218 57514 644454
rect 57750 644218 57792 644454
rect 57472 644134 57792 644218
rect 57472 643898 57514 644134
rect 57750 643898 57792 644134
rect 57472 643866 57792 643898
rect 79208 644454 79528 644486
rect 79208 644218 79250 644454
rect 79486 644218 79528 644454
rect 79208 644134 79528 644218
rect 79208 643898 79250 644134
rect 79486 643898 79528 644134
rect 79208 643866 79528 643898
rect 81390 634813 81450 657323
rect 82340 647829 82660 647861
rect 82340 647593 82382 647829
rect 82618 647593 82660 647829
rect 82340 647509 82660 647593
rect 82340 647273 82382 647509
rect 82618 647273 82660 647509
rect 82340 647241 82660 647273
rect 88604 647829 88924 647861
rect 88604 647593 88646 647829
rect 88882 647593 88924 647829
rect 88604 647509 88924 647593
rect 88604 647273 88646 647509
rect 88882 647273 88924 647509
rect 88604 647241 88924 647273
rect 104076 647829 104396 647861
rect 104076 647593 104118 647829
rect 104354 647593 104396 647829
rect 104076 647509 104396 647593
rect 104076 647273 104118 647509
rect 104354 647273 104396 647509
rect 104076 647241 104396 647273
rect 110340 647829 110660 647861
rect 110340 647593 110382 647829
rect 110618 647593 110660 647829
rect 110340 647509 110660 647593
rect 110340 647273 110382 647509
rect 110618 647273 110660 647509
rect 110340 647241 110660 647273
rect 116604 647829 116924 647861
rect 116604 647593 116646 647829
rect 116882 647593 116924 647829
rect 116604 647509 116924 647593
rect 116604 647273 116646 647509
rect 116882 647273 116924 647509
rect 116604 647241 116924 647273
rect 85472 644454 85792 644486
rect 85472 644218 85514 644454
rect 85750 644218 85792 644454
rect 85472 644134 85792 644218
rect 85472 643898 85514 644134
rect 85750 643898 85792 644134
rect 85472 643866 85792 643898
rect 107208 644454 107528 644486
rect 107208 644218 107250 644454
rect 107486 644218 107528 644454
rect 107208 644134 107528 644218
rect 107208 643898 107250 644134
rect 107486 643898 107528 644134
rect 107208 643866 107528 643898
rect 113472 644454 113792 644486
rect 113472 644218 113514 644454
rect 113750 644218 113792 644454
rect 113472 644134 113792 644218
rect 113472 643898 113514 644134
rect 113750 643898 113792 644134
rect 113472 643866 113792 643898
rect 128310 634813 128370 657323
rect 176331 656028 176397 656029
rect 176331 655964 176332 656028
rect 176396 655964 176397 656028
rect 176331 655963 176397 655964
rect 176334 648277 176394 655963
rect 176331 648276 176397 648277
rect 176331 648212 176332 648276
rect 176396 648212 176397 648276
rect 176331 648211 176397 648212
rect 132076 647829 132396 647861
rect 132076 647593 132118 647829
rect 132354 647593 132396 647829
rect 132076 647509 132396 647593
rect 132076 647273 132118 647509
rect 132354 647273 132396 647509
rect 132076 647241 132396 647273
rect 138340 647829 138660 647861
rect 138340 647593 138382 647829
rect 138618 647593 138660 647829
rect 138340 647509 138660 647593
rect 138340 647273 138382 647509
rect 138618 647273 138660 647509
rect 138340 647241 138660 647273
rect 144604 647829 144924 647861
rect 144604 647593 144646 647829
rect 144882 647593 144924 647829
rect 144604 647509 144924 647593
rect 144604 647273 144646 647509
rect 144882 647273 144924 647509
rect 144604 647241 144924 647273
rect 160076 647829 160396 647861
rect 160076 647593 160118 647829
rect 160354 647593 160396 647829
rect 160076 647509 160396 647593
rect 160076 647273 160118 647509
rect 160354 647273 160396 647509
rect 160076 647241 160396 647273
rect 166340 647829 166660 647861
rect 166340 647593 166382 647829
rect 166618 647593 166660 647829
rect 166340 647509 166660 647593
rect 166340 647273 166382 647509
rect 166618 647273 166660 647509
rect 166340 647241 166660 647273
rect 172604 647829 172924 647861
rect 172604 647593 172646 647829
rect 172882 647593 172924 647829
rect 172604 647509 172924 647593
rect 172604 647273 172646 647509
rect 172882 647273 172924 647509
rect 172604 647241 172924 647273
rect 188076 647829 188396 647861
rect 188076 647593 188118 647829
rect 188354 647593 188396 647829
rect 188076 647509 188396 647593
rect 188076 647273 188118 647509
rect 188354 647273 188396 647509
rect 188076 647241 188396 647273
rect 194340 647829 194660 647861
rect 194340 647593 194382 647829
rect 194618 647593 194660 647829
rect 194340 647509 194660 647593
rect 194340 647273 194382 647509
rect 194618 647273 194660 647509
rect 194340 647241 194660 647273
rect 135208 644454 135528 644486
rect 135208 644218 135250 644454
rect 135486 644218 135528 644454
rect 135208 644134 135528 644218
rect 135208 643898 135250 644134
rect 135486 643898 135528 644134
rect 135208 643866 135528 643898
rect 141472 644454 141792 644486
rect 141472 644218 141514 644454
rect 141750 644218 141792 644454
rect 141472 644134 141792 644218
rect 141472 643898 141514 644134
rect 141750 643898 141792 644134
rect 141472 643866 141792 643898
rect 163208 644454 163528 644486
rect 163208 644218 163250 644454
rect 163486 644218 163528 644454
rect 163208 644134 163528 644218
rect 163208 643898 163250 644134
rect 163486 643898 163528 644134
rect 163208 643866 163528 643898
rect 169472 644454 169792 644486
rect 169472 644218 169514 644454
rect 169750 644218 169792 644454
rect 169472 644134 169792 644218
rect 169472 643898 169514 644134
rect 169750 643898 169792 644134
rect 169472 643866 169792 643898
rect 191208 644454 191528 644486
rect 191208 644218 191250 644454
rect 191486 644218 191528 644454
rect 191208 644134 191528 644218
rect 191208 643898 191250 644134
rect 191486 643898 191528 644134
rect 191208 643866 191528 643898
rect 194734 634813 194794 657323
rect 277534 657250 277594 657323
rect 277166 657190 277594 657250
rect 200604 647829 200924 647861
rect 200604 647593 200646 647829
rect 200882 647593 200924 647829
rect 200604 647509 200924 647593
rect 200604 647273 200646 647509
rect 200882 647273 200924 647509
rect 200604 647241 200924 647273
rect 216076 647829 216396 647861
rect 216076 647593 216118 647829
rect 216354 647593 216396 647829
rect 216076 647509 216396 647593
rect 216076 647273 216118 647509
rect 216354 647273 216396 647509
rect 216076 647241 216396 647273
rect 222340 647829 222660 647861
rect 222340 647593 222382 647829
rect 222618 647593 222660 647829
rect 222340 647509 222660 647593
rect 222340 647273 222382 647509
rect 222618 647273 222660 647509
rect 222340 647241 222660 647273
rect 228604 647829 228924 647861
rect 228604 647593 228646 647829
rect 228882 647593 228924 647829
rect 228604 647509 228924 647593
rect 228604 647273 228646 647509
rect 228882 647273 228924 647509
rect 228604 647241 228924 647273
rect 244076 647829 244396 647861
rect 244076 647593 244118 647829
rect 244354 647593 244396 647829
rect 244076 647509 244396 647593
rect 244076 647273 244118 647509
rect 244354 647273 244396 647509
rect 244076 647241 244396 647273
rect 250340 647829 250660 647861
rect 250340 647593 250382 647829
rect 250618 647593 250660 647829
rect 250340 647509 250660 647593
rect 250340 647273 250382 647509
rect 250618 647273 250660 647509
rect 250340 647241 250660 647273
rect 256604 647829 256924 647861
rect 256604 647593 256646 647829
rect 256882 647593 256924 647829
rect 256604 647509 256924 647593
rect 256604 647273 256646 647509
rect 256882 647273 256924 647509
rect 256604 647241 256924 647273
rect 272076 647829 272396 647861
rect 272076 647593 272118 647829
rect 272354 647593 272396 647829
rect 272076 647509 272396 647593
rect 272076 647273 272118 647509
rect 272354 647273 272396 647509
rect 272076 647241 272396 647273
rect 197472 644454 197792 644486
rect 197472 644218 197514 644454
rect 197750 644218 197792 644454
rect 197472 644134 197792 644218
rect 197472 643898 197514 644134
rect 197750 643898 197792 644134
rect 197472 643866 197792 643898
rect 219208 644454 219528 644486
rect 219208 644218 219250 644454
rect 219486 644218 219528 644454
rect 219208 644134 219528 644218
rect 219208 643898 219250 644134
rect 219486 643898 219528 644134
rect 219208 643866 219528 643898
rect 225472 644454 225792 644486
rect 225472 644218 225514 644454
rect 225750 644218 225792 644454
rect 225472 644134 225792 644218
rect 225472 643898 225514 644134
rect 225750 643898 225792 644134
rect 225472 643866 225792 643898
rect 247208 644454 247528 644486
rect 247208 644218 247250 644454
rect 247486 644218 247528 644454
rect 247208 644134 247528 644218
rect 247208 643898 247250 644134
rect 247486 643898 247528 644134
rect 247208 643866 247528 643898
rect 253472 644454 253792 644486
rect 253472 644218 253514 644454
rect 253750 644218 253792 644454
rect 253472 644134 253792 644218
rect 253472 643898 253514 644134
rect 253750 643898 253792 644134
rect 253472 643866 253792 643898
rect 275208 644454 275528 644486
rect 275208 644218 275250 644454
rect 275486 644218 275528 644454
rect 275208 644134 275528 644218
rect 275208 643898 275250 644134
rect 275486 643898 275528 644134
rect 275208 643866 275528 643898
rect 277166 634813 277226 657190
rect 278340 647829 278660 647861
rect 278340 647593 278382 647829
rect 278618 647593 278660 647829
rect 278340 647509 278660 647593
rect 278340 647273 278382 647509
rect 278618 647273 278660 647509
rect 278340 647241 278660 647273
rect 284604 647829 284924 647861
rect 284604 647593 284646 647829
rect 284882 647593 284924 647829
rect 284604 647509 284924 647593
rect 284604 647273 284646 647509
rect 284882 647273 284924 647509
rect 284604 647241 284924 647273
rect 300076 647829 300396 647861
rect 300076 647593 300118 647829
rect 300354 647593 300396 647829
rect 300076 647509 300396 647593
rect 300076 647273 300118 647509
rect 300354 647273 300396 647509
rect 300076 647241 300396 647273
rect 306340 647829 306660 647861
rect 306340 647593 306382 647829
rect 306618 647593 306660 647829
rect 306340 647509 306660 647593
rect 306340 647273 306382 647509
rect 306618 647273 306660 647509
rect 306340 647241 306660 647273
rect 312604 647829 312924 647861
rect 312604 647593 312646 647829
rect 312882 647593 312924 647829
rect 312604 647509 312924 647593
rect 312604 647273 312646 647509
rect 312882 647273 312924 647509
rect 312604 647241 312924 647273
rect 328076 647829 328396 647861
rect 328076 647593 328118 647829
rect 328354 647593 328396 647829
rect 328076 647509 328396 647593
rect 328076 647273 328118 647509
rect 328354 647273 328396 647509
rect 328076 647241 328396 647273
rect 334340 647829 334660 647861
rect 334340 647593 334382 647829
rect 334618 647593 334660 647829
rect 334340 647509 334660 647593
rect 334340 647273 334382 647509
rect 334618 647273 334660 647509
rect 334340 647241 334660 647273
rect 340604 647829 340924 647861
rect 340604 647593 340646 647829
rect 340882 647593 340924 647829
rect 340604 647509 340924 647593
rect 340604 647273 340646 647509
rect 340882 647273 340924 647509
rect 340604 647241 340924 647273
rect 356076 647829 356396 647861
rect 356076 647593 356118 647829
rect 356354 647593 356396 647829
rect 356076 647509 356396 647593
rect 356076 647273 356118 647509
rect 356354 647273 356396 647509
rect 356076 647241 356396 647273
rect 362340 647829 362660 647861
rect 362340 647593 362382 647829
rect 362618 647593 362660 647829
rect 362340 647509 362660 647593
rect 362340 647273 362382 647509
rect 362618 647273 362660 647509
rect 362340 647241 362660 647273
rect 368604 647829 368924 647861
rect 368604 647593 368646 647829
rect 368882 647593 368924 647829
rect 368604 647509 368924 647593
rect 368604 647273 368646 647509
rect 368882 647273 368924 647509
rect 368604 647241 368924 647273
rect 384076 647829 384396 647861
rect 384076 647593 384118 647829
rect 384354 647593 384396 647829
rect 384076 647509 384396 647593
rect 384076 647273 384118 647509
rect 384354 647273 384396 647509
rect 384076 647241 384396 647273
rect 390340 647829 390660 647861
rect 390340 647593 390382 647829
rect 390618 647593 390660 647829
rect 390340 647509 390660 647593
rect 390340 647273 390382 647509
rect 390618 647273 390660 647509
rect 390340 647241 390660 647273
rect 281472 644454 281792 644486
rect 281472 644218 281514 644454
rect 281750 644218 281792 644454
rect 281472 644134 281792 644218
rect 281472 643898 281514 644134
rect 281750 643898 281792 644134
rect 281472 643866 281792 643898
rect 303208 644454 303528 644486
rect 303208 644218 303250 644454
rect 303486 644218 303528 644454
rect 303208 644134 303528 644218
rect 303208 643898 303250 644134
rect 303486 643898 303528 644134
rect 303208 643866 303528 643898
rect 309472 644454 309792 644486
rect 309472 644218 309514 644454
rect 309750 644218 309792 644454
rect 309472 644134 309792 644218
rect 309472 643898 309514 644134
rect 309750 643898 309792 644134
rect 309472 643866 309792 643898
rect 331208 644454 331528 644486
rect 331208 644218 331250 644454
rect 331486 644218 331528 644454
rect 331208 644134 331528 644218
rect 331208 643898 331250 644134
rect 331486 643898 331528 644134
rect 331208 643866 331528 643898
rect 337472 644454 337792 644486
rect 337472 644218 337514 644454
rect 337750 644218 337792 644454
rect 337472 644134 337792 644218
rect 337472 643898 337514 644134
rect 337750 643898 337792 644134
rect 337472 643866 337792 643898
rect 359208 644454 359528 644486
rect 359208 644218 359250 644454
rect 359486 644218 359528 644454
rect 359208 644134 359528 644218
rect 359208 643898 359250 644134
rect 359486 643898 359528 644134
rect 359208 643866 359528 643898
rect 365472 644454 365792 644486
rect 365472 644218 365514 644454
rect 365750 644218 365792 644454
rect 365472 644134 365792 644218
rect 365472 643898 365514 644134
rect 365750 643898 365792 644134
rect 365472 643866 365792 643898
rect 387208 644454 387528 644486
rect 387208 644218 387250 644454
rect 387486 644218 387528 644454
rect 387208 644134 387528 644218
rect 387208 643898 387250 644134
rect 387486 643898 387528 644134
rect 387208 643866 387528 643898
rect 390878 634813 390938 657323
rect 456379 656028 456445 656029
rect 456379 655964 456380 656028
rect 456444 655964 456445 656028
rect 456379 655963 456445 655964
rect 456382 648277 456442 655963
rect 456379 648276 456445 648277
rect 456379 648212 456380 648276
rect 456444 648212 456445 648276
rect 456379 648211 456445 648212
rect 396604 647829 396924 647861
rect 396604 647593 396646 647829
rect 396882 647593 396924 647829
rect 396604 647509 396924 647593
rect 396604 647273 396646 647509
rect 396882 647273 396924 647509
rect 396604 647241 396924 647273
rect 412076 647829 412396 647861
rect 412076 647593 412118 647829
rect 412354 647593 412396 647829
rect 412076 647509 412396 647593
rect 412076 647273 412118 647509
rect 412354 647273 412396 647509
rect 412076 647241 412396 647273
rect 418340 647829 418660 647861
rect 418340 647593 418382 647829
rect 418618 647593 418660 647829
rect 418340 647509 418660 647593
rect 418340 647273 418382 647509
rect 418618 647273 418660 647509
rect 418340 647241 418660 647273
rect 424604 647829 424924 647861
rect 424604 647593 424646 647829
rect 424882 647593 424924 647829
rect 424604 647509 424924 647593
rect 424604 647273 424646 647509
rect 424882 647273 424924 647509
rect 424604 647241 424924 647273
rect 440076 647829 440396 647861
rect 440076 647593 440118 647829
rect 440354 647593 440396 647829
rect 440076 647509 440396 647593
rect 440076 647273 440118 647509
rect 440354 647273 440396 647509
rect 440076 647241 440396 647273
rect 446340 647829 446660 647861
rect 446340 647593 446382 647829
rect 446618 647593 446660 647829
rect 446340 647509 446660 647593
rect 446340 647273 446382 647509
rect 446618 647273 446660 647509
rect 446340 647241 446660 647273
rect 452604 647829 452924 647861
rect 452604 647593 452646 647829
rect 452882 647593 452924 647829
rect 452604 647509 452924 647593
rect 452604 647273 452646 647509
rect 452882 647273 452924 647509
rect 452604 647241 452924 647273
rect 468076 647829 468396 647861
rect 468076 647593 468118 647829
rect 468354 647593 468396 647829
rect 468076 647509 468396 647593
rect 468076 647273 468118 647509
rect 468354 647273 468396 647509
rect 468076 647241 468396 647273
rect 393472 644454 393792 644486
rect 393472 644218 393514 644454
rect 393750 644218 393792 644454
rect 393472 644134 393792 644218
rect 393472 643898 393514 644134
rect 393750 643898 393792 644134
rect 393472 643866 393792 643898
rect 415208 644454 415528 644486
rect 415208 644218 415250 644454
rect 415486 644218 415528 644454
rect 415208 644134 415528 644218
rect 415208 643898 415250 644134
rect 415486 643898 415528 644134
rect 415208 643866 415528 643898
rect 421472 644454 421792 644486
rect 421472 644218 421514 644454
rect 421750 644218 421792 644454
rect 421472 644134 421792 644218
rect 421472 643898 421514 644134
rect 421750 643898 421792 644134
rect 421472 643866 421792 643898
rect 443208 644454 443528 644486
rect 443208 644218 443250 644454
rect 443486 644218 443528 644454
rect 443208 644134 443528 644218
rect 443208 643898 443250 644134
rect 443486 643898 443528 644134
rect 443208 643866 443528 643898
rect 449472 644454 449792 644486
rect 449472 644218 449514 644454
rect 449750 644218 449792 644454
rect 449472 644134 449792 644218
rect 449472 643898 449514 644134
rect 449750 643898 449792 644134
rect 449472 643866 449792 643898
rect 471208 644454 471528 644486
rect 471208 644218 471250 644454
rect 471486 644218 471528 644454
rect 471208 644134 471528 644218
rect 471208 643898 471250 644134
rect 471486 643898 471528 644134
rect 471208 643866 471528 643898
rect 473494 634813 473554 657323
rect 520227 657252 520293 657253
rect 520227 657188 520228 657252
rect 520292 657188 520293 657252
rect 520227 657187 520293 657188
rect 474340 647829 474660 647861
rect 474340 647593 474382 647829
rect 474618 647593 474660 647829
rect 474340 647509 474660 647593
rect 474340 647273 474382 647509
rect 474618 647273 474660 647509
rect 474340 647241 474660 647273
rect 480604 647829 480924 647861
rect 480604 647593 480646 647829
rect 480882 647593 480924 647829
rect 480604 647509 480924 647593
rect 480604 647273 480646 647509
rect 480882 647273 480924 647509
rect 480604 647241 480924 647273
rect 496076 647829 496396 647861
rect 496076 647593 496118 647829
rect 496354 647593 496396 647829
rect 496076 647509 496396 647593
rect 496076 647273 496118 647509
rect 496354 647273 496396 647509
rect 496076 647241 496396 647273
rect 502340 647829 502660 647861
rect 502340 647593 502382 647829
rect 502618 647593 502660 647829
rect 502340 647509 502660 647593
rect 502340 647273 502382 647509
rect 502618 647273 502660 647509
rect 502340 647241 502660 647273
rect 508604 647829 508924 647861
rect 508604 647593 508646 647829
rect 508882 647593 508924 647829
rect 508604 647509 508924 647593
rect 508604 647273 508646 647509
rect 508882 647273 508924 647509
rect 508604 647241 508924 647273
rect 477472 644454 477792 644486
rect 477472 644218 477514 644454
rect 477750 644218 477792 644454
rect 477472 644134 477792 644218
rect 477472 643898 477514 644134
rect 477750 643898 477792 644134
rect 477472 643866 477792 643898
rect 499208 644454 499528 644486
rect 499208 644218 499250 644454
rect 499486 644218 499528 644454
rect 499208 644134 499528 644218
rect 499208 643898 499250 644134
rect 499486 643898 499528 644134
rect 499208 643866 499528 643898
rect 505472 644454 505792 644486
rect 505472 644218 505514 644454
rect 505750 644218 505792 644454
rect 505472 644134 505792 644218
rect 505472 643898 505514 644134
rect 505750 643898 505792 644134
rect 505472 643866 505792 643898
rect 520230 634813 520290 657187
rect 568435 656028 568501 656029
rect 568435 655964 568436 656028
rect 568500 655964 568501 656028
rect 568435 655963 568501 655964
rect 568438 648277 568498 655963
rect 568435 648276 568501 648277
rect 568435 648212 568436 648276
rect 568500 648212 568501 648276
rect 568435 648211 568501 648212
rect 524076 647829 524396 647861
rect 524076 647593 524118 647829
rect 524354 647593 524396 647829
rect 524076 647509 524396 647593
rect 524076 647273 524118 647509
rect 524354 647273 524396 647509
rect 524076 647241 524396 647273
rect 530340 647829 530660 647861
rect 530340 647593 530382 647829
rect 530618 647593 530660 647829
rect 530340 647509 530660 647593
rect 530340 647273 530382 647509
rect 530618 647273 530660 647509
rect 530340 647241 530660 647273
rect 536604 647829 536924 647861
rect 536604 647593 536646 647829
rect 536882 647593 536924 647829
rect 536604 647509 536924 647593
rect 536604 647273 536646 647509
rect 536882 647273 536924 647509
rect 536604 647241 536924 647273
rect 552076 647829 552396 647861
rect 552076 647593 552118 647829
rect 552354 647593 552396 647829
rect 552076 647509 552396 647593
rect 552076 647273 552118 647509
rect 552354 647273 552396 647509
rect 552076 647241 552396 647273
rect 558340 647829 558660 647861
rect 558340 647593 558382 647829
rect 558618 647593 558660 647829
rect 558340 647509 558660 647593
rect 558340 647273 558382 647509
rect 558618 647273 558660 647509
rect 558340 647241 558660 647273
rect 564604 647829 564924 647861
rect 564604 647593 564646 647829
rect 564882 647593 564924 647829
rect 564604 647509 564924 647593
rect 564604 647273 564646 647509
rect 564882 647273 564924 647509
rect 564604 647241 564924 647273
rect 573494 647829 574114 674273
rect 573494 647593 573526 647829
rect 573762 647593 573846 647829
rect 574082 647593 574114 647829
rect 573494 647509 574114 647593
rect 573494 647273 573526 647509
rect 573762 647273 573846 647509
rect 574082 647273 574114 647509
rect 527208 644454 527528 644486
rect 527208 644218 527250 644454
rect 527486 644218 527528 644454
rect 527208 644134 527528 644218
rect 527208 643898 527250 644134
rect 527486 643898 527528 644134
rect 527208 643866 527528 643898
rect 533472 644454 533792 644486
rect 533472 644218 533514 644454
rect 533750 644218 533792 644454
rect 533472 644134 533792 644218
rect 533472 643898 533514 644134
rect 533750 643898 533792 644134
rect 533472 643866 533792 643898
rect 555208 644454 555528 644486
rect 555208 644218 555250 644454
rect 555486 644218 555528 644454
rect 555208 644134 555528 644218
rect 555208 643898 555250 644134
rect 555486 643898 555528 644134
rect 555208 643866 555528 643898
rect 561472 644454 561792 644486
rect 561472 644218 561514 644454
rect 561750 644218 561792 644454
rect 561472 644134 561792 644218
rect 561472 643898 561514 644134
rect 561750 643898 561792 644134
rect 561472 643866 561792 643898
rect 81387 634812 81453 634813
rect 81387 634748 81388 634812
rect 81452 634748 81453 634812
rect 81387 634747 81453 634748
rect 128307 634812 128373 634813
rect 128307 634748 128308 634812
rect 128372 634748 128373 634812
rect 128307 634747 128373 634748
rect 194731 634812 194797 634813
rect 194731 634748 194732 634812
rect 194796 634748 194797 634812
rect 194731 634747 194797 634748
rect 277163 634812 277229 634813
rect 277163 634748 277164 634812
rect 277228 634748 277229 634812
rect 277163 634747 277229 634748
rect 390875 634812 390941 634813
rect 390875 634748 390876 634812
rect 390940 634748 390941 634812
rect 390875 634747 390941 634748
rect 473491 634812 473557 634813
rect 473491 634748 473492 634812
rect 473556 634748 473557 634812
rect 473491 634747 473557 634748
rect 520227 634812 520293 634813
rect 520227 634748 520228 634812
rect 520292 634748 520293 634812
rect 520227 634747 520293 634748
rect 165659 630460 165725 630461
rect 165659 630396 165660 630460
rect 165724 630396 165725 630460
rect 165659 630395 165725 630396
rect 259499 630460 259565 630461
rect 259499 630396 259500 630460
rect 259564 630396 259565 630460
rect 259499 630395 259565 630396
rect 361619 630460 361685 630461
rect 361619 630396 361620 630460
rect 361684 630396 361685 630460
rect 361619 630395 361685 630396
rect 445707 630460 445773 630461
rect 445707 630396 445708 630460
rect 445772 630396 445773 630460
rect 445707 630395 445773 630396
rect 557579 630460 557645 630461
rect 557579 630396 557580 630460
rect 557644 630396 557645 630460
rect 557579 630395 557645 630396
rect -2006 620593 -1974 620829
rect -1738 620593 -1654 620829
rect -1418 620593 -1386 620829
rect -2006 620509 -1386 620593
rect -2006 620273 -1974 620509
rect -1738 620273 -1654 620509
rect -1418 620273 -1386 620509
rect -2006 593829 -1386 620273
rect 20076 620829 20396 620861
rect 20076 620593 20118 620829
rect 20354 620593 20396 620829
rect 20076 620509 20396 620593
rect 20076 620273 20118 620509
rect 20354 620273 20396 620509
rect 20076 620241 20396 620273
rect 26340 620829 26660 620861
rect 26340 620593 26382 620829
rect 26618 620593 26660 620829
rect 26340 620509 26660 620593
rect 26340 620273 26382 620509
rect 26618 620273 26660 620509
rect 26340 620241 26660 620273
rect 32604 620829 32924 620861
rect 32604 620593 32646 620829
rect 32882 620593 32924 620829
rect 32604 620509 32924 620593
rect 32604 620273 32646 620509
rect 32882 620273 32924 620509
rect 32604 620241 32924 620273
rect 48076 620829 48396 620861
rect 48076 620593 48118 620829
rect 48354 620593 48396 620829
rect 48076 620509 48396 620593
rect 48076 620273 48118 620509
rect 48354 620273 48396 620509
rect 48076 620241 48396 620273
rect 54340 620829 54660 620861
rect 54340 620593 54382 620829
rect 54618 620593 54660 620829
rect 54340 620509 54660 620593
rect 54340 620273 54382 620509
rect 54618 620273 54660 620509
rect 54340 620241 54660 620273
rect 60604 620829 60924 620861
rect 60604 620593 60646 620829
rect 60882 620593 60924 620829
rect 60604 620509 60924 620593
rect 60604 620273 60646 620509
rect 60882 620273 60924 620509
rect 60604 620241 60924 620273
rect 76076 620829 76396 620861
rect 76076 620593 76118 620829
rect 76354 620593 76396 620829
rect 76076 620509 76396 620593
rect 76076 620273 76118 620509
rect 76354 620273 76396 620509
rect 76076 620241 76396 620273
rect 82340 620829 82660 620861
rect 82340 620593 82382 620829
rect 82618 620593 82660 620829
rect 82340 620509 82660 620593
rect 82340 620273 82382 620509
rect 82618 620273 82660 620509
rect 82340 620241 82660 620273
rect 88604 620829 88924 620861
rect 88604 620593 88646 620829
rect 88882 620593 88924 620829
rect 88604 620509 88924 620593
rect 88604 620273 88646 620509
rect 88882 620273 88924 620509
rect 88604 620241 88924 620273
rect 104076 620829 104396 620861
rect 104076 620593 104118 620829
rect 104354 620593 104396 620829
rect 104076 620509 104396 620593
rect 104076 620273 104118 620509
rect 104354 620273 104396 620509
rect 104076 620241 104396 620273
rect 110340 620829 110660 620861
rect 110340 620593 110382 620829
rect 110618 620593 110660 620829
rect 110340 620509 110660 620593
rect 110340 620273 110382 620509
rect 110618 620273 110660 620509
rect 110340 620241 110660 620273
rect 116604 620829 116924 620861
rect 116604 620593 116646 620829
rect 116882 620593 116924 620829
rect 116604 620509 116924 620593
rect 116604 620273 116646 620509
rect 116882 620273 116924 620509
rect 116604 620241 116924 620273
rect 132076 620829 132396 620861
rect 132076 620593 132118 620829
rect 132354 620593 132396 620829
rect 132076 620509 132396 620593
rect 132076 620273 132118 620509
rect 132354 620273 132396 620509
rect 132076 620241 132396 620273
rect 138340 620829 138660 620861
rect 138340 620593 138382 620829
rect 138618 620593 138660 620829
rect 138340 620509 138660 620593
rect 138340 620273 138382 620509
rect 138618 620273 138660 620509
rect 138340 620241 138660 620273
rect 144604 620829 144924 620861
rect 144604 620593 144646 620829
rect 144882 620593 144924 620829
rect 144604 620509 144924 620593
rect 144604 620273 144646 620509
rect 144882 620273 144924 620509
rect 144604 620241 144924 620273
rect 160076 620829 160396 620861
rect 160076 620593 160118 620829
rect 160354 620593 160396 620829
rect 160076 620509 160396 620593
rect 160076 620273 160118 620509
rect 160354 620273 160396 620509
rect 160076 620241 160396 620273
rect 23208 617454 23528 617486
rect 23208 617218 23250 617454
rect 23486 617218 23528 617454
rect 23208 617134 23528 617218
rect 23208 616898 23250 617134
rect 23486 616898 23528 617134
rect 23208 616866 23528 616898
rect 29472 617454 29792 617486
rect 29472 617218 29514 617454
rect 29750 617218 29792 617454
rect 29472 617134 29792 617218
rect 29472 616898 29514 617134
rect 29750 616898 29792 617134
rect 29472 616866 29792 616898
rect 51208 617454 51528 617486
rect 51208 617218 51250 617454
rect 51486 617218 51528 617454
rect 51208 617134 51528 617218
rect 51208 616898 51250 617134
rect 51486 616898 51528 617134
rect 51208 616866 51528 616898
rect 57472 617454 57792 617486
rect 57472 617218 57514 617454
rect 57750 617218 57792 617454
rect 57472 617134 57792 617218
rect 57472 616898 57514 617134
rect 57750 616898 57792 617134
rect 57472 616866 57792 616898
rect 79208 617454 79528 617486
rect 79208 617218 79250 617454
rect 79486 617218 79528 617454
rect 79208 617134 79528 617218
rect 79208 616898 79250 617134
rect 79486 616898 79528 617134
rect 79208 616866 79528 616898
rect 85472 617454 85792 617486
rect 85472 617218 85514 617454
rect 85750 617218 85792 617454
rect 85472 617134 85792 617218
rect 85472 616898 85514 617134
rect 85750 616898 85792 617134
rect 85472 616866 85792 616898
rect 107208 617454 107528 617486
rect 107208 617218 107250 617454
rect 107486 617218 107528 617454
rect 107208 617134 107528 617218
rect 107208 616898 107250 617134
rect 107486 616898 107528 617134
rect 107208 616866 107528 616898
rect 113472 617454 113792 617486
rect 113472 617218 113514 617454
rect 113750 617218 113792 617454
rect 113472 617134 113792 617218
rect 113472 616898 113514 617134
rect 113750 616898 113792 617134
rect 113472 616866 113792 616898
rect 135208 617454 135528 617486
rect 135208 617218 135250 617454
rect 135486 617218 135528 617454
rect 135208 617134 135528 617218
rect 135208 616898 135250 617134
rect 135486 616898 135528 617134
rect 135208 616866 135528 616898
rect 141472 617454 141792 617486
rect 141472 617218 141514 617454
rect 141750 617218 141792 617454
rect 141472 617134 141792 617218
rect 141472 616898 141514 617134
rect 141750 616898 141792 617134
rect 141472 616866 141792 616898
rect 163208 617454 163528 617486
rect 163208 617218 163250 617454
rect 163486 617218 163528 617454
rect 163208 617134 163528 617218
rect 163208 616898 163250 617134
rect 163486 616898 163528 617134
rect 163208 616866 163528 616898
rect 165662 608565 165722 630395
rect 166340 620829 166660 620861
rect 166340 620593 166382 620829
rect 166618 620593 166660 620829
rect 166340 620509 166660 620593
rect 166340 620273 166382 620509
rect 166618 620273 166660 620509
rect 166340 620241 166660 620273
rect 172604 620829 172924 620861
rect 172604 620593 172646 620829
rect 172882 620593 172924 620829
rect 172604 620509 172924 620593
rect 172604 620273 172646 620509
rect 172882 620273 172924 620509
rect 172604 620241 172924 620273
rect 188076 620829 188396 620861
rect 188076 620593 188118 620829
rect 188354 620593 188396 620829
rect 188076 620509 188396 620593
rect 188076 620273 188118 620509
rect 188354 620273 188396 620509
rect 188076 620241 188396 620273
rect 194340 620829 194660 620861
rect 194340 620593 194382 620829
rect 194618 620593 194660 620829
rect 194340 620509 194660 620593
rect 194340 620273 194382 620509
rect 194618 620273 194660 620509
rect 194340 620241 194660 620273
rect 200604 620829 200924 620861
rect 200604 620593 200646 620829
rect 200882 620593 200924 620829
rect 200604 620509 200924 620593
rect 200604 620273 200646 620509
rect 200882 620273 200924 620509
rect 200604 620241 200924 620273
rect 216076 620829 216396 620861
rect 216076 620593 216118 620829
rect 216354 620593 216396 620829
rect 216076 620509 216396 620593
rect 216076 620273 216118 620509
rect 216354 620273 216396 620509
rect 216076 620241 216396 620273
rect 222340 620829 222660 620861
rect 222340 620593 222382 620829
rect 222618 620593 222660 620829
rect 222340 620509 222660 620593
rect 222340 620273 222382 620509
rect 222618 620273 222660 620509
rect 222340 620241 222660 620273
rect 228604 620829 228924 620861
rect 228604 620593 228646 620829
rect 228882 620593 228924 620829
rect 228604 620509 228924 620593
rect 228604 620273 228646 620509
rect 228882 620273 228924 620509
rect 228604 620241 228924 620273
rect 244076 620829 244396 620861
rect 244076 620593 244118 620829
rect 244354 620593 244396 620829
rect 244076 620509 244396 620593
rect 244076 620273 244118 620509
rect 244354 620273 244396 620509
rect 244076 620241 244396 620273
rect 250340 620829 250660 620861
rect 250340 620593 250382 620829
rect 250618 620593 250660 620829
rect 250340 620509 250660 620593
rect 250340 620273 250382 620509
rect 250618 620273 250660 620509
rect 250340 620241 250660 620273
rect 256604 620829 256924 620861
rect 256604 620593 256646 620829
rect 256882 620593 256924 620829
rect 256604 620509 256924 620593
rect 256604 620273 256646 620509
rect 256882 620273 256924 620509
rect 256604 620241 256924 620273
rect 169472 617454 169792 617486
rect 169472 617218 169514 617454
rect 169750 617218 169792 617454
rect 169472 617134 169792 617218
rect 169472 616898 169514 617134
rect 169750 616898 169792 617134
rect 169472 616866 169792 616898
rect 191208 617454 191528 617486
rect 191208 617218 191250 617454
rect 191486 617218 191528 617454
rect 191208 617134 191528 617218
rect 191208 616898 191250 617134
rect 191486 616898 191528 617134
rect 191208 616866 191528 616898
rect 197472 617454 197792 617486
rect 197472 617218 197514 617454
rect 197750 617218 197792 617454
rect 197472 617134 197792 617218
rect 197472 616898 197514 617134
rect 197750 616898 197792 617134
rect 197472 616866 197792 616898
rect 219208 617454 219528 617486
rect 219208 617218 219250 617454
rect 219486 617218 219528 617454
rect 219208 617134 219528 617218
rect 219208 616898 219250 617134
rect 219486 616898 219528 617134
rect 219208 616866 219528 616898
rect 225472 617454 225792 617486
rect 225472 617218 225514 617454
rect 225750 617218 225792 617454
rect 225472 617134 225792 617218
rect 225472 616898 225514 617134
rect 225750 616898 225792 617134
rect 225472 616866 225792 616898
rect 247208 617454 247528 617486
rect 247208 617218 247250 617454
rect 247486 617218 247528 617454
rect 247208 617134 247528 617218
rect 247208 616898 247250 617134
rect 247486 616898 247528 617134
rect 247208 616866 247528 616898
rect 253472 617454 253792 617486
rect 253472 617218 253514 617454
rect 253750 617218 253792 617454
rect 253472 617134 253792 617218
rect 253472 616898 253514 617134
rect 253750 616898 253792 617134
rect 253472 616866 253792 616898
rect 259502 608565 259562 630395
rect 272076 620829 272396 620861
rect 272076 620593 272118 620829
rect 272354 620593 272396 620829
rect 272076 620509 272396 620593
rect 272076 620273 272118 620509
rect 272354 620273 272396 620509
rect 272076 620241 272396 620273
rect 278340 620829 278660 620861
rect 278340 620593 278382 620829
rect 278618 620593 278660 620829
rect 278340 620509 278660 620593
rect 278340 620273 278382 620509
rect 278618 620273 278660 620509
rect 278340 620241 278660 620273
rect 284604 620829 284924 620861
rect 284604 620593 284646 620829
rect 284882 620593 284924 620829
rect 284604 620509 284924 620593
rect 284604 620273 284646 620509
rect 284882 620273 284924 620509
rect 284604 620241 284924 620273
rect 300076 620829 300396 620861
rect 300076 620593 300118 620829
rect 300354 620593 300396 620829
rect 300076 620509 300396 620593
rect 300076 620273 300118 620509
rect 300354 620273 300396 620509
rect 300076 620241 300396 620273
rect 306340 620829 306660 620861
rect 306340 620593 306382 620829
rect 306618 620593 306660 620829
rect 306340 620509 306660 620593
rect 306340 620273 306382 620509
rect 306618 620273 306660 620509
rect 306340 620241 306660 620273
rect 312604 620829 312924 620861
rect 312604 620593 312646 620829
rect 312882 620593 312924 620829
rect 312604 620509 312924 620593
rect 312604 620273 312646 620509
rect 312882 620273 312924 620509
rect 312604 620241 312924 620273
rect 328076 620829 328396 620861
rect 328076 620593 328118 620829
rect 328354 620593 328396 620829
rect 328076 620509 328396 620593
rect 328076 620273 328118 620509
rect 328354 620273 328396 620509
rect 328076 620241 328396 620273
rect 334340 620829 334660 620861
rect 334340 620593 334382 620829
rect 334618 620593 334660 620829
rect 334340 620509 334660 620593
rect 334340 620273 334382 620509
rect 334618 620273 334660 620509
rect 334340 620241 334660 620273
rect 340604 620829 340924 620861
rect 340604 620593 340646 620829
rect 340882 620593 340924 620829
rect 340604 620509 340924 620593
rect 340604 620273 340646 620509
rect 340882 620273 340924 620509
rect 340604 620241 340924 620273
rect 356076 620829 356396 620861
rect 356076 620593 356118 620829
rect 356354 620593 356396 620829
rect 356076 620509 356396 620593
rect 356076 620273 356118 620509
rect 356354 620273 356396 620509
rect 356076 620241 356396 620273
rect 275208 617454 275528 617486
rect 275208 617218 275250 617454
rect 275486 617218 275528 617454
rect 275208 617134 275528 617218
rect 275208 616898 275250 617134
rect 275486 616898 275528 617134
rect 275208 616866 275528 616898
rect 281472 617454 281792 617486
rect 281472 617218 281514 617454
rect 281750 617218 281792 617454
rect 281472 617134 281792 617218
rect 281472 616898 281514 617134
rect 281750 616898 281792 617134
rect 281472 616866 281792 616898
rect 303208 617454 303528 617486
rect 303208 617218 303250 617454
rect 303486 617218 303528 617454
rect 303208 617134 303528 617218
rect 303208 616898 303250 617134
rect 303486 616898 303528 617134
rect 303208 616866 303528 616898
rect 309472 617454 309792 617486
rect 309472 617218 309514 617454
rect 309750 617218 309792 617454
rect 309472 617134 309792 617218
rect 309472 616898 309514 617134
rect 309750 616898 309792 617134
rect 309472 616866 309792 616898
rect 331208 617454 331528 617486
rect 331208 617218 331250 617454
rect 331486 617218 331528 617454
rect 331208 617134 331528 617218
rect 331208 616898 331250 617134
rect 331486 616898 331528 617134
rect 331208 616866 331528 616898
rect 337472 617454 337792 617486
rect 337472 617218 337514 617454
rect 337750 617218 337792 617454
rect 337472 617134 337792 617218
rect 337472 616898 337514 617134
rect 337750 616898 337792 617134
rect 337472 616866 337792 616898
rect 359208 617454 359528 617486
rect 359208 617218 359250 617454
rect 359486 617218 359528 617454
rect 359208 617134 359528 617218
rect 359208 616898 359250 617134
rect 359486 616898 359528 617134
rect 359208 616866 359528 616898
rect 361622 608565 361682 630395
rect 362340 620829 362660 620861
rect 362340 620593 362382 620829
rect 362618 620593 362660 620829
rect 362340 620509 362660 620593
rect 362340 620273 362382 620509
rect 362618 620273 362660 620509
rect 362340 620241 362660 620273
rect 368604 620829 368924 620861
rect 368604 620593 368646 620829
rect 368882 620593 368924 620829
rect 368604 620509 368924 620593
rect 368604 620273 368646 620509
rect 368882 620273 368924 620509
rect 368604 620241 368924 620273
rect 384076 620829 384396 620861
rect 384076 620593 384118 620829
rect 384354 620593 384396 620829
rect 384076 620509 384396 620593
rect 384076 620273 384118 620509
rect 384354 620273 384396 620509
rect 384076 620241 384396 620273
rect 390340 620829 390660 620861
rect 390340 620593 390382 620829
rect 390618 620593 390660 620829
rect 390340 620509 390660 620593
rect 390340 620273 390382 620509
rect 390618 620273 390660 620509
rect 390340 620241 390660 620273
rect 396604 620829 396924 620861
rect 396604 620593 396646 620829
rect 396882 620593 396924 620829
rect 396604 620509 396924 620593
rect 396604 620273 396646 620509
rect 396882 620273 396924 620509
rect 396604 620241 396924 620273
rect 412076 620829 412396 620861
rect 412076 620593 412118 620829
rect 412354 620593 412396 620829
rect 412076 620509 412396 620593
rect 412076 620273 412118 620509
rect 412354 620273 412396 620509
rect 412076 620241 412396 620273
rect 418340 620829 418660 620861
rect 418340 620593 418382 620829
rect 418618 620593 418660 620829
rect 418340 620509 418660 620593
rect 418340 620273 418382 620509
rect 418618 620273 418660 620509
rect 418340 620241 418660 620273
rect 424604 620829 424924 620861
rect 424604 620593 424646 620829
rect 424882 620593 424924 620829
rect 424604 620509 424924 620593
rect 424604 620273 424646 620509
rect 424882 620273 424924 620509
rect 424604 620241 424924 620273
rect 440076 620829 440396 620861
rect 440076 620593 440118 620829
rect 440354 620593 440396 620829
rect 440076 620509 440396 620593
rect 440076 620273 440118 620509
rect 440354 620273 440396 620509
rect 440076 620241 440396 620273
rect 365472 617454 365792 617486
rect 365472 617218 365514 617454
rect 365750 617218 365792 617454
rect 365472 617134 365792 617218
rect 365472 616898 365514 617134
rect 365750 616898 365792 617134
rect 365472 616866 365792 616898
rect 387208 617454 387528 617486
rect 387208 617218 387250 617454
rect 387486 617218 387528 617454
rect 387208 617134 387528 617218
rect 387208 616898 387250 617134
rect 387486 616898 387528 617134
rect 387208 616866 387528 616898
rect 393472 617454 393792 617486
rect 393472 617218 393514 617454
rect 393750 617218 393792 617454
rect 393472 617134 393792 617218
rect 393472 616898 393514 617134
rect 393750 616898 393792 617134
rect 393472 616866 393792 616898
rect 415208 617454 415528 617486
rect 415208 617218 415250 617454
rect 415486 617218 415528 617454
rect 415208 617134 415528 617218
rect 415208 616898 415250 617134
rect 415486 616898 415528 617134
rect 415208 616866 415528 616898
rect 421472 617454 421792 617486
rect 421472 617218 421514 617454
rect 421750 617218 421792 617454
rect 421472 617134 421792 617218
rect 421472 616898 421514 617134
rect 421750 616898 421792 617134
rect 421472 616866 421792 616898
rect 443208 617454 443528 617486
rect 443208 617218 443250 617454
rect 443486 617218 443528 617454
rect 443208 617134 443528 617218
rect 443208 616898 443250 617134
rect 443486 616898 443528 617134
rect 443208 616866 443528 616898
rect 445710 608565 445770 630395
rect 446340 620829 446660 620861
rect 446340 620593 446382 620829
rect 446618 620593 446660 620829
rect 446340 620509 446660 620593
rect 446340 620273 446382 620509
rect 446618 620273 446660 620509
rect 446340 620241 446660 620273
rect 452604 620829 452924 620861
rect 452604 620593 452646 620829
rect 452882 620593 452924 620829
rect 452604 620509 452924 620593
rect 452604 620273 452646 620509
rect 452882 620273 452924 620509
rect 452604 620241 452924 620273
rect 468076 620829 468396 620861
rect 468076 620593 468118 620829
rect 468354 620593 468396 620829
rect 468076 620509 468396 620593
rect 468076 620273 468118 620509
rect 468354 620273 468396 620509
rect 468076 620241 468396 620273
rect 474340 620829 474660 620861
rect 474340 620593 474382 620829
rect 474618 620593 474660 620829
rect 474340 620509 474660 620593
rect 474340 620273 474382 620509
rect 474618 620273 474660 620509
rect 474340 620241 474660 620273
rect 480604 620829 480924 620861
rect 480604 620593 480646 620829
rect 480882 620593 480924 620829
rect 480604 620509 480924 620593
rect 480604 620273 480646 620509
rect 480882 620273 480924 620509
rect 480604 620241 480924 620273
rect 496076 620829 496396 620861
rect 496076 620593 496118 620829
rect 496354 620593 496396 620829
rect 496076 620509 496396 620593
rect 496076 620273 496118 620509
rect 496354 620273 496396 620509
rect 496076 620241 496396 620273
rect 502340 620829 502660 620861
rect 502340 620593 502382 620829
rect 502618 620593 502660 620829
rect 502340 620509 502660 620593
rect 502340 620273 502382 620509
rect 502618 620273 502660 620509
rect 502340 620241 502660 620273
rect 508604 620829 508924 620861
rect 508604 620593 508646 620829
rect 508882 620593 508924 620829
rect 508604 620509 508924 620593
rect 508604 620273 508646 620509
rect 508882 620273 508924 620509
rect 508604 620241 508924 620273
rect 524076 620829 524396 620861
rect 524076 620593 524118 620829
rect 524354 620593 524396 620829
rect 524076 620509 524396 620593
rect 524076 620273 524118 620509
rect 524354 620273 524396 620509
rect 524076 620241 524396 620273
rect 530340 620829 530660 620861
rect 530340 620593 530382 620829
rect 530618 620593 530660 620829
rect 530340 620509 530660 620593
rect 530340 620273 530382 620509
rect 530618 620273 530660 620509
rect 530340 620241 530660 620273
rect 536604 620829 536924 620861
rect 536604 620593 536646 620829
rect 536882 620593 536924 620829
rect 536604 620509 536924 620593
rect 536604 620273 536646 620509
rect 536882 620273 536924 620509
rect 536604 620241 536924 620273
rect 552076 620829 552396 620861
rect 552076 620593 552118 620829
rect 552354 620593 552396 620829
rect 552076 620509 552396 620593
rect 552076 620273 552118 620509
rect 552354 620273 552396 620509
rect 552076 620241 552396 620273
rect 449472 617454 449792 617486
rect 449472 617218 449514 617454
rect 449750 617218 449792 617454
rect 449472 617134 449792 617218
rect 449472 616898 449514 617134
rect 449750 616898 449792 617134
rect 449472 616866 449792 616898
rect 471208 617454 471528 617486
rect 471208 617218 471250 617454
rect 471486 617218 471528 617454
rect 471208 617134 471528 617218
rect 471208 616898 471250 617134
rect 471486 616898 471528 617134
rect 471208 616866 471528 616898
rect 477472 617454 477792 617486
rect 477472 617218 477514 617454
rect 477750 617218 477792 617454
rect 477472 617134 477792 617218
rect 477472 616898 477514 617134
rect 477750 616898 477792 617134
rect 477472 616866 477792 616898
rect 499208 617454 499528 617486
rect 499208 617218 499250 617454
rect 499486 617218 499528 617454
rect 499208 617134 499528 617218
rect 499208 616898 499250 617134
rect 499486 616898 499528 617134
rect 499208 616866 499528 616898
rect 505472 617454 505792 617486
rect 505472 617218 505514 617454
rect 505750 617218 505792 617454
rect 505472 617134 505792 617218
rect 505472 616898 505514 617134
rect 505750 616898 505792 617134
rect 505472 616866 505792 616898
rect 527208 617454 527528 617486
rect 527208 617218 527250 617454
rect 527486 617218 527528 617454
rect 527208 617134 527528 617218
rect 527208 616898 527250 617134
rect 527486 616898 527528 617134
rect 527208 616866 527528 616898
rect 533472 617454 533792 617486
rect 533472 617218 533514 617454
rect 533750 617218 533792 617454
rect 533472 617134 533792 617218
rect 533472 616898 533514 617134
rect 533750 616898 533792 617134
rect 533472 616866 533792 616898
rect 555208 617454 555528 617486
rect 555208 617218 555250 617454
rect 555486 617218 555528 617454
rect 555208 617134 555528 617218
rect 555208 616898 555250 617134
rect 555486 616898 555528 617134
rect 555208 616866 555528 616898
rect 557582 608565 557642 630395
rect 558340 620829 558660 620861
rect 558340 620593 558382 620829
rect 558618 620593 558660 620829
rect 558340 620509 558660 620593
rect 558340 620273 558382 620509
rect 558618 620273 558660 620509
rect 558340 620241 558660 620273
rect 564604 620829 564924 620861
rect 564604 620593 564646 620829
rect 564882 620593 564924 620829
rect 564604 620509 564924 620593
rect 564604 620273 564646 620509
rect 564882 620273 564924 620509
rect 564604 620241 564924 620273
rect 573494 620829 574114 647273
rect 573494 620593 573526 620829
rect 573762 620593 573846 620829
rect 574082 620593 574114 620829
rect 573494 620509 574114 620593
rect 573494 620273 573526 620509
rect 573762 620273 573846 620509
rect 574082 620273 574114 620509
rect 561472 617454 561792 617486
rect 561472 617218 561514 617454
rect 561750 617218 561792 617454
rect 561472 617134 561792 617218
rect 561472 616898 561514 617134
rect 561750 616898 561792 617134
rect 561472 616866 561792 616898
rect 165659 608564 165725 608565
rect 165659 608500 165660 608564
rect 165724 608500 165725 608564
rect 165659 608499 165725 608500
rect 259499 608564 259565 608565
rect 259499 608500 259500 608564
rect 259564 608500 259565 608564
rect 259499 608499 259565 608500
rect 361619 608564 361685 608565
rect 361619 608500 361620 608564
rect 361684 608500 361685 608564
rect 361619 608499 361685 608500
rect 445707 608564 445773 608565
rect 445707 608500 445708 608564
rect 445772 608500 445773 608564
rect 445707 608499 445773 608500
rect 557579 608564 557645 608565
rect 557579 608500 557580 608564
rect 557644 608500 557645 608564
rect 557579 608499 557645 608500
rect 128307 603396 128373 603397
rect 128307 603332 128308 603396
rect 128372 603332 128373 603396
rect 128307 603331 128373 603332
rect 194731 603396 194797 603397
rect 194731 603332 194732 603396
rect 194796 603332 194797 603396
rect 194731 603331 194797 603332
rect 390875 603396 390941 603397
rect 390875 603332 390876 603396
rect 390940 603332 390941 603396
rect 390875 603331 390941 603332
rect 92427 602172 92493 602173
rect 92427 602108 92428 602172
rect 92492 602108 92493 602172
rect 92427 602107 92493 602108
rect 64459 602036 64525 602037
rect 64459 601972 64460 602036
rect 64524 601972 64525 602036
rect 64459 601971 64525 601972
rect 64462 594285 64522 601971
rect 92430 594285 92490 602107
rect 64459 594284 64525 594285
rect 64459 594220 64460 594284
rect 64524 594220 64525 594284
rect 64459 594219 64525 594220
rect 92427 594284 92493 594285
rect 92427 594220 92428 594284
rect 92492 594220 92493 594284
rect 92427 594219 92493 594220
rect -2006 593593 -1974 593829
rect -1738 593593 -1654 593829
rect -1418 593593 -1386 593829
rect -2006 593509 -1386 593593
rect -2006 593273 -1974 593509
rect -1738 593273 -1654 593509
rect -1418 593273 -1386 593509
rect -2006 566829 -1386 593273
rect 20076 593829 20396 593861
rect 20076 593593 20118 593829
rect 20354 593593 20396 593829
rect 20076 593509 20396 593593
rect 20076 593273 20118 593509
rect 20354 593273 20396 593509
rect 20076 593241 20396 593273
rect 26340 593829 26660 593861
rect 26340 593593 26382 593829
rect 26618 593593 26660 593829
rect 26340 593509 26660 593593
rect 26340 593273 26382 593509
rect 26618 593273 26660 593509
rect 26340 593241 26660 593273
rect 32604 593829 32924 593861
rect 32604 593593 32646 593829
rect 32882 593593 32924 593829
rect 32604 593509 32924 593593
rect 32604 593273 32646 593509
rect 32882 593273 32924 593509
rect 32604 593241 32924 593273
rect 48076 593829 48396 593861
rect 48076 593593 48118 593829
rect 48354 593593 48396 593829
rect 48076 593509 48396 593593
rect 48076 593273 48118 593509
rect 48354 593273 48396 593509
rect 48076 593241 48396 593273
rect 54340 593829 54660 593861
rect 54340 593593 54382 593829
rect 54618 593593 54660 593829
rect 54340 593509 54660 593593
rect 54340 593273 54382 593509
rect 54618 593273 54660 593509
rect 54340 593241 54660 593273
rect 60604 593829 60924 593861
rect 60604 593593 60646 593829
rect 60882 593593 60924 593829
rect 60604 593509 60924 593593
rect 60604 593273 60646 593509
rect 60882 593273 60924 593509
rect 60604 593241 60924 593273
rect 76076 593829 76396 593861
rect 76076 593593 76118 593829
rect 76354 593593 76396 593829
rect 76076 593509 76396 593593
rect 76076 593273 76118 593509
rect 76354 593273 76396 593509
rect 76076 593241 76396 593273
rect 82340 593829 82660 593861
rect 82340 593593 82382 593829
rect 82618 593593 82660 593829
rect 82340 593509 82660 593593
rect 82340 593273 82382 593509
rect 82618 593273 82660 593509
rect 82340 593241 82660 593273
rect 88604 593829 88924 593861
rect 88604 593593 88646 593829
rect 88882 593593 88924 593829
rect 88604 593509 88924 593593
rect 88604 593273 88646 593509
rect 88882 593273 88924 593509
rect 88604 593241 88924 593273
rect 104076 593829 104396 593861
rect 104076 593593 104118 593829
rect 104354 593593 104396 593829
rect 104076 593509 104396 593593
rect 104076 593273 104118 593509
rect 104354 593273 104396 593509
rect 104076 593241 104396 593273
rect 110340 593829 110660 593861
rect 110340 593593 110382 593829
rect 110618 593593 110660 593829
rect 110340 593509 110660 593593
rect 110340 593273 110382 593509
rect 110618 593273 110660 593509
rect 110340 593241 110660 593273
rect 116604 593829 116924 593861
rect 116604 593593 116646 593829
rect 116882 593593 116924 593829
rect 116604 593509 116924 593593
rect 116604 593273 116646 593509
rect 116882 593273 116924 593509
rect 116604 593241 116924 593273
rect 23208 590454 23528 590486
rect 23208 590218 23250 590454
rect 23486 590218 23528 590454
rect 23208 590134 23528 590218
rect 23208 589898 23250 590134
rect 23486 589898 23528 590134
rect 23208 589866 23528 589898
rect 29472 590454 29792 590486
rect 29472 590218 29514 590454
rect 29750 590218 29792 590454
rect 29472 590134 29792 590218
rect 29472 589898 29514 590134
rect 29750 589898 29792 590134
rect 29472 589866 29792 589898
rect 51208 590454 51528 590486
rect 51208 590218 51250 590454
rect 51486 590218 51528 590454
rect 51208 590134 51528 590218
rect 51208 589898 51250 590134
rect 51486 589898 51528 590134
rect 51208 589866 51528 589898
rect 57472 590454 57792 590486
rect 57472 590218 57514 590454
rect 57750 590218 57792 590454
rect 57472 590134 57792 590218
rect 57472 589898 57514 590134
rect 57750 589898 57792 590134
rect 57472 589866 57792 589898
rect 79208 590454 79528 590486
rect 79208 590218 79250 590454
rect 79486 590218 79528 590454
rect 79208 590134 79528 590218
rect 79208 589898 79250 590134
rect 79486 589898 79528 590134
rect 79208 589866 79528 589898
rect 85472 590454 85792 590486
rect 85472 590218 85514 590454
rect 85750 590218 85792 590454
rect 85472 590134 85792 590218
rect 85472 589898 85514 590134
rect 85750 589898 85792 590134
rect 85472 589866 85792 589898
rect 107208 590454 107528 590486
rect 107208 590218 107250 590454
rect 107486 590218 107528 590454
rect 107208 590134 107528 590218
rect 107208 589898 107250 590134
rect 107486 589898 107528 590134
rect 107208 589866 107528 589898
rect 113472 590454 113792 590486
rect 113472 590218 113514 590454
rect 113750 590218 113792 590454
rect 113472 590134 113792 590218
rect 113472 589898 113514 590134
rect 113750 589898 113792 590134
rect 113472 589866 113792 589898
rect 128310 582390 128370 603331
rect 148363 602172 148429 602173
rect 148363 602108 148364 602172
rect 148428 602108 148429 602172
rect 148363 602107 148429 602108
rect 148366 594285 148426 602107
rect 176331 602036 176397 602037
rect 176331 601972 176332 602036
rect 176396 601972 176397 602036
rect 176331 601971 176397 601972
rect 176334 594285 176394 601971
rect 148363 594284 148429 594285
rect 148363 594220 148364 594284
rect 148428 594220 148429 594284
rect 148363 594219 148429 594220
rect 176331 594284 176397 594285
rect 176331 594220 176332 594284
rect 176396 594220 176397 594284
rect 176331 594219 176397 594220
rect 132076 593829 132396 593861
rect 132076 593593 132118 593829
rect 132354 593593 132396 593829
rect 132076 593509 132396 593593
rect 132076 593273 132118 593509
rect 132354 593273 132396 593509
rect 132076 593241 132396 593273
rect 138340 593829 138660 593861
rect 138340 593593 138382 593829
rect 138618 593593 138660 593829
rect 138340 593509 138660 593593
rect 138340 593273 138382 593509
rect 138618 593273 138660 593509
rect 138340 593241 138660 593273
rect 144604 593829 144924 593861
rect 144604 593593 144646 593829
rect 144882 593593 144924 593829
rect 144604 593509 144924 593593
rect 144604 593273 144646 593509
rect 144882 593273 144924 593509
rect 144604 593241 144924 593273
rect 160076 593829 160396 593861
rect 160076 593593 160118 593829
rect 160354 593593 160396 593829
rect 160076 593509 160396 593593
rect 160076 593273 160118 593509
rect 160354 593273 160396 593509
rect 160076 593241 160396 593273
rect 166340 593829 166660 593861
rect 166340 593593 166382 593829
rect 166618 593593 166660 593829
rect 166340 593509 166660 593593
rect 166340 593273 166382 593509
rect 166618 593273 166660 593509
rect 166340 593241 166660 593273
rect 172604 593829 172924 593861
rect 172604 593593 172646 593829
rect 172882 593593 172924 593829
rect 172604 593509 172924 593593
rect 172604 593273 172646 593509
rect 172882 593273 172924 593509
rect 172604 593241 172924 593273
rect 188076 593829 188396 593861
rect 188076 593593 188118 593829
rect 188354 593593 188396 593829
rect 188076 593509 188396 593593
rect 188076 593273 188118 593509
rect 188354 593273 188396 593509
rect 188076 593241 188396 593273
rect 194340 593829 194660 593861
rect 194340 593593 194382 593829
rect 194618 593593 194660 593829
rect 194340 593509 194660 593593
rect 194340 593273 194382 593509
rect 194618 593273 194660 593509
rect 194340 593241 194660 593273
rect 135208 590454 135528 590486
rect 135208 590218 135250 590454
rect 135486 590218 135528 590454
rect 135208 590134 135528 590218
rect 135208 589898 135250 590134
rect 135486 589898 135528 590134
rect 135208 589866 135528 589898
rect 141472 590454 141792 590486
rect 141472 590218 141514 590454
rect 141750 590218 141792 590454
rect 141472 590134 141792 590218
rect 141472 589898 141514 590134
rect 141750 589898 141792 590134
rect 141472 589866 141792 589898
rect 163208 590454 163528 590486
rect 163208 590218 163250 590454
rect 163486 590218 163528 590454
rect 163208 590134 163528 590218
rect 163208 589898 163250 590134
rect 163486 589898 163528 590134
rect 163208 589866 163528 589898
rect 169472 590454 169792 590486
rect 169472 590218 169514 590454
rect 169750 590218 169792 590454
rect 169472 590134 169792 590218
rect 169472 589898 169514 590134
rect 169750 589898 169792 590134
rect 169472 589866 169792 589898
rect 191208 590454 191528 590486
rect 191208 590218 191250 590454
rect 191486 590218 191528 590454
rect 191208 590134 191528 590218
rect 191208 589898 191250 590134
rect 191486 589898 191528 590134
rect 191208 589866 191528 589898
rect 128126 582330 128370 582390
rect 128126 580957 128186 582330
rect 194734 580957 194794 603331
rect 288387 602308 288453 602309
rect 288387 602244 288388 602308
rect 288452 602244 288453 602308
rect 288387 602243 288453 602244
rect 260419 602172 260485 602173
rect 260419 602108 260420 602172
rect 260484 602108 260485 602172
rect 260419 602107 260485 602108
rect 260422 594285 260482 602107
rect 288390 594285 288450 602243
rect 344323 602172 344389 602173
rect 344323 602108 344324 602172
rect 344388 602108 344389 602172
rect 344323 602107 344389 602108
rect 344326 594285 344386 602107
rect 372291 602036 372357 602037
rect 372291 601972 372292 602036
rect 372356 601972 372357 602036
rect 372291 601971 372357 601972
rect 372294 594285 372354 601971
rect 260419 594284 260485 594285
rect 260419 594220 260420 594284
rect 260484 594220 260485 594284
rect 260419 594219 260485 594220
rect 288387 594284 288453 594285
rect 288387 594220 288388 594284
rect 288452 594220 288453 594284
rect 288387 594219 288453 594220
rect 344323 594284 344389 594285
rect 344323 594220 344324 594284
rect 344388 594220 344389 594284
rect 344323 594219 344389 594220
rect 372291 594284 372357 594285
rect 372291 594220 372292 594284
rect 372356 594220 372357 594284
rect 372291 594219 372357 594220
rect 200604 593829 200924 593861
rect 200604 593593 200646 593829
rect 200882 593593 200924 593829
rect 200604 593509 200924 593593
rect 200604 593273 200646 593509
rect 200882 593273 200924 593509
rect 200604 593241 200924 593273
rect 216076 593829 216396 593861
rect 216076 593593 216118 593829
rect 216354 593593 216396 593829
rect 216076 593509 216396 593593
rect 216076 593273 216118 593509
rect 216354 593273 216396 593509
rect 216076 593241 216396 593273
rect 222340 593829 222660 593861
rect 222340 593593 222382 593829
rect 222618 593593 222660 593829
rect 222340 593509 222660 593593
rect 222340 593273 222382 593509
rect 222618 593273 222660 593509
rect 222340 593241 222660 593273
rect 228604 593829 228924 593861
rect 228604 593593 228646 593829
rect 228882 593593 228924 593829
rect 228604 593509 228924 593593
rect 228604 593273 228646 593509
rect 228882 593273 228924 593509
rect 228604 593241 228924 593273
rect 244076 593829 244396 593861
rect 244076 593593 244118 593829
rect 244354 593593 244396 593829
rect 244076 593509 244396 593593
rect 244076 593273 244118 593509
rect 244354 593273 244396 593509
rect 244076 593241 244396 593273
rect 250340 593829 250660 593861
rect 250340 593593 250382 593829
rect 250618 593593 250660 593829
rect 250340 593509 250660 593593
rect 250340 593273 250382 593509
rect 250618 593273 250660 593509
rect 250340 593241 250660 593273
rect 256604 593829 256924 593861
rect 256604 593593 256646 593829
rect 256882 593593 256924 593829
rect 256604 593509 256924 593593
rect 256604 593273 256646 593509
rect 256882 593273 256924 593509
rect 256604 593241 256924 593273
rect 272076 593829 272396 593861
rect 272076 593593 272118 593829
rect 272354 593593 272396 593829
rect 272076 593509 272396 593593
rect 272076 593273 272118 593509
rect 272354 593273 272396 593509
rect 272076 593241 272396 593273
rect 278340 593829 278660 593861
rect 278340 593593 278382 593829
rect 278618 593593 278660 593829
rect 278340 593509 278660 593593
rect 278340 593273 278382 593509
rect 278618 593273 278660 593509
rect 278340 593241 278660 593273
rect 284604 593829 284924 593861
rect 284604 593593 284646 593829
rect 284882 593593 284924 593829
rect 284604 593509 284924 593593
rect 284604 593273 284646 593509
rect 284882 593273 284924 593509
rect 284604 593241 284924 593273
rect 300076 593829 300396 593861
rect 300076 593593 300118 593829
rect 300354 593593 300396 593829
rect 300076 593509 300396 593593
rect 300076 593273 300118 593509
rect 300354 593273 300396 593509
rect 300076 593241 300396 593273
rect 306340 593829 306660 593861
rect 306340 593593 306382 593829
rect 306618 593593 306660 593829
rect 306340 593509 306660 593593
rect 306340 593273 306382 593509
rect 306618 593273 306660 593509
rect 306340 593241 306660 593273
rect 312604 593829 312924 593861
rect 312604 593593 312646 593829
rect 312882 593593 312924 593829
rect 312604 593509 312924 593593
rect 312604 593273 312646 593509
rect 312882 593273 312924 593509
rect 312604 593241 312924 593273
rect 328076 593829 328396 593861
rect 328076 593593 328118 593829
rect 328354 593593 328396 593829
rect 328076 593509 328396 593593
rect 328076 593273 328118 593509
rect 328354 593273 328396 593509
rect 328076 593241 328396 593273
rect 334340 593829 334660 593861
rect 334340 593593 334382 593829
rect 334618 593593 334660 593829
rect 334340 593509 334660 593593
rect 334340 593273 334382 593509
rect 334618 593273 334660 593509
rect 334340 593241 334660 593273
rect 340604 593829 340924 593861
rect 340604 593593 340646 593829
rect 340882 593593 340924 593829
rect 340604 593509 340924 593593
rect 340604 593273 340646 593509
rect 340882 593273 340924 593509
rect 340604 593241 340924 593273
rect 356076 593829 356396 593861
rect 356076 593593 356118 593829
rect 356354 593593 356396 593829
rect 356076 593509 356396 593593
rect 356076 593273 356118 593509
rect 356354 593273 356396 593509
rect 356076 593241 356396 593273
rect 362340 593829 362660 593861
rect 362340 593593 362382 593829
rect 362618 593593 362660 593829
rect 362340 593509 362660 593593
rect 362340 593273 362382 593509
rect 362618 593273 362660 593509
rect 362340 593241 362660 593273
rect 368604 593829 368924 593861
rect 368604 593593 368646 593829
rect 368882 593593 368924 593829
rect 368604 593509 368924 593593
rect 368604 593273 368646 593509
rect 368882 593273 368924 593509
rect 368604 593241 368924 593273
rect 384076 593829 384396 593861
rect 384076 593593 384118 593829
rect 384354 593593 384396 593829
rect 384076 593509 384396 593593
rect 384076 593273 384118 593509
rect 384354 593273 384396 593509
rect 384076 593241 384396 593273
rect 390340 593829 390660 593861
rect 390340 593593 390382 593829
rect 390618 593593 390660 593829
rect 390340 593509 390660 593593
rect 390340 593273 390382 593509
rect 390618 593273 390660 593509
rect 390340 593241 390660 593273
rect 197472 590454 197792 590486
rect 197472 590218 197514 590454
rect 197750 590218 197792 590454
rect 197472 590134 197792 590218
rect 197472 589898 197514 590134
rect 197750 589898 197792 590134
rect 197472 589866 197792 589898
rect 219208 590454 219528 590486
rect 219208 590218 219250 590454
rect 219486 590218 219528 590454
rect 219208 590134 219528 590218
rect 219208 589898 219250 590134
rect 219486 589898 219528 590134
rect 219208 589866 219528 589898
rect 225472 590454 225792 590486
rect 225472 590218 225514 590454
rect 225750 590218 225792 590454
rect 225472 590134 225792 590218
rect 225472 589898 225514 590134
rect 225750 589898 225792 590134
rect 225472 589866 225792 589898
rect 247208 590454 247528 590486
rect 247208 590218 247250 590454
rect 247486 590218 247528 590454
rect 247208 590134 247528 590218
rect 247208 589898 247250 590134
rect 247486 589898 247528 590134
rect 247208 589866 247528 589898
rect 253472 590454 253792 590486
rect 253472 590218 253514 590454
rect 253750 590218 253792 590454
rect 253472 590134 253792 590218
rect 253472 589898 253514 590134
rect 253750 589898 253792 590134
rect 253472 589866 253792 589898
rect 275208 590454 275528 590486
rect 275208 590218 275250 590454
rect 275486 590218 275528 590454
rect 275208 590134 275528 590218
rect 275208 589898 275250 590134
rect 275486 589898 275528 590134
rect 275208 589866 275528 589898
rect 281472 590454 281792 590486
rect 281472 590218 281514 590454
rect 281750 590218 281792 590454
rect 281472 590134 281792 590218
rect 281472 589898 281514 590134
rect 281750 589898 281792 590134
rect 281472 589866 281792 589898
rect 303208 590454 303528 590486
rect 303208 590218 303250 590454
rect 303486 590218 303528 590454
rect 303208 590134 303528 590218
rect 303208 589898 303250 590134
rect 303486 589898 303528 590134
rect 303208 589866 303528 589898
rect 309472 590454 309792 590486
rect 309472 590218 309514 590454
rect 309750 590218 309792 590454
rect 309472 590134 309792 590218
rect 309472 589898 309514 590134
rect 309750 589898 309792 590134
rect 309472 589866 309792 589898
rect 331208 590454 331528 590486
rect 331208 590218 331250 590454
rect 331486 590218 331528 590454
rect 331208 590134 331528 590218
rect 331208 589898 331250 590134
rect 331486 589898 331528 590134
rect 331208 589866 331528 589898
rect 337472 590454 337792 590486
rect 337472 590218 337514 590454
rect 337750 590218 337792 590454
rect 337472 590134 337792 590218
rect 337472 589898 337514 590134
rect 337750 589898 337792 590134
rect 337472 589866 337792 589898
rect 359208 590454 359528 590486
rect 359208 590218 359250 590454
rect 359486 590218 359528 590454
rect 359208 590134 359528 590218
rect 359208 589898 359250 590134
rect 359486 589898 359528 590134
rect 359208 589866 359528 589898
rect 365472 590454 365792 590486
rect 365472 590218 365514 590454
rect 365750 590218 365792 590454
rect 365472 590134 365792 590218
rect 365472 589898 365514 590134
rect 365750 589898 365792 590134
rect 365472 589866 365792 589898
rect 387208 590454 387528 590486
rect 387208 590218 387250 590454
rect 387486 590218 387528 590454
rect 387208 590134 387528 590218
rect 387208 589898 387250 590134
rect 387486 589898 387528 590134
rect 387208 589866 387528 589898
rect 390878 580957 390938 603331
rect 484347 602308 484413 602309
rect 484347 602244 484348 602308
rect 484412 602244 484413 602308
rect 484347 602243 484413 602244
rect 456379 602172 456445 602173
rect 456379 602108 456380 602172
rect 456444 602108 456445 602172
rect 456379 602107 456445 602108
rect 456382 594285 456442 602107
rect 484350 594285 484410 602243
rect 492811 602172 492877 602173
rect 492811 602108 492812 602172
rect 492876 602108 492877 602172
rect 492811 602107 492877 602108
rect 492814 596190 492874 602107
rect 520595 602036 520661 602037
rect 520595 601972 520596 602036
rect 520660 601972 520661 602036
rect 520595 601971 520661 601972
rect 492630 596130 492874 596190
rect 492630 594285 492690 596130
rect 520598 594285 520658 601971
rect 456379 594284 456445 594285
rect 456379 594220 456380 594284
rect 456444 594220 456445 594284
rect 456379 594219 456445 594220
rect 484347 594284 484413 594285
rect 484347 594220 484348 594284
rect 484412 594220 484413 594284
rect 484347 594219 484413 594220
rect 492627 594284 492693 594285
rect 492627 594220 492628 594284
rect 492692 594220 492693 594284
rect 492627 594219 492693 594220
rect 520595 594284 520661 594285
rect 520595 594220 520596 594284
rect 520660 594220 520661 594284
rect 520595 594219 520661 594220
rect 396604 593829 396924 593861
rect 396604 593593 396646 593829
rect 396882 593593 396924 593829
rect 396604 593509 396924 593593
rect 396604 593273 396646 593509
rect 396882 593273 396924 593509
rect 396604 593241 396924 593273
rect 412076 593829 412396 593861
rect 412076 593593 412118 593829
rect 412354 593593 412396 593829
rect 412076 593509 412396 593593
rect 412076 593273 412118 593509
rect 412354 593273 412396 593509
rect 412076 593241 412396 593273
rect 418340 593829 418660 593861
rect 418340 593593 418382 593829
rect 418618 593593 418660 593829
rect 418340 593509 418660 593593
rect 418340 593273 418382 593509
rect 418618 593273 418660 593509
rect 418340 593241 418660 593273
rect 424604 593829 424924 593861
rect 424604 593593 424646 593829
rect 424882 593593 424924 593829
rect 424604 593509 424924 593593
rect 424604 593273 424646 593509
rect 424882 593273 424924 593509
rect 424604 593241 424924 593273
rect 440076 593829 440396 593861
rect 440076 593593 440118 593829
rect 440354 593593 440396 593829
rect 440076 593509 440396 593593
rect 440076 593273 440118 593509
rect 440354 593273 440396 593509
rect 440076 593241 440396 593273
rect 446340 593829 446660 593861
rect 446340 593593 446382 593829
rect 446618 593593 446660 593829
rect 446340 593509 446660 593593
rect 446340 593273 446382 593509
rect 446618 593273 446660 593509
rect 446340 593241 446660 593273
rect 452604 593829 452924 593861
rect 452604 593593 452646 593829
rect 452882 593593 452924 593829
rect 452604 593509 452924 593593
rect 452604 593273 452646 593509
rect 452882 593273 452924 593509
rect 452604 593241 452924 593273
rect 468076 593829 468396 593861
rect 468076 593593 468118 593829
rect 468354 593593 468396 593829
rect 468076 593509 468396 593593
rect 468076 593273 468118 593509
rect 468354 593273 468396 593509
rect 468076 593241 468396 593273
rect 474340 593829 474660 593861
rect 474340 593593 474382 593829
rect 474618 593593 474660 593829
rect 474340 593509 474660 593593
rect 474340 593273 474382 593509
rect 474618 593273 474660 593509
rect 474340 593241 474660 593273
rect 480604 593829 480924 593861
rect 480604 593593 480646 593829
rect 480882 593593 480924 593829
rect 480604 593509 480924 593593
rect 480604 593273 480646 593509
rect 480882 593273 480924 593509
rect 480604 593241 480924 593273
rect 496076 593829 496396 593861
rect 496076 593593 496118 593829
rect 496354 593593 496396 593829
rect 496076 593509 496396 593593
rect 496076 593273 496118 593509
rect 496354 593273 496396 593509
rect 496076 593241 496396 593273
rect 502340 593829 502660 593861
rect 502340 593593 502382 593829
rect 502618 593593 502660 593829
rect 502340 593509 502660 593593
rect 502340 593273 502382 593509
rect 502618 593273 502660 593509
rect 502340 593241 502660 593273
rect 508604 593829 508924 593861
rect 508604 593593 508646 593829
rect 508882 593593 508924 593829
rect 508604 593509 508924 593593
rect 508604 593273 508646 593509
rect 508882 593273 508924 593509
rect 508604 593241 508924 593273
rect 524076 593829 524396 593861
rect 524076 593593 524118 593829
rect 524354 593593 524396 593829
rect 524076 593509 524396 593593
rect 524076 593273 524118 593509
rect 524354 593273 524396 593509
rect 524076 593241 524396 593273
rect 530340 593829 530660 593861
rect 530340 593593 530382 593829
rect 530618 593593 530660 593829
rect 530340 593509 530660 593593
rect 530340 593273 530382 593509
rect 530618 593273 530660 593509
rect 530340 593241 530660 593273
rect 536604 593829 536924 593861
rect 536604 593593 536646 593829
rect 536882 593593 536924 593829
rect 536604 593509 536924 593593
rect 536604 593273 536646 593509
rect 536882 593273 536924 593509
rect 536604 593241 536924 593273
rect 552076 593829 552396 593861
rect 552076 593593 552118 593829
rect 552354 593593 552396 593829
rect 552076 593509 552396 593593
rect 552076 593273 552118 593509
rect 552354 593273 552396 593509
rect 552076 593241 552396 593273
rect 558340 593829 558660 593861
rect 558340 593593 558382 593829
rect 558618 593593 558660 593829
rect 558340 593509 558660 593593
rect 558340 593273 558382 593509
rect 558618 593273 558660 593509
rect 558340 593241 558660 593273
rect 564604 593829 564924 593861
rect 564604 593593 564646 593829
rect 564882 593593 564924 593829
rect 564604 593509 564924 593593
rect 564604 593273 564646 593509
rect 564882 593273 564924 593509
rect 564604 593241 564924 593273
rect 573494 593829 574114 620273
rect 573494 593593 573526 593829
rect 573762 593593 573846 593829
rect 574082 593593 574114 593829
rect 573494 593509 574114 593593
rect 573494 593273 573526 593509
rect 573762 593273 573846 593509
rect 574082 593273 574114 593509
rect 393472 590454 393792 590486
rect 393472 590218 393514 590454
rect 393750 590218 393792 590454
rect 393472 590134 393792 590218
rect 393472 589898 393514 590134
rect 393750 589898 393792 590134
rect 393472 589866 393792 589898
rect 415208 590454 415528 590486
rect 415208 590218 415250 590454
rect 415486 590218 415528 590454
rect 415208 590134 415528 590218
rect 415208 589898 415250 590134
rect 415486 589898 415528 590134
rect 415208 589866 415528 589898
rect 421472 590454 421792 590486
rect 421472 590218 421514 590454
rect 421750 590218 421792 590454
rect 421472 590134 421792 590218
rect 421472 589898 421514 590134
rect 421750 589898 421792 590134
rect 421472 589866 421792 589898
rect 443208 590454 443528 590486
rect 443208 590218 443250 590454
rect 443486 590218 443528 590454
rect 443208 590134 443528 590218
rect 443208 589898 443250 590134
rect 443486 589898 443528 590134
rect 443208 589866 443528 589898
rect 449472 590454 449792 590486
rect 449472 590218 449514 590454
rect 449750 590218 449792 590454
rect 449472 590134 449792 590218
rect 449472 589898 449514 590134
rect 449750 589898 449792 590134
rect 449472 589866 449792 589898
rect 471208 590454 471528 590486
rect 471208 590218 471250 590454
rect 471486 590218 471528 590454
rect 471208 590134 471528 590218
rect 471208 589898 471250 590134
rect 471486 589898 471528 590134
rect 471208 589866 471528 589898
rect 477472 590454 477792 590486
rect 477472 590218 477514 590454
rect 477750 590218 477792 590454
rect 477472 590134 477792 590218
rect 477472 589898 477514 590134
rect 477750 589898 477792 590134
rect 477472 589866 477792 589898
rect 499208 590454 499528 590486
rect 499208 590218 499250 590454
rect 499486 590218 499528 590454
rect 499208 590134 499528 590218
rect 499208 589898 499250 590134
rect 499486 589898 499528 590134
rect 499208 589866 499528 589898
rect 505472 590454 505792 590486
rect 505472 590218 505514 590454
rect 505750 590218 505792 590454
rect 505472 590134 505792 590218
rect 505472 589898 505514 590134
rect 505750 589898 505792 590134
rect 505472 589866 505792 589898
rect 527208 590454 527528 590486
rect 527208 590218 527250 590454
rect 527486 590218 527528 590454
rect 527208 590134 527528 590218
rect 527208 589898 527250 590134
rect 527486 589898 527528 590134
rect 527208 589866 527528 589898
rect 533472 590454 533792 590486
rect 533472 590218 533514 590454
rect 533750 590218 533792 590454
rect 533472 590134 533792 590218
rect 533472 589898 533514 590134
rect 533750 589898 533792 590134
rect 533472 589866 533792 589898
rect 555208 590454 555528 590486
rect 555208 590218 555250 590454
rect 555486 590218 555528 590454
rect 555208 590134 555528 590218
rect 555208 589898 555250 590134
rect 555486 589898 555528 590134
rect 555208 589866 555528 589898
rect 561472 590454 561792 590486
rect 561472 590218 561514 590454
rect 561750 590218 561792 590454
rect 561472 590134 561792 590218
rect 561472 589898 561514 590134
rect 561750 589898 561792 590134
rect 561472 589866 561792 589898
rect 128123 580956 128189 580957
rect 128123 580892 128124 580956
rect 128188 580892 128189 580956
rect 128123 580891 128189 580892
rect 194731 580956 194797 580957
rect 194731 580892 194732 580956
rect 194796 580892 194797 580956
rect 194731 580891 194797 580892
rect 390875 580956 390941 580957
rect 390875 580892 390876 580956
rect 390940 580892 390941 580956
rect 390875 580891 390941 580892
rect 165659 576468 165725 576469
rect 165659 576404 165660 576468
rect 165724 576404 165725 576468
rect 165659 576403 165725 576404
rect 259499 576468 259565 576469
rect 259499 576404 259500 576468
rect 259564 576404 259565 576468
rect 259499 576403 259565 576404
rect 361619 576468 361685 576469
rect 361619 576404 361620 576468
rect 361684 576404 361685 576468
rect 361619 576403 361685 576404
rect 445707 576468 445773 576469
rect 445707 576404 445708 576468
rect 445772 576404 445773 576468
rect 445707 576403 445773 576404
rect 557579 576468 557645 576469
rect 557579 576404 557580 576468
rect 557644 576404 557645 576468
rect 557579 576403 557645 576404
rect -2006 566593 -1974 566829
rect -1738 566593 -1654 566829
rect -1418 566593 -1386 566829
rect -2006 566509 -1386 566593
rect -2006 566273 -1974 566509
rect -1738 566273 -1654 566509
rect -1418 566273 -1386 566509
rect -2006 539829 -1386 566273
rect 20076 566829 20396 566861
rect 20076 566593 20118 566829
rect 20354 566593 20396 566829
rect 20076 566509 20396 566593
rect 20076 566273 20118 566509
rect 20354 566273 20396 566509
rect 20076 566241 20396 566273
rect 26340 566829 26660 566861
rect 26340 566593 26382 566829
rect 26618 566593 26660 566829
rect 26340 566509 26660 566593
rect 26340 566273 26382 566509
rect 26618 566273 26660 566509
rect 26340 566241 26660 566273
rect 32604 566829 32924 566861
rect 32604 566593 32646 566829
rect 32882 566593 32924 566829
rect 32604 566509 32924 566593
rect 32604 566273 32646 566509
rect 32882 566273 32924 566509
rect 32604 566241 32924 566273
rect 48076 566829 48396 566861
rect 48076 566593 48118 566829
rect 48354 566593 48396 566829
rect 48076 566509 48396 566593
rect 48076 566273 48118 566509
rect 48354 566273 48396 566509
rect 48076 566241 48396 566273
rect 54340 566829 54660 566861
rect 54340 566593 54382 566829
rect 54618 566593 54660 566829
rect 54340 566509 54660 566593
rect 54340 566273 54382 566509
rect 54618 566273 54660 566509
rect 54340 566241 54660 566273
rect 60604 566829 60924 566861
rect 60604 566593 60646 566829
rect 60882 566593 60924 566829
rect 60604 566509 60924 566593
rect 60604 566273 60646 566509
rect 60882 566273 60924 566509
rect 60604 566241 60924 566273
rect 76076 566829 76396 566861
rect 76076 566593 76118 566829
rect 76354 566593 76396 566829
rect 76076 566509 76396 566593
rect 76076 566273 76118 566509
rect 76354 566273 76396 566509
rect 76076 566241 76396 566273
rect 82340 566829 82660 566861
rect 82340 566593 82382 566829
rect 82618 566593 82660 566829
rect 82340 566509 82660 566593
rect 82340 566273 82382 566509
rect 82618 566273 82660 566509
rect 82340 566241 82660 566273
rect 88604 566829 88924 566861
rect 88604 566593 88646 566829
rect 88882 566593 88924 566829
rect 88604 566509 88924 566593
rect 88604 566273 88646 566509
rect 88882 566273 88924 566509
rect 88604 566241 88924 566273
rect 104076 566829 104396 566861
rect 104076 566593 104118 566829
rect 104354 566593 104396 566829
rect 104076 566509 104396 566593
rect 104076 566273 104118 566509
rect 104354 566273 104396 566509
rect 104076 566241 104396 566273
rect 110340 566829 110660 566861
rect 110340 566593 110382 566829
rect 110618 566593 110660 566829
rect 110340 566509 110660 566593
rect 110340 566273 110382 566509
rect 110618 566273 110660 566509
rect 110340 566241 110660 566273
rect 116604 566829 116924 566861
rect 116604 566593 116646 566829
rect 116882 566593 116924 566829
rect 116604 566509 116924 566593
rect 116604 566273 116646 566509
rect 116882 566273 116924 566509
rect 116604 566241 116924 566273
rect 132076 566829 132396 566861
rect 132076 566593 132118 566829
rect 132354 566593 132396 566829
rect 132076 566509 132396 566593
rect 132076 566273 132118 566509
rect 132354 566273 132396 566509
rect 132076 566241 132396 566273
rect 138340 566829 138660 566861
rect 138340 566593 138382 566829
rect 138618 566593 138660 566829
rect 138340 566509 138660 566593
rect 138340 566273 138382 566509
rect 138618 566273 138660 566509
rect 138340 566241 138660 566273
rect 144604 566829 144924 566861
rect 144604 566593 144646 566829
rect 144882 566593 144924 566829
rect 144604 566509 144924 566593
rect 144604 566273 144646 566509
rect 144882 566273 144924 566509
rect 144604 566241 144924 566273
rect 160076 566829 160396 566861
rect 160076 566593 160118 566829
rect 160354 566593 160396 566829
rect 160076 566509 160396 566593
rect 160076 566273 160118 566509
rect 160354 566273 160396 566509
rect 160076 566241 160396 566273
rect 23208 563454 23528 563486
rect 23208 563218 23250 563454
rect 23486 563218 23528 563454
rect 23208 563134 23528 563218
rect 23208 562898 23250 563134
rect 23486 562898 23528 563134
rect 23208 562866 23528 562898
rect 29472 563454 29792 563486
rect 29472 563218 29514 563454
rect 29750 563218 29792 563454
rect 29472 563134 29792 563218
rect 29472 562898 29514 563134
rect 29750 562898 29792 563134
rect 29472 562866 29792 562898
rect 51208 563454 51528 563486
rect 51208 563218 51250 563454
rect 51486 563218 51528 563454
rect 51208 563134 51528 563218
rect 51208 562898 51250 563134
rect 51486 562898 51528 563134
rect 51208 562866 51528 562898
rect 57472 563454 57792 563486
rect 57472 563218 57514 563454
rect 57750 563218 57792 563454
rect 57472 563134 57792 563218
rect 57472 562898 57514 563134
rect 57750 562898 57792 563134
rect 57472 562866 57792 562898
rect 79208 563454 79528 563486
rect 79208 563218 79250 563454
rect 79486 563218 79528 563454
rect 79208 563134 79528 563218
rect 79208 562898 79250 563134
rect 79486 562898 79528 563134
rect 79208 562866 79528 562898
rect 85472 563454 85792 563486
rect 85472 563218 85514 563454
rect 85750 563218 85792 563454
rect 85472 563134 85792 563218
rect 85472 562898 85514 563134
rect 85750 562898 85792 563134
rect 85472 562866 85792 562898
rect 107208 563454 107528 563486
rect 107208 563218 107250 563454
rect 107486 563218 107528 563454
rect 107208 563134 107528 563218
rect 107208 562898 107250 563134
rect 107486 562898 107528 563134
rect 107208 562866 107528 562898
rect 113472 563454 113792 563486
rect 113472 563218 113514 563454
rect 113750 563218 113792 563454
rect 113472 563134 113792 563218
rect 113472 562898 113514 563134
rect 113750 562898 113792 563134
rect 113472 562866 113792 562898
rect 135208 563454 135528 563486
rect 135208 563218 135250 563454
rect 135486 563218 135528 563454
rect 135208 563134 135528 563218
rect 135208 562898 135250 563134
rect 135486 562898 135528 563134
rect 135208 562866 135528 562898
rect 141472 563454 141792 563486
rect 141472 563218 141514 563454
rect 141750 563218 141792 563454
rect 141472 563134 141792 563218
rect 141472 562898 141514 563134
rect 141750 562898 141792 563134
rect 141472 562866 141792 562898
rect 163208 563454 163528 563486
rect 163208 563218 163250 563454
rect 163486 563218 163528 563454
rect 163208 563134 163528 563218
rect 163208 562898 163250 563134
rect 163486 562898 163528 563134
rect 163208 562866 163528 562898
rect 165662 554709 165722 576403
rect 166340 566829 166660 566861
rect 166340 566593 166382 566829
rect 166618 566593 166660 566829
rect 166340 566509 166660 566593
rect 166340 566273 166382 566509
rect 166618 566273 166660 566509
rect 166340 566241 166660 566273
rect 172604 566829 172924 566861
rect 172604 566593 172646 566829
rect 172882 566593 172924 566829
rect 172604 566509 172924 566593
rect 172604 566273 172646 566509
rect 172882 566273 172924 566509
rect 172604 566241 172924 566273
rect 188076 566829 188396 566861
rect 188076 566593 188118 566829
rect 188354 566593 188396 566829
rect 188076 566509 188396 566593
rect 188076 566273 188118 566509
rect 188354 566273 188396 566509
rect 188076 566241 188396 566273
rect 194340 566829 194660 566861
rect 194340 566593 194382 566829
rect 194618 566593 194660 566829
rect 194340 566509 194660 566593
rect 194340 566273 194382 566509
rect 194618 566273 194660 566509
rect 194340 566241 194660 566273
rect 200604 566829 200924 566861
rect 200604 566593 200646 566829
rect 200882 566593 200924 566829
rect 200604 566509 200924 566593
rect 200604 566273 200646 566509
rect 200882 566273 200924 566509
rect 200604 566241 200924 566273
rect 216076 566829 216396 566861
rect 216076 566593 216118 566829
rect 216354 566593 216396 566829
rect 216076 566509 216396 566593
rect 216076 566273 216118 566509
rect 216354 566273 216396 566509
rect 216076 566241 216396 566273
rect 222340 566829 222660 566861
rect 222340 566593 222382 566829
rect 222618 566593 222660 566829
rect 222340 566509 222660 566593
rect 222340 566273 222382 566509
rect 222618 566273 222660 566509
rect 222340 566241 222660 566273
rect 228604 566829 228924 566861
rect 228604 566593 228646 566829
rect 228882 566593 228924 566829
rect 228604 566509 228924 566593
rect 228604 566273 228646 566509
rect 228882 566273 228924 566509
rect 228604 566241 228924 566273
rect 244076 566829 244396 566861
rect 244076 566593 244118 566829
rect 244354 566593 244396 566829
rect 244076 566509 244396 566593
rect 244076 566273 244118 566509
rect 244354 566273 244396 566509
rect 244076 566241 244396 566273
rect 250340 566829 250660 566861
rect 250340 566593 250382 566829
rect 250618 566593 250660 566829
rect 250340 566509 250660 566593
rect 250340 566273 250382 566509
rect 250618 566273 250660 566509
rect 250340 566241 250660 566273
rect 256604 566829 256924 566861
rect 256604 566593 256646 566829
rect 256882 566593 256924 566829
rect 256604 566509 256924 566593
rect 256604 566273 256646 566509
rect 256882 566273 256924 566509
rect 256604 566241 256924 566273
rect 169472 563454 169792 563486
rect 169472 563218 169514 563454
rect 169750 563218 169792 563454
rect 169472 563134 169792 563218
rect 169472 562898 169514 563134
rect 169750 562898 169792 563134
rect 169472 562866 169792 562898
rect 191208 563454 191528 563486
rect 191208 563218 191250 563454
rect 191486 563218 191528 563454
rect 191208 563134 191528 563218
rect 191208 562898 191250 563134
rect 191486 562898 191528 563134
rect 191208 562866 191528 562898
rect 197472 563454 197792 563486
rect 197472 563218 197514 563454
rect 197750 563218 197792 563454
rect 197472 563134 197792 563218
rect 197472 562898 197514 563134
rect 197750 562898 197792 563134
rect 197472 562866 197792 562898
rect 219208 563454 219528 563486
rect 219208 563218 219250 563454
rect 219486 563218 219528 563454
rect 219208 563134 219528 563218
rect 219208 562898 219250 563134
rect 219486 562898 219528 563134
rect 219208 562866 219528 562898
rect 225472 563454 225792 563486
rect 225472 563218 225514 563454
rect 225750 563218 225792 563454
rect 225472 563134 225792 563218
rect 225472 562898 225514 563134
rect 225750 562898 225792 563134
rect 225472 562866 225792 562898
rect 247208 563454 247528 563486
rect 247208 563218 247250 563454
rect 247486 563218 247528 563454
rect 247208 563134 247528 563218
rect 247208 562898 247250 563134
rect 247486 562898 247528 563134
rect 247208 562866 247528 562898
rect 253472 563454 253792 563486
rect 253472 563218 253514 563454
rect 253750 563218 253792 563454
rect 253472 563134 253792 563218
rect 253472 562898 253514 563134
rect 253750 562898 253792 563134
rect 253472 562866 253792 562898
rect 259502 554709 259562 576403
rect 272076 566829 272396 566861
rect 272076 566593 272118 566829
rect 272354 566593 272396 566829
rect 272076 566509 272396 566593
rect 272076 566273 272118 566509
rect 272354 566273 272396 566509
rect 272076 566241 272396 566273
rect 278340 566829 278660 566861
rect 278340 566593 278382 566829
rect 278618 566593 278660 566829
rect 278340 566509 278660 566593
rect 278340 566273 278382 566509
rect 278618 566273 278660 566509
rect 278340 566241 278660 566273
rect 284604 566829 284924 566861
rect 284604 566593 284646 566829
rect 284882 566593 284924 566829
rect 284604 566509 284924 566593
rect 284604 566273 284646 566509
rect 284882 566273 284924 566509
rect 284604 566241 284924 566273
rect 300076 566829 300396 566861
rect 300076 566593 300118 566829
rect 300354 566593 300396 566829
rect 300076 566509 300396 566593
rect 300076 566273 300118 566509
rect 300354 566273 300396 566509
rect 300076 566241 300396 566273
rect 306340 566829 306660 566861
rect 306340 566593 306382 566829
rect 306618 566593 306660 566829
rect 306340 566509 306660 566593
rect 306340 566273 306382 566509
rect 306618 566273 306660 566509
rect 306340 566241 306660 566273
rect 312604 566829 312924 566861
rect 312604 566593 312646 566829
rect 312882 566593 312924 566829
rect 312604 566509 312924 566593
rect 312604 566273 312646 566509
rect 312882 566273 312924 566509
rect 312604 566241 312924 566273
rect 328076 566829 328396 566861
rect 328076 566593 328118 566829
rect 328354 566593 328396 566829
rect 328076 566509 328396 566593
rect 328076 566273 328118 566509
rect 328354 566273 328396 566509
rect 328076 566241 328396 566273
rect 334340 566829 334660 566861
rect 334340 566593 334382 566829
rect 334618 566593 334660 566829
rect 334340 566509 334660 566593
rect 334340 566273 334382 566509
rect 334618 566273 334660 566509
rect 334340 566241 334660 566273
rect 340604 566829 340924 566861
rect 340604 566593 340646 566829
rect 340882 566593 340924 566829
rect 340604 566509 340924 566593
rect 340604 566273 340646 566509
rect 340882 566273 340924 566509
rect 340604 566241 340924 566273
rect 356076 566829 356396 566861
rect 356076 566593 356118 566829
rect 356354 566593 356396 566829
rect 356076 566509 356396 566593
rect 356076 566273 356118 566509
rect 356354 566273 356396 566509
rect 356076 566241 356396 566273
rect 275208 563454 275528 563486
rect 275208 563218 275250 563454
rect 275486 563218 275528 563454
rect 275208 563134 275528 563218
rect 275208 562898 275250 563134
rect 275486 562898 275528 563134
rect 275208 562866 275528 562898
rect 281472 563454 281792 563486
rect 281472 563218 281514 563454
rect 281750 563218 281792 563454
rect 281472 563134 281792 563218
rect 281472 562898 281514 563134
rect 281750 562898 281792 563134
rect 281472 562866 281792 562898
rect 303208 563454 303528 563486
rect 303208 563218 303250 563454
rect 303486 563218 303528 563454
rect 303208 563134 303528 563218
rect 303208 562898 303250 563134
rect 303486 562898 303528 563134
rect 303208 562866 303528 562898
rect 309472 563454 309792 563486
rect 309472 563218 309514 563454
rect 309750 563218 309792 563454
rect 309472 563134 309792 563218
rect 309472 562898 309514 563134
rect 309750 562898 309792 563134
rect 309472 562866 309792 562898
rect 331208 563454 331528 563486
rect 331208 563218 331250 563454
rect 331486 563218 331528 563454
rect 331208 563134 331528 563218
rect 331208 562898 331250 563134
rect 331486 562898 331528 563134
rect 331208 562866 331528 562898
rect 337472 563454 337792 563486
rect 337472 563218 337514 563454
rect 337750 563218 337792 563454
rect 337472 563134 337792 563218
rect 337472 562898 337514 563134
rect 337750 562898 337792 563134
rect 337472 562866 337792 562898
rect 359208 563454 359528 563486
rect 359208 563218 359250 563454
rect 359486 563218 359528 563454
rect 359208 563134 359528 563218
rect 359208 562898 359250 563134
rect 359486 562898 359528 563134
rect 359208 562866 359528 562898
rect 361622 554709 361682 576403
rect 362340 566829 362660 566861
rect 362340 566593 362382 566829
rect 362618 566593 362660 566829
rect 362340 566509 362660 566593
rect 362340 566273 362382 566509
rect 362618 566273 362660 566509
rect 362340 566241 362660 566273
rect 368604 566829 368924 566861
rect 368604 566593 368646 566829
rect 368882 566593 368924 566829
rect 368604 566509 368924 566593
rect 368604 566273 368646 566509
rect 368882 566273 368924 566509
rect 368604 566241 368924 566273
rect 384076 566829 384396 566861
rect 384076 566593 384118 566829
rect 384354 566593 384396 566829
rect 384076 566509 384396 566593
rect 384076 566273 384118 566509
rect 384354 566273 384396 566509
rect 384076 566241 384396 566273
rect 390340 566829 390660 566861
rect 390340 566593 390382 566829
rect 390618 566593 390660 566829
rect 390340 566509 390660 566593
rect 390340 566273 390382 566509
rect 390618 566273 390660 566509
rect 390340 566241 390660 566273
rect 396604 566829 396924 566861
rect 396604 566593 396646 566829
rect 396882 566593 396924 566829
rect 396604 566509 396924 566593
rect 396604 566273 396646 566509
rect 396882 566273 396924 566509
rect 396604 566241 396924 566273
rect 412076 566829 412396 566861
rect 412076 566593 412118 566829
rect 412354 566593 412396 566829
rect 412076 566509 412396 566593
rect 412076 566273 412118 566509
rect 412354 566273 412396 566509
rect 412076 566241 412396 566273
rect 418340 566829 418660 566861
rect 418340 566593 418382 566829
rect 418618 566593 418660 566829
rect 418340 566509 418660 566593
rect 418340 566273 418382 566509
rect 418618 566273 418660 566509
rect 418340 566241 418660 566273
rect 424604 566829 424924 566861
rect 424604 566593 424646 566829
rect 424882 566593 424924 566829
rect 424604 566509 424924 566593
rect 424604 566273 424646 566509
rect 424882 566273 424924 566509
rect 424604 566241 424924 566273
rect 440076 566829 440396 566861
rect 440076 566593 440118 566829
rect 440354 566593 440396 566829
rect 440076 566509 440396 566593
rect 440076 566273 440118 566509
rect 440354 566273 440396 566509
rect 440076 566241 440396 566273
rect 365472 563454 365792 563486
rect 365472 563218 365514 563454
rect 365750 563218 365792 563454
rect 365472 563134 365792 563218
rect 365472 562898 365514 563134
rect 365750 562898 365792 563134
rect 365472 562866 365792 562898
rect 387208 563454 387528 563486
rect 387208 563218 387250 563454
rect 387486 563218 387528 563454
rect 387208 563134 387528 563218
rect 387208 562898 387250 563134
rect 387486 562898 387528 563134
rect 387208 562866 387528 562898
rect 393472 563454 393792 563486
rect 393472 563218 393514 563454
rect 393750 563218 393792 563454
rect 393472 563134 393792 563218
rect 393472 562898 393514 563134
rect 393750 562898 393792 563134
rect 393472 562866 393792 562898
rect 415208 563454 415528 563486
rect 415208 563218 415250 563454
rect 415486 563218 415528 563454
rect 415208 563134 415528 563218
rect 415208 562898 415250 563134
rect 415486 562898 415528 563134
rect 415208 562866 415528 562898
rect 421472 563454 421792 563486
rect 421472 563218 421514 563454
rect 421750 563218 421792 563454
rect 421472 563134 421792 563218
rect 421472 562898 421514 563134
rect 421750 562898 421792 563134
rect 421472 562866 421792 562898
rect 443208 563454 443528 563486
rect 443208 563218 443250 563454
rect 443486 563218 443528 563454
rect 443208 563134 443528 563218
rect 443208 562898 443250 563134
rect 443486 562898 443528 563134
rect 443208 562866 443528 562898
rect 445710 554709 445770 576403
rect 446340 566829 446660 566861
rect 446340 566593 446382 566829
rect 446618 566593 446660 566829
rect 446340 566509 446660 566593
rect 446340 566273 446382 566509
rect 446618 566273 446660 566509
rect 446340 566241 446660 566273
rect 452604 566829 452924 566861
rect 452604 566593 452646 566829
rect 452882 566593 452924 566829
rect 452604 566509 452924 566593
rect 452604 566273 452646 566509
rect 452882 566273 452924 566509
rect 452604 566241 452924 566273
rect 468076 566829 468396 566861
rect 468076 566593 468118 566829
rect 468354 566593 468396 566829
rect 468076 566509 468396 566593
rect 468076 566273 468118 566509
rect 468354 566273 468396 566509
rect 468076 566241 468396 566273
rect 474340 566829 474660 566861
rect 474340 566593 474382 566829
rect 474618 566593 474660 566829
rect 474340 566509 474660 566593
rect 474340 566273 474382 566509
rect 474618 566273 474660 566509
rect 474340 566241 474660 566273
rect 480604 566829 480924 566861
rect 480604 566593 480646 566829
rect 480882 566593 480924 566829
rect 480604 566509 480924 566593
rect 480604 566273 480646 566509
rect 480882 566273 480924 566509
rect 480604 566241 480924 566273
rect 496076 566829 496396 566861
rect 496076 566593 496118 566829
rect 496354 566593 496396 566829
rect 496076 566509 496396 566593
rect 496076 566273 496118 566509
rect 496354 566273 496396 566509
rect 496076 566241 496396 566273
rect 502340 566829 502660 566861
rect 502340 566593 502382 566829
rect 502618 566593 502660 566829
rect 502340 566509 502660 566593
rect 502340 566273 502382 566509
rect 502618 566273 502660 566509
rect 502340 566241 502660 566273
rect 508604 566829 508924 566861
rect 508604 566593 508646 566829
rect 508882 566593 508924 566829
rect 508604 566509 508924 566593
rect 508604 566273 508646 566509
rect 508882 566273 508924 566509
rect 508604 566241 508924 566273
rect 524076 566829 524396 566861
rect 524076 566593 524118 566829
rect 524354 566593 524396 566829
rect 524076 566509 524396 566593
rect 524076 566273 524118 566509
rect 524354 566273 524396 566509
rect 524076 566241 524396 566273
rect 530340 566829 530660 566861
rect 530340 566593 530382 566829
rect 530618 566593 530660 566829
rect 530340 566509 530660 566593
rect 530340 566273 530382 566509
rect 530618 566273 530660 566509
rect 530340 566241 530660 566273
rect 536604 566829 536924 566861
rect 536604 566593 536646 566829
rect 536882 566593 536924 566829
rect 536604 566509 536924 566593
rect 536604 566273 536646 566509
rect 536882 566273 536924 566509
rect 536604 566241 536924 566273
rect 552076 566829 552396 566861
rect 552076 566593 552118 566829
rect 552354 566593 552396 566829
rect 552076 566509 552396 566593
rect 552076 566273 552118 566509
rect 552354 566273 552396 566509
rect 552076 566241 552396 566273
rect 449472 563454 449792 563486
rect 449472 563218 449514 563454
rect 449750 563218 449792 563454
rect 449472 563134 449792 563218
rect 449472 562898 449514 563134
rect 449750 562898 449792 563134
rect 449472 562866 449792 562898
rect 471208 563454 471528 563486
rect 471208 563218 471250 563454
rect 471486 563218 471528 563454
rect 471208 563134 471528 563218
rect 471208 562898 471250 563134
rect 471486 562898 471528 563134
rect 471208 562866 471528 562898
rect 477472 563454 477792 563486
rect 477472 563218 477514 563454
rect 477750 563218 477792 563454
rect 477472 563134 477792 563218
rect 477472 562898 477514 563134
rect 477750 562898 477792 563134
rect 477472 562866 477792 562898
rect 499208 563454 499528 563486
rect 499208 563218 499250 563454
rect 499486 563218 499528 563454
rect 499208 563134 499528 563218
rect 499208 562898 499250 563134
rect 499486 562898 499528 563134
rect 499208 562866 499528 562898
rect 505472 563454 505792 563486
rect 505472 563218 505514 563454
rect 505750 563218 505792 563454
rect 505472 563134 505792 563218
rect 505472 562898 505514 563134
rect 505750 562898 505792 563134
rect 505472 562866 505792 562898
rect 527208 563454 527528 563486
rect 527208 563218 527250 563454
rect 527486 563218 527528 563454
rect 527208 563134 527528 563218
rect 527208 562898 527250 563134
rect 527486 562898 527528 563134
rect 527208 562866 527528 562898
rect 533472 563454 533792 563486
rect 533472 563218 533514 563454
rect 533750 563218 533792 563454
rect 533472 563134 533792 563218
rect 533472 562898 533514 563134
rect 533750 562898 533792 563134
rect 533472 562866 533792 562898
rect 555208 563454 555528 563486
rect 555208 563218 555250 563454
rect 555486 563218 555528 563454
rect 555208 563134 555528 563218
rect 555208 562898 555250 563134
rect 555486 562898 555528 563134
rect 555208 562866 555528 562898
rect 557582 554709 557642 576403
rect 558340 566829 558660 566861
rect 558340 566593 558382 566829
rect 558618 566593 558660 566829
rect 558340 566509 558660 566593
rect 558340 566273 558382 566509
rect 558618 566273 558660 566509
rect 558340 566241 558660 566273
rect 564604 566829 564924 566861
rect 564604 566593 564646 566829
rect 564882 566593 564924 566829
rect 564604 566509 564924 566593
rect 564604 566273 564646 566509
rect 564882 566273 564924 566509
rect 564604 566241 564924 566273
rect 573494 566829 574114 593273
rect 573494 566593 573526 566829
rect 573762 566593 573846 566829
rect 574082 566593 574114 566829
rect 573494 566509 574114 566593
rect 573494 566273 573526 566509
rect 573762 566273 573846 566509
rect 574082 566273 574114 566509
rect 561472 563454 561792 563486
rect 561472 563218 561514 563454
rect 561750 563218 561792 563454
rect 561472 563134 561792 563218
rect 561472 562898 561514 563134
rect 561750 562898 561792 563134
rect 561472 562866 561792 562898
rect 165659 554708 165725 554709
rect 165659 554644 165660 554708
rect 165724 554644 165725 554708
rect 165659 554643 165725 554644
rect 259499 554708 259565 554709
rect 259499 554644 259500 554708
rect 259564 554644 259565 554708
rect 259499 554643 259565 554644
rect 361619 554708 361685 554709
rect 361619 554644 361620 554708
rect 361684 554644 361685 554708
rect 361619 554643 361685 554644
rect 445707 554708 445773 554709
rect 445707 554644 445708 554708
rect 445772 554644 445773 554708
rect 445707 554643 445773 554644
rect 557579 554708 557645 554709
rect 557579 554644 557580 554708
rect 557644 554644 557645 554708
rect 557579 554643 557645 554644
rect 128307 549404 128373 549405
rect 128307 549340 128308 549404
rect 128372 549340 128373 549404
rect 128307 549339 128373 549340
rect 194731 549404 194797 549405
rect 194731 549340 194732 549404
rect 194796 549340 194797 549404
rect 194731 549339 194797 549340
rect 390875 549404 390941 549405
rect 390875 549340 390876 549404
rect 390940 549340 390941 549404
rect 390875 549339 390941 549340
rect 92427 548180 92493 548181
rect 92427 548116 92428 548180
rect 92492 548116 92493 548180
rect 92427 548115 92493 548116
rect 64459 548044 64525 548045
rect 64459 547980 64460 548044
rect 64524 547980 64525 548044
rect 64459 547979 64525 547980
rect 64462 540293 64522 547979
rect 92430 540293 92490 548115
rect 64459 540292 64525 540293
rect 64459 540228 64460 540292
rect 64524 540228 64525 540292
rect 64459 540227 64525 540228
rect 92427 540292 92493 540293
rect 92427 540228 92428 540292
rect 92492 540228 92493 540292
rect 92427 540227 92493 540228
rect -2006 539593 -1974 539829
rect -1738 539593 -1654 539829
rect -1418 539593 -1386 539829
rect -2006 539509 -1386 539593
rect -2006 539273 -1974 539509
rect -1738 539273 -1654 539509
rect -1418 539273 -1386 539509
rect -2006 512829 -1386 539273
rect 20076 539829 20396 539861
rect 20076 539593 20118 539829
rect 20354 539593 20396 539829
rect 20076 539509 20396 539593
rect 20076 539273 20118 539509
rect 20354 539273 20396 539509
rect 20076 539241 20396 539273
rect 26340 539829 26660 539861
rect 26340 539593 26382 539829
rect 26618 539593 26660 539829
rect 26340 539509 26660 539593
rect 26340 539273 26382 539509
rect 26618 539273 26660 539509
rect 26340 539241 26660 539273
rect 32604 539829 32924 539861
rect 32604 539593 32646 539829
rect 32882 539593 32924 539829
rect 32604 539509 32924 539593
rect 32604 539273 32646 539509
rect 32882 539273 32924 539509
rect 32604 539241 32924 539273
rect 48076 539829 48396 539861
rect 48076 539593 48118 539829
rect 48354 539593 48396 539829
rect 48076 539509 48396 539593
rect 48076 539273 48118 539509
rect 48354 539273 48396 539509
rect 48076 539241 48396 539273
rect 54340 539829 54660 539861
rect 54340 539593 54382 539829
rect 54618 539593 54660 539829
rect 54340 539509 54660 539593
rect 54340 539273 54382 539509
rect 54618 539273 54660 539509
rect 54340 539241 54660 539273
rect 60604 539829 60924 539861
rect 60604 539593 60646 539829
rect 60882 539593 60924 539829
rect 60604 539509 60924 539593
rect 60604 539273 60646 539509
rect 60882 539273 60924 539509
rect 60604 539241 60924 539273
rect 76076 539829 76396 539861
rect 76076 539593 76118 539829
rect 76354 539593 76396 539829
rect 76076 539509 76396 539593
rect 76076 539273 76118 539509
rect 76354 539273 76396 539509
rect 76076 539241 76396 539273
rect 82340 539829 82660 539861
rect 82340 539593 82382 539829
rect 82618 539593 82660 539829
rect 82340 539509 82660 539593
rect 82340 539273 82382 539509
rect 82618 539273 82660 539509
rect 82340 539241 82660 539273
rect 88604 539829 88924 539861
rect 88604 539593 88646 539829
rect 88882 539593 88924 539829
rect 88604 539509 88924 539593
rect 88604 539273 88646 539509
rect 88882 539273 88924 539509
rect 88604 539241 88924 539273
rect 104076 539829 104396 539861
rect 104076 539593 104118 539829
rect 104354 539593 104396 539829
rect 104076 539509 104396 539593
rect 104076 539273 104118 539509
rect 104354 539273 104396 539509
rect 104076 539241 104396 539273
rect 110340 539829 110660 539861
rect 110340 539593 110382 539829
rect 110618 539593 110660 539829
rect 110340 539509 110660 539593
rect 110340 539273 110382 539509
rect 110618 539273 110660 539509
rect 110340 539241 110660 539273
rect 116604 539829 116924 539861
rect 116604 539593 116646 539829
rect 116882 539593 116924 539829
rect 116604 539509 116924 539593
rect 116604 539273 116646 539509
rect 116882 539273 116924 539509
rect 116604 539241 116924 539273
rect 23208 536454 23528 536486
rect 23208 536218 23250 536454
rect 23486 536218 23528 536454
rect 23208 536134 23528 536218
rect 23208 535898 23250 536134
rect 23486 535898 23528 536134
rect 23208 535866 23528 535898
rect 29472 536454 29792 536486
rect 29472 536218 29514 536454
rect 29750 536218 29792 536454
rect 29472 536134 29792 536218
rect 29472 535898 29514 536134
rect 29750 535898 29792 536134
rect 29472 535866 29792 535898
rect 51208 536454 51528 536486
rect 51208 536218 51250 536454
rect 51486 536218 51528 536454
rect 51208 536134 51528 536218
rect 51208 535898 51250 536134
rect 51486 535898 51528 536134
rect 51208 535866 51528 535898
rect 57472 536454 57792 536486
rect 57472 536218 57514 536454
rect 57750 536218 57792 536454
rect 57472 536134 57792 536218
rect 57472 535898 57514 536134
rect 57750 535898 57792 536134
rect 57472 535866 57792 535898
rect 79208 536454 79528 536486
rect 79208 536218 79250 536454
rect 79486 536218 79528 536454
rect 79208 536134 79528 536218
rect 79208 535898 79250 536134
rect 79486 535898 79528 536134
rect 79208 535866 79528 535898
rect 85472 536454 85792 536486
rect 85472 536218 85514 536454
rect 85750 536218 85792 536454
rect 85472 536134 85792 536218
rect 85472 535898 85514 536134
rect 85750 535898 85792 536134
rect 85472 535866 85792 535898
rect 107208 536454 107528 536486
rect 107208 536218 107250 536454
rect 107486 536218 107528 536454
rect 107208 536134 107528 536218
rect 107208 535898 107250 536134
rect 107486 535898 107528 536134
rect 107208 535866 107528 535898
rect 113472 536454 113792 536486
rect 113472 536218 113514 536454
rect 113750 536218 113792 536454
rect 113472 536134 113792 536218
rect 113472 535898 113514 536134
rect 113750 535898 113792 536134
rect 113472 535866 113792 535898
rect 128310 527101 128370 549339
rect 148363 548180 148429 548181
rect 148363 548116 148364 548180
rect 148428 548116 148429 548180
rect 148363 548115 148429 548116
rect 148366 540293 148426 548115
rect 176331 548044 176397 548045
rect 176331 547980 176332 548044
rect 176396 547980 176397 548044
rect 176331 547979 176397 547980
rect 176334 540293 176394 547979
rect 148363 540292 148429 540293
rect 148363 540228 148364 540292
rect 148428 540228 148429 540292
rect 148363 540227 148429 540228
rect 176331 540292 176397 540293
rect 176331 540228 176332 540292
rect 176396 540228 176397 540292
rect 176331 540227 176397 540228
rect 132076 539829 132396 539861
rect 132076 539593 132118 539829
rect 132354 539593 132396 539829
rect 132076 539509 132396 539593
rect 132076 539273 132118 539509
rect 132354 539273 132396 539509
rect 132076 539241 132396 539273
rect 138340 539829 138660 539861
rect 138340 539593 138382 539829
rect 138618 539593 138660 539829
rect 138340 539509 138660 539593
rect 138340 539273 138382 539509
rect 138618 539273 138660 539509
rect 138340 539241 138660 539273
rect 144604 539829 144924 539861
rect 144604 539593 144646 539829
rect 144882 539593 144924 539829
rect 144604 539509 144924 539593
rect 144604 539273 144646 539509
rect 144882 539273 144924 539509
rect 144604 539241 144924 539273
rect 160076 539829 160396 539861
rect 160076 539593 160118 539829
rect 160354 539593 160396 539829
rect 160076 539509 160396 539593
rect 160076 539273 160118 539509
rect 160354 539273 160396 539509
rect 160076 539241 160396 539273
rect 166340 539829 166660 539861
rect 166340 539593 166382 539829
rect 166618 539593 166660 539829
rect 166340 539509 166660 539593
rect 166340 539273 166382 539509
rect 166618 539273 166660 539509
rect 166340 539241 166660 539273
rect 172604 539829 172924 539861
rect 172604 539593 172646 539829
rect 172882 539593 172924 539829
rect 172604 539509 172924 539593
rect 172604 539273 172646 539509
rect 172882 539273 172924 539509
rect 172604 539241 172924 539273
rect 188076 539829 188396 539861
rect 188076 539593 188118 539829
rect 188354 539593 188396 539829
rect 188076 539509 188396 539593
rect 188076 539273 188118 539509
rect 188354 539273 188396 539509
rect 188076 539241 188396 539273
rect 194340 539829 194660 539861
rect 194340 539593 194382 539829
rect 194618 539593 194660 539829
rect 194340 539509 194660 539593
rect 194340 539273 194382 539509
rect 194618 539273 194660 539509
rect 194340 539241 194660 539273
rect 135208 536454 135528 536486
rect 135208 536218 135250 536454
rect 135486 536218 135528 536454
rect 135208 536134 135528 536218
rect 135208 535898 135250 536134
rect 135486 535898 135528 536134
rect 135208 535866 135528 535898
rect 141472 536454 141792 536486
rect 141472 536218 141514 536454
rect 141750 536218 141792 536454
rect 141472 536134 141792 536218
rect 141472 535898 141514 536134
rect 141750 535898 141792 536134
rect 141472 535866 141792 535898
rect 163208 536454 163528 536486
rect 163208 536218 163250 536454
rect 163486 536218 163528 536454
rect 163208 536134 163528 536218
rect 163208 535898 163250 536134
rect 163486 535898 163528 536134
rect 163208 535866 163528 535898
rect 169472 536454 169792 536486
rect 169472 536218 169514 536454
rect 169750 536218 169792 536454
rect 169472 536134 169792 536218
rect 169472 535898 169514 536134
rect 169750 535898 169792 536134
rect 169472 535866 169792 535898
rect 191208 536454 191528 536486
rect 191208 536218 191250 536454
rect 191486 536218 191528 536454
rect 191208 536134 191528 536218
rect 191208 535898 191250 536134
rect 191486 535898 191528 536134
rect 191208 535866 191528 535898
rect 194734 527101 194794 549339
rect 288387 548316 288453 548317
rect 288387 548252 288388 548316
rect 288452 548252 288453 548316
rect 288387 548251 288453 548252
rect 372291 548316 372357 548317
rect 372291 548252 372292 548316
rect 372356 548252 372357 548316
rect 372291 548251 372357 548252
rect 212579 548180 212645 548181
rect 212579 548116 212580 548180
rect 212644 548116 212645 548180
rect 212579 548115 212645 548116
rect 212582 540293 212642 548115
rect 288390 540293 288450 548251
rect 296851 548180 296917 548181
rect 296851 548116 296852 548180
rect 296916 548116 296917 548180
rect 296851 548115 296917 548116
rect 296854 540990 296914 548115
rect 296486 540930 296914 540990
rect 296486 540293 296546 540930
rect 372294 540293 372354 548251
rect 212579 540292 212645 540293
rect 212579 540228 212580 540292
rect 212644 540228 212645 540292
rect 212579 540227 212645 540228
rect 288387 540292 288453 540293
rect 288387 540228 288388 540292
rect 288452 540228 288453 540292
rect 288387 540227 288453 540228
rect 296483 540292 296549 540293
rect 296483 540228 296484 540292
rect 296548 540228 296549 540292
rect 296483 540227 296549 540228
rect 372291 540292 372357 540293
rect 372291 540228 372292 540292
rect 372356 540228 372357 540292
rect 372291 540227 372357 540228
rect 200604 539829 200924 539861
rect 200604 539593 200646 539829
rect 200882 539593 200924 539829
rect 200604 539509 200924 539593
rect 200604 539273 200646 539509
rect 200882 539273 200924 539509
rect 200604 539241 200924 539273
rect 216076 539829 216396 539861
rect 216076 539593 216118 539829
rect 216354 539593 216396 539829
rect 216076 539509 216396 539593
rect 216076 539273 216118 539509
rect 216354 539273 216396 539509
rect 216076 539241 216396 539273
rect 222340 539829 222660 539861
rect 222340 539593 222382 539829
rect 222618 539593 222660 539829
rect 222340 539509 222660 539593
rect 222340 539273 222382 539509
rect 222618 539273 222660 539509
rect 222340 539241 222660 539273
rect 228604 539829 228924 539861
rect 228604 539593 228646 539829
rect 228882 539593 228924 539829
rect 228604 539509 228924 539593
rect 228604 539273 228646 539509
rect 228882 539273 228924 539509
rect 228604 539241 228924 539273
rect 244076 539829 244396 539861
rect 244076 539593 244118 539829
rect 244354 539593 244396 539829
rect 244076 539509 244396 539593
rect 244076 539273 244118 539509
rect 244354 539273 244396 539509
rect 244076 539241 244396 539273
rect 250340 539829 250660 539861
rect 250340 539593 250382 539829
rect 250618 539593 250660 539829
rect 250340 539509 250660 539593
rect 250340 539273 250382 539509
rect 250618 539273 250660 539509
rect 250340 539241 250660 539273
rect 256604 539829 256924 539861
rect 256604 539593 256646 539829
rect 256882 539593 256924 539829
rect 256604 539509 256924 539593
rect 256604 539273 256646 539509
rect 256882 539273 256924 539509
rect 256604 539241 256924 539273
rect 272076 539829 272396 539861
rect 272076 539593 272118 539829
rect 272354 539593 272396 539829
rect 272076 539509 272396 539593
rect 272076 539273 272118 539509
rect 272354 539273 272396 539509
rect 272076 539241 272396 539273
rect 278340 539829 278660 539861
rect 278340 539593 278382 539829
rect 278618 539593 278660 539829
rect 278340 539509 278660 539593
rect 278340 539273 278382 539509
rect 278618 539273 278660 539509
rect 278340 539241 278660 539273
rect 284604 539829 284924 539861
rect 284604 539593 284646 539829
rect 284882 539593 284924 539829
rect 284604 539509 284924 539593
rect 284604 539273 284646 539509
rect 284882 539273 284924 539509
rect 284604 539241 284924 539273
rect 300076 539829 300396 539861
rect 300076 539593 300118 539829
rect 300354 539593 300396 539829
rect 300076 539509 300396 539593
rect 300076 539273 300118 539509
rect 300354 539273 300396 539509
rect 300076 539241 300396 539273
rect 306340 539829 306660 539861
rect 306340 539593 306382 539829
rect 306618 539593 306660 539829
rect 306340 539509 306660 539593
rect 306340 539273 306382 539509
rect 306618 539273 306660 539509
rect 306340 539241 306660 539273
rect 312604 539829 312924 539861
rect 312604 539593 312646 539829
rect 312882 539593 312924 539829
rect 312604 539509 312924 539593
rect 312604 539273 312646 539509
rect 312882 539273 312924 539509
rect 312604 539241 312924 539273
rect 328076 539829 328396 539861
rect 328076 539593 328118 539829
rect 328354 539593 328396 539829
rect 328076 539509 328396 539593
rect 328076 539273 328118 539509
rect 328354 539273 328396 539509
rect 328076 539241 328396 539273
rect 334340 539829 334660 539861
rect 334340 539593 334382 539829
rect 334618 539593 334660 539829
rect 334340 539509 334660 539593
rect 334340 539273 334382 539509
rect 334618 539273 334660 539509
rect 334340 539241 334660 539273
rect 340604 539829 340924 539861
rect 340604 539593 340646 539829
rect 340882 539593 340924 539829
rect 340604 539509 340924 539593
rect 340604 539273 340646 539509
rect 340882 539273 340924 539509
rect 340604 539241 340924 539273
rect 356076 539829 356396 539861
rect 356076 539593 356118 539829
rect 356354 539593 356396 539829
rect 356076 539509 356396 539593
rect 356076 539273 356118 539509
rect 356354 539273 356396 539509
rect 356076 539241 356396 539273
rect 362340 539829 362660 539861
rect 362340 539593 362382 539829
rect 362618 539593 362660 539829
rect 362340 539509 362660 539593
rect 362340 539273 362382 539509
rect 362618 539273 362660 539509
rect 362340 539241 362660 539273
rect 368604 539829 368924 539861
rect 368604 539593 368646 539829
rect 368882 539593 368924 539829
rect 368604 539509 368924 539593
rect 368604 539273 368646 539509
rect 368882 539273 368924 539509
rect 368604 539241 368924 539273
rect 384076 539829 384396 539861
rect 384076 539593 384118 539829
rect 384354 539593 384396 539829
rect 384076 539509 384396 539593
rect 384076 539273 384118 539509
rect 384354 539273 384396 539509
rect 384076 539241 384396 539273
rect 390340 539829 390660 539861
rect 390340 539593 390382 539829
rect 390618 539593 390660 539829
rect 390340 539509 390660 539593
rect 390340 539273 390382 539509
rect 390618 539273 390660 539509
rect 390340 539241 390660 539273
rect 197472 536454 197792 536486
rect 197472 536218 197514 536454
rect 197750 536218 197792 536454
rect 197472 536134 197792 536218
rect 197472 535898 197514 536134
rect 197750 535898 197792 536134
rect 197472 535866 197792 535898
rect 219208 536454 219528 536486
rect 219208 536218 219250 536454
rect 219486 536218 219528 536454
rect 219208 536134 219528 536218
rect 219208 535898 219250 536134
rect 219486 535898 219528 536134
rect 219208 535866 219528 535898
rect 225472 536454 225792 536486
rect 225472 536218 225514 536454
rect 225750 536218 225792 536454
rect 225472 536134 225792 536218
rect 225472 535898 225514 536134
rect 225750 535898 225792 536134
rect 225472 535866 225792 535898
rect 247208 536454 247528 536486
rect 247208 536218 247250 536454
rect 247486 536218 247528 536454
rect 247208 536134 247528 536218
rect 247208 535898 247250 536134
rect 247486 535898 247528 536134
rect 247208 535866 247528 535898
rect 253472 536454 253792 536486
rect 253472 536218 253514 536454
rect 253750 536218 253792 536454
rect 253472 536134 253792 536218
rect 253472 535898 253514 536134
rect 253750 535898 253792 536134
rect 253472 535866 253792 535898
rect 275208 536454 275528 536486
rect 275208 536218 275250 536454
rect 275486 536218 275528 536454
rect 275208 536134 275528 536218
rect 275208 535898 275250 536134
rect 275486 535898 275528 536134
rect 275208 535866 275528 535898
rect 281472 536454 281792 536486
rect 281472 536218 281514 536454
rect 281750 536218 281792 536454
rect 281472 536134 281792 536218
rect 281472 535898 281514 536134
rect 281750 535898 281792 536134
rect 281472 535866 281792 535898
rect 303208 536454 303528 536486
rect 303208 536218 303250 536454
rect 303486 536218 303528 536454
rect 303208 536134 303528 536218
rect 303208 535898 303250 536134
rect 303486 535898 303528 536134
rect 303208 535866 303528 535898
rect 309472 536454 309792 536486
rect 309472 536218 309514 536454
rect 309750 536218 309792 536454
rect 309472 536134 309792 536218
rect 309472 535898 309514 536134
rect 309750 535898 309792 536134
rect 309472 535866 309792 535898
rect 331208 536454 331528 536486
rect 331208 536218 331250 536454
rect 331486 536218 331528 536454
rect 331208 536134 331528 536218
rect 331208 535898 331250 536134
rect 331486 535898 331528 536134
rect 331208 535866 331528 535898
rect 337472 536454 337792 536486
rect 337472 536218 337514 536454
rect 337750 536218 337792 536454
rect 337472 536134 337792 536218
rect 337472 535898 337514 536134
rect 337750 535898 337792 536134
rect 337472 535866 337792 535898
rect 359208 536454 359528 536486
rect 359208 536218 359250 536454
rect 359486 536218 359528 536454
rect 359208 536134 359528 536218
rect 359208 535898 359250 536134
rect 359486 535898 359528 536134
rect 359208 535866 359528 535898
rect 365472 536454 365792 536486
rect 365472 536218 365514 536454
rect 365750 536218 365792 536454
rect 365472 536134 365792 536218
rect 365472 535898 365514 536134
rect 365750 535898 365792 536134
rect 365472 535866 365792 535898
rect 387208 536454 387528 536486
rect 387208 536218 387250 536454
rect 387486 536218 387528 536454
rect 387208 536134 387528 536218
rect 387208 535898 387250 536134
rect 387486 535898 387528 536134
rect 387208 535866 387528 535898
rect 390878 527101 390938 549339
rect 484347 548180 484413 548181
rect 484347 548116 484348 548180
rect 484412 548116 484413 548180
rect 484347 548115 484413 548116
rect 540467 548180 540533 548181
rect 540467 548116 540468 548180
rect 540532 548116 540533 548180
rect 540467 548115 540533 548116
rect 408539 548044 408605 548045
rect 408539 547980 408540 548044
rect 408604 547980 408605 548044
rect 408539 547979 408605 547980
rect 408542 540293 408602 547979
rect 484350 540293 484410 548115
rect 520595 548044 520661 548045
rect 520595 547980 520596 548044
rect 520660 547980 520661 548044
rect 520595 547979 520661 547980
rect 520598 540293 520658 547979
rect 540470 540293 540530 548115
rect 408539 540292 408605 540293
rect 408539 540228 408540 540292
rect 408604 540228 408605 540292
rect 408539 540227 408605 540228
rect 484347 540292 484413 540293
rect 484347 540228 484348 540292
rect 484412 540228 484413 540292
rect 484347 540227 484413 540228
rect 520595 540292 520661 540293
rect 520595 540228 520596 540292
rect 520660 540228 520661 540292
rect 520595 540227 520661 540228
rect 540467 540292 540533 540293
rect 540467 540228 540468 540292
rect 540532 540228 540533 540292
rect 540467 540227 540533 540228
rect 396604 539829 396924 539861
rect 396604 539593 396646 539829
rect 396882 539593 396924 539829
rect 396604 539509 396924 539593
rect 396604 539273 396646 539509
rect 396882 539273 396924 539509
rect 396604 539241 396924 539273
rect 412076 539829 412396 539861
rect 412076 539593 412118 539829
rect 412354 539593 412396 539829
rect 412076 539509 412396 539593
rect 412076 539273 412118 539509
rect 412354 539273 412396 539509
rect 412076 539241 412396 539273
rect 418340 539829 418660 539861
rect 418340 539593 418382 539829
rect 418618 539593 418660 539829
rect 418340 539509 418660 539593
rect 418340 539273 418382 539509
rect 418618 539273 418660 539509
rect 418340 539241 418660 539273
rect 424604 539829 424924 539861
rect 424604 539593 424646 539829
rect 424882 539593 424924 539829
rect 424604 539509 424924 539593
rect 424604 539273 424646 539509
rect 424882 539273 424924 539509
rect 424604 539241 424924 539273
rect 440076 539829 440396 539861
rect 440076 539593 440118 539829
rect 440354 539593 440396 539829
rect 440076 539509 440396 539593
rect 440076 539273 440118 539509
rect 440354 539273 440396 539509
rect 440076 539241 440396 539273
rect 446340 539829 446660 539861
rect 446340 539593 446382 539829
rect 446618 539593 446660 539829
rect 446340 539509 446660 539593
rect 446340 539273 446382 539509
rect 446618 539273 446660 539509
rect 446340 539241 446660 539273
rect 452604 539829 452924 539861
rect 452604 539593 452646 539829
rect 452882 539593 452924 539829
rect 452604 539509 452924 539593
rect 452604 539273 452646 539509
rect 452882 539273 452924 539509
rect 452604 539241 452924 539273
rect 468076 539829 468396 539861
rect 468076 539593 468118 539829
rect 468354 539593 468396 539829
rect 468076 539509 468396 539593
rect 468076 539273 468118 539509
rect 468354 539273 468396 539509
rect 468076 539241 468396 539273
rect 474340 539829 474660 539861
rect 474340 539593 474382 539829
rect 474618 539593 474660 539829
rect 474340 539509 474660 539593
rect 474340 539273 474382 539509
rect 474618 539273 474660 539509
rect 474340 539241 474660 539273
rect 480604 539829 480924 539861
rect 480604 539593 480646 539829
rect 480882 539593 480924 539829
rect 480604 539509 480924 539593
rect 480604 539273 480646 539509
rect 480882 539273 480924 539509
rect 480604 539241 480924 539273
rect 496076 539829 496396 539861
rect 496076 539593 496118 539829
rect 496354 539593 496396 539829
rect 496076 539509 496396 539593
rect 496076 539273 496118 539509
rect 496354 539273 496396 539509
rect 496076 539241 496396 539273
rect 502340 539829 502660 539861
rect 502340 539593 502382 539829
rect 502618 539593 502660 539829
rect 502340 539509 502660 539593
rect 502340 539273 502382 539509
rect 502618 539273 502660 539509
rect 502340 539241 502660 539273
rect 508604 539829 508924 539861
rect 508604 539593 508646 539829
rect 508882 539593 508924 539829
rect 508604 539509 508924 539593
rect 508604 539273 508646 539509
rect 508882 539273 508924 539509
rect 508604 539241 508924 539273
rect 524076 539829 524396 539861
rect 524076 539593 524118 539829
rect 524354 539593 524396 539829
rect 524076 539509 524396 539593
rect 524076 539273 524118 539509
rect 524354 539273 524396 539509
rect 524076 539241 524396 539273
rect 530340 539829 530660 539861
rect 530340 539593 530382 539829
rect 530618 539593 530660 539829
rect 530340 539509 530660 539593
rect 530340 539273 530382 539509
rect 530618 539273 530660 539509
rect 530340 539241 530660 539273
rect 536604 539829 536924 539861
rect 536604 539593 536646 539829
rect 536882 539593 536924 539829
rect 536604 539509 536924 539593
rect 536604 539273 536646 539509
rect 536882 539273 536924 539509
rect 536604 539241 536924 539273
rect 552076 539829 552396 539861
rect 552076 539593 552118 539829
rect 552354 539593 552396 539829
rect 552076 539509 552396 539593
rect 552076 539273 552118 539509
rect 552354 539273 552396 539509
rect 552076 539241 552396 539273
rect 558340 539829 558660 539861
rect 558340 539593 558382 539829
rect 558618 539593 558660 539829
rect 558340 539509 558660 539593
rect 558340 539273 558382 539509
rect 558618 539273 558660 539509
rect 558340 539241 558660 539273
rect 564604 539829 564924 539861
rect 564604 539593 564646 539829
rect 564882 539593 564924 539829
rect 564604 539509 564924 539593
rect 564604 539273 564646 539509
rect 564882 539273 564924 539509
rect 564604 539241 564924 539273
rect 573494 539829 574114 566273
rect 573494 539593 573526 539829
rect 573762 539593 573846 539829
rect 574082 539593 574114 539829
rect 573494 539509 574114 539593
rect 573494 539273 573526 539509
rect 573762 539273 573846 539509
rect 574082 539273 574114 539509
rect 393472 536454 393792 536486
rect 393472 536218 393514 536454
rect 393750 536218 393792 536454
rect 393472 536134 393792 536218
rect 393472 535898 393514 536134
rect 393750 535898 393792 536134
rect 393472 535866 393792 535898
rect 415208 536454 415528 536486
rect 415208 536218 415250 536454
rect 415486 536218 415528 536454
rect 415208 536134 415528 536218
rect 415208 535898 415250 536134
rect 415486 535898 415528 536134
rect 415208 535866 415528 535898
rect 421472 536454 421792 536486
rect 421472 536218 421514 536454
rect 421750 536218 421792 536454
rect 421472 536134 421792 536218
rect 421472 535898 421514 536134
rect 421750 535898 421792 536134
rect 421472 535866 421792 535898
rect 443208 536454 443528 536486
rect 443208 536218 443250 536454
rect 443486 536218 443528 536454
rect 443208 536134 443528 536218
rect 443208 535898 443250 536134
rect 443486 535898 443528 536134
rect 443208 535866 443528 535898
rect 449472 536454 449792 536486
rect 449472 536218 449514 536454
rect 449750 536218 449792 536454
rect 449472 536134 449792 536218
rect 449472 535898 449514 536134
rect 449750 535898 449792 536134
rect 449472 535866 449792 535898
rect 471208 536454 471528 536486
rect 471208 536218 471250 536454
rect 471486 536218 471528 536454
rect 471208 536134 471528 536218
rect 471208 535898 471250 536134
rect 471486 535898 471528 536134
rect 471208 535866 471528 535898
rect 477472 536454 477792 536486
rect 477472 536218 477514 536454
rect 477750 536218 477792 536454
rect 477472 536134 477792 536218
rect 477472 535898 477514 536134
rect 477750 535898 477792 536134
rect 477472 535866 477792 535898
rect 499208 536454 499528 536486
rect 499208 536218 499250 536454
rect 499486 536218 499528 536454
rect 499208 536134 499528 536218
rect 499208 535898 499250 536134
rect 499486 535898 499528 536134
rect 499208 535866 499528 535898
rect 505472 536454 505792 536486
rect 505472 536218 505514 536454
rect 505750 536218 505792 536454
rect 505472 536134 505792 536218
rect 505472 535898 505514 536134
rect 505750 535898 505792 536134
rect 505472 535866 505792 535898
rect 527208 536454 527528 536486
rect 527208 536218 527250 536454
rect 527486 536218 527528 536454
rect 527208 536134 527528 536218
rect 527208 535898 527250 536134
rect 527486 535898 527528 536134
rect 527208 535866 527528 535898
rect 533472 536454 533792 536486
rect 533472 536218 533514 536454
rect 533750 536218 533792 536454
rect 533472 536134 533792 536218
rect 533472 535898 533514 536134
rect 533750 535898 533792 536134
rect 533472 535866 533792 535898
rect 555208 536454 555528 536486
rect 555208 536218 555250 536454
rect 555486 536218 555528 536454
rect 555208 536134 555528 536218
rect 555208 535898 555250 536134
rect 555486 535898 555528 536134
rect 555208 535866 555528 535898
rect 561472 536454 561792 536486
rect 561472 536218 561514 536454
rect 561750 536218 561792 536454
rect 561472 536134 561792 536218
rect 561472 535898 561514 536134
rect 561750 535898 561792 536134
rect 561472 535866 561792 535898
rect 128307 527100 128373 527101
rect 128307 527036 128308 527100
rect 128372 527036 128373 527100
rect 128307 527035 128373 527036
rect 194731 527100 194797 527101
rect 194731 527036 194732 527100
rect 194796 527036 194797 527100
rect 194731 527035 194797 527036
rect 390875 527100 390941 527101
rect 390875 527036 390876 527100
rect 390940 527036 390941 527100
rect 390875 527035 390941 527036
rect 165659 522476 165725 522477
rect 165659 522412 165660 522476
rect 165724 522412 165725 522476
rect 165659 522411 165725 522412
rect 259499 522476 259565 522477
rect 259499 522412 259500 522476
rect 259564 522412 259565 522476
rect 259499 522411 259565 522412
rect 361619 522476 361685 522477
rect 361619 522412 361620 522476
rect 361684 522412 361685 522476
rect 361619 522411 361685 522412
rect 445707 522476 445773 522477
rect 445707 522412 445708 522476
rect 445772 522412 445773 522476
rect 445707 522411 445773 522412
rect 557579 522476 557645 522477
rect 557579 522412 557580 522476
rect 557644 522412 557645 522476
rect 557579 522411 557645 522412
rect 44587 520980 44653 520981
rect 44587 520916 44588 520980
rect 44652 520916 44653 520980
rect 44587 520915 44653 520916
rect -2006 512593 -1974 512829
rect -1738 512593 -1654 512829
rect -1418 512593 -1386 512829
rect -2006 512509 -1386 512593
rect -2006 512273 -1974 512509
rect -1738 512273 -1654 512509
rect -1418 512273 -1386 512509
rect -2006 485829 -1386 512273
rect 20076 512829 20396 512861
rect 20076 512593 20118 512829
rect 20354 512593 20396 512829
rect 20076 512509 20396 512593
rect 20076 512273 20118 512509
rect 20354 512273 20396 512509
rect 20076 512241 20396 512273
rect 26340 512829 26660 512861
rect 26340 512593 26382 512829
rect 26618 512593 26660 512829
rect 26340 512509 26660 512593
rect 26340 512273 26382 512509
rect 26618 512273 26660 512509
rect 26340 512241 26660 512273
rect 32604 512829 32924 512861
rect 32604 512593 32646 512829
rect 32882 512593 32924 512829
rect 44590 512821 44650 520915
rect 48076 512829 48396 512861
rect 44587 512820 44653 512821
rect 44587 512756 44588 512820
rect 44652 512756 44653 512820
rect 44587 512755 44653 512756
rect 32604 512509 32924 512593
rect 32604 512273 32646 512509
rect 32882 512273 32924 512509
rect 32604 512241 32924 512273
rect 48076 512593 48118 512829
rect 48354 512593 48396 512829
rect 48076 512509 48396 512593
rect 48076 512273 48118 512509
rect 48354 512273 48396 512509
rect 48076 512241 48396 512273
rect 54340 512829 54660 512861
rect 54340 512593 54382 512829
rect 54618 512593 54660 512829
rect 54340 512509 54660 512593
rect 54340 512273 54382 512509
rect 54618 512273 54660 512509
rect 54340 512241 54660 512273
rect 60604 512829 60924 512861
rect 60604 512593 60646 512829
rect 60882 512593 60924 512829
rect 60604 512509 60924 512593
rect 60604 512273 60646 512509
rect 60882 512273 60924 512509
rect 60604 512241 60924 512273
rect 76076 512829 76396 512861
rect 76076 512593 76118 512829
rect 76354 512593 76396 512829
rect 76076 512509 76396 512593
rect 76076 512273 76118 512509
rect 76354 512273 76396 512509
rect 76076 512241 76396 512273
rect 82340 512829 82660 512861
rect 82340 512593 82382 512829
rect 82618 512593 82660 512829
rect 82340 512509 82660 512593
rect 82340 512273 82382 512509
rect 82618 512273 82660 512509
rect 82340 512241 82660 512273
rect 88604 512829 88924 512861
rect 88604 512593 88646 512829
rect 88882 512593 88924 512829
rect 88604 512509 88924 512593
rect 88604 512273 88646 512509
rect 88882 512273 88924 512509
rect 88604 512241 88924 512273
rect 104076 512829 104396 512861
rect 104076 512593 104118 512829
rect 104354 512593 104396 512829
rect 104076 512509 104396 512593
rect 104076 512273 104118 512509
rect 104354 512273 104396 512509
rect 104076 512241 104396 512273
rect 110340 512829 110660 512861
rect 110340 512593 110382 512829
rect 110618 512593 110660 512829
rect 110340 512509 110660 512593
rect 110340 512273 110382 512509
rect 110618 512273 110660 512509
rect 110340 512241 110660 512273
rect 116604 512829 116924 512861
rect 116604 512593 116646 512829
rect 116882 512593 116924 512829
rect 116604 512509 116924 512593
rect 116604 512273 116646 512509
rect 116882 512273 116924 512509
rect 116604 512241 116924 512273
rect 132076 512829 132396 512861
rect 132076 512593 132118 512829
rect 132354 512593 132396 512829
rect 132076 512509 132396 512593
rect 132076 512273 132118 512509
rect 132354 512273 132396 512509
rect 132076 512241 132396 512273
rect 138340 512829 138660 512861
rect 138340 512593 138382 512829
rect 138618 512593 138660 512829
rect 138340 512509 138660 512593
rect 138340 512273 138382 512509
rect 138618 512273 138660 512509
rect 138340 512241 138660 512273
rect 144604 512829 144924 512861
rect 144604 512593 144646 512829
rect 144882 512593 144924 512829
rect 144604 512509 144924 512593
rect 144604 512273 144646 512509
rect 144882 512273 144924 512509
rect 144604 512241 144924 512273
rect 160076 512829 160396 512861
rect 160076 512593 160118 512829
rect 160354 512593 160396 512829
rect 160076 512509 160396 512593
rect 160076 512273 160118 512509
rect 160354 512273 160396 512509
rect 160076 512241 160396 512273
rect 23208 509454 23528 509486
rect 23208 509218 23250 509454
rect 23486 509218 23528 509454
rect 23208 509134 23528 509218
rect 23208 508898 23250 509134
rect 23486 508898 23528 509134
rect 23208 508866 23528 508898
rect 29472 509454 29792 509486
rect 29472 509218 29514 509454
rect 29750 509218 29792 509454
rect 29472 509134 29792 509218
rect 29472 508898 29514 509134
rect 29750 508898 29792 509134
rect 29472 508866 29792 508898
rect 51208 509454 51528 509486
rect 51208 509218 51250 509454
rect 51486 509218 51528 509454
rect 51208 509134 51528 509218
rect 51208 508898 51250 509134
rect 51486 508898 51528 509134
rect 51208 508866 51528 508898
rect 57472 509454 57792 509486
rect 57472 509218 57514 509454
rect 57750 509218 57792 509454
rect 57472 509134 57792 509218
rect 57472 508898 57514 509134
rect 57750 508898 57792 509134
rect 57472 508866 57792 508898
rect 79208 509454 79528 509486
rect 79208 509218 79250 509454
rect 79486 509218 79528 509454
rect 79208 509134 79528 509218
rect 79208 508898 79250 509134
rect 79486 508898 79528 509134
rect 79208 508866 79528 508898
rect 85472 509454 85792 509486
rect 85472 509218 85514 509454
rect 85750 509218 85792 509454
rect 85472 509134 85792 509218
rect 85472 508898 85514 509134
rect 85750 508898 85792 509134
rect 85472 508866 85792 508898
rect 107208 509454 107528 509486
rect 107208 509218 107250 509454
rect 107486 509218 107528 509454
rect 107208 509134 107528 509218
rect 107208 508898 107250 509134
rect 107486 508898 107528 509134
rect 107208 508866 107528 508898
rect 113472 509454 113792 509486
rect 113472 509218 113514 509454
rect 113750 509218 113792 509454
rect 113472 509134 113792 509218
rect 113472 508898 113514 509134
rect 113750 508898 113792 509134
rect 113472 508866 113792 508898
rect 135208 509454 135528 509486
rect 135208 509218 135250 509454
rect 135486 509218 135528 509454
rect 135208 509134 135528 509218
rect 135208 508898 135250 509134
rect 135486 508898 135528 509134
rect 135208 508866 135528 508898
rect 141472 509454 141792 509486
rect 141472 509218 141514 509454
rect 141750 509218 141792 509454
rect 141472 509134 141792 509218
rect 141472 508898 141514 509134
rect 141750 508898 141792 509134
rect 141472 508866 141792 508898
rect 163208 509454 163528 509486
rect 163208 509218 163250 509454
rect 163486 509218 163528 509454
rect 163208 509134 163528 509218
rect 163208 508898 163250 509134
rect 163486 508898 163528 509134
rect 163208 508866 163528 508898
rect 165662 500853 165722 522411
rect 176331 520980 176397 520981
rect 176331 520916 176332 520980
rect 176396 520916 176397 520980
rect 176331 520915 176397 520916
rect 166340 512829 166660 512861
rect 166340 512593 166382 512829
rect 166618 512593 166660 512829
rect 166340 512509 166660 512593
rect 166340 512273 166382 512509
rect 166618 512273 166660 512509
rect 166340 512241 166660 512273
rect 172604 512829 172924 512861
rect 172604 512593 172646 512829
rect 172882 512593 172924 512829
rect 176334 512821 176394 520915
rect 212579 520844 212645 520845
rect 212579 520780 212580 520844
rect 212644 520780 212645 520844
rect 212579 520779 212645 520780
rect 188076 512829 188396 512861
rect 176331 512820 176397 512821
rect 176331 512756 176332 512820
rect 176396 512756 176397 512820
rect 176331 512755 176397 512756
rect 172604 512509 172924 512593
rect 172604 512273 172646 512509
rect 172882 512273 172924 512509
rect 172604 512241 172924 512273
rect 188076 512593 188118 512829
rect 188354 512593 188396 512829
rect 188076 512509 188396 512593
rect 188076 512273 188118 512509
rect 188354 512273 188396 512509
rect 188076 512241 188396 512273
rect 194340 512829 194660 512861
rect 194340 512593 194382 512829
rect 194618 512593 194660 512829
rect 194340 512509 194660 512593
rect 194340 512273 194382 512509
rect 194618 512273 194660 512509
rect 194340 512241 194660 512273
rect 200604 512829 200924 512861
rect 200604 512593 200646 512829
rect 200882 512593 200924 512829
rect 212582 512821 212642 520779
rect 216076 512829 216396 512861
rect 212579 512820 212645 512821
rect 212579 512756 212580 512820
rect 212644 512756 212645 512820
rect 212579 512755 212645 512756
rect 200604 512509 200924 512593
rect 200604 512273 200646 512509
rect 200882 512273 200924 512509
rect 200604 512241 200924 512273
rect 216076 512593 216118 512829
rect 216354 512593 216396 512829
rect 216076 512509 216396 512593
rect 216076 512273 216118 512509
rect 216354 512273 216396 512509
rect 216076 512241 216396 512273
rect 222340 512829 222660 512861
rect 222340 512593 222382 512829
rect 222618 512593 222660 512829
rect 222340 512509 222660 512593
rect 222340 512273 222382 512509
rect 222618 512273 222660 512509
rect 222340 512241 222660 512273
rect 228604 512829 228924 512861
rect 228604 512593 228646 512829
rect 228882 512593 228924 512829
rect 228604 512509 228924 512593
rect 228604 512273 228646 512509
rect 228882 512273 228924 512509
rect 228604 512241 228924 512273
rect 244076 512829 244396 512861
rect 244076 512593 244118 512829
rect 244354 512593 244396 512829
rect 244076 512509 244396 512593
rect 244076 512273 244118 512509
rect 244354 512273 244396 512509
rect 244076 512241 244396 512273
rect 250340 512829 250660 512861
rect 250340 512593 250382 512829
rect 250618 512593 250660 512829
rect 250340 512509 250660 512593
rect 250340 512273 250382 512509
rect 250618 512273 250660 512509
rect 250340 512241 250660 512273
rect 256604 512829 256924 512861
rect 256604 512593 256646 512829
rect 256882 512593 256924 512829
rect 256604 512509 256924 512593
rect 256604 512273 256646 512509
rect 256882 512273 256924 512509
rect 256604 512241 256924 512273
rect 169472 509454 169792 509486
rect 169472 509218 169514 509454
rect 169750 509218 169792 509454
rect 169472 509134 169792 509218
rect 169472 508898 169514 509134
rect 169750 508898 169792 509134
rect 169472 508866 169792 508898
rect 191208 509454 191528 509486
rect 191208 509218 191250 509454
rect 191486 509218 191528 509454
rect 191208 509134 191528 509218
rect 191208 508898 191250 509134
rect 191486 508898 191528 509134
rect 191208 508866 191528 508898
rect 197472 509454 197792 509486
rect 197472 509218 197514 509454
rect 197750 509218 197792 509454
rect 197472 509134 197792 509218
rect 197472 508898 197514 509134
rect 197750 508898 197792 509134
rect 197472 508866 197792 508898
rect 219208 509454 219528 509486
rect 219208 509218 219250 509454
rect 219486 509218 219528 509454
rect 219208 509134 219528 509218
rect 219208 508898 219250 509134
rect 219486 508898 219528 509134
rect 219208 508866 219528 508898
rect 225472 509454 225792 509486
rect 225472 509218 225514 509454
rect 225750 509218 225792 509454
rect 225472 509134 225792 509218
rect 225472 508898 225514 509134
rect 225750 508898 225792 509134
rect 225472 508866 225792 508898
rect 247208 509454 247528 509486
rect 247208 509218 247250 509454
rect 247486 509218 247528 509454
rect 247208 509134 247528 509218
rect 247208 508898 247250 509134
rect 247486 508898 247528 509134
rect 247208 508866 247528 508898
rect 253472 509454 253792 509486
rect 253472 509218 253514 509454
rect 253750 509218 253792 509454
rect 253472 509134 253792 509218
rect 253472 508898 253514 509134
rect 253750 508898 253792 509134
rect 253472 508866 253792 508898
rect 259502 500853 259562 522411
rect 288387 520980 288453 520981
rect 288387 520916 288388 520980
rect 288452 520916 288453 520980
rect 288387 520915 288453 520916
rect 272076 512829 272396 512861
rect 272076 512593 272118 512829
rect 272354 512593 272396 512829
rect 272076 512509 272396 512593
rect 272076 512273 272118 512509
rect 272354 512273 272396 512509
rect 272076 512241 272396 512273
rect 278340 512829 278660 512861
rect 278340 512593 278382 512829
rect 278618 512593 278660 512829
rect 278340 512509 278660 512593
rect 278340 512273 278382 512509
rect 278618 512273 278660 512509
rect 278340 512241 278660 512273
rect 284604 512829 284924 512861
rect 284604 512593 284646 512829
rect 284882 512593 284924 512829
rect 288390 512821 288450 520915
rect 296851 520844 296917 520845
rect 296851 520780 296852 520844
rect 296916 520780 296917 520844
rect 296851 520779 296917 520780
rect 296854 520570 296914 520779
rect 296486 520510 296914 520570
rect 296486 512821 296546 520510
rect 300076 512829 300396 512861
rect 288387 512820 288453 512821
rect 288387 512756 288388 512820
rect 288452 512756 288453 512820
rect 288387 512755 288453 512756
rect 296483 512820 296549 512821
rect 296483 512756 296484 512820
rect 296548 512756 296549 512820
rect 296483 512755 296549 512756
rect 284604 512509 284924 512593
rect 284604 512273 284646 512509
rect 284882 512273 284924 512509
rect 284604 512241 284924 512273
rect 300076 512593 300118 512829
rect 300354 512593 300396 512829
rect 300076 512509 300396 512593
rect 300076 512273 300118 512509
rect 300354 512273 300396 512509
rect 300076 512241 300396 512273
rect 306340 512829 306660 512861
rect 306340 512593 306382 512829
rect 306618 512593 306660 512829
rect 306340 512509 306660 512593
rect 306340 512273 306382 512509
rect 306618 512273 306660 512509
rect 306340 512241 306660 512273
rect 312604 512829 312924 512861
rect 312604 512593 312646 512829
rect 312882 512593 312924 512829
rect 312604 512509 312924 512593
rect 312604 512273 312646 512509
rect 312882 512273 312924 512509
rect 312604 512241 312924 512273
rect 328076 512829 328396 512861
rect 328076 512593 328118 512829
rect 328354 512593 328396 512829
rect 328076 512509 328396 512593
rect 328076 512273 328118 512509
rect 328354 512273 328396 512509
rect 328076 512241 328396 512273
rect 334340 512829 334660 512861
rect 334340 512593 334382 512829
rect 334618 512593 334660 512829
rect 334340 512509 334660 512593
rect 334340 512273 334382 512509
rect 334618 512273 334660 512509
rect 334340 512241 334660 512273
rect 340604 512829 340924 512861
rect 340604 512593 340646 512829
rect 340882 512593 340924 512829
rect 340604 512509 340924 512593
rect 340604 512273 340646 512509
rect 340882 512273 340924 512509
rect 340604 512241 340924 512273
rect 356076 512829 356396 512861
rect 356076 512593 356118 512829
rect 356354 512593 356396 512829
rect 356076 512509 356396 512593
rect 356076 512273 356118 512509
rect 356354 512273 356396 512509
rect 356076 512241 356396 512273
rect 275208 509454 275528 509486
rect 275208 509218 275250 509454
rect 275486 509218 275528 509454
rect 275208 509134 275528 509218
rect 275208 508898 275250 509134
rect 275486 508898 275528 509134
rect 275208 508866 275528 508898
rect 281472 509454 281792 509486
rect 281472 509218 281514 509454
rect 281750 509218 281792 509454
rect 281472 509134 281792 509218
rect 281472 508898 281514 509134
rect 281750 508898 281792 509134
rect 281472 508866 281792 508898
rect 303208 509454 303528 509486
rect 303208 509218 303250 509454
rect 303486 509218 303528 509454
rect 303208 509134 303528 509218
rect 303208 508898 303250 509134
rect 303486 508898 303528 509134
rect 303208 508866 303528 508898
rect 309472 509454 309792 509486
rect 309472 509218 309514 509454
rect 309750 509218 309792 509454
rect 309472 509134 309792 509218
rect 309472 508898 309514 509134
rect 309750 508898 309792 509134
rect 309472 508866 309792 508898
rect 331208 509454 331528 509486
rect 331208 509218 331250 509454
rect 331486 509218 331528 509454
rect 331208 509134 331528 509218
rect 331208 508898 331250 509134
rect 331486 508898 331528 509134
rect 331208 508866 331528 508898
rect 337472 509454 337792 509486
rect 337472 509218 337514 509454
rect 337750 509218 337792 509454
rect 337472 509134 337792 509218
rect 337472 508898 337514 509134
rect 337750 508898 337792 509134
rect 337472 508866 337792 508898
rect 359208 509454 359528 509486
rect 359208 509218 359250 509454
rect 359486 509218 359528 509454
rect 359208 509134 359528 509218
rect 359208 508898 359250 509134
rect 359486 508898 359528 509134
rect 359208 508866 359528 508898
rect 361622 500853 361682 522411
rect 408539 520844 408605 520845
rect 408539 520780 408540 520844
rect 408604 520780 408605 520844
rect 408539 520779 408605 520780
rect 372291 520708 372357 520709
rect 372291 520644 372292 520708
rect 372356 520644 372357 520708
rect 372291 520643 372357 520644
rect 362340 512829 362660 512861
rect 362340 512593 362382 512829
rect 362618 512593 362660 512829
rect 362340 512509 362660 512593
rect 362340 512273 362382 512509
rect 362618 512273 362660 512509
rect 362340 512241 362660 512273
rect 368604 512829 368924 512861
rect 368604 512593 368646 512829
rect 368882 512593 368924 512829
rect 372294 512821 372354 520643
rect 384076 512829 384396 512861
rect 372291 512820 372357 512821
rect 372291 512756 372292 512820
rect 372356 512756 372357 512820
rect 372291 512755 372357 512756
rect 368604 512509 368924 512593
rect 368604 512273 368646 512509
rect 368882 512273 368924 512509
rect 368604 512241 368924 512273
rect 384076 512593 384118 512829
rect 384354 512593 384396 512829
rect 384076 512509 384396 512593
rect 384076 512273 384118 512509
rect 384354 512273 384396 512509
rect 384076 512241 384396 512273
rect 390340 512829 390660 512861
rect 390340 512593 390382 512829
rect 390618 512593 390660 512829
rect 390340 512509 390660 512593
rect 390340 512273 390382 512509
rect 390618 512273 390660 512509
rect 390340 512241 390660 512273
rect 396604 512829 396924 512861
rect 396604 512593 396646 512829
rect 396882 512593 396924 512829
rect 408542 512821 408602 520779
rect 412076 512829 412396 512861
rect 408539 512820 408605 512821
rect 408539 512756 408540 512820
rect 408604 512756 408605 512820
rect 408539 512755 408605 512756
rect 396604 512509 396924 512593
rect 396604 512273 396646 512509
rect 396882 512273 396924 512509
rect 396604 512241 396924 512273
rect 412076 512593 412118 512829
rect 412354 512593 412396 512829
rect 412076 512509 412396 512593
rect 412076 512273 412118 512509
rect 412354 512273 412396 512509
rect 412076 512241 412396 512273
rect 418340 512829 418660 512861
rect 418340 512593 418382 512829
rect 418618 512593 418660 512829
rect 418340 512509 418660 512593
rect 418340 512273 418382 512509
rect 418618 512273 418660 512509
rect 418340 512241 418660 512273
rect 424604 512829 424924 512861
rect 424604 512593 424646 512829
rect 424882 512593 424924 512829
rect 424604 512509 424924 512593
rect 424604 512273 424646 512509
rect 424882 512273 424924 512509
rect 424604 512241 424924 512273
rect 440076 512829 440396 512861
rect 440076 512593 440118 512829
rect 440354 512593 440396 512829
rect 440076 512509 440396 512593
rect 440076 512273 440118 512509
rect 440354 512273 440396 512509
rect 440076 512241 440396 512273
rect 365472 509454 365792 509486
rect 365472 509218 365514 509454
rect 365750 509218 365792 509454
rect 365472 509134 365792 509218
rect 365472 508898 365514 509134
rect 365750 508898 365792 509134
rect 365472 508866 365792 508898
rect 387208 509454 387528 509486
rect 387208 509218 387250 509454
rect 387486 509218 387528 509454
rect 387208 509134 387528 509218
rect 387208 508898 387250 509134
rect 387486 508898 387528 509134
rect 387208 508866 387528 508898
rect 393472 509454 393792 509486
rect 393472 509218 393514 509454
rect 393750 509218 393792 509454
rect 393472 509134 393792 509218
rect 393472 508898 393514 509134
rect 393750 508898 393792 509134
rect 393472 508866 393792 508898
rect 415208 509454 415528 509486
rect 415208 509218 415250 509454
rect 415486 509218 415528 509454
rect 415208 509134 415528 509218
rect 415208 508898 415250 509134
rect 415486 508898 415528 509134
rect 415208 508866 415528 508898
rect 421472 509454 421792 509486
rect 421472 509218 421514 509454
rect 421750 509218 421792 509454
rect 421472 509134 421792 509218
rect 421472 508898 421514 509134
rect 421750 508898 421792 509134
rect 421472 508866 421792 508898
rect 443208 509454 443528 509486
rect 443208 509218 443250 509454
rect 443486 509218 443528 509454
rect 443208 509134 443528 509218
rect 443208 508898 443250 509134
rect 443486 508898 443528 509134
rect 443208 508866 443528 508898
rect 445710 500853 445770 522411
rect 484347 520980 484413 520981
rect 484347 520916 484348 520980
rect 484412 520916 484413 520980
rect 484347 520915 484413 520916
rect 446340 512829 446660 512861
rect 446340 512593 446382 512829
rect 446618 512593 446660 512829
rect 446340 512509 446660 512593
rect 446340 512273 446382 512509
rect 446618 512273 446660 512509
rect 446340 512241 446660 512273
rect 452604 512829 452924 512861
rect 452604 512593 452646 512829
rect 452882 512593 452924 512829
rect 452604 512509 452924 512593
rect 452604 512273 452646 512509
rect 452882 512273 452924 512509
rect 452604 512241 452924 512273
rect 468076 512829 468396 512861
rect 468076 512593 468118 512829
rect 468354 512593 468396 512829
rect 468076 512509 468396 512593
rect 468076 512273 468118 512509
rect 468354 512273 468396 512509
rect 468076 512241 468396 512273
rect 474340 512829 474660 512861
rect 474340 512593 474382 512829
rect 474618 512593 474660 512829
rect 474340 512509 474660 512593
rect 474340 512273 474382 512509
rect 474618 512273 474660 512509
rect 474340 512241 474660 512273
rect 480604 512829 480924 512861
rect 480604 512593 480646 512829
rect 480882 512593 480924 512829
rect 484350 512821 484410 520915
rect 492811 520844 492877 520845
rect 492811 520780 492812 520844
rect 492876 520780 492877 520844
rect 492811 520779 492877 520780
rect 492814 518910 492874 520779
rect 520595 520708 520661 520709
rect 520595 520644 520596 520708
rect 520660 520644 520661 520708
rect 520595 520643 520661 520644
rect 492630 518850 492874 518910
rect 492630 512821 492690 518850
rect 496076 512829 496396 512861
rect 484347 512820 484413 512821
rect 484347 512756 484348 512820
rect 484412 512756 484413 512820
rect 484347 512755 484413 512756
rect 492627 512820 492693 512821
rect 492627 512756 492628 512820
rect 492692 512756 492693 512820
rect 492627 512755 492693 512756
rect 480604 512509 480924 512593
rect 480604 512273 480646 512509
rect 480882 512273 480924 512509
rect 480604 512241 480924 512273
rect 496076 512593 496118 512829
rect 496354 512593 496396 512829
rect 496076 512509 496396 512593
rect 496076 512273 496118 512509
rect 496354 512273 496396 512509
rect 496076 512241 496396 512273
rect 502340 512829 502660 512861
rect 502340 512593 502382 512829
rect 502618 512593 502660 512829
rect 502340 512509 502660 512593
rect 502340 512273 502382 512509
rect 502618 512273 502660 512509
rect 502340 512241 502660 512273
rect 508604 512829 508924 512861
rect 508604 512593 508646 512829
rect 508882 512593 508924 512829
rect 520598 512821 520658 520643
rect 524076 512829 524396 512861
rect 520595 512820 520661 512821
rect 520595 512756 520596 512820
rect 520660 512756 520661 512820
rect 520595 512755 520661 512756
rect 508604 512509 508924 512593
rect 508604 512273 508646 512509
rect 508882 512273 508924 512509
rect 508604 512241 508924 512273
rect 524076 512593 524118 512829
rect 524354 512593 524396 512829
rect 524076 512509 524396 512593
rect 524076 512273 524118 512509
rect 524354 512273 524396 512509
rect 524076 512241 524396 512273
rect 530340 512829 530660 512861
rect 530340 512593 530382 512829
rect 530618 512593 530660 512829
rect 530340 512509 530660 512593
rect 530340 512273 530382 512509
rect 530618 512273 530660 512509
rect 530340 512241 530660 512273
rect 536604 512829 536924 512861
rect 536604 512593 536646 512829
rect 536882 512593 536924 512829
rect 536604 512509 536924 512593
rect 536604 512273 536646 512509
rect 536882 512273 536924 512509
rect 536604 512241 536924 512273
rect 552076 512829 552396 512861
rect 552076 512593 552118 512829
rect 552354 512593 552396 512829
rect 552076 512509 552396 512593
rect 552076 512273 552118 512509
rect 552354 512273 552396 512509
rect 552076 512241 552396 512273
rect 449472 509454 449792 509486
rect 449472 509218 449514 509454
rect 449750 509218 449792 509454
rect 449472 509134 449792 509218
rect 449472 508898 449514 509134
rect 449750 508898 449792 509134
rect 449472 508866 449792 508898
rect 471208 509454 471528 509486
rect 471208 509218 471250 509454
rect 471486 509218 471528 509454
rect 471208 509134 471528 509218
rect 471208 508898 471250 509134
rect 471486 508898 471528 509134
rect 471208 508866 471528 508898
rect 477472 509454 477792 509486
rect 477472 509218 477514 509454
rect 477750 509218 477792 509454
rect 477472 509134 477792 509218
rect 477472 508898 477514 509134
rect 477750 508898 477792 509134
rect 477472 508866 477792 508898
rect 499208 509454 499528 509486
rect 499208 509218 499250 509454
rect 499486 509218 499528 509454
rect 499208 509134 499528 509218
rect 499208 508898 499250 509134
rect 499486 508898 499528 509134
rect 499208 508866 499528 508898
rect 505472 509454 505792 509486
rect 505472 509218 505514 509454
rect 505750 509218 505792 509454
rect 505472 509134 505792 509218
rect 505472 508898 505514 509134
rect 505750 508898 505792 509134
rect 505472 508866 505792 508898
rect 527208 509454 527528 509486
rect 527208 509218 527250 509454
rect 527486 509218 527528 509454
rect 527208 509134 527528 509218
rect 527208 508898 527250 509134
rect 527486 508898 527528 509134
rect 527208 508866 527528 508898
rect 533472 509454 533792 509486
rect 533472 509218 533514 509454
rect 533750 509218 533792 509454
rect 533472 509134 533792 509218
rect 533472 508898 533514 509134
rect 533750 508898 533792 509134
rect 533472 508866 533792 508898
rect 555208 509454 555528 509486
rect 555208 509218 555250 509454
rect 555486 509218 555528 509454
rect 555208 509134 555528 509218
rect 555208 508898 555250 509134
rect 555486 508898 555528 509134
rect 555208 508866 555528 508898
rect 557582 500853 557642 522411
rect 558340 512829 558660 512861
rect 558340 512593 558382 512829
rect 558618 512593 558660 512829
rect 558340 512509 558660 512593
rect 558340 512273 558382 512509
rect 558618 512273 558660 512509
rect 558340 512241 558660 512273
rect 564604 512829 564924 512861
rect 564604 512593 564646 512829
rect 564882 512593 564924 512829
rect 564604 512509 564924 512593
rect 564604 512273 564646 512509
rect 564882 512273 564924 512509
rect 564604 512241 564924 512273
rect 573494 512829 574114 539273
rect 573494 512593 573526 512829
rect 573762 512593 573846 512829
rect 574082 512593 574114 512829
rect 573494 512509 574114 512593
rect 573494 512273 573526 512509
rect 573762 512273 573846 512509
rect 574082 512273 574114 512509
rect 561472 509454 561792 509486
rect 561472 509218 561514 509454
rect 561750 509218 561792 509454
rect 561472 509134 561792 509218
rect 561472 508898 561514 509134
rect 561750 508898 561792 509134
rect 561472 508866 561792 508898
rect 165659 500852 165725 500853
rect 165659 500788 165660 500852
rect 165724 500788 165725 500852
rect 165659 500787 165725 500788
rect 259499 500852 259565 500853
rect 259499 500788 259500 500852
rect 259564 500788 259565 500852
rect 259499 500787 259565 500788
rect 361619 500852 361685 500853
rect 361619 500788 361620 500852
rect 361684 500788 361685 500852
rect 361619 500787 361685 500788
rect 445707 500852 445773 500853
rect 445707 500788 445708 500852
rect 445772 500788 445773 500852
rect 445707 500787 445773 500788
rect 557579 500852 557645 500853
rect 557579 500788 557580 500852
rect 557644 500788 557645 500852
rect 557579 500787 557645 500788
rect 194731 495548 194797 495549
rect 194731 495484 194732 495548
rect 194796 495484 194797 495548
rect 194731 495483 194797 495484
rect 390875 495548 390941 495549
rect 390875 495484 390876 495548
rect 390940 495484 390941 495548
rect 390875 495483 390941 495484
rect 128307 495276 128373 495277
rect 128307 495212 128308 495276
rect 128372 495212 128373 495276
rect 128307 495211 128373 495212
rect -2006 485593 -1974 485829
rect -1738 485593 -1654 485829
rect -1418 485593 -1386 485829
rect -2006 485509 -1386 485593
rect -2006 485273 -1974 485509
rect -1738 485273 -1654 485509
rect -1418 485273 -1386 485509
rect -2006 458829 -1386 485273
rect 20076 485829 20396 485861
rect 20076 485593 20118 485829
rect 20354 485593 20396 485829
rect 20076 485509 20396 485593
rect 20076 485273 20118 485509
rect 20354 485273 20396 485509
rect 20076 485241 20396 485273
rect 26340 485829 26660 485861
rect 26340 485593 26382 485829
rect 26618 485593 26660 485829
rect 26340 485509 26660 485593
rect 26340 485273 26382 485509
rect 26618 485273 26660 485509
rect 26340 485241 26660 485273
rect 32604 485829 32924 485861
rect 32604 485593 32646 485829
rect 32882 485593 32924 485829
rect 32604 485509 32924 485593
rect 32604 485273 32646 485509
rect 32882 485273 32924 485509
rect 32604 485241 32924 485273
rect 48076 485829 48396 485861
rect 48076 485593 48118 485829
rect 48354 485593 48396 485829
rect 48076 485509 48396 485593
rect 48076 485273 48118 485509
rect 48354 485273 48396 485509
rect 48076 485241 48396 485273
rect 54340 485829 54660 485861
rect 54340 485593 54382 485829
rect 54618 485593 54660 485829
rect 54340 485509 54660 485593
rect 54340 485273 54382 485509
rect 54618 485273 54660 485509
rect 54340 485241 54660 485273
rect 60604 485829 60924 485861
rect 60604 485593 60646 485829
rect 60882 485593 60924 485829
rect 60604 485509 60924 485593
rect 60604 485273 60646 485509
rect 60882 485273 60924 485509
rect 60604 485241 60924 485273
rect 76076 485829 76396 485861
rect 76076 485593 76118 485829
rect 76354 485593 76396 485829
rect 76076 485509 76396 485593
rect 76076 485273 76118 485509
rect 76354 485273 76396 485509
rect 76076 485241 76396 485273
rect 82340 485829 82660 485861
rect 82340 485593 82382 485829
rect 82618 485593 82660 485829
rect 82340 485509 82660 485593
rect 82340 485273 82382 485509
rect 82618 485273 82660 485509
rect 82340 485241 82660 485273
rect 88604 485829 88924 485861
rect 88604 485593 88646 485829
rect 88882 485593 88924 485829
rect 88604 485509 88924 485593
rect 88604 485273 88646 485509
rect 88882 485273 88924 485509
rect 88604 485241 88924 485273
rect 104076 485829 104396 485861
rect 104076 485593 104118 485829
rect 104354 485593 104396 485829
rect 104076 485509 104396 485593
rect 104076 485273 104118 485509
rect 104354 485273 104396 485509
rect 104076 485241 104396 485273
rect 110340 485829 110660 485861
rect 110340 485593 110382 485829
rect 110618 485593 110660 485829
rect 110340 485509 110660 485593
rect 110340 485273 110382 485509
rect 110618 485273 110660 485509
rect 110340 485241 110660 485273
rect 116604 485829 116924 485861
rect 116604 485593 116646 485829
rect 116882 485593 116924 485829
rect 116604 485509 116924 485593
rect 116604 485273 116646 485509
rect 116882 485273 116924 485509
rect 116604 485241 116924 485273
rect 64459 485212 64525 485213
rect 64459 485148 64460 485212
rect 64524 485148 64525 485212
rect 64459 485147 64525 485148
rect 92427 485212 92493 485213
rect 92427 485148 92428 485212
rect 92492 485148 92493 485212
rect 92427 485147 92493 485148
rect 23208 482454 23528 482486
rect 23208 482218 23250 482454
rect 23486 482218 23528 482454
rect 23208 482134 23528 482218
rect 23208 481898 23250 482134
rect 23486 481898 23528 482134
rect 23208 481866 23528 481898
rect 29472 482454 29792 482486
rect 29472 482218 29514 482454
rect 29750 482218 29792 482454
rect 29472 482134 29792 482218
rect 29472 481898 29514 482134
rect 29750 481898 29792 482134
rect 29472 481866 29792 481898
rect 51208 482454 51528 482486
rect 51208 482218 51250 482454
rect 51486 482218 51528 482454
rect 51208 482134 51528 482218
rect 51208 481898 51250 482134
rect 51486 481898 51528 482134
rect 51208 481866 51528 481898
rect 57472 482454 57792 482486
rect 57472 482218 57514 482454
rect 57750 482218 57792 482454
rect 57472 482134 57792 482218
rect 57472 481898 57514 482134
rect 57750 481898 57792 482134
rect 57472 481866 57792 481898
rect 64462 477325 64522 485147
rect 79208 482454 79528 482486
rect 79208 482218 79250 482454
rect 79486 482218 79528 482454
rect 79208 482134 79528 482218
rect 79208 481898 79250 482134
rect 79486 481898 79528 482134
rect 79208 481866 79528 481898
rect 85472 482454 85792 482486
rect 85472 482218 85514 482454
rect 85750 482218 85792 482454
rect 85472 482134 85792 482218
rect 85472 481898 85514 482134
rect 85750 481898 85792 482134
rect 85472 481866 85792 481898
rect 64459 477324 64525 477325
rect 64459 477260 64460 477324
rect 64524 477260 64525 477324
rect 64459 477259 64525 477260
rect 92430 477189 92490 485147
rect 107208 482454 107528 482486
rect 107208 482218 107250 482454
rect 107486 482218 107528 482454
rect 107208 482134 107528 482218
rect 107208 481898 107250 482134
rect 107486 481898 107528 482134
rect 107208 481866 107528 481898
rect 113472 482454 113792 482486
rect 113472 482218 113514 482454
rect 113750 482218 113792 482454
rect 113472 482134 113792 482218
rect 113472 481898 113514 482134
rect 113750 481898 113792 482134
rect 113472 481866 113792 481898
rect 92427 477188 92493 477189
rect 92427 477124 92428 477188
rect 92492 477124 92493 477188
rect 92427 477123 92493 477124
rect 128310 473245 128370 495211
rect 132076 485829 132396 485861
rect 132076 485593 132118 485829
rect 132354 485593 132396 485829
rect 132076 485509 132396 485593
rect 132076 485273 132118 485509
rect 132354 485273 132396 485509
rect 132076 485241 132396 485273
rect 138340 485829 138660 485861
rect 138340 485593 138382 485829
rect 138618 485593 138660 485829
rect 138340 485509 138660 485593
rect 138340 485273 138382 485509
rect 138618 485273 138660 485509
rect 138340 485241 138660 485273
rect 144604 485829 144924 485861
rect 144604 485593 144646 485829
rect 144882 485593 144924 485829
rect 144604 485509 144924 485593
rect 144604 485273 144646 485509
rect 144882 485273 144924 485509
rect 144604 485241 144924 485273
rect 160076 485829 160396 485861
rect 160076 485593 160118 485829
rect 160354 485593 160396 485829
rect 160076 485509 160396 485593
rect 160076 485273 160118 485509
rect 160354 485273 160396 485509
rect 160076 485241 160396 485273
rect 166340 485829 166660 485861
rect 166340 485593 166382 485829
rect 166618 485593 166660 485829
rect 166340 485509 166660 485593
rect 166340 485273 166382 485509
rect 166618 485273 166660 485509
rect 166340 485241 166660 485273
rect 172604 485829 172924 485861
rect 172604 485593 172646 485829
rect 172882 485593 172924 485829
rect 172604 485509 172924 485593
rect 172604 485273 172646 485509
rect 172882 485273 172924 485509
rect 172604 485241 172924 485273
rect 188076 485829 188396 485861
rect 188076 485593 188118 485829
rect 188354 485593 188396 485829
rect 188076 485509 188396 485593
rect 188076 485273 188118 485509
rect 188354 485273 188396 485509
rect 188076 485241 188396 485273
rect 194340 485829 194660 485861
rect 194340 485593 194382 485829
rect 194618 485593 194660 485829
rect 194340 485509 194660 485593
rect 194340 485273 194382 485509
rect 194618 485273 194660 485509
rect 194340 485241 194660 485273
rect 148363 485212 148429 485213
rect 148363 485148 148364 485212
rect 148428 485148 148429 485212
rect 148363 485147 148429 485148
rect 176331 485212 176397 485213
rect 176331 485148 176332 485212
rect 176396 485148 176397 485212
rect 176331 485147 176397 485148
rect 135208 482454 135528 482486
rect 135208 482218 135250 482454
rect 135486 482218 135528 482454
rect 135208 482134 135528 482218
rect 135208 481898 135250 482134
rect 135486 481898 135528 482134
rect 135208 481866 135528 481898
rect 141472 482454 141792 482486
rect 141472 482218 141514 482454
rect 141750 482218 141792 482454
rect 141472 482134 141792 482218
rect 141472 481898 141514 482134
rect 141750 481898 141792 482134
rect 141472 481866 141792 481898
rect 148366 477189 148426 485147
rect 163208 482454 163528 482486
rect 163208 482218 163250 482454
rect 163486 482218 163528 482454
rect 163208 482134 163528 482218
rect 163208 481898 163250 482134
rect 163486 481898 163528 482134
rect 163208 481866 163528 481898
rect 169472 482454 169792 482486
rect 169472 482218 169514 482454
rect 169750 482218 169792 482454
rect 169472 482134 169792 482218
rect 169472 481898 169514 482134
rect 169750 481898 169792 482134
rect 169472 481866 169792 481898
rect 176334 477325 176394 485147
rect 191208 482454 191528 482486
rect 191208 482218 191250 482454
rect 191486 482218 191528 482454
rect 191208 482134 191528 482218
rect 191208 481898 191250 482134
rect 191486 481898 191528 482134
rect 191208 481866 191528 481898
rect 176331 477324 176397 477325
rect 176331 477260 176332 477324
rect 176396 477260 176397 477324
rect 176331 477259 176397 477260
rect 148363 477188 148429 477189
rect 148363 477124 148364 477188
rect 148428 477124 148429 477188
rect 148363 477123 148429 477124
rect 194734 473245 194794 495483
rect 200604 485829 200924 485861
rect 200604 485593 200646 485829
rect 200882 485593 200924 485829
rect 200604 485509 200924 485593
rect 200604 485273 200646 485509
rect 200882 485273 200924 485509
rect 200604 485241 200924 485273
rect 216076 485829 216396 485861
rect 216076 485593 216118 485829
rect 216354 485593 216396 485829
rect 216076 485509 216396 485593
rect 216076 485273 216118 485509
rect 216354 485273 216396 485509
rect 216076 485241 216396 485273
rect 222340 485829 222660 485861
rect 222340 485593 222382 485829
rect 222618 485593 222660 485829
rect 222340 485509 222660 485593
rect 222340 485273 222382 485509
rect 222618 485273 222660 485509
rect 222340 485241 222660 485273
rect 228604 485829 228924 485861
rect 228604 485593 228646 485829
rect 228882 485593 228924 485829
rect 228604 485509 228924 485593
rect 228604 485273 228646 485509
rect 228882 485273 228924 485509
rect 228604 485241 228924 485273
rect 244076 485829 244396 485861
rect 244076 485593 244118 485829
rect 244354 485593 244396 485829
rect 244076 485509 244396 485593
rect 244076 485273 244118 485509
rect 244354 485273 244396 485509
rect 244076 485241 244396 485273
rect 250340 485829 250660 485861
rect 250340 485593 250382 485829
rect 250618 485593 250660 485829
rect 250340 485509 250660 485593
rect 250340 485273 250382 485509
rect 250618 485273 250660 485509
rect 250340 485241 250660 485273
rect 256604 485829 256924 485861
rect 256604 485593 256646 485829
rect 256882 485593 256924 485829
rect 256604 485509 256924 485593
rect 256604 485273 256646 485509
rect 256882 485273 256924 485509
rect 256604 485241 256924 485273
rect 272076 485829 272396 485861
rect 272076 485593 272118 485829
rect 272354 485593 272396 485829
rect 272076 485509 272396 485593
rect 272076 485273 272118 485509
rect 272354 485273 272396 485509
rect 272076 485241 272396 485273
rect 278340 485829 278660 485861
rect 278340 485593 278382 485829
rect 278618 485593 278660 485829
rect 278340 485509 278660 485593
rect 278340 485273 278382 485509
rect 278618 485273 278660 485509
rect 278340 485241 278660 485273
rect 284604 485829 284924 485861
rect 284604 485593 284646 485829
rect 284882 485593 284924 485829
rect 284604 485509 284924 485593
rect 284604 485273 284646 485509
rect 284882 485273 284924 485509
rect 284604 485241 284924 485273
rect 300076 485829 300396 485861
rect 300076 485593 300118 485829
rect 300354 485593 300396 485829
rect 300076 485509 300396 485593
rect 300076 485273 300118 485509
rect 300354 485273 300396 485509
rect 300076 485241 300396 485273
rect 306340 485829 306660 485861
rect 306340 485593 306382 485829
rect 306618 485593 306660 485829
rect 306340 485509 306660 485593
rect 306340 485273 306382 485509
rect 306618 485273 306660 485509
rect 306340 485241 306660 485273
rect 312604 485829 312924 485861
rect 312604 485593 312646 485829
rect 312882 485593 312924 485829
rect 312604 485509 312924 485593
rect 312604 485273 312646 485509
rect 312882 485273 312924 485509
rect 312604 485241 312924 485273
rect 328076 485829 328396 485861
rect 328076 485593 328118 485829
rect 328354 485593 328396 485829
rect 328076 485509 328396 485593
rect 328076 485273 328118 485509
rect 328354 485273 328396 485509
rect 328076 485241 328396 485273
rect 334340 485829 334660 485861
rect 334340 485593 334382 485829
rect 334618 485593 334660 485829
rect 334340 485509 334660 485593
rect 334340 485273 334382 485509
rect 334618 485273 334660 485509
rect 334340 485241 334660 485273
rect 340604 485829 340924 485861
rect 340604 485593 340646 485829
rect 340882 485593 340924 485829
rect 340604 485509 340924 485593
rect 340604 485273 340646 485509
rect 340882 485273 340924 485509
rect 340604 485241 340924 485273
rect 356076 485829 356396 485861
rect 356076 485593 356118 485829
rect 356354 485593 356396 485829
rect 356076 485509 356396 485593
rect 356076 485273 356118 485509
rect 356354 485273 356396 485509
rect 356076 485241 356396 485273
rect 362340 485829 362660 485861
rect 362340 485593 362382 485829
rect 362618 485593 362660 485829
rect 362340 485509 362660 485593
rect 362340 485273 362382 485509
rect 362618 485273 362660 485509
rect 362340 485241 362660 485273
rect 368604 485829 368924 485861
rect 368604 485593 368646 485829
rect 368882 485593 368924 485829
rect 368604 485509 368924 485593
rect 368604 485273 368646 485509
rect 368882 485273 368924 485509
rect 368604 485241 368924 485273
rect 384076 485829 384396 485861
rect 384076 485593 384118 485829
rect 384354 485593 384396 485829
rect 384076 485509 384396 485593
rect 384076 485273 384118 485509
rect 384354 485273 384396 485509
rect 384076 485241 384396 485273
rect 390340 485829 390660 485861
rect 390340 485593 390382 485829
rect 390618 485593 390660 485829
rect 390340 485509 390660 485593
rect 390340 485273 390382 485509
rect 390618 485273 390660 485509
rect 390340 485241 390660 485273
rect 212579 485212 212645 485213
rect 212579 485148 212580 485212
rect 212644 485148 212645 485212
rect 212579 485147 212645 485148
rect 288387 485212 288453 485213
rect 288387 485148 288388 485212
rect 288452 485148 288453 485212
rect 288387 485147 288453 485148
rect 296483 485212 296549 485213
rect 296483 485148 296484 485212
rect 296548 485148 296549 485212
rect 296483 485147 296549 485148
rect 372291 485212 372357 485213
rect 372291 485148 372292 485212
rect 372356 485148 372357 485212
rect 372291 485147 372357 485148
rect 197472 482454 197792 482486
rect 197472 482218 197514 482454
rect 197750 482218 197792 482454
rect 197472 482134 197792 482218
rect 197472 481898 197514 482134
rect 197750 481898 197792 482134
rect 197472 481866 197792 481898
rect 212582 477189 212642 485147
rect 219208 482454 219528 482486
rect 219208 482218 219250 482454
rect 219486 482218 219528 482454
rect 219208 482134 219528 482218
rect 219208 481898 219250 482134
rect 219486 481898 219528 482134
rect 219208 481866 219528 481898
rect 225472 482454 225792 482486
rect 225472 482218 225514 482454
rect 225750 482218 225792 482454
rect 225472 482134 225792 482218
rect 225472 481898 225514 482134
rect 225750 481898 225792 482134
rect 225472 481866 225792 481898
rect 247208 482454 247528 482486
rect 247208 482218 247250 482454
rect 247486 482218 247528 482454
rect 247208 482134 247528 482218
rect 247208 481898 247250 482134
rect 247486 481898 247528 482134
rect 247208 481866 247528 481898
rect 253472 482454 253792 482486
rect 253472 482218 253514 482454
rect 253750 482218 253792 482454
rect 253472 482134 253792 482218
rect 253472 481898 253514 482134
rect 253750 481898 253792 482134
rect 253472 481866 253792 481898
rect 275208 482454 275528 482486
rect 275208 482218 275250 482454
rect 275486 482218 275528 482454
rect 275208 482134 275528 482218
rect 275208 481898 275250 482134
rect 275486 481898 275528 482134
rect 275208 481866 275528 481898
rect 281472 482454 281792 482486
rect 281472 482218 281514 482454
rect 281750 482218 281792 482454
rect 281472 482134 281792 482218
rect 281472 481898 281514 482134
rect 281750 481898 281792 482134
rect 281472 481866 281792 481898
rect 212579 477188 212645 477189
rect 212579 477124 212580 477188
rect 212644 477124 212645 477188
rect 212579 477123 212645 477124
rect 288390 477053 288450 485147
rect 296486 483030 296546 485147
rect 296486 482970 296914 483030
rect 296854 477189 296914 482970
rect 303208 482454 303528 482486
rect 303208 482218 303250 482454
rect 303486 482218 303528 482454
rect 303208 482134 303528 482218
rect 303208 481898 303250 482134
rect 303486 481898 303528 482134
rect 303208 481866 303528 481898
rect 309472 482454 309792 482486
rect 309472 482218 309514 482454
rect 309750 482218 309792 482454
rect 309472 482134 309792 482218
rect 309472 481898 309514 482134
rect 309750 481898 309792 482134
rect 309472 481866 309792 481898
rect 331208 482454 331528 482486
rect 331208 482218 331250 482454
rect 331486 482218 331528 482454
rect 331208 482134 331528 482218
rect 331208 481898 331250 482134
rect 331486 481898 331528 482134
rect 331208 481866 331528 481898
rect 337472 482454 337792 482486
rect 337472 482218 337514 482454
rect 337750 482218 337792 482454
rect 337472 482134 337792 482218
rect 337472 481898 337514 482134
rect 337750 481898 337792 482134
rect 337472 481866 337792 481898
rect 359208 482454 359528 482486
rect 359208 482218 359250 482454
rect 359486 482218 359528 482454
rect 359208 482134 359528 482218
rect 359208 481898 359250 482134
rect 359486 481898 359528 482134
rect 359208 481866 359528 481898
rect 365472 482454 365792 482486
rect 365472 482218 365514 482454
rect 365750 482218 365792 482454
rect 365472 482134 365792 482218
rect 365472 481898 365514 482134
rect 365750 481898 365792 482134
rect 365472 481866 365792 481898
rect 296851 477188 296917 477189
rect 296851 477124 296852 477188
rect 296916 477124 296917 477188
rect 296851 477123 296917 477124
rect 372294 477053 372354 485147
rect 387208 482454 387528 482486
rect 387208 482218 387250 482454
rect 387486 482218 387528 482454
rect 387208 482134 387528 482218
rect 387208 481898 387250 482134
rect 387486 481898 387528 482134
rect 387208 481866 387528 481898
rect 288387 477052 288453 477053
rect 288387 476988 288388 477052
rect 288452 476988 288453 477052
rect 288387 476987 288453 476988
rect 372291 477052 372357 477053
rect 372291 476988 372292 477052
rect 372356 476988 372357 477052
rect 372291 476987 372357 476988
rect 390878 473245 390938 495483
rect 396604 485829 396924 485861
rect 396604 485593 396646 485829
rect 396882 485593 396924 485829
rect 396604 485509 396924 485593
rect 396604 485273 396646 485509
rect 396882 485273 396924 485509
rect 396604 485241 396924 485273
rect 412076 485829 412396 485861
rect 412076 485593 412118 485829
rect 412354 485593 412396 485829
rect 412076 485509 412396 485593
rect 412076 485273 412118 485509
rect 412354 485273 412396 485509
rect 412076 485241 412396 485273
rect 418340 485829 418660 485861
rect 418340 485593 418382 485829
rect 418618 485593 418660 485829
rect 418340 485509 418660 485593
rect 418340 485273 418382 485509
rect 418618 485273 418660 485509
rect 418340 485241 418660 485273
rect 424604 485829 424924 485861
rect 424604 485593 424646 485829
rect 424882 485593 424924 485829
rect 424604 485509 424924 485593
rect 424604 485273 424646 485509
rect 424882 485273 424924 485509
rect 424604 485241 424924 485273
rect 440076 485829 440396 485861
rect 440076 485593 440118 485829
rect 440354 485593 440396 485829
rect 440076 485509 440396 485593
rect 440076 485273 440118 485509
rect 440354 485273 440396 485509
rect 440076 485241 440396 485273
rect 446340 485829 446660 485861
rect 446340 485593 446382 485829
rect 446618 485593 446660 485829
rect 446340 485509 446660 485593
rect 446340 485273 446382 485509
rect 446618 485273 446660 485509
rect 446340 485241 446660 485273
rect 452604 485829 452924 485861
rect 452604 485593 452646 485829
rect 452882 485593 452924 485829
rect 452604 485509 452924 485593
rect 452604 485273 452646 485509
rect 452882 485273 452924 485509
rect 452604 485241 452924 485273
rect 468076 485829 468396 485861
rect 468076 485593 468118 485829
rect 468354 485593 468396 485829
rect 468076 485509 468396 485593
rect 468076 485273 468118 485509
rect 468354 485273 468396 485509
rect 468076 485241 468396 485273
rect 474340 485829 474660 485861
rect 474340 485593 474382 485829
rect 474618 485593 474660 485829
rect 474340 485509 474660 485593
rect 474340 485273 474382 485509
rect 474618 485273 474660 485509
rect 474340 485241 474660 485273
rect 480604 485829 480924 485861
rect 480604 485593 480646 485829
rect 480882 485593 480924 485829
rect 480604 485509 480924 485593
rect 480604 485273 480646 485509
rect 480882 485273 480924 485509
rect 480604 485241 480924 485273
rect 496076 485829 496396 485861
rect 496076 485593 496118 485829
rect 496354 485593 496396 485829
rect 496076 485509 496396 485593
rect 496076 485273 496118 485509
rect 496354 485273 496396 485509
rect 496076 485241 496396 485273
rect 502340 485829 502660 485861
rect 502340 485593 502382 485829
rect 502618 485593 502660 485829
rect 502340 485509 502660 485593
rect 502340 485273 502382 485509
rect 502618 485273 502660 485509
rect 502340 485241 502660 485273
rect 508604 485829 508924 485861
rect 508604 485593 508646 485829
rect 508882 485593 508924 485829
rect 508604 485509 508924 485593
rect 508604 485273 508646 485509
rect 508882 485273 508924 485509
rect 508604 485241 508924 485273
rect 524076 485829 524396 485861
rect 524076 485593 524118 485829
rect 524354 485593 524396 485829
rect 524076 485509 524396 485593
rect 524076 485273 524118 485509
rect 524354 485273 524396 485509
rect 524076 485241 524396 485273
rect 530340 485829 530660 485861
rect 530340 485593 530382 485829
rect 530618 485593 530660 485829
rect 530340 485509 530660 485593
rect 530340 485273 530382 485509
rect 530618 485273 530660 485509
rect 530340 485241 530660 485273
rect 536604 485829 536924 485861
rect 536604 485593 536646 485829
rect 536882 485593 536924 485829
rect 536604 485509 536924 485593
rect 536604 485273 536646 485509
rect 536882 485273 536924 485509
rect 536604 485241 536924 485273
rect 552076 485829 552396 485861
rect 552076 485593 552118 485829
rect 552354 485593 552396 485829
rect 552076 485509 552396 485593
rect 552076 485273 552118 485509
rect 552354 485273 552396 485509
rect 552076 485241 552396 485273
rect 558340 485829 558660 485861
rect 558340 485593 558382 485829
rect 558618 485593 558660 485829
rect 558340 485509 558660 485593
rect 558340 485273 558382 485509
rect 558618 485273 558660 485509
rect 558340 485241 558660 485273
rect 564604 485829 564924 485861
rect 564604 485593 564646 485829
rect 564882 485593 564924 485829
rect 564604 485509 564924 485593
rect 564604 485273 564646 485509
rect 564882 485273 564924 485509
rect 564604 485241 564924 485273
rect 573494 485829 574114 512273
rect 573494 485593 573526 485829
rect 573762 485593 573846 485829
rect 574082 485593 574114 485829
rect 573494 485509 574114 485593
rect 573494 485273 573526 485509
rect 573762 485273 573846 485509
rect 574082 485273 574114 485509
rect 408539 485212 408605 485213
rect 408539 485148 408540 485212
rect 408604 485148 408605 485212
rect 408539 485147 408605 485148
rect 484347 485212 484413 485213
rect 484347 485148 484348 485212
rect 484412 485148 484413 485212
rect 484347 485147 484413 485148
rect 520595 485212 520661 485213
rect 520595 485148 520596 485212
rect 520660 485148 520661 485212
rect 520595 485147 520661 485148
rect 540467 485212 540533 485213
rect 540467 485148 540468 485212
rect 540532 485148 540533 485212
rect 540467 485147 540533 485148
rect 393472 482454 393792 482486
rect 393472 482218 393514 482454
rect 393750 482218 393792 482454
rect 393472 482134 393792 482218
rect 393472 481898 393514 482134
rect 393750 481898 393792 482134
rect 393472 481866 393792 481898
rect 408542 477325 408602 485147
rect 415208 482454 415528 482486
rect 415208 482218 415250 482454
rect 415486 482218 415528 482454
rect 415208 482134 415528 482218
rect 415208 481898 415250 482134
rect 415486 481898 415528 482134
rect 415208 481866 415528 481898
rect 421472 482454 421792 482486
rect 421472 482218 421514 482454
rect 421750 482218 421792 482454
rect 421472 482134 421792 482218
rect 421472 481898 421514 482134
rect 421750 481898 421792 482134
rect 421472 481866 421792 481898
rect 443208 482454 443528 482486
rect 443208 482218 443250 482454
rect 443486 482218 443528 482454
rect 443208 482134 443528 482218
rect 443208 481898 443250 482134
rect 443486 481898 443528 482134
rect 443208 481866 443528 481898
rect 449472 482454 449792 482486
rect 449472 482218 449514 482454
rect 449750 482218 449792 482454
rect 449472 482134 449792 482218
rect 449472 481898 449514 482134
rect 449750 481898 449792 482134
rect 449472 481866 449792 481898
rect 471208 482454 471528 482486
rect 471208 482218 471250 482454
rect 471486 482218 471528 482454
rect 471208 482134 471528 482218
rect 471208 481898 471250 482134
rect 471486 481898 471528 482134
rect 471208 481866 471528 481898
rect 477472 482454 477792 482486
rect 477472 482218 477514 482454
rect 477750 482218 477792 482454
rect 477472 482134 477792 482218
rect 477472 481898 477514 482134
rect 477750 481898 477792 482134
rect 477472 481866 477792 481898
rect 408539 477324 408605 477325
rect 408539 477260 408540 477324
rect 408604 477260 408605 477324
rect 408539 477259 408605 477260
rect 484350 477189 484410 485147
rect 499208 482454 499528 482486
rect 499208 482218 499250 482454
rect 499486 482218 499528 482454
rect 499208 482134 499528 482218
rect 499208 481898 499250 482134
rect 499486 481898 499528 482134
rect 499208 481866 499528 481898
rect 505472 482454 505792 482486
rect 505472 482218 505514 482454
rect 505750 482218 505792 482454
rect 505472 482134 505792 482218
rect 505472 481898 505514 482134
rect 505750 481898 505792 482134
rect 505472 481866 505792 481898
rect 520598 477325 520658 485147
rect 527208 482454 527528 482486
rect 527208 482218 527250 482454
rect 527486 482218 527528 482454
rect 527208 482134 527528 482218
rect 527208 481898 527250 482134
rect 527486 481898 527528 482134
rect 527208 481866 527528 481898
rect 533472 482454 533792 482486
rect 533472 482218 533514 482454
rect 533750 482218 533792 482454
rect 533472 482134 533792 482218
rect 533472 481898 533514 482134
rect 533750 481898 533792 482134
rect 533472 481866 533792 481898
rect 520595 477324 520661 477325
rect 520595 477260 520596 477324
rect 520660 477260 520661 477324
rect 520595 477259 520661 477260
rect 540470 477189 540530 485147
rect 555208 482454 555528 482486
rect 555208 482218 555250 482454
rect 555486 482218 555528 482454
rect 555208 482134 555528 482218
rect 555208 481898 555250 482134
rect 555486 481898 555528 482134
rect 555208 481866 555528 481898
rect 561472 482454 561792 482486
rect 561472 482218 561514 482454
rect 561750 482218 561792 482454
rect 561472 482134 561792 482218
rect 561472 481898 561514 482134
rect 561750 481898 561792 482134
rect 561472 481866 561792 481898
rect 484347 477188 484413 477189
rect 484347 477124 484348 477188
rect 484412 477124 484413 477188
rect 484347 477123 484413 477124
rect 540467 477188 540533 477189
rect 540467 477124 540468 477188
rect 540532 477124 540533 477188
rect 540467 477123 540533 477124
rect 128307 473244 128373 473245
rect 128307 473180 128308 473244
rect 128372 473180 128373 473244
rect 128307 473179 128373 473180
rect 194731 473244 194797 473245
rect 194731 473180 194732 473244
rect 194796 473180 194797 473244
rect 194731 473179 194797 473180
rect 390875 473244 390941 473245
rect 390875 473180 390876 473244
rect 390940 473180 390941 473244
rect 390875 473179 390941 473180
rect 81387 468484 81453 468485
rect 81387 468420 81388 468484
rect 81452 468420 81453 468484
rect 81387 468419 81453 468420
rect 165659 468484 165725 468485
rect 165659 468420 165660 468484
rect 165724 468420 165725 468484
rect 165659 468419 165725 468420
rect 259499 468484 259565 468485
rect 259499 468420 259500 468484
rect 259564 468420 259565 468484
rect 259499 468419 259565 468420
rect 361619 468484 361685 468485
rect 361619 468420 361620 468484
rect 361684 468420 361685 468484
rect 361619 468419 361685 468420
rect 445707 468484 445773 468485
rect 445707 468420 445708 468484
rect 445772 468420 445773 468484
rect 445707 468419 445773 468420
rect 455459 468484 455525 468485
rect 455459 468420 455460 468484
rect 455524 468420 455525 468484
rect 455459 468419 455525 468420
rect 557579 468484 557645 468485
rect 557579 468420 557580 468484
rect 557644 468420 557645 468484
rect 557579 468419 557645 468420
rect 44587 466852 44653 466853
rect 44587 466788 44588 466852
rect 44652 466788 44653 466852
rect 44587 466787 44653 466788
rect -2006 458593 -1974 458829
rect -1738 458593 -1654 458829
rect -1418 458593 -1386 458829
rect -2006 458509 -1386 458593
rect -2006 458273 -1974 458509
rect -1738 458273 -1654 458509
rect -1418 458273 -1386 458509
rect -2006 431829 -1386 458273
rect 20076 458829 20396 458861
rect 20076 458593 20118 458829
rect 20354 458593 20396 458829
rect 20076 458509 20396 458593
rect 20076 458273 20118 458509
rect 20354 458273 20396 458509
rect 20076 458241 20396 458273
rect 26340 458829 26660 458861
rect 26340 458593 26382 458829
rect 26618 458593 26660 458829
rect 26340 458509 26660 458593
rect 26340 458273 26382 458509
rect 26618 458273 26660 458509
rect 26340 458241 26660 458273
rect 32604 458829 32924 458861
rect 44590 458829 44650 466787
rect 48076 458829 48396 458861
rect 32604 458593 32646 458829
rect 32882 458593 32924 458829
rect 44587 458828 44653 458829
rect 44587 458764 44588 458828
rect 44652 458764 44653 458828
rect 44587 458763 44653 458764
rect 32604 458509 32924 458593
rect 32604 458273 32646 458509
rect 32882 458273 32924 458509
rect 32604 458241 32924 458273
rect 48076 458593 48118 458829
rect 48354 458593 48396 458829
rect 48076 458509 48396 458593
rect 48076 458273 48118 458509
rect 48354 458273 48396 458509
rect 48076 458241 48396 458273
rect 54340 458829 54660 458861
rect 54340 458593 54382 458829
rect 54618 458593 54660 458829
rect 54340 458509 54660 458593
rect 54340 458273 54382 458509
rect 54618 458273 54660 458509
rect 54340 458241 54660 458273
rect 60604 458829 60924 458861
rect 60604 458593 60646 458829
rect 60882 458593 60924 458829
rect 60604 458509 60924 458593
rect 60604 458273 60646 458509
rect 60882 458273 60924 458509
rect 60604 458241 60924 458273
rect 76076 458829 76396 458861
rect 76076 458593 76118 458829
rect 76354 458593 76396 458829
rect 76076 458509 76396 458593
rect 76076 458273 76118 458509
rect 76354 458273 76396 458509
rect 76076 458241 76396 458273
rect 23208 455454 23528 455486
rect 23208 455218 23250 455454
rect 23486 455218 23528 455454
rect 23208 455134 23528 455218
rect 23208 454898 23250 455134
rect 23486 454898 23528 455134
rect 23208 454866 23528 454898
rect 29472 455454 29792 455486
rect 29472 455218 29514 455454
rect 29750 455218 29792 455454
rect 29472 455134 29792 455218
rect 29472 454898 29514 455134
rect 29750 454898 29792 455134
rect 29472 454866 29792 454898
rect 51208 455454 51528 455486
rect 51208 455218 51250 455454
rect 51486 455218 51528 455454
rect 51208 455134 51528 455218
rect 51208 454898 51250 455134
rect 51486 454898 51528 455134
rect 51208 454866 51528 454898
rect 57472 455454 57792 455486
rect 57472 455218 57514 455454
rect 57750 455218 57792 455454
rect 57472 455134 57792 455218
rect 57472 454898 57514 455134
rect 57750 454898 57792 455134
rect 57472 454866 57792 454898
rect 79208 455454 79528 455486
rect 79208 455218 79250 455454
rect 79486 455218 79528 455454
rect 79208 455134 79528 455218
rect 79208 454898 79250 455134
rect 79486 454898 79528 455134
rect 79208 454866 79528 454898
rect 81390 445637 81450 468419
rect 128491 466716 128557 466717
rect 128491 466652 128492 466716
rect 128556 466652 128557 466716
rect 128491 466651 128557 466652
rect 82340 458829 82660 458861
rect 82340 458593 82382 458829
rect 82618 458593 82660 458829
rect 82340 458509 82660 458593
rect 82340 458273 82382 458509
rect 82618 458273 82660 458509
rect 82340 458241 82660 458273
rect 88604 458829 88924 458861
rect 88604 458593 88646 458829
rect 88882 458593 88924 458829
rect 88604 458509 88924 458593
rect 88604 458273 88646 458509
rect 88882 458273 88924 458509
rect 88604 458241 88924 458273
rect 104076 458829 104396 458861
rect 104076 458593 104118 458829
rect 104354 458593 104396 458829
rect 104076 458509 104396 458593
rect 104076 458273 104118 458509
rect 104354 458273 104396 458509
rect 104076 458241 104396 458273
rect 110340 458829 110660 458861
rect 110340 458593 110382 458829
rect 110618 458593 110660 458829
rect 110340 458509 110660 458593
rect 110340 458273 110382 458509
rect 110618 458273 110660 458509
rect 110340 458241 110660 458273
rect 116604 458829 116924 458861
rect 128494 458829 128554 466651
rect 132076 458829 132396 458861
rect 116604 458593 116646 458829
rect 116882 458593 116924 458829
rect 128491 458828 128557 458829
rect 128491 458764 128492 458828
rect 128556 458764 128557 458828
rect 128491 458763 128557 458764
rect 116604 458509 116924 458593
rect 116604 458273 116646 458509
rect 116882 458273 116924 458509
rect 116604 458241 116924 458273
rect 132076 458593 132118 458829
rect 132354 458593 132396 458829
rect 132076 458509 132396 458593
rect 132076 458273 132118 458509
rect 132354 458273 132396 458509
rect 132076 458241 132396 458273
rect 138340 458829 138660 458861
rect 138340 458593 138382 458829
rect 138618 458593 138660 458829
rect 138340 458509 138660 458593
rect 138340 458273 138382 458509
rect 138618 458273 138660 458509
rect 138340 458241 138660 458273
rect 144604 458829 144924 458861
rect 144604 458593 144646 458829
rect 144882 458593 144924 458829
rect 144604 458509 144924 458593
rect 144604 458273 144646 458509
rect 144882 458273 144924 458509
rect 144604 458241 144924 458273
rect 160076 458829 160396 458861
rect 160076 458593 160118 458829
rect 160354 458593 160396 458829
rect 160076 458509 160396 458593
rect 160076 458273 160118 458509
rect 160354 458273 160396 458509
rect 160076 458241 160396 458273
rect 85472 455454 85792 455486
rect 85472 455218 85514 455454
rect 85750 455218 85792 455454
rect 85472 455134 85792 455218
rect 85472 454898 85514 455134
rect 85750 454898 85792 455134
rect 85472 454866 85792 454898
rect 107208 455454 107528 455486
rect 107208 455218 107250 455454
rect 107486 455218 107528 455454
rect 107208 455134 107528 455218
rect 107208 454898 107250 455134
rect 107486 454898 107528 455134
rect 107208 454866 107528 454898
rect 113472 455454 113792 455486
rect 113472 455218 113514 455454
rect 113750 455218 113792 455454
rect 113472 455134 113792 455218
rect 113472 454898 113514 455134
rect 113750 454898 113792 455134
rect 113472 454866 113792 454898
rect 135208 455454 135528 455486
rect 135208 455218 135250 455454
rect 135486 455218 135528 455454
rect 135208 455134 135528 455218
rect 135208 454898 135250 455134
rect 135486 454898 135528 455134
rect 135208 454866 135528 454898
rect 141472 455454 141792 455486
rect 141472 455218 141514 455454
rect 141750 455218 141792 455454
rect 141472 455134 141792 455218
rect 141472 454898 141514 455134
rect 141750 454898 141792 455134
rect 141472 454866 141792 454898
rect 163208 455454 163528 455486
rect 163208 455218 163250 455454
rect 163486 455218 163528 455454
rect 163208 455134 163528 455218
rect 163208 454898 163250 455134
rect 163486 454898 163528 455134
rect 163208 454866 163528 454898
rect 165662 445637 165722 468419
rect 212579 466988 212645 466989
rect 212579 466924 212580 466988
rect 212644 466924 212645 466988
rect 212579 466923 212645 466924
rect 166340 458829 166660 458861
rect 166340 458593 166382 458829
rect 166618 458593 166660 458829
rect 166340 458509 166660 458593
rect 166340 458273 166382 458509
rect 166618 458273 166660 458509
rect 166340 458241 166660 458273
rect 172604 458829 172924 458861
rect 172604 458593 172646 458829
rect 172882 458593 172924 458829
rect 172604 458509 172924 458593
rect 172604 458273 172646 458509
rect 172882 458273 172924 458509
rect 172604 458241 172924 458273
rect 188076 458829 188396 458861
rect 188076 458593 188118 458829
rect 188354 458593 188396 458829
rect 188076 458509 188396 458593
rect 188076 458273 188118 458509
rect 188354 458273 188396 458509
rect 188076 458241 188396 458273
rect 194340 458829 194660 458861
rect 194340 458593 194382 458829
rect 194618 458593 194660 458829
rect 194340 458509 194660 458593
rect 194340 458273 194382 458509
rect 194618 458273 194660 458509
rect 194340 458241 194660 458273
rect 200604 458829 200924 458861
rect 212582 458829 212642 466923
rect 240547 466852 240613 466853
rect 240547 466788 240548 466852
rect 240612 466788 240613 466852
rect 240547 466787 240613 466788
rect 216076 458829 216396 458861
rect 200604 458593 200646 458829
rect 200882 458593 200924 458829
rect 212579 458828 212645 458829
rect 212579 458764 212580 458828
rect 212644 458764 212645 458828
rect 212579 458763 212645 458764
rect 200604 458509 200924 458593
rect 200604 458273 200646 458509
rect 200882 458273 200924 458509
rect 200604 458241 200924 458273
rect 216076 458593 216118 458829
rect 216354 458593 216396 458829
rect 216076 458509 216396 458593
rect 216076 458273 216118 458509
rect 216354 458273 216396 458509
rect 216076 458241 216396 458273
rect 222340 458829 222660 458861
rect 222340 458593 222382 458829
rect 222618 458593 222660 458829
rect 222340 458509 222660 458593
rect 222340 458273 222382 458509
rect 222618 458273 222660 458509
rect 222340 458241 222660 458273
rect 228604 458829 228924 458861
rect 240550 458829 240610 466787
rect 244076 458829 244396 458861
rect 228604 458593 228646 458829
rect 228882 458593 228924 458829
rect 240547 458828 240613 458829
rect 240547 458764 240548 458828
rect 240612 458764 240613 458828
rect 240547 458763 240613 458764
rect 228604 458509 228924 458593
rect 228604 458273 228646 458509
rect 228882 458273 228924 458509
rect 228604 458241 228924 458273
rect 244076 458593 244118 458829
rect 244354 458593 244396 458829
rect 244076 458509 244396 458593
rect 244076 458273 244118 458509
rect 244354 458273 244396 458509
rect 244076 458241 244396 458273
rect 250340 458829 250660 458861
rect 250340 458593 250382 458829
rect 250618 458593 250660 458829
rect 250340 458509 250660 458593
rect 250340 458273 250382 458509
rect 250618 458273 250660 458509
rect 250340 458241 250660 458273
rect 256604 458829 256924 458861
rect 256604 458593 256646 458829
rect 256882 458593 256924 458829
rect 256604 458509 256924 458593
rect 256604 458273 256646 458509
rect 256882 458273 256924 458509
rect 256604 458241 256924 458273
rect 169472 455454 169792 455486
rect 169472 455218 169514 455454
rect 169750 455218 169792 455454
rect 169472 455134 169792 455218
rect 169472 454898 169514 455134
rect 169750 454898 169792 455134
rect 169472 454866 169792 454898
rect 191208 455454 191528 455486
rect 191208 455218 191250 455454
rect 191486 455218 191528 455454
rect 191208 455134 191528 455218
rect 191208 454898 191250 455134
rect 191486 454898 191528 455134
rect 191208 454866 191528 454898
rect 197472 455454 197792 455486
rect 197472 455218 197514 455454
rect 197750 455218 197792 455454
rect 197472 455134 197792 455218
rect 197472 454898 197514 455134
rect 197750 454898 197792 455134
rect 197472 454866 197792 454898
rect 219208 455454 219528 455486
rect 219208 455218 219250 455454
rect 219486 455218 219528 455454
rect 219208 455134 219528 455218
rect 219208 454898 219250 455134
rect 219486 454898 219528 455134
rect 219208 454866 219528 454898
rect 225472 455454 225792 455486
rect 225472 455218 225514 455454
rect 225750 455218 225792 455454
rect 225472 455134 225792 455218
rect 225472 454898 225514 455134
rect 225750 454898 225792 455134
rect 225472 454866 225792 454898
rect 247208 455454 247528 455486
rect 247208 455218 247250 455454
rect 247486 455218 247528 455454
rect 247208 455134 247528 455218
rect 247208 454898 247250 455134
rect 247486 454898 247528 455134
rect 247208 454866 247528 454898
rect 253472 455454 253792 455486
rect 253472 455218 253514 455454
rect 253750 455218 253792 455454
rect 253472 455134 253792 455218
rect 253472 454898 253514 455134
rect 253750 454898 253792 455134
rect 253472 454866 253792 454898
rect 259502 445637 259562 468419
rect 296851 466852 296917 466853
rect 296851 466788 296852 466852
rect 296916 466788 296917 466852
rect 296851 466787 296917 466788
rect 296854 463710 296914 466787
rect 324635 466716 324701 466717
rect 324635 466652 324636 466716
rect 324700 466652 324701 466716
rect 324635 466651 324701 466652
rect 296486 463650 296914 463710
rect 272076 458829 272396 458861
rect 272076 458593 272118 458829
rect 272354 458593 272396 458829
rect 272076 458509 272396 458593
rect 272076 458273 272118 458509
rect 272354 458273 272396 458509
rect 272076 458241 272396 458273
rect 278340 458829 278660 458861
rect 278340 458593 278382 458829
rect 278618 458593 278660 458829
rect 278340 458509 278660 458593
rect 278340 458273 278382 458509
rect 278618 458273 278660 458509
rect 278340 458241 278660 458273
rect 284604 458829 284924 458861
rect 296486 458829 296546 463650
rect 300076 458829 300396 458861
rect 284604 458593 284646 458829
rect 284882 458593 284924 458829
rect 296483 458828 296549 458829
rect 296483 458764 296484 458828
rect 296548 458764 296549 458828
rect 296483 458763 296549 458764
rect 284604 458509 284924 458593
rect 284604 458273 284646 458509
rect 284882 458273 284924 458509
rect 284604 458241 284924 458273
rect 300076 458593 300118 458829
rect 300354 458593 300396 458829
rect 300076 458509 300396 458593
rect 300076 458273 300118 458509
rect 300354 458273 300396 458509
rect 300076 458241 300396 458273
rect 306340 458829 306660 458861
rect 306340 458593 306382 458829
rect 306618 458593 306660 458829
rect 306340 458509 306660 458593
rect 306340 458273 306382 458509
rect 306618 458273 306660 458509
rect 306340 458241 306660 458273
rect 312604 458829 312924 458861
rect 324638 458829 324698 466651
rect 328076 458829 328396 458861
rect 312604 458593 312646 458829
rect 312882 458593 312924 458829
rect 324635 458828 324701 458829
rect 324635 458764 324636 458828
rect 324700 458764 324701 458828
rect 324635 458763 324701 458764
rect 312604 458509 312924 458593
rect 312604 458273 312646 458509
rect 312882 458273 312924 458509
rect 312604 458241 312924 458273
rect 328076 458593 328118 458829
rect 328354 458593 328396 458829
rect 328076 458509 328396 458593
rect 328076 458273 328118 458509
rect 328354 458273 328396 458509
rect 328076 458241 328396 458273
rect 334340 458829 334660 458861
rect 334340 458593 334382 458829
rect 334618 458593 334660 458829
rect 334340 458509 334660 458593
rect 334340 458273 334382 458509
rect 334618 458273 334660 458509
rect 334340 458241 334660 458273
rect 340604 458829 340924 458861
rect 340604 458593 340646 458829
rect 340882 458593 340924 458829
rect 340604 458509 340924 458593
rect 340604 458273 340646 458509
rect 340882 458273 340924 458509
rect 340604 458241 340924 458273
rect 356076 458829 356396 458861
rect 356076 458593 356118 458829
rect 356354 458593 356396 458829
rect 356076 458509 356396 458593
rect 356076 458273 356118 458509
rect 356354 458273 356396 458509
rect 356076 458241 356396 458273
rect 275208 455454 275528 455486
rect 275208 455218 275250 455454
rect 275486 455218 275528 455454
rect 275208 455134 275528 455218
rect 275208 454898 275250 455134
rect 275486 454898 275528 455134
rect 275208 454866 275528 454898
rect 281472 455454 281792 455486
rect 281472 455218 281514 455454
rect 281750 455218 281792 455454
rect 281472 455134 281792 455218
rect 281472 454898 281514 455134
rect 281750 454898 281792 455134
rect 281472 454866 281792 454898
rect 303208 455454 303528 455486
rect 303208 455218 303250 455454
rect 303486 455218 303528 455454
rect 303208 455134 303528 455218
rect 303208 454898 303250 455134
rect 303486 454898 303528 455134
rect 303208 454866 303528 454898
rect 309472 455454 309792 455486
rect 309472 455218 309514 455454
rect 309750 455218 309792 455454
rect 309472 455134 309792 455218
rect 309472 454898 309514 455134
rect 309750 454898 309792 455134
rect 309472 454866 309792 454898
rect 331208 455454 331528 455486
rect 331208 455218 331250 455454
rect 331486 455218 331528 455454
rect 331208 455134 331528 455218
rect 331208 454898 331250 455134
rect 331486 454898 331528 455134
rect 331208 454866 331528 454898
rect 337472 455454 337792 455486
rect 337472 455218 337514 455454
rect 337750 455218 337792 455454
rect 337472 455134 337792 455218
rect 337472 454898 337514 455134
rect 337750 454898 337792 455134
rect 337472 454866 337792 454898
rect 359208 455454 359528 455486
rect 359208 455218 359250 455454
rect 359486 455218 359528 455454
rect 359208 455134 359528 455218
rect 359208 454898 359250 455134
rect 359486 454898 359528 455134
rect 359208 454866 359528 454898
rect 361622 445637 361682 468419
rect 408539 466988 408605 466989
rect 408539 466924 408540 466988
rect 408604 466924 408605 466988
rect 408539 466923 408605 466924
rect 362340 458829 362660 458861
rect 362340 458593 362382 458829
rect 362618 458593 362660 458829
rect 362340 458509 362660 458593
rect 362340 458273 362382 458509
rect 362618 458273 362660 458509
rect 362340 458241 362660 458273
rect 368604 458829 368924 458861
rect 368604 458593 368646 458829
rect 368882 458593 368924 458829
rect 368604 458509 368924 458593
rect 368604 458273 368646 458509
rect 368882 458273 368924 458509
rect 368604 458241 368924 458273
rect 384076 458829 384396 458861
rect 384076 458593 384118 458829
rect 384354 458593 384396 458829
rect 384076 458509 384396 458593
rect 384076 458273 384118 458509
rect 384354 458273 384396 458509
rect 384076 458241 384396 458273
rect 390340 458829 390660 458861
rect 390340 458593 390382 458829
rect 390618 458593 390660 458829
rect 390340 458509 390660 458593
rect 390340 458273 390382 458509
rect 390618 458273 390660 458509
rect 390340 458241 390660 458273
rect 396604 458829 396924 458861
rect 408542 458829 408602 466923
rect 436507 466852 436573 466853
rect 436507 466788 436508 466852
rect 436572 466788 436573 466852
rect 436507 466787 436573 466788
rect 412076 458829 412396 458861
rect 396604 458593 396646 458829
rect 396882 458593 396924 458829
rect 408539 458828 408605 458829
rect 408539 458764 408540 458828
rect 408604 458764 408605 458828
rect 408539 458763 408605 458764
rect 396604 458509 396924 458593
rect 396604 458273 396646 458509
rect 396882 458273 396924 458509
rect 396604 458241 396924 458273
rect 412076 458593 412118 458829
rect 412354 458593 412396 458829
rect 412076 458509 412396 458593
rect 412076 458273 412118 458509
rect 412354 458273 412396 458509
rect 412076 458241 412396 458273
rect 418340 458829 418660 458861
rect 418340 458593 418382 458829
rect 418618 458593 418660 458829
rect 418340 458509 418660 458593
rect 418340 458273 418382 458509
rect 418618 458273 418660 458509
rect 418340 458241 418660 458273
rect 424604 458829 424924 458861
rect 436510 458829 436570 466787
rect 440076 458829 440396 458861
rect 424604 458593 424646 458829
rect 424882 458593 424924 458829
rect 436507 458828 436573 458829
rect 436507 458764 436508 458828
rect 436572 458764 436573 458828
rect 436507 458763 436573 458764
rect 424604 458509 424924 458593
rect 424604 458273 424646 458509
rect 424882 458273 424924 458509
rect 424604 458241 424924 458273
rect 440076 458593 440118 458829
rect 440354 458593 440396 458829
rect 440076 458509 440396 458593
rect 440076 458273 440118 458509
rect 440354 458273 440396 458509
rect 440076 458241 440396 458273
rect 365472 455454 365792 455486
rect 365472 455218 365514 455454
rect 365750 455218 365792 455454
rect 365472 455134 365792 455218
rect 365472 454898 365514 455134
rect 365750 454898 365792 455134
rect 365472 454866 365792 454898
rect 387208 455454 387528 455486
rect 387208 455218 387250 455454
rect 387486 455218 387528 455454
rect 387208 455134 387528 455218
rect 387208 454898 387250 455134
rect 387486 454898 387528 455134
rect 387208 454866 387528 454898
rect 393472 455454 393792 455486
rect 393472 455218 393514 455454
rect 393750 455218 393792 455454
rect 393472 455134 393792 455218
rect 393472 454898 393514 455134
rect 393750 454898 393792 455134
rect 393472 454866 393792 454898
rect 415208 455454 415528 455486
rect 415208 455218 415250 455454
rect 415486 455218 415528 455454
rect 415208 455134 415528 455218
rect 415208 454898 415250 455134
rect 415486 454898 415528 455134
rect 415208 454866 415528 454898
rect 421472 455454 421792 455486
rect 421472 455218 421514 455454
rect 421750 455218 421792 455454
rect 421472 455134 421792 455218
rect 421472 454898 421514 455134
rect 421750 454898 421792 455134
rect 421472 454866 421792 454898
rect 443208 455454 443528 455486
rect 443208 455218 443250 455454
rect 443486 455218 443528 455454
rect 443208 455134 443528 455218
rect 443208 454898 443250 455134
rect 443486 454898 443528 455134
rect 443208 454866 443528 454898
rect 81387 445636 81453 445637
rect 81387 445572 81388 445636
rect 81452 445572 81453 445636
rect 81387 445571 81453 445572
rect 165659 445636 165725 445637
rect 165659 445572 165660 445636
rect 165724 445572 165725 445636
rect 165659 445571 165725 445572
rect 259499 445636 259565 445637
rect 259499 445572 259500 445636
rect 259564 445572 259565 445636
rect 259499 445571 259565 445572
rect 361619 445636 361685 445637
rect 361619 445572 361620 445636
rect 361684 445572 361685 445636
rect 361619 445571 361685 445572
rect 445710 445501 445770 468419
rect 446340 458829 446660 458861
rect 446340 458593 446382 458829
rect 446618 458593 446660 458829
rect 446340 458509 446660 458593
rect 446340 458273 446382 458509
rect 446618 458273 446660 458509
rect 446340 458241 446660 458273
rect 452604 458829 452924 458861
rect 452604 458593 452646 458829
rect 452882 458593 452924 458829
rect 452604 458509 452924 458593
rect 452604 458273 452646 458509
rect 452882 458273 452924 458509
rect 452604 458241 452924 458273
rect 449472 455454 449792 455486
rect 449472 455218 449514 455454
rect 449750 455218 449792 455454
rect 449472 455134 449792 455218
rect 449472 454898 449514 455134
rect 449750 454898 449792 455134
rect 449472 454866 449792 454898
rect 455462 445637 455522 468419
rect 492811 466852 492877 466853
rect 492811 466788 492812 466852
rect 492876 466788 492877 466852
rect 492811 466787 492877 466788
rect 492814 460950 492874 466787
rect 520595 466716 520661 466717
rect 520595 466652 520596 466716
rect 520660 466652 520661 466716
rect 520595 466651 520661 466652
rect 492630 460890 492874 460950
rect 468076 458829 468396 458861
rect 468076 458593 468118 458829
rect 468354 458593 468396 458829
rect 468076 458509 468396 458593
rect 468076 458273 468118 458509
rect 468354 458273 468396 458509
rect 468076 458241 468396 458273
rect 474340 458829 474660 458861
rect 474340 458593 474382 458829
rect 474618 458593 474660 458829
rect 474340 458509 474660 458593
rect 474340 458273 474382 458509
rect 474618 458273 474660 458509
rect 474340 458241 474660 458273
rect 480604 458829 480924 458861
rect 492630 458829 492690 460890
rect 496076 458829 496396 458861
rect 480604 458593 480646 458829
rect 480882 458593 480924 458829
rect 492627 458828 492693 458829
rect 492627 458764 492628 458828
rect 492692 458764 492693 458828
rect 492627 458763 492693 458764
rect 480604 458509 480924 458593
rect 480604 458273 480646 458509
rect 480882 458273 480924 458509
rect 480604 458241 480924 458273
rect 496076 458593 496118 458829
rect 496354 458593 496396 458829
rect 496076 458509 496396 458593
rect 496076 458273 496118 458509
rect 496354 458273 496396 458509
rect 496076 458241 496396 458273
rect 502340 458829 502660 458861
rect 502340 458593 502382 458829
rect 502618 458593 502660 458829
rect 502340 458509 502660 458593
rect 502340 458273 502382 458509
rect 502618 458273 502660 458509
rect 502340 458241 502660 458273
rect 508604 458829 508924 458861
rect 520598 458829 520658 466651
rect 524076 458829 524396 458861
rect 508604 458593 508646 458829
rect 508882 458593 508924 458829
rect 520595 458828 520661 458829
rect 520595 458764 520596 458828
rect 520660 458764 520661 458828
rect 520595 458763 520661 458764
rect 508604 458509 508924 458593
rect 508604 458273 508646 458509
rect 508882 458273 508924 458509
rect 508604 458241 508924 458273
rect 524076 458593 524118 458829
rect 524354 458593 524396 458829
rect 524076 458509 524396 458593
rect 524076 458273 524118 458509
rect 524354 458273 524396 458509
rect 524076 458241 524396 458273
rect 530340 458829 530660 458861
rect 530340 458593 530382 458829
rect 530618 458593 530660 458829
rect 530340 458509 530660 458593
rect 530340 458273 530382 458509
rect 530618 458273 530660 458509
rect 530340 458241 530660 458273
rect 536604 458829 536924 458861
rect 536604 458593 536646 458829
rect 536882 458593 536924 458829
rect 536604 458509 536924 458593
rect 536604 458273 536646 458509
rect 536882 458273 536924 458509
rect 536604 458241 536924 458273
rect 552076 458829 552396 458861
rect 552076 458593 552118 458829
rect 552354 458593 552396 458829
rect 552076 458509 552396 458593
rect 552076 458273 552118 458509
rect 552354 458273 552396 458509
rect 552076 458241 552396 458273
rect 471208 455454 471528 455486
rect 471208 455218 471250 455454
rect 471486 455218 471528 455454
rect 471208 455134 471528 455218
rect 471208 454898 471250 455134
rect 471486 454898 471528 455134
rect 471208 454866 471528 454898
rect 477472 455454 477792 455486
rect 477472 455218 477514 455454
rect 477750 455218 477792 455454
rect 477472 455134 477792 455218
rect 477472 454898 477514 455134
rect 477750 454898 477792 455134
rect 477472 454866 477792 454898
rect 499208 455454 499528 455486
rect 499208 455218 499250 455454
rect 499486 455218 499528 455454
rect 499208 455134 499528 455218
rect 499208 454898 499250 455134
rect 499486 454898 499528 455134
rect 499208 454866 499528 454898
rect 505472 455454 505792 455486
rect 505472 455218 505514 455454
rect 505750 455218 505792 455454
rect 505472 455134 505792 455218
rect 505472 454898 505514 455134
rect 505750 454898 505792 455134
rect 505472 454866 505792 454898
rect 527208 455454 527528 455486
rect 527208 455218 527250 455454
rect 527486 455218 527528 455454
rect 527208 455134 527528 455218
rect 527208 454898 527250 455134
rect 527486 454898 527528 455134
rect 527208 454866 527528 454898
rect 533472 455454 533792 455486
rect 533472 455218 533514 455454
rect 533750 455218 533792 455454
rect 533472 455134 533792 455218
rect 533472 454898 533514 455134
rect 533750 454898 533792 455134
rect 533472 454866 533792 454898
rect 555208 455454 555528 455486
rect 555208 455218 555250 455454
rect 555486 455218 555528 455454
rect 555208 455134 555528 455218
rect 555208 454898 555250 455134
rect 555486 454898 555528 455134
rect 555208 454866 555528 454898
rect 557582 445637 557642 468419
rect 558340 458829 558660 458861
rect 558340 458593 558382 458829
rect 558618 458593 558660 458829
rect 558340 458509 558660 458593
rect 558340 458273 558382 458509
rect 558618 458273 558660 458509
rect 558340 458241 558660 458273
rect 564604 458829 564924 458861
rect 564604 458593 564646 458829
rect 564882 458593 564924 458829
rect 564604 458509 564924 458593
rect 564604 458273 564646 458509
rect 564882 458273 564924 458509
rect 564604 458241 564924 458273
rect 573494 458829 574114 485273
rect 573494 458593 573526 458829
rect 573762 458593 573846 458829
rect 574082 458593 574114 458829
rect 573494 458509 574114 458593
rect 573494 458273 573526 458509
rect 573762 458273 573846 458509
rect 574082 458273 574114 458509
rect 561472 455454 561792 455486
rect 561472 455218 561514 455454
rect 561750 455218 561792 455454
rect 561472 455134 561792 455218
rect 561472 454898 561514 455134
rect 561750 454898 561792 455134
rect 561472 454866 561792 454898
rect 455459 445636 455525 445637
rect 455459 445572 455460 445636
rect 455524 445572 455525 445636
rect 455459 445571 455525 445572
rect 557579 445636 557645 445637
rect 557579 445572 557580 445636
rect 557644 445572 557645 445636
rect 557579 445571 557645 445572
rect 445707 445500 445773 445501
rect 445707 445436 445708 445500
rect 445772 445436 445773 445500
rect 445707 445435 445773 445436
rect 128307 441692 128373 441693
rect 128307 441628 128308 441692
rect 128372 441628 128373 441692
rect 128307 441627 128373 441628
rect 194731 441692 194797 441693
rect 194731 441628 194732 441692
rect 194796 441628 194797 441692
rect 194731 441627 194797 441628
rect 390875 441692 390941 441693
rect 390875 441628 390876 441692
rect 390940 441628 390941 441692
rect 390875 441627 390941 441628
rect -2006 431593 -1974 431829
rect -1738 431593 -1654 431829
rect -1418 431593 -1386 431829
rect -2006 431509 -1386 431593
rect -2006 431273 -1974 431509
rect -1738 431273 -1654 431509
rect -1418 431273 -1386 431509
rect -2006 404829 -1386 431273
rect 20076 431829 20396 431861
rect 20076 431593 20118 431829
rect 20354 431593 20396 431829
rect 20076 431509 20396 431593
rect 20076 431273 20118 431509
rect 20354 431273 20396 431509
rect 20076 431241 20396 431273
rect 26340 431829 26660 431861
rect 26340 431593 26382 431829
rect 26618 431593 26660 431829
rect 26340 431509 26660 431593
rect 26340 431273 26382 431509
rect 26618 431273 26660 431509
rect 26340 431241 26660 431273
rect 32604 431829 32924 431861
rect 32604 431593 32646 431829
rect 32882 431593 32924 431829
rect 32604 431509 32924 431593
rect 32604 431273 32646 431509
rect 32882 431273 32924 431509
rect 32604 431241 32924 431273
rect 48076 431829 48396 431861
rect 48076 431593 48118 431829
rect 48354 431593 48396 431829
rect 48076 431509 48396 431593
rect 48076 431273 48118 431509
rect 48354 431273 48396 431509
rect 48076 431241 48396 431273
rect 54340 431829 54660 431861
rect 54340 431593 54382 431829
rect 54618 431593 54660 431829
rect 54340 431509 54660 431593
rect 54340 431273 54382 431509
rect 54618 431273 54660 431509
rect 54340 431241 54660 431273
rect 60604 431829 60924 431861
rect 60604 431593 60646 431829
rect 60882 431593 60924 431829
rect 60604 431509 60924 431593
rect 60604 431273 60646 431509
rect 60882 431273 60924 431509
rect 60604 431241 60924 431273
rect 76076 431829 76396 431861
rect 76076 431593 76118 431829
rect 76354 431593 76396 431829
rect 76076 431509 76396 431593
rect 76076 431273 76118 431509
rect 76354 431273 76396 431509
rect 76076 431241 76396 431273
rect 82340 431829 82660 431861
rect 82340 431593 82382 431829
rect 82618 431593 82660 431829
rect 82340 431509 82660 431593
rect 82340 431273 82382 431509
rect 82618 431273 82660 431509
rect 82340 431241 82660 431273
rect 88604 431829 88924 431861
rect 88604 431593 88646 431829
rect 88882 431593 88924 431829
rect 88604 431509 88924 431593
rect 88604 431273 88646 431509
rect 88882 431273 88924 431509
rect 88604 431241 88924 431273
rect 104076 431829 104396 431861
rect 104076 431593 104118 431829
rect 104354 431593 104396 431829
rect 104076 431509 104396 431593
rect 104076 431273 104118 431509
rect 104354 431273 104396 431509
rect 104076 431241 104396 431273
rect 110340 431829 110660 431861
rect 110340 431593 110382 431829
rect 110618 431593 110660 431829
rect 110340 431509 110660 431593
rect 110340 431273 110382 431509
rect 110618 431273 110660 431509
rect 110340 431241 110660 431273
rect 116604 431829 116924 431861
rect 116604 431593 116646 431829
rect 116882 431593 116924 431829
rect 116604 431509 116924 431593
rect 116604 431273 116646 431509
rect 116882 431273 116924 431509
rect 116604 431241 116924 431273
rect 64459 431220 64525 431221
rect 64459 431156 64460 431220
rect 64524 431156 64525 431220
rect 64459 431155 64525 431156
rect 92427 431220 92493 431221
rect 92427 431156 92428 431220
rect 92492 431156 92493 431220
rect 92427 431155 92493 431156
rect 23208 428454 23528 428486
rect 23208 428218 23250 428454
rect 23486 428218 23528 428454
rect 23208 428134 23528 428218
rect 23208 427898 23250 428134
rect 23486 427898 23528 428134
rect 23208 427866 23528 427898
rect 29472 428454 29792 428486
rect 29472 428218 29514 428454
rect 29750 428218 29792 428454
rect 29472 428134 29792 428218
rect 29472 427898 29514 428134
rect 29750 427898 29792 428134
rect 29472 427866 29792 427898
rect 51208 428454 51528 428486
rect 51208 428218 51250 428454
rect 51486 428218 51528 428454
rect 51208 428134 51528 428218
rect 51208 427898 51250 428134
rect 51486 427898 51528 428134
rect 51208 427866 51528 427898
rect 57472 428454 57792 428486
rect 57472 428218 57514 428454
rect 57750 428218 57792 428454
rect 57472 428134 57792 428218
rect 57472 427898 57514 428134
rect 57750 427898 57792 428134
rect 57472 427866 57792 427898
rect 64462 423333 64522 431155
rect 79208 428454 79528 428486
rect 79208 428218 79250 428454
rect 79486 428218 79528 428454
rect 79208 428134 79528 428218
rect 79208 427898 79250 428134
rect 79486 427898 79528 428134
rect 79208 427866 79528 427898
rect 85472 428454 85792 428486
rect 85472 428218 85514 428454
rect 85750 428218 85792 428454
rect 85472 428134 85792 428218
rect 85472 427898 85514 428134
rect 85750 427898 85792 428134
rect 85472 427866 85792 427898
rect 64459 423332 64525 423333
rect 64459 423268 64460 423332
rect 64524 423268 64525 423332
rect 64459 423267 64525 423268
rect 92430 423197 92490 431155
rect 107208 428454 107528 428486
rect 107208 428218 107250 428454
rect 107486 428218 107528 428454
rect 107208 428134 107528 428218
rect 107208 427898 107250 428134
rect 107486 427898 107528 428134
rect 107208 427866 107528 427898
rect 113472 428454 113792 428486
rect 113472 428218 113514 428454
rect 113750 428218 113792 428454
rect 113472 428134 113792 428218
rect 113472 427898 113514 428134
rect 113750 427898 113792 428134
rect 113472 427866 113792 427898
rect 92427 423196 92493 423197
rect 92427 423132 92428 423196
rect 92492 423132 92493 423196
rect 92427 423131 92493 423132
rect 128310 419525 128370 441627
rect 132076 431829 132396 431861
rect 132076 431593 132118 431829
rect 132354 431593 132396 431829
rect 132076 431509 132396 431593
rect 132076 431273 132118 431509
rect 132354 431273 132396 431509
rect 132076 431241 132396 431273
rect 138340 431829 138660 431861
rect 138340 431593 138382 431829
rect 138618 431593 138660 431829
rect 138340 431509 138660 431593
rect 138340 431273 138382 431509
rect 138618 431273 138660 431509
rect 138340 431241 138660 431273
rect 144604 431829 144924 431861
rect 144604 431593 144646 431829
rect 144882 431593 144924 431829
rect 144604 431509 144924 431593
rect 144604 431273 144646 431509
rect 144882 431273 144924 431509
rect 144604 431241 144924 431273
rect 160076 431829 160396 431861
rect 160076 431593 160118 431829
rect 160354 431593 160396 431829
rect 160076 431509 160396 431593
rect 160076 431273 160118 431509
rect 160354 431273 160396 431509
rect 160076 431241 160396 431273
rect 166340 431829 166660 431861
rect 166340 431593 166382 431829
rect 166618 431593 166660 431829
rect 166340 431509 166660 431593
rect 166340 431273 166382 431509
rect 166618 431273 166660 431509
rect 166340 431241 166660 431273
rect 172604 431829 172924 431861
rect 172604 431593 172646 431829
rect 172882 431593 172924 431829
rect 172604 431509 172924 431593
rect 172604 431273 172646 431509
rect 172882 431273 172924 431509
rect 172604 431241 172924 431273
rect 188076 431829 188396 431861
rect 188076 431593 188118 431829
rect 188354 431593 188396 431829
rect 188076 431509 188396 431593
rect 188076 431273 188118 431509
rect 188354 431273 188396 431509
rect 188076 431241 188396 431273
rect 194340 431829 194660 431861
rect 194340 431593 194382 431829
rect 194618 431593 194660 431829
rect 194340 431509 194660 431593
rect 194340 431273 194382 431509
rect 194618 431273 194660 431509
rect 194340 431241 194660 431273
rect 148363 431220 148429 431221
rect 148363 431156 148364 431220
rect 148428 431156 148429 431220
rect 148363 431155 148429 431156
rect 176331 431220 176397 431221
rect 176331 431156 176332 431220
rect 176396 431156 176397 431220
rect 176331 431155 176397 431156
rect 135208 428454 135528 428486
rect 135208 428218 135250 428454
rect 135486 428218 135528 428454
rect 135208 428134 135528 428218
rect 135208 427898 135250 428134
rect 135486 427898 135528 428134
rect 135208 427866 135528 427898
rect 141472 428454 141792 428486
rect 141472 428218 141514 428454
rect 141750 428218 141792 428454
rect 141472 428134 141792 428218
rect 141472 427898 141514 428134
rect 141750 427898 141792 428134
rect 141472 427866 141792 427898
rect 148366 423197 148426 431155
rect 163208 428454 163528 428486
rect 163208 428218 163250 428454
rect 163486 428218 163528 428454
rect 163208 428134 163528 428218
rect 163208 427898 163250 428134
rect 163486 427898 163528 428134
rect 163208 427866 163528 427898
rect 169472 428454 169792 428486
rect 169472 428218 169514 428454
rect 169750 428218 169792 428454
rect 169472 428134 169792 428218
rect 169472 427898 169514 428134
rect 169750 427898 169792 428134
rect 169472 427866 169792 427898
rect 176334 423333 176394 431155
rect 191208 428454 191528 428486
rect 191208 428218 191250 428454
rect 191486 428218 191528 428454
rect 191208 428134 191528 428218
rect 191208 427898 191250 428134
rect 191486 427898 191528 428134
rect 191208 427866 191528 427898
rect 176331 423332 176397 423333
rect 176331 423268 176332 423332
rect 176396 423268 176397 423332
rect 176331 423267 176397 423268
rect 148363 423196 148429 423197
rect 148363 423132 148364 423196
rect 148428 423132 148429 423196
rect 148363 423131 148429 423132
rect 194734 419525 194794 441627
rect 200604 431829 200924 431861
rect 200604 431593 200646 431829
rect 200882 431593 200924 431829
rect 200604 431509 200924 431593
rect 200604 431273 200646 431509
rect 200882 431273 200924 431509
rect 200604 431241 200924 431273
rect 216076 431829 216396 431861
rect 216076 431593 216118 431829
rect 216354 431593 216396 431829
rect 216076 431509 216396 431593
rect 216076 431273 216118 431509
rect 216354 431273 216396 431509
rect 216076 431241 216396 431273
rect 222340 431829 222660 431861
rect 222340 431593 222382 431829
rect 222618 431593 222660 431829
rect 222340 431509 222660 431593
rect 222340 431273 222382 431509
rect 222618 431273 222660 431509
rect 222340 431241 222660 431273
rect 228604 431829 228924 431861
rect 228604 431593 228646 431829
rect 228882 431593 228924 431829
rect 228604 431509 228924 431593
rect 228604 431273 228646 431509
rect 228882 431273 228924 431509
rect 228604 431241 228924 431273
rect 244076 431829 244396 431861
rect 244076 431593 244118 431829
rect 244354 431593 244396 431829
rect 244076 431509 244396 431593
rect 244076 431273 244118 431509
rect 244354 431273 244396 431509
rect 244076 431241 244396 431273
rect 250340 431829 250660 431861
rect 250340 431593 250382 431829
rect 250618 431593 250660 431829
rect 250340 431509 250660 431593
rect 250340 431273 250382 431509
rect 250618 431273 250660 431509
rect 250340 431241 250660 431273
rect 256604 431829 256924 431861
rect 256604 431593 256646 431829
rect 256882 431593 256924 431829
rect 256604 431509 256924 431593
rect 256604 431273 256646 431509
rect 256882 431273 256924 431509
rect 256604 431241 256924 431273
rect 272076 431829 272396 431861
rect 272076 431593 272118 431829
rect 272354 431593 272396 431829
rect 272076 431509 272396 431593
rect 272076 431273 272118 431509
rect 272354 431273 272396 431509
rect 272076 431241 272396 431273
rect 278340 431829 278660 431861
rect 278340 431593 278382 431829
rect 278618 431593 278660 431829
rect 278340 431509 278660 431593
rect 278340 431273 278382 431509
rect 278618 431273 278660 431509
rect 278340 431241 278660 431273
rect 284604 431829 284924 431861
rect 284604 431593 284646 431829
rect 284882 431593 284924 431829
rect 284604 431509 284924 431593
rect 284604 431273 284646 431509
rect 284882 431273 284924 431509
rect 284604 431241 284924 431273
rect 300076 431829 300396 431861
rect 300076 431593 300118 431829
rect 300354 431593 300396 431829
rect 300076 431509 300396 431593
rect 300076 431273 300118 431509
rect 300354 431273 300396 431509
rect 300076 431241 300396 431273
rect 306340 431829 306660 431861
rect 306340 431593 306382 431829
rect 306618 431593 306660 431829
rect 306340 431509 306660 431593
rect 306340 431273 306382 431509
rect 306618 431273 306660 431509
rect 306340 431241 306660 431273
rect 312604 431829 312924 431861
rect 312604 431593 312646 431829
rect 312882 431593 312924 431829
rect 312604 431509 312924 431593
rect 312604 431273 312646 431509
rect 312882 431273 312924 431509
rect 312604 431241 312924 431273
rect 328076 431829 328396 431861
rect 328076 431593 328118 431829
rect 328354 431593 328396 431829
rect 328076 431509 328396 431593
rect 328076 431273 328118 431509
rect 328354 431273 328396 431509
rect 328076 431241 328396 431273
rect 334340 431829 334660 431861
rect 334340 431593 334382 431829
rect 334618 431593 334660 431829
rect 334340 431509 334660 431593
rect 334340 431273 334382 431509
rect 334618 431273 334660 431509
rect 334340 431241 334660 431273
rect 340604 431829 340924 431861
rect 340604 431593 340646 431829
rect 340882 431593 340924 431829
rect 340604 431509 340924 431593
rect 340604 431273 340646 431509
rect 340882 431273 340924 431509
rect 340604 431241 340924 431273
rect 356076 431829 356396 431861
rect 356076 431593 356118 431829
rect 356354 431593 356396 431829
rect 356076 431509 356396 431593
rect 356076 431273 356118 431509
rect 356354 431273 356396 431509
rect 356076 431241 356396 431273
rect 362340 431829 362660 431861
rect 362340 431593 362382 431829
rect 362618 431593 362660 431829
rect 362340 431509 362660 431593
rect 362340 431273 362382 431509
rect 362618 431273 362660 431509
rect 362340 431241 362660 431273
rect 368604 431829 368924 431861
rect 368604 431593 368646 431829
rect 368882 431593 368924 431829
rect 368604 431509 368924 431593
rect 368604 431273 368646 431509
rect 368882 431273 368924 431509
rect 368604 431241 368924 431273
rect 384076 431829 384396 431861
rect 384076 431593 384118 431829
rect 384354 431593 384396 431829
rect 384076 431509 384396 431593
rect 384076 431273 384118 431509
rect 384354 431273 384396 431509
rect 384076 431241 384396 431273
rect 390340 431829 390660 431861
rect 390340 431593 390382 431829
rect 390618 431593 390660 431829
rect 390340 431509 390660 431593
rect 390340 431273 390382 431509
rect 390618 431273 390660 431509
rect 390340 431241 390660 431273
rect 260419 431220 260485 431221
rect 260419 431156 260420 431220
rect 260484 431156 260485 431220
rect 260419 431155 260485 431156
rect 288387 431220 288453 431221
rect 288387 431156 288388 431220
rect 288452 431156 288453 431220
rect 288387 431155 288453 431156
rect 344323 431220 344389 431221
rect 344323 431156 344324 431220
rect 344388 431156 344389 431220
rect 344323 431155 344389 431156
rect 372291 431220 372357 431221
rect 372291 431156 372292 431220
rect 372356 431156 372357 431220
rect 372291 431155 372357 431156
rect 197472 428454 197792 428486
rect 197472 428218 197514 428454
rect 197750 428218 197792 428454
rect 197472 428134 197792 428218
rect 197472 427898 197514 428134
rect 197750 427898 197792 428134
rect 197472 427866 197792 427898
rect 219208 428454 219528 428486
rect 219208 428218 219250 428454
rect 219486 428218 219528 428454
rect 219208 428134 219528 428218
rect 219208 427898 219250 428134
rect 219486 427898 219528 428134
rect 219208 427866 219528 427898
rect 225472 428454 225792 428486
rect 225472 428218 225514 428454
rect 225750 428218 225792 428454
rect 225472 428134 225792 428218
rect 225472 427898 225514 428134
rect 225750 427898 225792 428134
rect 225472 427866 225792 427898
rect 247208 428454 247528 428486
rect 247208 428218 247250 428454
rect 247486 428218 247528 428454
rect 247208 428134 247528 428218
rect 247208 427898 247250 428134
rect 247486 427898 247528 428134
rect 247208 427866 247528 427898
rect 253472 428454 253792 428486
rect 253472 428218 253514 428454
rect 253750 428218 253792 428454
rect 253472 428134 253792 428218
rect 253472 427898 253514 428134
rect 253750 427898 253792 428134
rect 253472 427866 253792 427898
rect 260422 423197 260482 431155
rect 275208 428454 275528 428486
rect 275208 428218 275250 428454
rect 275486 428218 275528 428454
rect 275208 428134 275528 428218
rect 275208 427898 275250 428134
rect 275486 427898 275528 428134
rect 275208 427866 275528 427898
rect 281472 428454 281792 428486
rect 281472 428218 281514 428454
rect 281750 428218 281792 428454
rect 281472 428134 281792 428218
rect 281472 427898 281514 428134
rect 281750 427898 281792 428134
rect 281472 427866 281792 427898
rect 260419 423196 260485 423197
rect 260419 423132 260420 423196
rect 260484 423132 260485 423196
rect 260419 423131 260485 423132
rect 288390 423061 288450 431155
rect 303208 428454 303528 428486
rect 303208 428218 303250 428454
rect 303486 428218 303528 428454
rect 303208 428134 303528 428218
rect 303208 427898 303250 428134
rect 303486 427898 303528 428134
rect 303208 427866 303528 427898
rect 309472 428454 309792 428486
rect 309472 428218 309514 428454
rect 309750 428218 309792 428454
rect 309472 428134 309792 428218
rect 309472 427898 309514 428134
rect 309750 427898 309792 428134
rect 309472 427866 309792 427898
rect 331208 428454 331528 428486
rect 331208 428218 331250 428454
rect 331486 428218 331528 428454
rect 331208 428134 331528 428218
rect 331208 427898 331250 428134
rect 331486 427898 331528 428134
rect 331208 427866 331528 427898
rect 337472 428454 337792 428486
rect 337472 428218 337514 428454
rect 337750 428218 337792 428454
rect 337472 428134 337792 428218
rect 337472 427898 337514 428134
rect 337750 427898 337792 428134
rect 337472 427866 337792 427898
rect 344326 423197 344386 431155
rect 359208 428454 359528 428486
rect 359208 428218 359250 428454
rect 359486 428218 359528 428454
rect 359208 428134 359528 428218
rect 359208 427898 359250 428134
rect 359486 427898 359528 428134
rect 359208 427866 359528 427898
rect 365472 428454 365792 428486
rect 365472 428218 365514 428454
rect 365750 428218 365792 428454
rect 365472 428134 365792 428218
rect 365472 427898 365514 428134
rect 365750 427898 365792 428134
rect 365472 427866 365792 427898
rect 372294 423333 372354 431155
rect 387208 428454 387528 428486
rect 387208 428218 387250 428454
rect 387486 428218 387528 428454
rect 387208 428134 387528 428218
rect 387208 427898 387250 428134
rect 387486 427898 387528 428134
rect 387208 427866 387528 427898
rect 372291 423332 372357 423333
rect 372291 423268 372292 423332
rect 372356 423268 372357 423332
rect 372291 423267 372357 423268
rect 344323 423196 344389 423197
rect 344323 423132 344324 423196
rect 344388 423132 344389 423196
rect 344323 423131 344389 423132
rect 288387 423060 288453 423061
rect 288387 422996 288388 423060
rect 288452 422996 288453 423060
rect 288387 422995 288453 422996
rect 390878 419525 390938 441627
rect 396604 431829 396924 431861
rect 396604 431593 396646 431829
rect 396882 431593 396924 431829
rect 396604 431509 396924 431593
rect 396604 431273 396646 431509
rect 396882 431273 396924 431509
rect 396604 431241 396924 431273
rect 412076 431829 412396 431861
rect 412076 431593 412118 431829
rect 412354 431593 412396 431829
rect 412076 431509 412396 431593
rect 412076 431273 412118 431509
rect 412354 431273 412396 431509
rect 412076 431241 412396 431273
rect 418340 431829 418660 431861
rect 418340 431593 418382 431829
rect 418618 431593 418660 431829
rect 418340 431509 418660 431593
rect 418340 431273 418382 431509
rect 418618 431273 418660 431509
rect 418340 431241 418660 431273
rect 424604 431829 424924 431861
rect 424604 431593 424646 431829
rect 424882 431593 424924 431829
rect 424604 431509 424924 431593
rect 424604 431273 424646 431509
rect 424882 431273 424924 431509
rect 424604 431241 424924 431273
rect 440076 431829 440396 431861
rect 440076 431593 440118 431829
rect 440354 431593 440396 431829
rect 440076 431509 440396 431593
rect 440076 431273 440118 431509
rect 440354 431273 440396 431509
rect 440076 431241 440396 431273
rect 446340 431829 446660 431861
rect 446340 431593 446382 431829
rect 446618 431593 446660 431829
rect 446340 431509 446660 431593
rect 446340 431273 446382 431509
rect 446618 431273 446660 431509
rect 446340 431241 446660 431273
rect 452604 431829 452924 431861
rect 452604 431593 452646 431829
rect 452882 431593 452924 431829
rect 452604 431509 452924 431593
rect 452604 431273 452646 431509
rect 452882 431273 452924 431509
rect 452604 431241 452924 431273
rect 468076 431829 468396 431861
rect 468076 431593 468118 431829
rect 468354 431593 468396 431829
rect 468076 431509 468396 431593
rect 468076 431273 468118 431509
rect 468354 431273 468396 431509
rect 468076 431241 468396 431273
rect 474340 431829 474660 431861
rect 474340 431593 474382 431829
rect 474618 431593 474660 431829
rect 474340 431509 474660 431593
rect 474340 431273 474382 431509
rect 474618 431273 474660 431509
rect 474340 431241 474660 431273
rect 480604 431829 480924 431861
rect 480604 431593 480646 431829
rect 480882 431593 480924 431829
rect 480604 431509 480924 431593
rect 480604 431273 480646 431509
rect 480882 431273 480924 431509
rect 480604 431241 480924 431273
rect 496076 431829 496396 431861
rect 496076 431593 496118 431829
rect 496354 431593 496396 431829
rect 496076 431509 496396 431593
rect 496076 431273 496118 431509
rect 496354 431273 496396 431509
rect 496076 431241 496396 431273
rect 502340 431829 502660 431861
rect 502340 431593 502382 431829
rect 502618 431593 502660 431829
rect 502340 431509 502660 431593
rect 502340 431273 502382 431509
rect 502618 431273 502660 431509
rect 502340 431241 502660 431273
rect 508604 431829 508924 431861
rect 508604 431593 508646 431829
rect 508882 431593 508924 431829
rect 508604 431509 508924 431593
rect 508604 431273 508646 431509
rect 508882 431273 508924 431509
rect 508604 431241 508924 431273
rect 524076 431829 524396 431861
rect 524076 431593 524118 431829
rect 524354 431593 524396 431829
rect 524076 431509 524396 431593
rect 524076 431273 524118 431509
rect 524354 431273 524396 431509
rect 524076 431241 524396 431273
rect 530340 431829 530660 431861
rect 530340 431593 530382 431829
rect 530618 431593 530660 431829
rect 530340 431509 530660 431593
rect 530340 431273 530382 431509
rect 530618 431273 530660 431509
rect 530340 431241 530660 431273
rect 536604 431829 536924 431861
rect 536604 431593 536646 431829
rect 536882 431593 536924 431829
rect 536604 431509 536924 431593
rect 536604 431273 536646 431509
rect 536882 431273 536924 431509
rect 536604 431241 536924 431273
rect 552076 431829 552396 431861
rect 552076 431593 552118 431829
rect 552354 431593 552396 431829
rect 552076 431509 552396 431593
rect 552076 431273 552118 431509
rect 552354 431273 552396 431509
rect 552076 431241 552396 431273
rect 558340 431829 558660 431861
rect 558340 431593 558382 431829
rect 558618 431593 558660 431829
rect 558340 431509 558660 431593
rect 558340 431273 558382 431509
rect 558618 431273 558660 431509
rect 558340 431241 558660 431273
rect 564604 431829 564924 431861
rect 564604 431593 564646 431829
rect 564882 431593 564924 431829
rect 564604 431509 564924 431593
rect 564604 431273 564646 431509
rect 564882 431273 564924 431509
rect 564604 431241 564924 431273
rect 573494 431829 574114 458273
rect 573494 431593 573526 431829
rect 573762 431593 573846 431829
rect 574082 431593 574114 431829
rect 573494 431509 574114 431593
rect 573494 431273 573526 431509
rect 573762 431273 573846 431509
rect 574082 431273 574114 431509
rect 456379 431220 456445 431221
rect 456379 431156 456380 431220
rect 456444 431156 456445 431220
rect 456379 431155 456445 431156
rect 484347 431220 484413 431221
rect 484347 431156 484348 431220
rect 484412 431156 484413 431220
rect 484347 431155 484413 431156
rect 492627 431220 492693 431221
rect 492627 431156 492628 431220
rect 492692 431156 492693 431220
rect 492627 431155 492693 431156
rect 520595 431220 520661 431221
rect 520595 431156 520596 431220
rect 520660 431156 520661 431220
rect 520595 431155 520661 431156
rect 393472 428454 393792 428486
rect 393472 428218 393514 428454
rect 393750 428218 393792 428454
rect 393472 428134 393792 428218
rect 393472 427898 393514 428134
rect 393750 427898 393792 428134
rect 393472 427866 393792 427898
rect 415208 428454 415528 428486
rect 415208 428218 415250 428454
rect 415486 428218 415528 428454
rect 415208 428134 415528 428218
rect 415208 427898 415250 428134
rect 415486 427898 415528 428134
rect 415208 427866 415528 427898
rect 421472 428454 421792 428486
rect 421472 428218 421514 428454
rect 421750 428218 421792 428454
rect 421472 428134 421792 428218
rect 421472 427898 421514 428134
rect 421750 427898 421792 428134
rect 421472 427866 421792 427898
rect 443208 428454 443528 428486
rect 443208 428218 443250 428454
rect 443486 428218 443528 428454
rect 443208 428134 443528 428218
rect 443208 427898 443250 428134
rect 443486 427898 443528 428134
rect 443208 427866 443528 427898
rect 449472 428454 449792 428486
rect 449472 428218 449514 428454
rect 449750 428218 449792 428454
rect 449472 428134 449792 428218
rect 449472 427898 449514 428134
rect 449750 427898 449792 428134
rect 449472 427866 449792 427898
rect 456382 423197 456442 431155
rect 471208 428454 471528 428486
rect 471208 428218 471250 428454
rect 471486 428218 471528 428454
rect 471208 428134 471528 428218
rect 471208 427898 471250 428134
rect 471486 427898 471528 428134
rect 471208 427866 471528 427898
rect 477472 428454 477792 428486
rect 477472 428218 477514 428454
rect 477750 428218 477792 428454
rect 477472 428134 477792 428218
rect 477472 427898 477514 428134
rect 477750 427898 477792 428134
rect 477472 427866 477792 427898
rect 456379 423196 456445 423197
rect 456379 423132 456380 423196
rect 456444 423132 456445 423196
rect 456379 423131 456445 423132
rect 484350 423061 484410 431155
rect 492630 423197 492690 431155
rect 499208 428454 499528 428486
rect 499208 428218 499250 428454
rect 499486 428218 499528 428454
rect 499208 428134 499528 428218
rect 499208 427898 499250 428134
rect 499486 427898 499528 428134
rect 499208 427866 499528 427898
rect 505472 428454 505792 428486
rect 505472 428218 505514 428454
rect 505750 428218 505792 428454
rect 505472 428134 505792 428218
rect 505472 427898 505514 428134
rect 505750 427898 505792 428134
rect 505472 427866 505792 427898
rect 520598 423333 520658 431155
rect 527208 428454 527528 428486
rect 527208 428218 527250 428454
rect 527486 428218 527528 428454
rect 527208 428134 527528 428218
rect 527208 427898 527250 428134
rect 527486 427898 527528 428134
rect 527208 427866 527528 427898
rect 533472 428454 533792 428486
rect 533472 428218 533514 428454
rect 533750 428218 533792 428454
rect 533472 428134 533792 428218
rect 533472 427898 533514 428134
rect 533750 427898 533792 428134
rect 533472 427866 533792 427898
rect 555208 428454 555528 428486
rect 555208 428218 555250 428454
rect 555486 428218 555528 428454
rect 555208 428134 555528 428218
rect 555208 427898 555250 428134
rect 555486 427898 555528 428134
rect 555208 427866 555528 427898
rect 561472 428454 561792 428486
rect 561472 428218 561514 428454
rect 561750 428218 561792 428454
rect 561472 428134 561792 428218
rect 561472 427898 561514 428134
rect 561750 427898 561792 428134
rect 561472 427866 561792 427898
rect 520595 423332 520661 423333
rect 520595 423268 520596 423332
rect 520660 423268 520661 423332
rect 520595 423267 520661 423268
rect 492627 423196 492693 423197
rect 492627 423132 492628 423196
rect 492692 423132 492693 423196
rect 492627 423131 492693 423132
rect 484347 423060 484413 423061
rect 484347 422996 484348 423060
rect 484412 422996 484413 423060
rect 484347 422995 484413 422996
rect 128307 419524 128373 419525
rect 128307 419460 128308 419524
rect 128372 419460 128373 419524
rect 128307 419459 128373 419460
rect 194731 419524 194797 419525
rect 194731 419460 194732 419524
rect 194796 419460 194797 419524
rect 194731 419459 194797 419460
rect 390875 419524 390941 419525
rect 390875 419460 390876 419524
rect 390940 419460 390941 419524
rect 390875 419459 390941 419460
rect 81387 414492 81453 414493
rect 81387 414428 81388 414492
rect 81452 414428 81453 414492
rect 81387 414427 81453 414428
rect 165659 414492 165725 414493
rect 165659 414428 165660 414492
rect 165724 414428 165725 414492
rect 165659 414427 165725 414428
rect 259499 414492 259565 414493
rect 259499 414428 259500 414492
rect 259564 414428 259565 414492
rect 259499 414427 259565 414428
rect 361619 414492 361685 414493
rect 361619 414428 361620 414492
rect 361684 414428 361685 414492
rect 361619 414427 361685 414428
rect 445707 414492 445773 414493
rect 445707 414428 445708 414492
rect 445772 414428 445773 414492
rect 445707 414427 445773 414428
rect 455459 414492 455525 414493
rect 455459 414428 455460 414492
rect 455524 414428 455525 414492
rect 455459 414427 455525 414428
rect 557579 414492 557645 414493
rect 557579 414428 557580 414492
rect 557644 414428 557645 414492
rect 557579 414427 557645 414428
rect -2006 404593 -1974 404829
rect -1738 404593 -1654 404829
rect -1418 404593 -1386 404829
rect -2006 404509 -1386 404593
rect -2006 404273 -1974 404509
rect -1738 404273 -1654 404509
rect -1418 404273 -1386 404509
rect -2006 377829 -1386 404273
rect 20076 404829 20396 404861
rect 20076 404593 20118 404829
rect 20354 404593 20396 404829
rect 20076 404509 20396 404593
rect 20076 404273 20118 404509
rect 20354 404273 20396 404509
rect 20076 404241 20396 404273
rect 26340 404829 26660 404861
rect 26340 404593 26382 404829
rect 26618 404593 26660 404829
rect 26340 404509 26660 404593
rect 26340 404273 26382 404509
rect 26618 404273 26660 404509
rect 26340 404241 26660 404273
rect 32604 404829 32924 404861
rect 32604 404593 32646 404829
rect 32882 404593 32924 404829
rect 32604 404509 32924 404593
rect 32604 404273 32646 404509
rect 32882 404273 32924 404509
rect 32604 404241 32924 404273
rect 48076 404829 48396 404861
rect 48076 404593 48118 404829
rect 48354 404593 48396 404829
rect 48076 404509 48396 404593
rect 48076 404273 48118 404509
rect 48354 404273 48396 404509
rect 48076 404241 48396 404273
rect 54340 404829 54660 404861
rect 54340 404593 54382 404829
rect 54618 404593 54660 404829
rect 54340 404509 54660 404593
rect 54340 404273 54382 404509
rect 54618 404273 54660 404509
rect 54340 404241 54660 404273
rect 60604 404829 60924 404861
rect 60604 404593 60646 404829
rect 60882 404593 60924 404829
rect 60604 404509 60924 404593
rect 60604 404273 60646 404509
rect 60882 404273 60924 404509
rect 60604 404241 60924 404273
rect 76076 404829 76396 404861
rect 76076 404593 76118 404829
rect 76354 404593 76396 404829
rect 76076 404509 76396 404593
rect 76076 404273 76118 404509
rect 76354 404273 76396 404509
rect 76076 404241 76396 404273
rect 44587 403748 44653 403749
rect 44587 403684 44588 403748
rect 44652 403684 44653 403748
rect 44587 403683 44653 403684
rect 23208 401454 23528 401486
rect 23208 401218 23250 401454
rect 23486 401218 23528 401454
rect 23208 401134 23528 401218
rect 23208 400898 23250 401134
rect 23486 400898 23528 401134
rect 23208 400866 23528 400898
rect 29472 401454 29792 401486
rect 29472 401218 29514 401454
rect 29750 401218 29792 401454
rect 29472 401134 29792 401218
rect 29472 400898 29514 401134
rect 29750 400898 29792 401134
rect 29472 400866 29792 400898
rect 44590 395861 44650 403683
rect 51208 401454 51528 401486
rect 51208 401218 51250 401454
rect 51486 401218 51528 401454
rect 51208 401134 51528 401218
rect 51208 400898 51250 401134
rect 51486 400898 51528 401134
rect 51208 400866 51528 400898
rect 57472 401454 57792 401486
rect 57472 401218 57514 401454
rect 57750 401218 57792 401454
rect 57472 401134 57792 401218
rect 57472 400898 57514 401134
rect 57750 400898 57792 401134
rect 57472 400866 57792 400898
rect 79208 401454 79528 401486
rect 79208 401218 79250 401454
rect 79486 401218 79528 401454
rect 79208 401134 79528 401218
rect 79208 400898 79250 401134
rect 79486 400898 79528 401134
rect 79208 400866 79528 400898
rect 44587 395860 44653 395861
rect 44587 395796 44588 395860
rect 44652 395796 44653 395860
rect 44587 395795 44653 395796
rect 81390 391917 81450 414427
rect 82340 404829 82660 404861
rect 82340 404593 82382 404829
rect 82618 404593 82660 404829
rect 82340 404509 82660 404593
rect 82340 404273 82382 404509
rect 82618 404273 82660 404509
rect 82340 404241 82660 404273
rect 88604 404829 88924 404861
rect 88604 404593 88646 404829
rect 88882 404593 88924 404829
rect 88604 404509 88924 404593
rect 88604 404273 88646 404509
rect 88882 404273 88924 404509
rect 88604 404241 88924 404273
rect 104076 404829 104396 404861
rect 104076 404593 104118 404829
rect 104354 404593 104396 404829
rect 104076 404509 104396 404593
rect 104076 404273 104118 404509
rect 104354 404273 104396 404509
rect 104076 404241 104396 404273
rect 110340 404829 110660 404861
rect 110340 404593 110382 404829
rect 110618 404593 110660 404829
rect 110340 404509 110660 404593
rect 110340 404273 110382 404509
rect 110618 404273 110660 404509
rect 110340 404241 110660 404273
rect 116604 404829 116924 404861
rect 116604 404593 116646 404829
rect 116882 404593 116924 404829
rect 116604 404509 116924 404593
rect 116604 404273 116646 404509
rect 116882 404273 116924 404509
rect 116604 404241 116924 404273
rect 132076 404829 132396 404861
rect 132076 404593 132118 404829
rect 132354 404593 132396 404829
rect 132076 404509 132396 404593
rect 132076 404273 132118 404509
rect 132354 404273 132396 404509
rect 132076 404241 132396 404273
rect 138340 404829 138660 404861
rect 138340 404593 138382 404829
rect 138618 404593 138660 404829
rect 138340 404509 138660 404593
rect 138340 404273 138382 404509
rect 138618 404273 138660 404509
rect 138340 404241 138660 404273
rect 144604 404829 144924 404861
rect 144604 404593 144646 404829
rect 144882 404593 144924 404829
rect 144604 404509 144924 404593
rect 144604 404273 144646 404509
rect 144882 404273 144924 404509
rect 144604 404241 144924 404273
rect 160076 404829 160396 404861
rect 160076 404593 160118 404829
rect 160354 404593 160396 404829
rect 160076 404509 160396 404593
rect 160076 404273 160118 404509
rect 160354 404273 160396 404509
rect 160076 404241 160396 404273
rect 128491 403748 128557 403749
rect 128491 403684 128492 403748
rect 128556 403684 128557 403748
rect 128491 403683 128557 403684
rect 85472 401454 85792 401486
rect 85472 401218 85514 401454
rect 85750 401218 85792 401454
rect 85472 401134 85792 401218
rect 85472 400898 85514 401134
rect 85750 400898 85792 401134
rect 85472 400866 85792 400898
rect 107208 401454 107528 401486
rect 107208 401218 107250 401454
rect 107486 401218 107528 401454
rect 107208 401134 107528 401218
rect 107208 400898 107250 401134
rect 107486 400898 107528 401134
rect 107208 400866 107528 400898
rect 113472 401454 113792 401486
rect 113472 401218 113514 401454
rect 113750 401218 113792 401454
rect 113472 401134 113792 401218
rect 113472 400898 113514 401134
rect 113750 400898 113792 401134
rect 113472 400866 113792 400898
rect 128494 395997 128554 403683
rect 135208 401454 135528 401486
rect 135208 401218 135250 401454
rect 135486 401218 135528 401454
rect 135208 401134 135528 401218
rect 135208 400898 135250 401134
rect 135486 400898 135528 401134
rect 135208 400866 135528 400898
rect 141472 401454 141792 401486
rect 141472 401218 141514 401454
rect 141750 401218 141792 401454
rect 141472 401134 141792 401218
rect 141472 400898 141514 401134
rect 141750 400898 141792 401134
rect 141472 400866 141792 400898
rect 163208 401454 163528 401486
rect 163208 401218 163250 401454
rect 163486 401218 163528 401454
rect 163208 401134 163528 401218
rect 163208 400898 163250 401134
rect 163486 400898 163528 401134
rect 163208 400866 163528 400898
rect 128491 395996 128557 395997
rect 128491 395932 128492 395996
rect 128556 395932 128557 395996
rect 128491 395931 128557 395932
rect 165662 391917 165722 414427
rect 166340 404829 166660 404861
rect 166340 404593 166382 404829
rect 166618 404593 166660 404829
rect 166340 404509 166660 404593
rect 166340 404273 166382 404509
rect 166618 404273 166660 404509
rect 166340 404241 166660 404273
rect 172604 404829 172924 404861
rect 172604 404593 172646 404829
rect 172882 404593 172924 404829
rect 172604 404509 172924 404593
rect 172604 404273 172646 404509
rect 172882 404273 172924 404509
rect 172604 404241 172924 404273
rect 188076 404829 188396 404861
rect 188076 404593 188118 404829
rect 188354 404593 188396 404829
rect 188076 404509 188396 404593
rect 188076 404273 188118 404509
rect 188354 404273 188396 404509
rect 188076 404241 188396 404273
rect 194340 404829 194660 404861
rect 194340 404593 194382 404829
rect 194618 404593 194660 404829
rect 194340 404509 194660 404593
rect 194340 404273 194382 404509
rect 194618 404273 194660 404509
rect 194340 404241 194660 404273
rect 200604 404829 200924 404861
rect 200604 404593 200646 404829
rect 200882 404593 200924 404829
rect 200604 404509 200924 404593
rect 200604 404273 200646 404509
rect 200882 404273 200924 404509
rect 200604 404241 200924 404273
rect 216076 404829 216396 404861
rect 216076 404593 216118 404829
rect 216354 404593 216396 404829
rect 216076 404509 216396 404593
rect 216076 404273 216118 404509
rect 216354 404273 216396 404509
rect 216076 404241 216396 404273
rect 222340 404829 222660 404861
rect 222340 404593 222382 404829
rect 222618 404593 222660 404829
rect 222340 404509 222660 404593
rect 222340 404273 222382 404509
rect 222618 404273 222660 404509
rect 222340 404241 222660 404273
rect 228604 404829 228924 404861
rect 228604 404593 228646 404829
rect 228882 404593 228924 404829
rect 228604 404509 228924 404593
rect 228604 404273 228646 404509
rect 228882 404273 228924 404509
rect 228604 404241 228924 404273
rect 244076 404829 244396 404861
rect 244076 404593 244118 404829
rect 244354 404593 244396 404829
rect 244076 404509 244396 404593
rect 244076 404273 244118 404509
rect 244354 404273 244396 404509
rect 244076 404241 244396 404273
rect 250340 404829 250660 404861
rect 250340 404593 250382 404829
rect 250618 404593 250660 404829
rect 250340 404509 250660 404593
rect 250340 404273 250382 404509
rect 250618 404273 250660 404509
rect 250340 404241 250660 404273
rect 256604 404829 256924 404861
rect 256604 404593 256646 404829
rect 256882 404593 256924 404829
rect 256604 404509 256924 404593
rect 256604 404273 256646 404509
rect 256882 404273 256924 404509
rect 256604 404241 256924 404273
rect 212579 403748 212645 403749
rect 212579 403684 212580 403748
rect 212644 403684 212645 403748
rect 212579 403683 212645 403684
rect 240547 403748 240613 403749
rect 240547 403684 240548 403748
rect 240612 403684 240613 403748
rect 240547 403683 240613 403684
rect 169472 401454 169792 401486
rect 169472 401218 169514 401454
rect 169750 401218 169792 401454
rect 169472 401134 169792 401218
rect 169472 400898 169514 401134
rect 169750 400898 169792 401134
rect 169472 400866 169792 400898
rect 191208 401454 191528 401486
rect 191208 401218 191250 401454
rect 191486 401218 191528 401454
rect 191208 401134 191528 401218
rect 191208 400898 191250 401134
rect 191486 400898 191528 401134
rect 191208 400866 191528 400898
rect 197472 401454 197792 401486
rect 197472 401218 197514 401454
rect 197750 401218 197792 401454
rect 197472 401134 197792 401218
rect 197472 400898 197514 401134
rect 197750 400898 197792 401134
rect 197472 400866 197792 400898
rect 212582 395725 212642 403683
rect 219208 401454 219528 401486
rect 219208 401218 219250 401454
rect 219486 401218 219528 401454
rect 219208 401134 219528 401218
rect 219208 400898 219250 401134
rect 219486 400898 219528 401134
rect 219208 400866 219528 400898
rect 225472 401454 225792 401486
rect 225472 401218 225514 401454
rect 225750 401218 225792 401454
rect 225472 401134 225792 401218
rect 225472 400898 225514 401134
rect 225750 400898 225792 401134
rect 225472 400866 225792 400898
rect 240550 395861 240610 403683
rect 247208 401454 247528 401486
rect 247208 401218 247250 401454
rect 247486 401218 247528 401454
rect 247208 401134 247528 401218
rect 247208 400898 247250 401134
rect 247486 400898 247528 401134
rect 247208 400866 247528 400898
rect 253472 401454 253792 401486
rect 253472 401218 253514 401454
rect 253750 401218 253792 401454
rect 253472 401134 253792 401218
rect 253472 400898 253514 401134
rect 253750 400898 253792 401134
rect 253472 400866 253792 400898
rect 240547 395860 240613 395861
rect 240547 395796 240548 395860
rect 240612 395796 240613 395860
rect 240547 395795 240613 395796
rect 212579 395724 212645 395725
rect 212579 395660 212580 395724
rect 212644 395660 212645 395724
rect 212579 395659 212645 395660
rect 259502 391917 259562 414427
rect 272076 404829 272396 404861
rect 272076 404593 272118 404829
rect 272354 404593 272396 404829
rect 272076 404509 272396 404593
rect 272076 404273 272118 404509
rect 272354 404273 272396 404509
rect 272076 404241 272396 404273
rect 278340 404829 278660 404861
rect 278340 404593 278382 404829
rect 278618 404593 278660 404829
rect 278340 404509 278660 404593
rect 278340 404273 278382 404509
rect 278618 404273 278660 404509
rect 278340 404241 278660 404273
rect 284604 404829 284924 404861
rect 284604 404593 284646 404829
rect 284882 404593 284924 404829
rect 284604 404509 284924 404593
rect 284604 404273 284646 404509
rect 284882 404273 284924 404509
rect 284604 404241 284924 404273
rect 300076 404829 300396 404861
rect 300076 404593 300118 404829
rect 300354 404593 300396 404829
rect 300076 404509 300396 404593
rect 300076 404273 300118 404509
rect 300354 404273 300396 404509
rect 300076 404241 300396 404273
rect 306340 404829 306660 404861
rect 306340 404593 306382 404829
rect 306618 404593 306660 404829
rect 306340 404509 306660 404593
rect 306340 404273 306382 404509
rect 306618 404273 306660 404509
rect 306340 404241 306660 404273
rect 312604 404829 312924 404861
rect 312604 404593 312646 404829
rect 312882 404593 312924 404829
rect 312604 404509 312924 404593
rect 312604 404273 312646 404509
rect 312882 404273 312924 404509
rect 312604 404241 312924 404273
rect 328076 404829 328396 404861
rect 328076 404593 328118 404829
rect 328354 404593 328396 404829
rect 328076 404509 328396 404593
rect 328076 404273 328118 404509
rect 328354 404273 328396 404509
rect 328076 404241 328396 404273
rect 334340 404829 334660 404861
rect 334340 404593 334382 404829
rect 334618 404593 334660 404829
rect 334340 404509 334660 404593
rect 334340 404273 334382 404509
rect 334618 404273 334660 404509
rect 334340 404241 334660 404273
rect 340604 404829 340924 404861
rect 340604 404593 340646 404829
rect 340882 404593 340924 404829
rect 340604 404509 340924 404593
rect 340604 404273 340646 404509
rect 340882 404273 340924 404509
rect 340604 404241 340924 404273
rect 356076 404829 356396 404861
rect 356076 404593 356118 404829
rect 356354 404593 356396 404829
rect 356076 404509 356396 404593
rect 356076 404273 356118 404509
rect 356354 404273 356396 404509
rect 356076 404241 356396 404273
rect 296483 403748 296549 403749
rect 296483 403684 296484 403748
rect 296548 403684 296549 403748
rect 296483 403683 296549 403684
rect 324635 403748 324701 403749
rect 324635 403684 324636 403748
rect 324700 403684 324701 403748
rect 324635 403683 324701 403684
rect 275208 401454 275528 401486
rect 275208 401218 275250 401454
rect 275486 401218 275528 401454
rect 275208 401134 275528 401218
rect 275208 400898 275250 401134
rect 275486 400898 275528 401134
rect 275208 400866 275528 400898
rect 281472 401454 281792 401486
rect 281472 401218 281514 401454
rect 281750 401218 281792 401454
rect 281472 401134 281792 401218
rect 281472 400898 281514 401134
rect 281750 400898 281792 401134
rect 281472 400866 281792 400898
rect 296486 396090 296546 403683
rect 303208 401454 303528 401486
rect 303208 401218 303250 401454
rect 303486 401218 303528 401454
rect 303208 401134 303528 401218
rect 303208 400898 303250 401134
rect 303486 400898 303528 401134
rect 303208 400866 303528 400898
rect 309472 401454 309792 401486
rect 309472 401218 309514 401454
rect 309750 401218 309792 401454
rect 309472 401134 309792 401218
rect 309472 400898 309514 401134
rect 309750 400898 309792 401134
rect 309472 400866 309792 400898
rect 296486 396030 296914 396090
rect 296854 395725 296914 396030
rect 324638 395861 324698 403683
rect 331208 401454 331528 401486
rect 331208 401218 331250 401454
rect 331486 401218 331528 401454
rect 331208 401134 331528 401218
rect 331208 400898 331250 401134
rect 331486 400898 331528 401134
rect 331208 400866 331528 400898
rect 337472 401454 337792 401486
rect 337472 401218 337514 401454
rect 337750 401218 337792 401454
rect 337472 401134 337792 401218
rect 337472 400898 337514 401134
rect 337750 400898 337792 401134
rect 337472 400866 337792 400898
rect 359208 401454 359528 401486
rect 359208 401218 359250 401454
rect 359486 401218 359528 401454
rect 359208 401134 359528 401218
rect 359208 400898 359250 401134
rect 359486 400898 359528 401134
rect 359208 400866 359528 400898
rect 324635 395860 324701 395861
rect 324635 395796 324636 395860
rect 324700 395796 324701 395860
rect 324635 395795 324701 395796
rect 296851 395724 296917 395725
rect 296851 395660 296852 395724
rect 296916 395660 296917 395724
rect 296851 395659 296917 395660
rect 361622 391917 361682 414427
rect 362340 404829 362660 404861
rect 362340 404593 362382 404829
rect 362618 404593 362660 404829
rect 362340 404509 362660 404593
rect 362340 404273 362382 404509
rect 362618 404273 362660 404509
rect 362340 404241 362660 404273
rect 368604 404829 368924 404861
rect 368604 404593 368646 404829
rect 368882 404593 368924 404829
rect 368604 404509 368924 404593
rect 368604 404273 368646 404509
rect 368882 404273 368924 404509
rect 368604 404241 368924 404273
rect 384076 404829 384396 404861
rect 384076 404593 384118 404829
rect 384354 404593 384396 404829
rect 384076 404509 384396 404593
rect 384076 404273 384118 404509
rect 384354 404273 384396 404509
rect 384076 404241 384396 404273
rect 390340 404829 390660 404861
rect 390340 404593 390382 404829
rect 390618 404593 390660 404829
rect 390340 404509 390660 404593
rect 390340 404273 390382 404509
rect 390618 404273 390660 404509
rect 390340 404241 390660 404273
rect 396604 404829 396924 404861
rect 396604 404593 396646 404829
rect 396882 404593 396924 404829
rect 396604 404509 396924 404593
rect 396604 404273 396646 404509
rect 396882 404273 396924 404509
rect 396604 404241 396924 404273
rect 412076 404829 412396 404861
rect 412076 404593 412118 404829
rect 412354 404593 412396 404829
rect 412076 404509 412396 404593
rect 412076 404273 412118 404509
rect 412354 404273 412396 404509
rect 412076 404241 412396 404273
rect 418340 404829 418660 404861
rect 418340 404593 418382 404829
rect 418618 404593 418660 404829
rect 418340 404509 418660 404593
rect 418340 404273 418382 404509
rect 418618 404273 418660 404509
rect 418340 404241 418660 404273
rect 424604 404829 424924 404861
rect 424604 404593 424646 404829
rect 424882 404593 424924 404829
rect 424604 404509 424924 404593
rect 424604 404273 424646 404509
rect 424882 404273 424924 404509
rect 424604 404241 424924 404273
rect 440076 404829 440396 404861
rect 440076 404593 440118 404829
rect 440354 404593 440396 404829
rect 440076 404509 440396 404593
rect 440076 404273 440118 404509
rect 440354 404273 440396 404509
rect 440076 404241 440396 404273
rect 408539 403748 408605 403749
rect 408539 403684 408540 403748
rect 408604 403684 408605 403748
rect 408539 403683 408605 403684
rect 436507 403748 436573 403749
rect 436507 403684 436508 403748
rect 436572 403684 436573 403748
rect 436507 403683 436573 403684
rect 365472 401454 365792 401486
rect 365472 401218 365514 401454
rect 365750 401218 365792 401454
rect 365472 401134 365792 401218
rect 365472 400898 365514 401134
rect 365750 400898 365792 401134
rect 365472 400866 365792 400898
rect 387208 401454 387528 401486
rect 387208 401218 387250 401454
rect 387486 401218 387528 401454
rect 387208 401134 387528 401218
rect 387208 400898 387250 401134
rect 387486 400898 387528 401134
rect 387208 400866 387528 400898
rect 393472 401454 393792 401486
rect 393472 401218 393514 401454
rect 393750 401218 393792 401454
rect 393472 401134 393792 401218
rect 393472 400898 393514 401134
rect 393750 400898 393792 401134
rect 393472 400866 393792 400898
rect 408542 395997 408602 403683
rect 415208 401454 415528 401486
rect 415208 401218 415250 401454
rect 415486 401218 415528 401454
rect 415208 401134 415528 401218
rect 415208 400898 415250 401134
rect 415486 400898 415528 401134
rect 415208 400866 415528 400898
rect 421472 401454 421792 401486
rect 421472 401218 421514 401454
rect 421750 401218 421792 401454
rect 421472 401134 421792 401218
rect 421472 400898 421514 401134
rect 421750 400898 421792 401134
rect 421472 400866 421792 400898
rect 408539 395996 408605 395997
rect 408539 395932 408540 395996
rect 408604 395932 408605 395996
rect 408539 395931 408605 395932
rect 436510 395861 436570 403683
rect 443208 401454 443528 401486
rect 443208 401218 443250 401454
rect 443486 401218 443528 401454
rect 443208 401134 443528 401218
rect 443208 400898 443250 401134
rect 443486 400898 443528 401134
rect 443208 400866 443528 400898
rect 436507 395860 436573 395861
rect 436507 395796 436508 395860
rect 436572 395796 436573 395860
rect 436507 395795 436573 395796
rect 81387 391916 81453 391917
rect 81387 391852 81388 391916
rect 81452 391852 81453 391916
rect 81387 391851 81453 391852
rect 165659 391916 165725 391917
rect 165659 391852 165660 391916
rect 165724 391852 165725 391916
rect 165659 391851 165725 391852
rect 259499 391916 259565 391917
rect 259499 391852 259500 391916
rect 259564 391852 259565 391916
rect 259499 391851 259565 391852
rect 361619 391916 361685 391917
rect 361619 391852 361620 391916
rect 361684 391852 361685 391916
rect 361619 391851 361685 391852
rect 445710 391781 445770 414427
rect 446340 404829 446660 404861
rect 446340 404593 446382 404829
rect 446618 404593 446660 404829
rect 446340 404509 446660 404593
rect 446340 404273 446382 404509
rect 446618 404273 446660 404509
rect 446340 404241 446660 404273
rect 452604 404829 452924 404861
rect 452604 404593 452646 404829
rect 452882 404593 452924 404829
rect 452604 404509 452924 404593
rect 452604 404273 452646 404509
rect 452882 404273 452924 404509
rect 452604 404241 452924 404273
rect 449472 401454 449792 401486
rect 449472 401218 449514 401454
rect 449750 401218 449792 401454
rect 449472 401134 449792 401218
rect 449472 400898 449514 401134
rect 449750 400898 449792 401134
rect 449472 400866 449792 400898
rect 455462 391917 455522 414427
rect 468076 404829 468396 404861
rect 468076 404593 468118 404829
rect 468354 404593 468396 404829
rect 468076 404509 468396 404593
rect 468076 404273 468118 404509
rect 468354 404273 468396 404509
rect 468076 404241 468396 404273
rect 474340 404829 474660 404861
rect 474340 404593 474382 404829
rect 474618 404593 474660 404829
rect 474340 404509 474660 404593
rect 474340 404273 474382 404509
rect 474618 404273 474660 404509
rect 474340 404241 474660 404273
rect 480604 404829 480924 404861
rect 480604 404593 480646 404829
rect 480882 404593 480924 404829
rect 480604 404509 480924 404593
rect 480604 404273 480646 404509
rect 480882 404273 480924 404509
rect 480604 404241 480924 404273
rect 496076 404829 496396 404861
rect 496076 404593 496118 404829
rect 496354 404593 496396 404829
rect 496076 404509 496396 404593
rect 496076 404273 496118 404509
rect 496354 404273 496396 404509
rect 496076 404241 496396 404273
rect 502340 404829 502660 404861
rect 502340 404593 502382 404829
rect 502618 404593 502660 404829
rect 502340 404509 502660 404593
rect 502340 404273 502382 404509
rect 502618 404273 502660 404509
rect 502340 404241 502660 404273
rect 508604 404829 508924 404861
rect 508604 404593 508646 404829
rect 508882 404593 508924 404829
rect 508604 404509 508924 404593
rect 508604 404273 508646 404509
rect 508882 404273 508924 404509
rect 508604 404241 508924 404273
rect 524076 404829 524396 404861
rect 524076 404593 524118 404829
rect 524354 404593 524396 404829
rect 524076 404509 524396 404593
rect 524076 404273 524118 404509
rect 524354 404273 524396 404509
rect 524076 404241 524396 404273
rect 530340 404829 530660 404861
rect 530340 404593 530382 404829
rect 530618 404593 530660 404829
rect 530340 404509 530660 404593
rect 530340 404273 530382 404509
rect 530618 404273 530660 404509
rect 530340 404241 530660 404273
rect 536604 404829 536924 404861
rect 536604 404593 536646 404829
rect 536882 404593 536924 404829
rect 536604 404509 536924 404593
rect 536604 404273 536646 404509
rect 536882 404273 536924 404509
rect 536604 404241 536924 404273
rect 552076 404829 552396 404861
rect 552076 404593 552118 404829
rect 552354 404593 552396 404829
rect 552076 404509 552396 404593
rect 552076 404273 552118 404509
rect 552354 404273 552396 404509
rect 552076 404241 552396 404273
rect 492627 403748 492693 403749
rect 492627 403684 492628 403748
rect 492692 403684 492693 403748
rect 492627 403683 492693 403684
rect 520595 403748 520661 403749
rect 520595 403684 520596 403748
rect 520660 403684 520661 403748
rect 520595 403683 520661 403684
rect 471208 401454 471528 401486
rect 471208 401218 471250 401454
rect 471486 401218 471528 401454
rect 471208 401134 471528 401218
rect 471208 400898 471250 401134
rect 471486 400898 471528 401134
rect 471208 400866 471528 400898
rect 477472 401454 477792 401486
rect 477472 401218 477514 401454
rect 477750 401218 477792 401454
rect 477472 401134 477792 401218
rect 477472 400898 477514 401134
rect 477750 400898 477792 401134
rect 477472 400866 477792 400898
rect 492630 395861 492690 403683
rect 499208 401454 499528 401486
rect 499208 401218 499250 401454
rect 499486 401218 499528 401454
rect 499208 401134 499528 401218
rect 499208 400898 499250 401134
rect 499486 400898 499528 401134
rect 499208 400866 499528 400898
rect 505472 401454 505792 401486
rect 505472 401218 505514 401454
rect 505750 401218 505792 401454
rect 505472 401134 505792 401218
rect 505472 400898 505514 401134
rect 505750 400898 505792 401134
rect 505472 400866 505792 400898
rect 520598 395997 520658 403683
rect 527208 401454 527528 401486
rect 527208 401218 527250 401454
rect 527486 401218 527528 401454
rect 527208 401134 527528 401218
rect 527208 400898 527250 401134
rect 527486 400898 527528 401134
rect 527208 400866 527528 400898
rect 533472 401454 533792 401486
rect 533472 401218 533514 401454
rect 533750 401218 533792 401454
rect 533472 401134 533792 401218
rect 533472 400898 533514 401134
rect 533750 400898 533792 401134
rect 533472 400866 533792 400898
rect 555208 401454 555528 401486
rect 555208 401218 555250 401454
rect 555486 401218 555528 401454
rect 555208 401134 555528 401218
rect 555208 400898 555250 401134
rect 555486 400898 555528 401134
rect 555208 400866 555528 400898
rect 520595 395996 520661 395997
rect 520595 395932 520596 395996
rect 520660 395932 520661 395996
rect 520595 395931 520661 395932
rect 492627 395860 492693 395861
rect 492627 395796 492628 395860
rect 492692 395796 492693 395860
rect 492627 395795 492693 395796
rect 557582 391917 557642 414427
rect 558340 404829 558660 404861
rect 558340 404593 558382 404829
rect 558618 404593 558660 404829
rect 558340 404509 558660 404593
rect 558340 404273 558382 404509
rect 558618 404273 558660 404509
rect 558340 404241 558660 404273
rect 564604 404829 564924 404861
rect 564604 404593 564646 404829
rect 564882 404593 564924 404829
rect 564604 404509 564924 404593
rect 564604 404273 564646 404509
rect 564882 404273 564924 404509
rect 564604 404241 564924 404273
rect 573494 404829 574114 431273
rect 573494 404593 573526 404829
rect 573762 404593 573846 404829
rect 574082 404593 574114 404829
rect 573494 404509 574114 404593
rect 573494 404273 573526 404509
rect 573762 404273 573846 404509
rect 574082 404273 574114 404509
rect 561472 401454 561792 401486
rect 561472 401218 561514 401454
rect 561750 401218 561792 401454
rect 561472 401134 561792 401218
rect 561472 400898 561514 401134
rect 561750 400898 561792 401134
rect 561472 400866 561792 400898
rect 455459 391916 455525 391917
rect 455459 391852 455460 391916
rect 455524 391852 455525 391916
rect 455459 391851 455525 391852
rect 557579 391916 557645 391917
rect 557579 391852 557580 391916
rect 557644 391852 557645 391916
rect 557579 391851 557645 391852
rect 445707 391780 445773 391781
rect 445707 391716 445708 391780
rect 445772 391716 445773 391780
rect 445707 391715 445773 391716
rect 128307 387428 128373 387429
rect 128307 387364 128308 387428
rect 128372 387364 128373 387428
rect 128307 387363 128373 387364
rect 194731 387428 194797 387429
rect 194731 387364 194732 387428
rect 194796 387364 194797 387428
rect 194731 387363 194797 387364
rect 390875 387428 390941 387429
rect 390875 387364 390876 387428
rect 390940 387364 390941 387428
rect 390875 387363 390941 387364
rect -2006 377593 -1974 377829
rect -1738 377593 -1654 377829
rect -1418 377593 -1386 377829
rect -2006 377509 -1386 377593
rect -2006 377273 -1974 377509
rect -1738 377273 -1654 377509
rect -1418 377273 -1386 377509
rect -2006 350829 -1386 377273
rect 20076 377829 20396 377861
rect 20076 377593 20118 377829
rect 20354 377593 20396 377829
rect 20076 377509 20396 377593
rect 20076 377273 20118 377509
rect 20354 377273 20396 377509
rect 20076 377241 20396 377273
rect 26340 377829 26660 377861
rect 26340 377593 26382 377829
rect 26618 377593 26660 377829
rect 26340 377509 26660 377593
rect 26340 377273 26382 377509
rect 26618 377273 26660 377509
rect 26340 377241 26660 377273
rect 32604 377829 32924 377861
rect 32604 377593 32646 377829
rect 32882 377593 32924 377829
rect 32604 377509 32924 377593
rect 32604 377273 32646 377509
rect 32882 377273 32924 377509
rect 32604 377241 32924 377273
rect 48076 377829 48396 377861
rect 48076 377593 48118 377829
rect 48354 377593 48396 377829
rect 48076 377509 48396 377593
rect 48076 377273 48118 377509
rect 48354 377273 48396 377509
rect 48076 377241 48396 377273
rect 54340 377829 54660 377861
rect 54340 377593 54382 377829
rect 54618 377593 54660 377829
rect 54340 377509 54660 377593
rect 54340 377273 54382 377509
rect 54618 377273 54660 377509
rect 54340 377241 54660 377273
rect 60604 377829 60924 377861
rect 60604 377593 60646 377829
rect 60882 377593 60924 377829
rect 60604 377509 60924 377593
rect 60604 377273 60646 377509
rect 60882 377273 60924 377509
rect 60604 377241 60924 377273
rect 76076 377829 76396 377861
rect 76076 377593 76118 377829
rect 76354 377593 76396 377829
rect 76076 377509 76396 377593
rect 76076 377273 76118 377509
rect 76354 377273 76396 377509
rect 76076 377241 76396 377273
rect 82340 377829 82660 377861
rect 82340 377593 82382 377829
rect 82618 377593 82660 377829
rect 82340 377509 82660 377593
rect 82340 377273 82382 377509
rect 82618 377273 82660 377509
rect 82340 377241 82660 377273
rect 88604 377829 88924 377861
rect 88604 377593 88646 377829
rect 88882 377593 88924 377829
rect 88604 377509 88924 377593
rect 88604 377273 88646 377509
rect 88882 377273 88924 377509
rect 88604 377241 88924 377273
rect 104076 377829 104396 377861
rect 104076 377593 104118 377829
rect 104354 377593 104396 377829
rect 104076 377509 104396 377593
rect 104076 377273 104118 377509
rect 104354 377273 104396 377509
rect 104076 377241 104396 377273
rect 110340 377829 110660 377861
rect 110340 377593 110382 377829
rect 110618 377593 110660 377829
rect 110340 377509 110660 377593
rect 110340 377273 110382 377509
rect 110618 377273 110660 377509
rect 110340 377241 110660 377273
rect 116604 377829 116924 377861
rect 116604 377593 116646 377829
rect 116882 377593 116924 377829
rect 116604 377509 116924 377593
rect 116604 377273 116646 377509
rect 116882 377273 116924 377509
rect 116604 377241 116924 377273
rect 23208 374454 23528 374486
rect 23208 374218 23250 374454
rect 23486 374218 23528 374454
rect 23208 374134 23528 374218
rect 23208 373898 23250 374134
rect 23486 373898 23528 374134
rect 23208 373866 23528 373898
rect 29472 374454 29792 374486
rect 29472 374218 29514 374454
rect 29750 374218 29792 374454
rect 29472 374134 29792 374218
rect 29472 373898 29514 374134
rect 29750 373898 29792 374134
rect 29472 373866 29792 373898
rect 51208 374454 51528 374486
rect 51208 374218 51250 374454
rect 51486 374218 51528 374454
rect 51208 374134 51528 374218
rect 51208 373898 51250 374134
rect 51486 373898 51528 374134
rect 51208 373866 51528 373898
rect 57472 374454 57792 374486
rect 57472 374218 57514 374454
rect 57750 374218 57792 374454
rect 57472 374134 57792 374218
rect 57472 373898 57514 374134
rect 57750 373898 57792 374134
rect 57472 373866 57792 373898
rect 79208 374454 79528 374486
rect 79208 374218 79250 374454
rect 79486 374218 79528 374454
rect 79208 374134 79528 374218
rect 79208 373898 79250 374134
rect 79486 373898 79528 374134
rect 79208 373866 79528 373898
rect 85472 374454 85792 374486
rect 85472 374218 85514 374454
rect 85750 374218 85792 374454
rect 85472 374134 85792 374218
rect 85472 373898 85514 374134
rect 85750 373898 85792 374134
rect 85472 373866 85792 373898
rect 107208 374454 107528 374486
rect 107208 374218 107250 374454
rect 107486 374218 107528 374454
rect 107208 374134 107528 374218
rect 107208 373898 107250 374134
rect 107486 373898 107528 374134
rect 107208 373866 107528 373898
rect 113472 374454 113792 374486
rect 113472 374218 113514 374454
rect 113750 374218 113792 374454
rect 113472 374134 113792 374218
rect 113472 373898 113514 374134
rect 113750 373898 113792 374134
rect 113472 373866 113792 373898
rect 128310 365669 128370 387363
rect 132076 377829 132396 377861
rect 132076 377593 132118 377829
rect 132354 377593 132396 377829
rect 132076 377509 132396 377593
rect 132076 377273 132118 377509
rect 132354 377273 132396 377509
rect 132076 377241 132396 377273
rect 138340 377829 138660 377861
rect 138340 377593 138382 377829
rect 138618 377593 138660 377829
rect 138340 377509 138660 377593
rect 138340 377273 138382 377509
rect 138618 377273 138660 377509
rect 138340 377241 138660 377273
rect 144604 377829 144924 377861
rect 144604 377593 144646 377829
rect 144882 377593 144924 377829
rect 144604 377509 144924 377593
rect 144604 377273 144646 377509
rect 144882 377273 144924 377509
rect 144604 377241 144924 377273
rect 160076 377829 160396 377861
rect 160076 377593 160118 377829
rect 160354 377593 160396 377829
rect 160076 377509 160396 377593
rect 160076 377273 160118 377509
rect 160354 377273 160396 377509
rect 160076 377241 160396 377273
rect 166340 377829 166660 377861
rect 166340 377593 166382 377829
rect 166618 377593 166660 377829
rect 166340 377509 166660 377593
rect 166340 377273 166382 377509
rect 166618 377273 166660 377509
rect 166340 377241 166660 377273
rect 172604 377829 172924 377861
rect 172604 377593 172646 377829
rect 172882 377593 172924 377829
rect 172604 377509 172924 377593
rect 172604 377273 172646 377509
rect 172882 377273 172924 377509
rect 172604 377241 172924 377273
rect 188076 377829 188396 377861
rect 188076 377593 188118 377829
rect 188354 377593 188396 377829
rect 188076 377509 188396 377593
rect 188076 377273 188118 377509
rect 188354 377273 188396 377509
rect 188076 377241 188396 377273
rect 194340 377829 194660 377861
rect 194340 377593 194382 377829
rect 194618 377593 194660 377829
rect 194340 377509 194660 377593
rect 194340 377273 194382 377509
rect 194618 377273 194660 377509
rect 194340 377241 194660 377273
rect 176331 377228 176397 377229
rect 176331 377164 176332 377228
rect 176396 377164 176397 377228
rect 176331 377163 176397 377164
rect 135208 374454 135528 374486
rect 135208 374218 135250 374454
rect 135486 374218 135528 374454
rect 135208 374134 135528 374218
rect 135208 373898 135250 374134
rect 135486 373898 135528 374134
rect 135208 373866 135528 373898
rect 141472 374454 141792 374486
rect 141472 374218 141514 374454
rect 141750 374218 141792 374454
rect 141472 374134 141792 374218
rect 141472 373898 141514 374134
rect 141750 373898 141792 374134
rect 141472 373866 141792 373898
rect 163208 374454 163528 374486
rect 163208 374218 163250 374454
rect 163486 374218 163528 374454
rect 163208 374134 163528 374218
rect 163208 373898 163250 374134
rect 163486 373898 163528 374134
rect 163208 373866 163528 373898
rect 169472 374454 169792 374486
rect 169472 374218 169514 374454
rect 169750 374218 169792 374454
rect 169472 374134 169792 374218
rect 169472 373898 169514 374134
rect 169750 373898 169792 374134
rect 176334 374010 176394 377163
rect 169472 373866 169792 373898
rect 175230 373950 176394 374010
rect 191208 374454 191528 374486
rect 191208 374218 191250 374454
rect 191486 374218 191528 374454
rect 191208 374134 191528 374218
rect 175230 369341 175290 373950
rect 191208 373898 191250 374134
rect 191486 373898 191528 374134
rect 191208 373866 191528 373898
rect 175227 369340 175293 369341
rect 175227 369276 175228 369340
rect 175292 369276 175293 369340
rect 175227 369275 175293 369276
rect 194734 365669 194794 387363
rect 200604 377829 200924 377861
rect 200604 377593 200646 377829
rect 200882 377593 200924 377829
rect 200604 377509 200924 377593
rect 200604 377273 200646 377509
rect 200882 377273 200924 377509
rect 200604 377241 200924 377273
rect 216076 377829 216396 377861
rect 216076 377593 216118 377829
rect 216354 377593 216396 377829
rect 216076 377509 216396 377593
rect 216076 377273 216118 377509
rect 216354 377273 216396 377509
rect 216076 377241 216396 377273
rect 222340 377829 222660 377861
rect 222340 377593 222382 377829
rect 222618 377593 222660 377829
rect 222340 377509 222660 377593
rect 222340 377273 222382 377509
rect 222618 377273 222660 377509
rect 222340 377241 222660 377273
rect 228604 377829 228924 377861
rect 228604 377593 228646 377829
rect 228882 377593 228924 377829
rect 228604 377509 228924 377593
rect 228604 377273 228646 377509
rect 228882 377273 228924 377509
rect 228604 377241 228924 377273
rect 244076 377829 244396 377861
rect 244076 377593 244118 377829
rect 244354 377593 244396 377829
rect 244076 377509 244396 377593
rect 244076 377273 244118 377509
rect 244354 377273 244396 377509
rect 244076 377241 244396 377273
rect 250340 377829 250660 377861
rect 250340 377593 250382 377829
rect 250618 377593 250660 377829
rect 250340 377509 250660 377593
rect 250340 377273 250382 377509
rect 250618 377273 250660 377509
rect 250340 377241 250660 377273
rect 256604 377829 256924 377861
rect 256604 377593 256646 377829
rect 256882 377593 256924 377829
rect 256604 377509 256924 377593
rect 256604 377273 256646 377509
rect 256882 377273 256924 377509
rect 256604 377241 256924 377273
rect 272076 377829 272396 377861
rect 272076 377593 272118 377829
rect 272354 377593 272396 377829
rect 272076 377509 272396 377593
rect 272076 377273 272118 377509
rect 272354 377273 272396 377509
rect 272076 377241 272396 377273
rect 278340 377829 278660 377861
rect 278340 377593 278382 377829
rect 278618 377593 278660 377829
rect 278340 377509 278660 377593
rect 278340 377273 278382 377509
rect 278618 377273 278660 377509
rect 278340 377241 278660 377273
rect 284604 377829 284924 377861
rect 284604 377593 284646 377829
rect 284882 377593 284924 377829
rect 284604 377509 284924 377593
rect 284604 377273 284646 377509
rect 284882 377273 284924 377509
rect 284604 377241 284924 377273
rect 300076 377829 300396 377861
rect 300076 377593 300118 377829
rect 300354 377593 300396 377829
rect 300076 377509 300396 377593
rect 300076 377273 300118 377509
rect 300354 377273 300396 377509
rect 300076 377241 300396 377273
rect 306340 377829 306660 377861
rect 306340 377593 306382 377829
rect 306618 377593 306660 377829
rect 306340 377509 306660 377593
rect 306340 377273 306382 377509
rect 306618 377273 306660 377509
rect 306340 377241 306660 377273
rect 312604 377829 312924 377861
rect 312604 377593 312646 377829
rect 312882 377593 312924 377829
rect 312604 377509 312924 377593
rect 312604 377273 312646 377509
rect 312882 377273 312924 377509
rect 312604 377241 312924 377273
rect 328076 377829 328396 377861
rect 328076 377593 328118 377829
rect 328354 377593 328396 377829
rect 328076 377509 328396 377593
rect 328076 377273 328118 377509
rect 328354 377273 328396 377509
rect 328076 377241 328396 377273
rect 334340 377829 334660 377861
rect 334340 377593 334382 377829
rect 334618 377593 334660 377829
rect 334340 377509 334660 377593
rect 334340 377273 334382 377509
rect 334618 377273 334660 377509
rect 334340 377241 334660 377273
rect 340604 377829 340924 377861
rect 340604 377593 340646 377829
rect 340882 377593 340924 377829
rect 340604 377509 340924 377593
rect 340604 377273 340646 377509
rect 340882 377273 340924 377509
rect 340604 377241 340924 377273
rect 356076 377829 356396 377861
rect 356076 377593 356118 377829
rect 356354 377593 356396 377829
rect 356076 377509 356396 377593
rect 356076 377273 356118 377509
rect 356354 377273 356396 377509
rect 356076 377241 356396 377273
rect 362340 377829 362660 377861
rect 362340 377593 362382 377829
rect 362618 377593 362660 377829
rect 362340 377509 362660 377593
rect 362340 377273 362382 377509
rect 362618 377273 362660 377509
rect 362340 377241 362660 377273
rect 368604 377829 368924 377861
rect 368604 377593 368646 377829
rect 368882 377593 368924 377829
rect 368604 377509 368924 377593
rect 368604 377273 368646 377509
rect 368882 377273 368924 377509
rect 368604 377241 368924 377273
rect 384076 377829 384396 377861
rect 384076 377593 384118 377829
rect 384354 377593 384396 377829
rect 384076 377509 384396 377593
rect 384076 377273 384118 377509
rect 384354 377273 384396 377509
rect 384076 377241 384396 377273
rect 390340 377829 390660 377861
rect 390340 377593 390382 377829
rect 390618 377593 390660 377829
rect 390340 377509 390660 377593
rect 390340 377273 390382 377509
rect 390618 377273 390660 377509
rect 390340 377241 390660 377273
rect 197472 374454 197792 374486
rect 197472 374218 197514 374454
rect 197750 374218 197792 374454
rect 197472 374134 197792 374218
rect 197472 373898 197514 374134
rect 197750 373898 197792 374134
rect 197472 373866 197792 373898
rect 219208 374454 219528 374486
rect 219208 374218 219250 374454
rect 219486 374218 219528 374454
rect 219208 374134 219528 374218
rect 219208 373898 219250 374134
rect 219486 373898 219528 374134
rect 219208 373866 219528 373898
rect 225472 374454 225792 374486
rect 225472 374218 225514 374454
rect 225750 374218 225792 374454
rect 225472 374134 225792 374218
rect 225472 373898 225514 374134
rect 225750 373898 225792 374134
rect 225472 373866 225792 373898
rect 247208 374454 247528 374486
rect 247208 374218 247250 374454
rect 247486 374218 247528 374454
rect 247208 374134 247528 374218
rect 247208 373898 247250 374134
rect 247486 373898 247528 374134
rect 247208 373866 247528 373898
rect 253472 374454 253792 374486
rect 253472 374218 253514 374454
rect 253750 374218 253792 374454
rect 253472 374134 253792 374218
rect 253472 373898 253514 374134
rect 253750 373898 253792 374134
rect 253472 373866 253792 373898
rect 275208 374454 275528 374486
rect 275208 374218 275250 374454
rect 275486 374218 275528 374454
rect 275208 374134 275528 374218
rect 275208 373898 275250 374134
rect 275486 373898 275528 374134
rect 275208 373866 275528 373898
rect 281472 374454 281792 374486
rect 281472 374218 281514 374454
rect 281750 374218 281792 374454
rect 281472 374134 281792 374218
rect 281472 373898 281514 374134
rect 281750 373898 281792 374134
rect 281472 373866 281792 373898
rect 303208 374454 303528 374486
rect 303208 374218 303250 374454
rect 303486 374218 303528 374454
rect 303208 374134 303528 374218
rect 303208 373898 303250 374134
rect 303486 373898 303528 374134
rect 303208 373866 303528 373898
rect 309472 374454 309792 374486
rect 309472 374218 309514 374454
rect 309750 374218 309792 374454
rect 309472 374134 309792 374218
rect 309472 373898 309514 374134
rect 309750 373898 309792 374134
rect 309472 373866 309792 373898
rect 331208 374454 331528 374486
rect 331208 374218 331250 374454
rect 331486 374218 331528 374454
rect 331208 374134 331528 374218
rect 331208 373898 331250 374134
rect 331486 373898 331528 374134
rect 331208 373866 331528 373898
rect 337472 374454 337792 374486
rect 337472 374218 337514 374454
rect 337750 374218 337792 374454
rect 337472 374134 337792 374218
rect 337472 373898 337514 374134
rect 337750 373898 337792 374134
rect 337472 373866 337792 373898
rect 359208 374454 359528 374486
rect 359208 374218 359250 374454
rect 359486 374218 359528 374454
rect 359208 374134 359528 374218
rect 359208 373898 359250 374134
rect 359486 373898 359528 374134
rect 359208 373866 359528 373898
rect 365472 374454 365792 374486
rect 365472 374218 365514 374454
rect 365750 374218 365792 374454
rect 365472 374134 365792 374218
rect 365472 373898 365514 374134
rect 365750 373898 365792 374134
rect 365472 373866 365792 373898
rect 387208 374454 387528 374486
rect 387208 374218 387250 374454
rect 387486 374218 387528 374454
rect 387208 374134 387528 374218
rect 387208 373898 387250 374134
rect 387486 373898 387528 374134
rect 387208 373866 387528 373898
rect 390878 365669 390938 387363
rect 396604 377829 396924 377861
rect 396604 377593 396646 377829
rect 396882 377593 396924 377829
rect 396604 377509 396924 377593
rect 396604 377273 396646 377509
rect 396882 377273 396924 377509
rect 396604 377241 396924 377273
rect 412076 377829 412396 377861
rect 412076 377593 412118 377829
rect 412354 377593 412396 377829
rect 412076 377509 412396 377593
rect 412076 377273 412118 377509
rect 412354 377273 412396 377509
rect 412076 377241 412396 377273
rect 418340 377829 418660 377861
rect 418340 377593 418382 377829
rect 418618 377593 418660 377829
rect 418340 377509 418660 377593
rect 418340 377273 418382 377509
rect 418618 377273 418660 377509
rect 418340 377241 418660 377273
rect 424604 377829 424924 377861
rect 424604 377593 424646 377829
rect 424882 377593 424924 377829
rect 424604 377509 424924 377593
rect 424604 377273 424646 377509
rect 424882 377273 424924 377509
rect 424604 377241 424924 377273
rect 440076 377829 440396 377861
rect 440076 377593 440118 377829
rect 440354 377593 440396 377829
rect 440076 377509 440396 377593
rect 440076 377273 440118 377509
rect 440354 377273 440396 377509
rect 440076 377241 440396 377273
rect 446340 377829 446660 377861
rect 446340 377593 446382 377829
rect 446618 377593 446660 377829
rect 446340 377509 446660 377593
rect 446340 377273 446382 377509
rect 446618 377273 446660 377509
rect 446340 377241 446660 377273
rect 452604 377829 452924 377861
rect 452604 377593 452646 377829
rect 452882 377593 452924 377829
rect 452604 377509 452924 377593
rect 452604 377273 452646 377509
rect 452882 377273 452924 377509
rect 452604 377241 452924 377273
rect 468076 377829 468396 377861
rect 468076 377593 468118 377829
rect 468354 377593 468396 377829
rect 468076 377509 468396 377593
rect 468076 377273 468118 377509
rect 468354 377273 468396 377509
rect 468076 377241 468396 377273
rect 474340 377829 474660 377861
rect 474340 377593 474382 377829
rect 474618 377593 474660 377829
rect 474340 377509 474660 377593
rect 474340 377273 474382 377509
rect 474618 377273 474660 377509
rect 474340 377241 474660 377273
rect 480604 377829 480924 377861
rect 480604 377593 480646 377829
rect 480882 377593 480924 377829
rect 480604 377509 480924 377593
rect 480604 377273 480646 377509
rect 480882 377273 480924 377509
rect 480604 377241 480924 377273
rect 496076 377829 496396 377861
rect 496076 377593 496118 377829
rect 496354 377593 496396 377829
rect 496076 377509 496396 377593
rect 496076 377273 496118 377509
rect 496354 377273 496396 377509
rect 496076 377241 496396 377273
rect 502340 377829 502660 377861
rect 502340 377593 502382 377829
rect 502618 377593 502660 377829
rect 502340 377509 502660 377593
rect 502340 377273 502382 377509
rect 502618 377273 502660 377509
rect 502340 377241 502660 377273
rect 508604 377829 508924 377861
rect 508604 377593 508646 377829
rect 508882 377593 508924 377829
rect 508604 377509 508924 377593
rect 508604 377273 508646 377509
rect 508882 377273 508924 377509
rect 508604 377241 508924 377273
rect 524076 377829 524396 377861
rect 524076 377593 524118 377829
rect 524354 377593 524396 377829
rect 524076 377509 524396 377593
rect 524076 377273 524118 377509
rect 524354 377273 524396 377509
rect 524076 377241 524396 377273
rect 530340 377829 530660 377861
rect 530340 377593 530382 377829
rect 530618 377593 530660 377829
rect 530340 377509 530660 377593
rect 530340 377273 530382 377509
rect 530618 377273 530660 377509
rect 530340 377241 530660 377273
rect 536604 377829 536924 377861
rect 536604 377593 536646 377829
rect 536882 377593 536924 377829
rect 536604 377509 536924 377593
rect 536604 377273 536646 377509
rect 536882 377273 536924 377509
rect 536604 377241 536924 377273
rect 552076 377829 552396 377861
rect 552076 377593 552118 377829
rect 552354 377593 552396 377829
rect 552076 377509 552396 377593
rect 552076 377273 552118 377509
rect 552354 377273 552396 377509
rect 552076 377241 552396 377273
rect 558340 377829 558660 377861
rect 558340 377593 558382 377829
rect 558618 377593 558660 377829
rect 558340 377509 558660 377593
rect 558340 377273 558382 377509
rect 558618 377273 558660 377509
rect 558340 377241 558660 377273
rect 564604 377829 564924 377861
rect 564604 377593 564646 377829
rect 564882 377593 564924 377829
rect 564604 377509 564924 377593
rect 564604 377273 564646 377509
rect 564882 377273 564924 377509
rect 564604 377241 564924 377273
rect 573494 377829 574114 404273
rect 573494 377593 573526 377829
rect 573762 377593 573846 377829
rect 574082 377593 574114 377829
rect 573494 377509 574114 377593
rect 573494 377273 573526 377509
rect 573762 377273 573846 377509
rect 574082 377273 574114 377509
rect 456379 377228 456445 377229
rect 456379 377164 456380 377228
rect 456444 377164 456445 377228
rect 456379 377163 456445 377164
rect 568435 377228 568501 377229
rect 568435 377164 568436 377228
rect 568500 377164 568501 377228
rect 568435 377163 568501 377164
rect 393472 374454 393792 374486
rect 393472 374218 393514 374454
rect 393750 374218 393792 374454
rect 393472 374134 393792 374218
rect 393472 373898 393514 374134
rect 393750 373898 393792 374134
rect 393472 373866 393792 373898
rect 415208 374454 415528 374486
rect 415208 374218 415250 374454
rect 415486 374218 415528 374454
rect 415208 374134 415528 374218
rect 415208 373898 415250 374134
rect 415486 373898 415528 374134
rect 415208 373866 415528 373898
rect 421472 374454 421792 374486
rect 421472 374218 421514 374454
rect 421750 374218 421792 374454
rect 421472 374134 421792 374218
rect 421472 373898 421514 374134
rect 421750 373898 421792 374134
rect 421472 373866 421792 373898
rect 443208 374454 443528 374486
rect 443208 374218 443250 374454
rect 443486 374218 443528 374454
rect 443208 374134 443528 374218
rect 443208 373898 443250 374134
rect 443486 373898 443528 374134
rect 443208 373866 443528 373898
rect 449472 374454 449792 374486
rect 449472 374218 449514 374454
rect 449750 374218 449792 374454
rect 449472 374134 449792 374218
rect 449472 373898 449514 374134
rect 449750 373898 449792 374134
rect 456382 374010 456442 377163
rect 568438 376770 568498 377163
rect 566966 376710 568498 376770
rect 449472 373866 449792 373898
rect 455462 373950 456442 374010
rect 471208 374454 471528 374486
rect 471208 374218 471250 374454
rect 471486 374218 471528 374454
rect 471208 374134 471528 374218
rect 455462 369341 455522 373950
rect 471208 373898 471250 374134
rect 471486 373898 471528 374134
rect 471208 373866 471528 373898
rect 477472 374454 477792 374486
rect 477472 374218 477514 374454
rect 477750 374218 477792 374454
rect 477472 374134 477792 374218
rect 477472 373898 477514 374134
rect 477750 373898 477792 374134
rect 477472 373866 477792 373898
rect 499208 374454 499528 374486
rect 499208 374218 499250 374454
rect 499486 374218 499528 374454
rect 499208 374134 499528 374218
rect 499208 373898 499250 374134
rect 499486 373898 499528 374134
rect 499208 373866 499528 373898
rect 505472 374454 505792 374486
rect 505472 374218 505514 374454
rect 505750 374218 505792 374454
rect 505472 374134 505792 374218
rect 505472 373898 505514 374134
rect 505750 373898 505792 374134
rect 505472 373866 505792 373898
rect 527208 374454 527528 374486
rect 527208 374218 527250 374454
rect 527486 374218 527528 374454
rect 527208 374134 527528 374218
rect 527208 373898 527250 374134
rect 527486 373898 527528 374134
rect 527208 373866 527528 373898
rect 533472 374454 533792 374486
rect 533472 374218 533514 374454
rect 533750 374218 533792 374454
rect 533472 374134 533792 374218
rect 533472 373898 533514 374134
rect 533750 373898 533792 374134
rect 533472 373866 533792 373898
rect 555208 374454 555528 374486
rect 555208 374218 555250 374454
rect 555486 374218 555528 374454
rect 555208 374134 555528 374218
rect 555208 373898 555250 374134
rect 555486 373898 555528 374134
rect 555208 373866 555528 373898
rect 561472 374454 561792 374486
rect 561472 374218 561514 374454
rect 561750 374218 561792 374454
rect 561472 374134 561792 374218
rect 561472 373898 561514 374134
rect 561750 373898 561792 374134
rect 561472 373866 561792 373898
rect 566966 369341 567026 376710
rect 455459 369340 455525 369341
rect 455459 369276 455460 369340
rect 455524 369276 455525 369340
rect 455459 369275 455525 369276
rect 566963 369340 567029 369341
rect 566963 369276 566964 369340
rect 567028 369276 567029 369340
rect 566963 369275 567029 369276
rect 128307 365668 128373 365669
rect 128307 365604 128308 365668
rect 128372 365604 128373 365668
rect 128307 365603 128373 365604
rect 194731 365668 194797 365669
rect 194731 365604 194732 365668
rect 194796 365604 194797 365668
rect 194731 365603 194797 365604
rect 390875 365668 390941 365669
rect 390875 365604 390876 365668
rect 390940 365604 390941 365668
rect 390875 365603 390941 365604
rect 165659 360500 165725 360501
rect 165659 360436 165660 360500
rect 165724 360436 165725 360500
rect 165659 360435 165725 360436
rect 259499 360500 259565 360501
rect 259499 360436 259500 360500
rect 259564 360436 259565 360500
rect 259499 360435 259565 360436
rect 361619 360500 361685 360501
rect 361619 360436 361620 360500
rect 361684 360436 361685 360500
rect 361619 360435 361685 360436
rect 445707 360500 445773 360501
rect 445707 360436 445708 360500
rect 445772 360436 445773 360500
rect 445707 360435 445773 360436
rect 557579 360500 557645 360501
rect 557579 360436 557580 360500
rect 557644 360436 557645 360500
rect 557579 360435 557645 360436
rect -2006 350593 -1974 350829
rect -1738 350593 -1654 350829
rect -1418 350593 -1386 350829
rect -2006 350509 -1386 350593
rect -2006 350273 -1974 350509
rect -1738 350273 -1654 350509
rect -1418 350273 -1386 350509
rect -2006 323829 -1386 350273
rect 20076 350829 20396 350861
rect 20076 350593 20118 350829
rect 20354 350593 20396 350829
rect 20076 350509 20396 350593
rect 20076 350273 20118 350509
rect 20354 350273 20396 350509
rect 20076 350241 20396 350273
rect 26340 350829 26660 350861
rect 26340 350593 26382 350829
rect 26618 350593 26660 350829
rect 26340 350509 26660 350593
rect 26340 350273 26382 350509
rect 26618 350273 26660 350509
rect 26340 350241 26660 350273
rect 32604 350829 32924 350861
rect 32604 350593 32646 350829
rect 32882 350593 32924 350829
rect 32604 350509 32924 350593
rect 32604 350273 32646 350509
rect 32882 350273 32924 350509
rect 32604 350241 32924 350273
rect 48076 350829 48396 350861
rect 48076 350593 48118 350829
rect 48354 350593 48396 350829
rect 48076 350509 48396 350593
rect 48076 350273 48118 350509
rect 48354 350273 48396 350509
rect 48076 350241 48396 350273
rect 54340 350829 54660 350861
rect 54340 350593 54382 350829
rect 54618 350593 54660 350829
rect 54340 350509 54660 350593
rect 54340 350273 54382 350509
rect 54618 350273 54660 350509
rect 54340 350241 54660 350273
rect 60604 350829 60924 350861
rect 60604 350593 60646 350829
rect 60882 350593 60924 350829
rect 60604 350509 60924 350593
rect 60604 350273 60646 350509
rect 60882 350273 60924 350509
rect 60604 350241 60924 350273
rect 76076 350829 76396 350861
rect 76076 350593 76118 350829
rect 76354 350593 76396 350829
rect 76076 350509 76396 350593
rect 76076 350273 76118 350509
rect 76354 350273 76396 350509
rect 76076 350241 76396 350273
rect 82340 350829 82660 350861
rect 82340 350593 82382 350829
rect 82618 350593 82660 350829
rect 82340 350509 82660 350593
rect 82340 350273 82382 350509
rect 82618 350273 82660 350509
rect 82340 350241 82660 350273
rect 88604 350829 88924 350861
rect 88604 350593 88646 350829
rect 88882 350593 88924 350829
rect 88604 350509 88924 350593
rect 88604 350273 88646 350509
rect 88882 350273 88924 350509
rect 88604 350241 88924 350273
rect 104076 350829 104396 350861
rect 104076 350593 104118 350829
rect 104354 350593 104396 350829
rect 104076 350509 104396 350593
rect 104076 350273 104118 350509
rect 104354 350273 104396 350509
rect 104076 350241 104396 350273
rect 110340 350829 110660 350861
rect 110340 350593 110382 350829
rect 110618 350593 110660 350829
rect 110340 350509 110660 350593
rect 110340 350273 110382 350509
rect 110618 350273 110660 350509
rect 110340 350241 110660 350273
rect 116604 350829 116924 350861
rect 116604 350593 116646 350829
rect 116882 350593 116924 350829
rect 116604 350509 116924 350593
rect 116604 350273 116646 350509
rect 116882 350273 116924 350509
rect 116604 350241 116924 350273
rect 132076 350829 132396 350861
rect 132076 350593 132118 350829
rect 132354 350593 132396 350829
rect 132076 350509 132396 350593
rect 132076 350273 132118 350509
rect 132354 350273 132396 350509
rect 132076 350241 132396 350273
rect 138340 350829 138660 350861
rect 138340 350593 138382 350829
rect 138618 350593 138660 350829
rect 138340 350509 138660 350593
rect 138340 350273 138382 350509
rect 138618 350273 138660 350509
rect 138340 350241 138660 350273
rect 144604 350829 144924 350861
rect 144604 350593 144646 350829
rect 144882 350593 144924 350829
rect 144604 350509 144924 350593
rect 144604 350273 144646 350509
rect 144882 350273 144924 350509
rect 144604 350241 144924 350273
rect 160076 350829 160396 350861
rect 160076 350593 160118 350829
rect 160354 350593 160396 350829
rect 160076 350509 160396 350593
rect 160076 350273 160118 350509
rect 160354 350273 160396 350509
rect 160076 350241 160396 350273
rect 44587 349756 44653 349757
rect 44587 349692 44588 349756
rect 44652 349692 44653 349756
rect 44587 349691 44653 349692
rect 128491 349756 128557 349757
rect 128491 349692 128492 349756
rect 128556 349692 128557 349756
rect 128491 349691 128557 349692
rect 23208 347454 23528 347486
rect 23208 347218 23250 347454
rect 23486 347218 23528 347454
rect 23208 347134 23528 347218
rect 23208 346898 23250 347134
rect 23486 346898 23528 347134
rect 23208 346866 23528 346898
rect 29472 347454 29792 347486
rect 29472 347218 29514 347454
rect 29750 347218 29792 347454
rect 29472 347134 29792 347218
rect 29472 346898 29514 347134
rect 29750 346898 29792 347134
rect 29472 346866 29792 346898
rect 44590 341733 44650 349691
rect 51208 347454 51528 347486
rect 51208 347218 51250 347454
rect 51486 347218 51528 347454
rect 51208 347134 51528 347218
rect 51208 346898 51250 347134
rect 51486 346898 51528 347134
rect 51208 346866 51528 346898
rect 57472 347454 57792 347486
rect 57472 347218 57514 347454
rect 57750 347218 57792 347454
rect 57472 347134 57792 347218
rect 57472 346898 57514 347134
rect 57750 346898 57792 347134
rect 57472 346866 57792 346898
rect 79208 347454 79528 347486
rect 79208 347218 79250 347454
rect 79486 347218 79528 347454
rect 79208 347134 79528 347218
rect 79208 346898 79250 347134
rect 79486 346898 79528 347134
rect 79208 346866 79528 346898
rect 85472 347454 85792 347486
rect 85472 347218 85514 347454
rect 85750 347218 85792 347454
rect 85472 347134 85792 347218
rect 85472 346898 85514 347134
rect 85750 346898 85792 347134
rect 85472 346866 85792 346898
rect 107208 347454 107528 347486
rect 107208 347218 107250 347454
rect 107486 347218 107528 347454
rect 107208 347134 107528 347218
rect 107208 346898 107250 347134
rect 107486 346898 107528 347134
rect 107208 346866 107528 346898
rect 113472 347454 113792 347486
rect 113472 347218 113514 347454
rect 113750 347218 113792 347454
rect 113472 347134 113792 347218
rect 113472 346898 113514 347134
rect 113750 346898 113792 347134
rect 113472 346866 113792 346898
rect 128494 341733 128554 349691
rect 135208 347454 135528 347486
rect 135208 347218 135250 347454
rect 135486 347218 135528 347454
rect 135208 347134 135528 347218
rect 135208 346898 135250 347134
rect 135486 346898 135528 347134
rect 135208 346866 135528 346898
rect 141472 347454 141792 347486
rect 141472 347218 141514 347454
rect 141750 347218 141792 347454
rect 141472 347134 141792 347218
rect 141472 346898 141514 347134
rect 141750 346898 141792 347134
rect 141472 346866 141792 346898
rect 163208 347454 163528 347486
rect 163208 347218 163250 347454
rect 163486 347218 163528 347454
rect 163208 347134 163528 347218
rect 163208 346898 163250 347134
rect 163486 346898 163528 347134
rect 163208 346866 163528 346898
rect 44587 341732 44653 341733
rect 44587 341668 44588 341732
rect 44652 341668 44653 341732
rect 44587 341667 44653 341668
rect 128491 341732 128557 341733
rect 128491 341668 128492 341732
rect 128556 341668 128557 341732
rect 128491 341667 128557 341668
rect 165662 338061 165722 360435
rect 166340 350829 166660 350861
rect 166340 350593 166382 350829
rect 166618 350593 166660 350829
rect 166340 350509 166660 350593
rect 166340 350273 166382 350509
rect 166618 350273 166660 350509
rect 166340 350241 166660 350273
rect 172604 350829 172924 350861
rect 172604 350593 172646 350829
rect 172882 350593 172924 350829
rect 172604 350509 172924 350593
rect 172604 350273 172646 350509
rect 172882 350273 172924 350509
rect 172604 350241 172924 350273
rect 188076 350829 188396 350861
rect 188076 350593 188118 350829
rect 188354 350593 188396 350829
rect 188076 350509 188396 350593
rect 188076 350273 188118 350509
rect 188354 350273 188396 350509
rect 188076 350241 188396 350273
rect 194340 350829 194660 350861
rect 194340 350593 194382 350829
rect 194618 350593 194660 350829
rect 194340 350509 194660 350593
rect 194340 350273 194382 350509
rect 194618 350273 194660 350509
rect 194340 350241 194660 350273
rect 200604 350829 200924 350861
rect 200604 350593 200646 350829
rect 200882 350593 200924 350829
rect 200604 350509 200924 350593
rect 200604 350273 200646 350509
rect 200882 350273 200924 350509
rect 200604 350241 200924 350273
rect 216076 350829 216396 350861
rect 216076 350593 216118 350829
rect 216354 350593 216396 350829
rect 216076 350509 216396 350593
rect 216076 350273 216118 350509
rect 216354 350273 216396 350509
rect 216076 350241 216396 350273
rect 222340 350829 222660 350861
rect 222340 350593 222382 350829
rect 222618 350593 222660 350829
rect 222340 350509 222660 350593
rect 222340 350273 222382 350509
rect 222618 350273 222660 350509
rect 222340 350241 222660 350273
rect 228604 350829 228924 350861
rect 228604 350593 228646 350829
rect 228882 350593 228924 350829
rect 228604 350509 228924 350593
rect 228604 350273 228646 350509
rect 228882 350273 228924 350509
rect 228604 350241 228924 350273
rect 244076 350829 244396 350861
rect 244076 350593 244118 350829
rect 244354 350593 244396 350829
rect 244076 350509 244396 350593
rect 244076 350273 244118 350509
rect 244354 350273 244396 350509
rect 244076 350241 244396 350273
rect 250340 350829 250660 350861
rect 250340 350593 250382 350829
rect 250618 350593 250660 350829
rect 250340 350509 250660 350593
rect 250340 350273 250382 350509
rect 250618 350273 250660 350509
rect 250340 350241 250660 350273
rect 256604 350829 256924 350861
rect 256604 350593 256646 350829
rect 256882 350593 256924 350829
rect 256604 350509 256924 350593
rect 256604 350273 256646 350509
rect 256882 350273 256924 350509
rect 256604 350241 256924 350273
rect 212579 349756 212645 349757
rect 212579 349692 212580 349756
rect 212644 349692 212645 349756
rect 212579 349691 212645 349692
rect 240547 349756 240613 349757
rect 240547 349692 240548 349756
rect 240612 349692 240613 349756
rect 240547 349691 240613 349692
rect 169472 347454 169792 347486
rect 169472 347218 169514 347454
rect 169750 347218 169792 347454
rect 169472 347134 169792 347218
rect 169472 346898 169514 347134
rect 169750 346898 169792 347134
rect 169472 346866 169792 346898
rect 191208 347454 191528 347486
rect 191208 347218 191250 347454
rect 191486 347218 191528 347454
rect 191208 347134 191528 347218
rect 191208 346898 191250 347134
rect 191486 346898 191528 347134
rect 191208 346866 191528 346898
rect 197472 347454 197792 347486
rect 197472 347218 197514 347454
rect 197750 347218 197792 347454
rect 197472 347134 197792 347218
rect 197472 346898 197514 347134
rect 197750 346898 197792 347134
rect 197472 346866 197792 346898
rect 212582 341733 212642 349691
rect 219208 347454 219528 347486
rect 219208 347218 219250 347454
rect 219486 347218 219528 347454
rect 219208 347134 219528 347218
rect 219208 346898 219250 347134
rect 219486 346898 219528 347134
rect 219208 346866 219528 346898
rect 225472 347454 225792 347486
rect 225472 347218 225514 347454
rect 225750 347218 225792 347454
rect 225472 347134 225792 347218
rect 225472 346898 225514 347134
rect 225750 346898 225792 347134
rect 225472 346866 225792 346898
rect 240550 341869 240610 349691
rect 247208 347454 247528 347486
rect 247208 347218 247250 347454
rect 247486 347218 247528 347454
rect 247208 347134 247528 347218
rect 247208 346898 247250 347134
rect 247486 346898 247528 347134
rect 247208 346866 247528 346898
rect 253472 347454 253792 347486
rect 253472 347218 253514 347454
rect 253750 347218 253792 347454
rect 253472 347134 253792 347218
rect 253472 346898 253514 347134
rect 253750 346898 253792 347134
rect 253472 346866 253792 346898
rect 240547 341868 240613 341869
rect 240547 341804 240548 341868
rect 240612 341804 240613 341868
rect 240547 341803 240613 341804
rect 212579 341732 212645 341733
rect 212579 341668 212580 341732
rect 212644 341668 212645 341732
rect 212579 341667 212645 341668
rect 259502 338061 259562 360435
rect 272076 350829 272396 350861
rect 272076 350593 272118 350829
rect 272354 350593 272396 350829
rect 272076 350509 272396 350593
rect 272076 350273 272118 350509
rect 272354 350273 272396 350509
rect 272076 350241 272396 350273
rect 278340 350829 278660 350861
rect 278340 350593 278382 350829
rect 278618 350593 278660 350829
rect 278340 350509 278660 350593
rect 278340 350273 278382 350509
rect 278618 350273 278660 350509
rect 278340 350241 278660 350273
rect 284604 350829 284924 350861
rect 284604 350593 284646 350829
rect 284882 350593 284924 350829
rect 284604 350509 284924 350593
rect 284604 350273 284646 350509
rect 284882 350273 284924 350509
rect 284604 350241 284924 350273
rect 300076 350829 300396 350861
rect 300076 350593 300118 350829
rect 300354 350593 300396 350829
rect 300076 350509 300396 350593
rect 300076 350273 300118 350509
rect 300354 350273 300396 350509
rect 300076 350241 300396 350273
rect 306340 350829 306660 350861
rect 306340 350593 306382 350829
rect 306618 350593 306660 350829
rect 306340 350509 306660 350593
rect 306340 350273 306382 350509
rect 306618 350273 306660 350509
rect 306340 350241 306660 350273
rect 312604 350829 312924 350861
rect 312604 350593 312646 350829
rect 312882 350593 312924 350829
rect 312604 350509 312924 350593
rect 312604 350273 312646 350509
rect 312882 350273 312924 350509
rect 312604 350241 312924 350273
rect 328076 350829 328396 350861
rect 328076 350593 328118 350829
rect 328354 350593 328396 350829
rect 328076 350509 328396 350593
rect 328076 350273 328118 350509
rect 328354 350273 328396 350509
rect 328076 350241 328396 350273
rect 334340 350829 334660 350861
rect 334340 350593 334382 350829
rect 334618 350593 334660 350829
rect 334340 350509 334660 350593
rect 334340 350273 334382 350509
rect 334618 350273 334660 350509
rect 334340 350241 334660 350273
rect 340604 350829 340924 350861
rect 340604 350593 340646 350829
rect 340882 350593 340924 350829
rect 340604 350509 340924 350593
rect 340604 350273 340646 350509
rect 340882 350273 340924 350509
rect 340604 350241 340924 350273
rect 356076 350829 356396 350861
rect 356076 350593 356118 350829
rect 356354 350593 356396 350829
rect 356076 350509 356396 350593
rect 356076 350273 356118 350509
rect 356354 350273 356396 350509
rect 356076 350241 356396 350273
rect 296483 349756 296549 349757
rect 296483 349692 296484 349756
rect 296548 349692 296549 349756
rect 296483 349691 296549 349692
rect 324635 349756 324701 349757
rect 324635 349692 324636 349756
rect 324700 349692 324701 349756
rect 324635 349691 324701 349692
rect 296486 347790 296546 349691
rect 296486 347730 296914 347790
rect 275208 347454 275528 347486
rect 275208 347218 275250 347454
rect 275486 347218 275528 347454
rect 275208 347134 275528 347218
rect 275208 346898 275250 347134
rect 275486 346898 275528 347134
rect 275208 346866 275528 346898
rect 281472 347454 281792 347486
rect 281472 347218 281514 347454
rect 281750 347218 281792 347454
rect 281472 347134 281792 347218
rect 281472 346898 281514 347134
rect 281750 346898 281792 347134
rect 281472 346866 281792 346898
rect 296854 341733 296914 347730
rect 303208 347454 303528 347486
rect 303208 347218 303250 347454
rect 303486 347218 303528 347454
rect 303208 347134 303528 347218
rect 303208 346898 303250 347134
rect 303486 346898 303528 347134
rect 303208 346866 303528 346898
rect 309472 347454 309792 347486
rect 309472 347218 309514 347454
rect 309750 347218 309792 347454
rect 309472 347134 309792 347218
rect 309472 346898 309514 347134
rect 309750 346898 309792 347134
rect 309472 346866 309792 346898
rect 324638 341869 324698 349691
rect 331208 347454 331528 347486
rect 331208 347218 331250 347454
rect 331486 347218 331528 347454
rect 331208 347134 331528 347218
rect 331208 346898 331250 347134
rect 331486 346898 331528 347134
rect 331208 346866 331528 346898
rect 337472 347454 337792 347486
rect 337472 347218 337514 347454
rect 337750 347218 337792 347454
rect 337472 347134 337792 347218
rect 337472 346898 337514 347134
rect 337750 346898 337792 347134
rect 337472 346866 337792 346898
rect 359208 347454 359528 347486
rect 359208 347218 359250 347454
rect 359486 347218 359528 347454
rect 359208 347134 359528 347218
rect 359208 346898 359250 347134
rect 359486 346898 359528 347134
rect 359208 346866 359528 346898
rect 324635 341868 324701 341869
rect 324635 341804 324636 341868
rect 324700 341804 324701 341868
rect 324635 341803 324701 341804
rect 296851 341732 296917 341733
rect 296851 341668 296852 341732
rect 296916 341668 296917 341732
rect 296851 341667 296917 341668
rect 361622 338061 361682 360435
rect 362340 350829 362660 350861
rect 362340 350593 362382 350829
rect 362618 350593 362660 350829
rect 362340 350509 362660 350593
rect 362340 350273 362382 350509
rect 362618 350273 362660 350509
rect 362340 350241 362660 350273
rect 368604 350829 368924 350861
rect 368604 350593 368646 350829
rect 368882 350593 368924 350829
rect 368604 350509 368924 350593
rect 368604 350273 368646 350509
rect 368882 350273 368924 350509
rect 368604 350241 368924 350273
rect 384076 350829 384396 350861
rect 384076 350593 384118 350829
rect 384354 350593 384396 350829
rect 384076 350509 384396 350593
rect 384076 350273 384118 350509
rect 384354 350273 384396 350509
rect 384076 350241 384396 350273
rect 390340 350829 390660 350861
rect 390340 350593 390382 350829
rect 390618 350593 390660 350829
rect 390340 350509 390660 350593
rect 390340 350273 390382 350509
rect 390618 350273 390660 350509
rect 390340 350241 390660 350273
rect 396604 350829 396924 350861
rect 396604 350593 396646 350829
rect 396882 350593 396924 350829
rect 396604 350509 396924 350593
rect 396604 350273 396646 350509
rect 396882 350273 396924 350509
rect 396604 350241 396924 350273
rect 412076 350829 412396 350861
rect 412076 350593 412118 350829
rect 412354 350593 412396 350829
rect 412076 350509 412396 350593
rect 412076 350273 412118 350509
rect 412354 350273 412396 350509
rect 412076 350241 412396 350273
rect 418340 350829 418660 350861
rect 418340 350593 418382 350829
rect 418618 350593 418660 350829
rect 418340 350509 418660 350593
rect 418340 350273 418382 350509
rect 418618 350273 418660 350509
rect 418340 350241 418660 350273
rect 424604 350829 424924 350861
rect 424604 350593 424646 350829
rect 424882 350593 424924 350829
rect 424604 350509 424924 350593
rect 424604 350273 424646 350509
rect 424882 350273 424924 350509
rect 424604 350241 424924 350273
rect 440076 350829 440396 350861
rect 440076 350593 440118 350829
rect 440354 350593 440396 350829
rect 440076 350509 440396 350593
rect 440076 350273 440118 350509
rect 440354 350273 440396 350509
rect 440076 350241 440396 350273
rect 408539 349756 408605 349757
rect 408539 349692 408540 349756
rect 408604 349692 408605 349756
rect 408539 349691 408605 349692
rect 436507 349756 436573 349757
rect 436507 349692 436508 349756
rect 436572 349692 436573 349756
rect 436507 349691 436573 349692
rect 365472 347454 365792 347486
rect 365472 347218 365514 347454
rect 365750 347218 365792 347454
rect 365472 347134 365792 347218
rect 365472 346898 365514 347134
rect 365750 346898 365792 347134
rect 365472 346866 365792 346898
rect 387208 347454 387528 347486
rect 387208 347218 387250 347454
rect 387486 347218 387528 347454
rect 387208 347134 387528 347218
rect 387208 346898 387250 347134
rect 387486 346898 387528 347134
rect 387208 346866 387528 346898
rect 393472 347454 393792 347486
rect 393472 347218 393514 347454
rect 393750 347218 393792 347454
rect 393472 347134 393792 347218
rect 393472 346898 393514 347134
rect 393750 346898 393792 347134
rect 393472 346866 393792 346898
rect 408542 342005 408602 349691
rect 415208 347454 415528 347486
rect 415208 347218 415250 347454
rect 415486 347218 415528 347454
rect 415208 347134 415528 347218
rect 415208 346898 415250 347134
rect 415486 346898 415528 347134
rect 415208 346866 415528 346898
rect 421472 347454 421792 347486
rect 421472 347218 421514 347454
rect 421750 347218 421792 347454
rect 421472 347134 421792 347218
rect 421472 346898 421514 347134
rect 421750 346898 421792 347134
rect 421472 346866 421792 346898
rect 408539 342004 408605 342005
rect 408539 341940 408540 342004
rect 408604 341940 408605 342004
rect 408539 341939 408605 341940
rect 436510 341869 436570 349691
rect 443208 347454 443528 347486
rect 443208 347218 443250 347454
rect 443486 347218 443528 347454
rect 443208 347134 443528 347218
rect 443208 346898 443250 347134
rect 443486 346898 443528 347134
rect 443208 346866 443528 346898
rect 436507 341868 436573 341869
rect 436507 341804 436508 341868
rect 436572 341804 436573 341868
rect 436507 341803 436573 341804
rect 445710 338061 445770 360435
rect 446340 350829 446660 350861
rect 446340 350593 446382 350829
rect 446618 350593 446660 350829
rect 446340 350509 446660 350593
rect 446340 350273 446382 350509
rect 446618 350273 446660 350509
rect 446340 350241 446660 350273
rect 452604 350829 452924 350861
rect 452604 350593 452646 350829
rect 452882 350593 452924 350829
rect 452604 350509 452924 350593
rect 452604 350273 452646 350509
rect 452882 350273 452924 350509
rect 452604 350241 452924 350273
rect 468076 350829 468396 350861
rect 468076 350593 468118 350829
rect 468354 350593 468396 350829
rect 468076 350509 468396 350593
rect 468076 350273 468118 350509
rect 468354 350273 468396 350509
rect 468076 350241 468396 350273
rect 474340 350829 474660 350861
rect 474340 350593 474382 350829
rect 474618 350593 474660 350829
rect 474340 350509 474660 350593
rect 474340 350273 474382 350509
rect 474618 350273 474660 350509
rect 474340 350241 474660 350273
rect 480604 350829 480924 350861
rect 480604 350593 480646 350829
rect 480882 350593 480924 350829
rect 480604 350509 480924 350593
rect 480604 350273 480646 350509
rect 480882 350273 480924 350509
rect 480604 350241 480924 350273
rect 496076 350829 496396 350861
rect 496076 350593 496118 350829
rect 496354 350593 496396 350829
rect 496076 350509 496396 350593
rect 496076 350273 496118 350509
rect 496354 350273 496396 350509
rect 496076 350241 496396 350273
rect 502340 350829 502660 350861
rect 502340 350593 502382 350829
rect 502618 350593 502660 350829
rect 502340 350509 502660 350593
rect 502340 350273 502382 350509
rect 502618 350273 502660 350509
rect 502340 350241 502660 350273
rect 508604 350829 508924 350861
rect 508604 350593 508646 350829
rect 508882 350593 508924 350829
rect 508604 350509 508924 350593
rect 508604 350273 508646 350509
rect 508882 350273 508924 350509
rect 508604 350241 508924 350273
rect 524076 350829 524396 350861
rect 524076 350593 524118 350829
rect 524354 350593 524396 350829
rect 524076 350509 524396 350593
rect 524076 350273 524118 350509
rect 524354 350273 524396 350509
rect 524076 350241 524396 350273
rect 530340 350829 530660 350861
rect 530340 350593 530382 350829
rect 530618 350593 530660 350829
rect 530340 350509 530660 350593
rect 530340 350273 530382 350509
rect 530618 350273 530660 350509
rect 530340 350241 530660 350273
rect 536604 350829 536924 350861
rect 536604 350593 536646 350829
rect 536882 350593 536924 350829
rect 536604 350509 536924 350593
rect 536604 350273 536646 350509
rect 536882 350273 536924 350509
rect 536604 350241 536924 350273
rect 552076 350829 552396 350861
rect 552076 350593 552118 350829
rect 552354 350593 552396 350829
rect 552076 350509 552396 350593
rect 552076 350273 552118 350509
rect 552354 350273 552396 350509
rect 552076 350241 552396 350273
rect 492627 349756 492693 349757
rect 492627 349692 492628 349756
rect 492692 349692 492693 349756
rect 492627 349691 492693 349692
rect 520595 349756 520661 349757
rect 520595 349692 520596 349756
rect 520660 349692 520661 349756
rect 520595 349691 520661 349692
rect 449472 347454 449792 347486
rect 449472 347218 449514 347454
rect 449750 347218 449792 347454
rect 449472 347134 449792 347218
rect 449472 346898 449514 347134
rect 449750 346898 449792 347134
rect 449472 346866 449792 346898
rect 471208 347454 471528 347486
rect 471208 347218 471250 347454
rect 471486 347218 471528 347454
rect 471208 347134 471528 347218
rect 471208 346898 471250 347134
rect 471486 346898 471528 347134
rect 471208 346866 471528 346898
rect 477472 347454 477792 347486
rect 477472 347218 477514 347454
rect 477750 347218 477792 347454
rect 477472 347134 477792 347218
rect 477472 346898 477514 347134
rect 477750 346898 477792 347134
rect 477472 346866 477792 346898
rect 492630 341869 492690 349691
rect 499208 347454 499528 347486
rect 499208 347218 499250 347454
rect 499486 347218 499528 347454
rect 499208 347134 499528 347218
rect 499208 346898 499250 347134
rect 499486 346898 499528 347134
rect 499208 346866 499528 346898
rect 505472 347454 505792 347486
rect 505472 347218 505514 347454
rect 505750 347218 505792 347454
rect 505472 347134 505792 347218
rect 505472 346898 505514 347134
rect 505750 346898 505792 347134
rect 505472 346866 505792 346898
rect 520598 342005 520658 349691
rect 527208 347454 527528 347486
rect 527208 347218 527250 347454
rect 527486 347218 527528 347454
rect 527208 347134 527528 347218
rect 527208 346898 527250 347134
rect 527486 346898 527528 347134
rect 527208 346866 527528 346898
rect 533472 347454 533792 347486
rect 533472 347218 533514 347454
rect 533750 347218 533792 347454
rect 533472 347134 533792 347218
rect 533472 346898 533514 347134
rect 533750 346898 533792 347134
rect 533472 346866 533792 346898
rect 555208 347454 555528 347486
rect 555208 347218 555250 347454
rect 555486 347218 555528 347454
rect 555208 347134 555528 347218
rect 555208 346898 555250 347134
rect 555486 346898 555528 347134
rect 555208 346866 555528 346898
rect 520595 342004 520661 342005
rect 520595 341940 520596 342004
rect 520660 341940 520661 342004
rect 520595 341939 520661 341940
rect 492627 341868 492693 341869
rect 492627 341804 492628 341868
rect 492692 341804 492693 341868
rect 492627 341803 492693 341804
rect 557582 338061 557642 360435
rect 558340 350829 558660 350861
rect 558340 350593 558382 350829
rect 558618 350593 558660 350829
rect 558340 350509 558660 350593
rect 558340 350273 558382 350509
rect 558618 350273 558660 350509
rect 558340 350241 558660 350273
rect 564604 350829 564924 350861
rect 564604 350593 564646 350829
rect 564882 350593 564924 350829
rect 564604 350509 564924 350593
rect 564604 350273 564646 350509
rect 564882 350273 564924 350509
rect 564604 350241 564924 350273
rect 573494 350829 574114 377273
rect 573494 350593 573526 350829
rect 573762 350593 573846 350829
rect 574082 350593 574114 350829
rect 573494 350509 574114 350593
rect 573494 350273 573526 350509
rect 573762 350273 573846 350509
rect 574082 350273 574114 350509
rect 561472 347454 561792 347486
rect 561472 347218 561514 347454
rect 561750 347218 561792 347454
rect 561472 347134 561792 347218
rect 561472 346898 561514 347134
rect 561750 346898 561792 347134
rect 561472 346866 561792 346898
rect 165659 338060 165725 338061
rect 165659 337996 165660 338060
rect 165724 337996 165725 338060
rect 165659 337995 165725 337996
rect 259499 338060 259565 338061
rect 259499 337996 259500 338060
rect 259564 337996 259565 338060
rect 259499 337995 259565 337996
rect 361619 338060 361685 338061
rect 361619 337996 361620 338060
rect 361684 337996 361685 338060
rect 361619 337995 361685 337996
rect 445707 338060 445773 338061
rect 445707 337996 445708 338060
rect 445772 337996 445773 338060
rect 445707 337995 445773 337996
rect 557579 338060 557645 338061
rect 557579 337996 557580 338060
rect 557644 337996 557645 338060
rect 557579 337995 557645 337996
rect 128307 333300 128373 333301
rect 128307 333236 128308 333300
rect 128372 333236 128373 333300
rect 128307 333235 128373 333236
rect 194731 333300 194797 333301
rect 194731 333236 194732 333300
rect 194796 333236 194797 333300
rect 194731 333235 194797 333236
rect 390875 333300 390941 333301
rect 390875 333236 390876 333300
rect 390940 333236 390941 333300
rect 390875 333235 390941 333236
rect -2006 323593 -1974 323829
rect -1738 323593 -1654 323829
rect -1418 323593 -1386 323829
rect -2006 323509 -1386 323593
rect -2006 323273 -1974 323509
rect -1738 323273 -1654 323509
rect -1418 323273 -1386 323509
rect -2006 296829 -1386 323273
rect 20076 323829 20396 323861
rect 20076 323593 20118 323829
rect 20354 323593 20396 323829
rect 20076 323509 20396 323593
rect 20076 323273 20118 323509
rect 20354 323273 20396 323509
rect 20076 323241 20396 323273
rect 26340 323829 26660 323861
rect 26340 323593 26382 323829
rect 26618 323593 26660 323829
rect 26340 323509 26660 323593
rect 26340 323273 26382 323509
rect 26618 323273 26660 323509
rect 26340 323241 26660 323273
rect 32604 323829 32924 323861
rect 32604 323593 32646 323829
rect 32882 323593 32924 323829
rect 32604 323509 32924 323593
rect 32604 323273 32646 323509
rect 32882 323273 32924 323509
rect 32604 323241 32924 323273
rect 48076 323829 48396 323861
rect 48076 323593 48118 323829
rect 48354 323593 48396 323829
rect 48076 323509 48396 323593
rect 48076 323273 48118 323509
rect 48354 323273 48396 323509
rect 48076 323241 48396 323273
rect 54340 323829 54660 323861
rect 54340 323593 54382 323829
rect 54618 323593 54660 323829
rect 54340 323509 54660 323593
rect 54340 323273 54382 323509
rect 54618 323273 54660 323509
rect 54340 323241 54660 323273
rect 60604 323829 60924 323861
rect 60604 323593 60646 323829
rect 60882 323593 60924 323829
rect 60604 323509 60924 323593
rect 60604 323273 60646 323509
rect 60882 323273 60924 323509
rect 60604 323241 60924 323273
rect 76076 323829 76396 323861
rect 76076 323593 76118 323829
rect 76354 323593 76396 323829
rect 76076 323509 76396 323593
rect 76076 323273 76118 323509
rect 76354 323273 76396 323509
rect 76076 323241 76396 323273
rect 82340 323829 82660 323861
rect 82340 323593 82382 323829
rect 82618 323593 82660 323829
rect 82340 323509 82660 323593
rect 82340 323273 82382 323509
rect 82618 323273 82660 323509
rect 82340 323241 82660 323273
rect 88604 323829 88924 323861
rect 88604 323593 88646 323829
rect 88882 323593 88924 323829
rect 88604 323509 88924 323593
rect 88604 323273 88646 323509
rect 88882 323273 88924 323509
rect 88604 323241 88924 323273
rect 104076 323829 104396 323861
rect 104076 323593 104118 323829
rect 104354 323593 104396 323829
rect 104076 323509 104396 323593
rect 104076 323273 104118 323509
rect 104354 323273 104396 323509
rect 104076 323241 104396 323273
rect 110340 323829 110660 323861
rect 110340 323593 110382 323829
rect 110618 323593 110660 323829
rect 110340 323509 110660 323593
rect 110340 323273 110382 323509
rect 110618 323273 110660 323509
rect 110340 323241 110660 323273
rect 116604 323829 116924 323861
rect 116604 323593 116646 323829
rect 116882 323593 116924 323829
rect 116604 323509 116924 323593
rect 116604 323273 116646 323509
rect 116882 323273 116924 323509
rect 116604 323241 116924 323273
rect 23208 320454 23528 320486
rect 23208 320218 23250 320454
rect 23486 320218 23528 320454
rect 23208 320134 23528 320218
rect 23208 319898 23250 320134
rect 23486 319898 23528 320134
rect 23208 319866 23528 319898
rect 29472 320454 29792 320486
rect 29472 320218 29514 320454
rect 29750 320218 29792 320454
rect 29472 320134 29792 320218
rect 29472 319898 29514 320134
rect 29750 319898 29792 320134
rect 29472 319866 29792 319898
rect 51208 320454 51528 320486
rect 51208 320218 51250 320454
rect 51486 320218 51528 320454
rect 51208 320134 51528 320218
rect 51208 319898 51250 320134
rect 51486 319898 51528 320134
rect 51208 319866 51528 319898
rect 57472 320454 57792 320486
rect 57472 320218 57514 320454
rect 57750 320218 57792 320454
rect 57472 320134 57792 320218
rect 57472 319898 57514 320134
rect 57750 319898 57792 320134
rect 57472 319866 57792 319898
rect 79208 320454 79528 320486
rect 79208 320218 79250 320454
rect 79486 320218 79528 320454
rect 79208 320134 79528 320218
rect 79208 319898 79250 320134
rect 79486 319898 79528 320134
rect 79208 319866 79528 319898
rect 85472 320454 85792 320486
rect 85472 320218 85514 320454
rect 85750 320218 85792 320454
rect 85472 320134 85792 320218
rect 85472 319898 85514 320134
rect 85750 319898 85792 320134
rect 85472 319866 85792 319898
rect 107208 320454 107528 320486
rect 107208 320218 107250 320454
rect 107486 320218 107528 320454
rect 107208 320134 107528 320218
rect 107208 319898 107250 320134
rect 107486 319898 107528 320134
rect 107208 319866 107528 319898
rect 113472 320454 113792 320486
rect 113472 320218 113514 320454
rect 113750 320218 113792 320454
rect 113472 320134 113792 320218
rect 113472 319898 113514 320134
rect 113750 319898 113792 320134
rect 113472 319866 113792 319898
rect 128310 311813 128370 333235
rect 132076 323829 132396 323861
rect 132076 323593 132118 323829
rect 132354 323593 132396 323829
rect 132076 323509 132396 323593
rect 132076 323273 132118 323509
rect 132354 323273 132396 323509
rect 132076 323241 132396 323273
rect 138340 323829 138660 323861
rect 138340 323593 138382 323829
rect 138618 323593 138660 323829
rect 138340 323509 138660 323593
rect 138340 323273 138382 323509
rect 138618 323273 138660 323509
rect 138340 323241 138660 323273
rect 144604 323829 144924 323861
rect 144604 323593 144646 323829
rect 144882 323593 144924 323829
rect 144604 323509 144924 323593
rect 144604 323273 144646 323509
rect 144882 323273 144924 323509
rect 144604 323241 144924 323273
rect 160076 323829 160396 323861
rect 160076 323593 160118 323829
rect 160354 323593 160396 323829
rect 160076 323509 160396 323593
rect 160076 323273 160118 323509
rect 160354 323273 160396 323509
rect 160076 323241 160396 323273
rect 166340 323829 166660 323861
rect 166340 323593 166382 323829
rect 166618 323593 166660 323829
rect 166340 323509 166660 323593
rect 166340 323273 166382 323509
rect 166618 323273 166660 323509
rect 166340 323241 166660 323273
rect 172604 323829 172924 323861
rect 172604 323593 172646 323829
rect 172882 323593 172924 323829
rect 172604 323509 172924 323593
rect 172604 323273 172646 323509
rect 172882 323273 172924 323509
rect 172604 323241 172924 323273
rect 188076 323829 188396 323861
rect 188076 323593 188118 323829
rect 188354 323593 188396 323829
rect 188076 323509 188396 323593
rect 188076 323273 188118 323509
rect 188354 323273 188396 323509
rect 188076 323241 188396 323273
rect 194340 323829 194660 323861
rect 194340 323593 194382 323829
rect 194618 323593 194660 323829
rect 194340 323509 194660 323593
rect 194340 323273 194382 323509
rect 194618 323273 194660 323509
rect 194340 323241 194660 323273
rect 176331 323236 176397 323237
rect 176331 323172 176332 323236
rect 176396 323172 176397 323236
rect 176331 323171 176397 323172
rect 135208 320454 135528 320486
rect 135208 320218 135250 320454
rect 135486 320218 135528 320454
rect 135208 320134 135528 320218
rect 135208 319898 135250 320134
rect 135486 319898 135528 320134
rect 135208 319866 135528 319898
rect 141472 320454 141792 320486
rect 141472 320218 141514 320454
rect 141750 320218 141792 320454
rect 141472 320134 141792 320218
rect 141472 319898 141514 320134
rect 141750 319898 141792 320134
rect 141472 319866 141792 319898
rect 163208 320454 163528 320486
rect 163208 320218 163250 320454
rect 163486 320218 163528 320454
rect 163208 320134 163528 320218
rect 163208 319898 163250 320134
rect 163486 319898 163528 320134
rect 163208 319866 163528 319898
rect 169472 320454 169792 320486
rect 169472 320218 169514 320454
rect 169750 320218 169792 320454
rect 169472 320134 169792 320218
rect 169472 319898 169514 320134
rect 169750 319898 169792 320134
rect 169472 319866 169792 319898
rect 176334 316050 176394 323171
rect 191208 320454 191528 320486
rect 191208 320218 191250 320454
rect 191486 320218 191528 320454
rect 191208 320134 191528 320218
rect 191208 319898 191250 320134
rect 191486 319898 191528 320134
rect 191208 319866 191528 319898
rect 175230 315990 176394 316050
rect 175230 315349 175290 315990
rect 175227 315348 175293 315349
rect 175227 315284 175228 315348
rect 175292 315284 175293 315348
rect 175227 315283 175293 315284
rect 194734 311813 194794 333235
rect 200604 323829 200924 323861
rect 200604 323593 200646 323829
rect 200882 323593 200924 323829
rect 200604 323509 200924 323593
rect 200604 323273 200646 323509
rect 200882 323273 200924 323509
rect 200604 323241 200924 323273
rect 216076 323829 216396 323861
rect 216076 323593 216118 323829
rect 216354 323593 216396 323829
rect 216076 323509 216396 323593
rect 216076 323273 216118 323509
rect 216354 323273 216396 323509
rect 216076 323241 216396 323273
rect 222340 323829 222660 323861
rect 222340 323593 222382 323829
rect 222618 323593 222660 323829
rect 222340 323509 222660 323593
rect 222340 323273 222382 323509
rect 222618 323273 222660 323509
rect 222340 323241 222660 323273
rect 228604 323829 228924 323861
rect 228604 323593 228646 323829
rect 228882 323593 228924 323829
rect 228604 323509 228924 323593
rect 228604 323273 228646 323509
rect 228882 323273 228924 323509
rect 228604 323241 228924 323273
rect 244076 323829 244396 323861
rect 244076 323593 244118 323829
rect 244354 323593 244396 323829
rect 244076 323509 244396 323593
rect 244076 323273 244118 323509
rect 244354 323273 244396 323509
rect 244076 323241 244396 323273
rect 250340 323829 250660 323861
rect 250340 323593 250382 323829
rect 250618 323593 250660 323829
rect 250340 323509 250660 323593
rect 250340 323273 250382 323509
rect 250618 323273 250660 323509
rect 250340 323241 250660 323273
rect 256604 323829 256924 323861
rect 256604 323593 256646 323829
rect 256882 323593 256924 323829
rect 256604 323509 256924 323593
rect 256604 323273 256646 323509
rect 256882 323273 256924 323509
rect 256604 323241 256924 323273
rect 272076 323829 272396 323861
rect 272076 323593 272118 323829
rect 272354 323593 272396 323829
rect 272076 323509 272396 323593
rect 272076 323273 272118 323509
rect 272354 323273 272396 323509
rect 272076 323241 272396 323273
rect 278340 323829 278660 323861
rect 278340 323593 278382 323829
rect 278618 323593 278660 323829
rect 278340 323509 278660 323593
rect 278340 323273 278382 323509
rect 278618 323273 278660 323509
rect 278340 323241 278660 323273
rect 284604 323829 284924 323861
rect 284604 323593 284646 323829
rect 284882 323593 284924 323829
rect 284604 323509 284924 323593
rect 284604 323273 284646 323509
rect 284882 323273 284924 323509
rect 284604 323241 284924 323273
rect 300076 323829 300396 323861
rect 300076 323593 300118 323829
rect 300354 323593 300396 323829
rect 300076 323509 300396 323593
rect 300076 323273 300118 323509
rect 300354 323273 300396 323509
rect 300076 323241 300396 323273
rect 306340 323829 306660 323861
rect 306340 323593 306382 323829
rect 306618 323593 306660 323829
rect 306340 323509 306660 323593
rect 306340 323273 306382 323509
rect 306618 323273 306660 323509
rect 306340 323241 306660 323273
rect 312604 323829 312924 323861
rect 312604 323593 312646 323829
rect 312882 323593 312924 323829
rect 312604 323509 312924 323593
rect 312604 323273 312646 323509
rect 312882 323273 312924 323509
rect 312604 323241 312924 323273
rect 328076 323829 328396 323861
rect 328076 323593 328118 323829
rect 328354 323593 328396 323829
rect 328076 323509 328396 323593
rect 328076 323273 328118 323509
rect 328354 323273 328396 323509
rect 328076 323241 328396 323273
rect 334340 323829 334660 323861
rect 334340 323593 334382 323829
rect 334618 323593 334660 323829
rect 334340 323509 334660 323593
rect 334340 323273 334382 323509
rect 334618 323273 334660 323509
rect 334340 323241 334660 323273
rect 340604 323829 340924 323861
rect 340604 323593 340646 323829
rect 340882 323593 340924 323829
rect 340604 323509 340924 323593
rect 340604 323273 340646 323509
rect 340882 323273 340924 323509
rect 340604 323241 340924 323273
rect 356076 323829 356396 323861
rect 356076 323593 356118 323829
rect 356354 323593 356396 323829
rect 356076 323509 356396 323593
rect 356076 323273 356118 323509
rect 356354 323273 356396 323509
rect 356076 323241 356396 323273
rect 362340 323829 362660 323861
rect 362340 323593 362382 323829
rect 362618 323593 362660 323829
rect 362340 323509 362660 323593
rect 362340 323273 362382 323509
rect 362618 323273 362660 323509
rect 362340 323241 362660 323273
rect 368604 323829 368924 323861
rect 368604 323593 368646 323829
rect 368882 323593 368924 323829
rect 368604 323509 368924 323593
rect 368604 323273 368646 323509
rect 368882 323273 368924 323509
rect 368604 323241 368924 323273
rect 384076 323829 384396 323861
rect 384076 323593 384118 323829
rect 384354 323593 384396 323829
rect 384076 323509 384396 323593
rect 384076 323273 384118 323509
rect 384354 323273 384396 323509
rect 384076 323241 384396 323273
rect 390340 323829 390660 323861
rect 390340 323593 390382 323829
rect 390618 323593 390660 323829
rect 390340 323509 390660 323593
rect 390340 323273 390382 323509
rect 390618 323273 390660 323509
rect 390340 323241 390660 323273
rect 197472 320454 197792 320486
rect 197472 320218 197514 320454
rect 197750 320218 197792 320454
rect 197472 320134 197792 320218
rect 197472 319898 197514 320134
rect 197750 319898 197792 320134
rect 197472 319866 197792 319898
rect 219208 320454 219528 320486
rect 219208 320218 219250 320454
rect 219486 320218 219528 320454
rect 219208 320134 219528 320218
rect 219208 319898 219250 320134
rect 219486 319898 219528 320134
rect 219208 319866 219528 319898
rect 225472 320454 225792 320486
rect 225472 320218 225514 320454
rect 225750 320218 225792 320454
rect 225472 320134 225792 320218
rect 225472 319898 225514 320134
rect 225750 319898 225792 320134
rect 225472 319866 225792 319898
rect 247208 320454 247528 320486
rect 247208 320218 247250 320454
rect 247486 320218 247528 320454
rect 247208 320134 247528 320218
rect 247208 319898 247250 320134
rect 247486 319898 247528 320134
rect 247208 319866 247528 319898
rect 253472 320454 253792 320486
rect 253472 320218 253514 320454
rect 253750 320218 253792 320454
rect 253472 320134 253792 320218
rect 253472 319898 253514 320134
rect 253750 319898 253792 320134
rect 253472 319866 253792 319898
rect 275208 320454 275528 320486
rect 275208 320218 275250 320454
rect 275486 320218 275528 320454
rect 275208 320134 275528 320218
rect 275208 319898 275250 320134
rect 275486 319898 275528 320134
rect 275208 319866 275528 319898
rect 281472 320454 281792 320486
rect 281472 320218 281514 320454
rect 281750 320218 281792 320454
rect 281472 320134 281792 320218
rect 281472 319898 281514 320134
rect 281750 319898 281792 320134
rect 281472 319866 281792 319898
rect 303208 320454 303528 320486
rect 303208 320218 303250 320454
rect 303486 320218 303528 320454
rect 303208 320134 303528 320218
rect 303208 319898 303250 320134
rect 303486 319898 303528 320134
rect 303208 319866 303528 319898
rect 309472 320454 309792 320486
rect 309472 320218 309514 320454
rect 309750 320218 309792 320454
rect 309472 320134 309792 320218
rect 309472 319898 309514 320134
rect 309750 319898 309792 320134
rect 309472 319866 309792 319898
rect 331208 320454 331528 320486
rect 331208 320218 331250 320454
rect 331486 320218 331528 320454
rect 331208 320134 331528 320218
rect 331208 319898 331250 320134
rect 331486 319898 331528 320134
rect 331208 319866 331528 319898
rect 337472 320454 337792 320486
rect 337472 320218 337514 320454
rect 337750 320218 337792 320454
rect 337472 320134 337792 320218
rect 337472 319898 337514 320134
rect 337750 319898 337792 320134
rect 337472 319866 337792 319898
rect 359208 320454 359528 320486
rect 359208 320218 359250 320454
rect 359486 320218 359528 320454
rect 359208 320134 359528 320218
rect 359208 319898 359250 320134
rect 359486 319898 359528 320134
rect 359208 319866 359528 319898
rect 365472 320454 365792 320486
rect 365472 320218 365514 320454
rect 365750 320218 365792 320454
rect 365472 320134 365792 320218
rect 365472 319898 365514 320134
rect 365750 319898 365792 320134
rect 365472 319866 365792 319898
rect 387208 320454 387528 320486
rect 387208 320218 387250 320454
rect 387486 320218 387528 320454
rect 387208 320134 387528 320218
rect 387208 319898 387250 320134
rect 387486 319898 387528 320134
rect 387208 319866 387528 319898
rect 390878 311813 390938 333235
rect 396604 323829 396924 323861
rect 396604 323593 396646 323829
rect 396882 323593 396924 323829
rect 396604 323509 396924 323593
rect 396604 323273 396646 323509
rect 396882 323273 396924 323509
rect 396604 323241 396924 323273
rect 412076 323829 412396 323861
rect 412076 323593 412118 323829
rect 412354 323593 412396 323829
rect 412076 323509 412396 323593
rect 412076 323273 412118 323509
rect 412354 323273 412396 323509
rect 412076 323241 412396 323273
rect 418340 323829 418660 323861
rect 418340 323593 418382 323829
rect 418618 323593 418660 323829
rect 418340 323509 418660 323593
rect 418340 323273 418382 323509
rect 418618 323273 418660 323509
rect 418340 323241 418660 323273
rect 424604 323829 424924 323861
rect 424604 323593 424646 323829
rect 424882 323593 424924 323829
rect 424604 323509 424924 323593
rect 424604 323273 424646 323509
rect 424882 323273 424924 323509
rect 424604 323241 424924 323273
rect 440076 323829 440396 323861
rect 440076 323593 440118 323829
rect 440354 323593 440396 323829
rect 440076 323509 440396 323593
rect 440076 323273 440118 323509
rect 440354 323273 440396 323509
rect 440076 323241 440396 323273
rect 446340 323829 446660 323861
rect 446340 323593 446382 323829
rect 446618 323593 446660 323829
rect 446340 323509 446660 323593
rect 446340 323273 446382 323509
rect 446618 323273 446660 323509
rect 446340 323241 446660 323273
rect 452604 323829 452924 323861
rect 452604 323593 452646 323829
rect 452882 323593 452924 323829
rect 452604 323509 452924 323593
rect 452604 323273 452646 323509
rect 452882 323273 452924 323509
rect 452604 323241 452924 323273
rect 468076 323829 468396 323861
rect 468076 323593 468118 323829
rect 468354 323593 468396 323829
rect 468076 323509 468396 323593
rect 468076 323273 468118 323509
rect 468354 323273 468396 323509
rect 468076 323241 468396 323273
rect 474340 323829 474660 323861
rect 474340 323593 474382 323829
rect 474618 323593 474660 323829
rect 474340 323509 474660 323593
rect 474340 323273 474382 323509
rect 474618 323273 474660 323509
rect 474340 323241 474660 323273
rect 480604 323829 480924 323861
rect 480604 323593 480646 323829
rect 480882 323593 480924 323829
rect 480604 323509 480924 323593
rect 480604 323273 480646 323509
rect 480882 323273 480924 323509
rect 480604 323241 480924 323273
rect 496076 323829 496396 323861
rect 496076 323593 496118 323829
rect 496354 323593 496396 323829
rect 496076 323509 496396 323593
rect 496076 323273 496118 323509
rect 496354 323273 496396 323509
rect 496076 323241 496396 323273
rect 502340 323829 502660 323861
rect 502340 323593 502382 323829
rect 502618 323593 502660 323829
rect 502340 323509 502660 323593
rect 502340 323273 502382 323509
rect 502618 323273 502660 323509
rect 502340 323241 502660 323273
rect 508604 323829 508924 323861
rect 508604 323593 508646 323829
rect 508882 323593 508924 323829
rect 508604 323509 508924 323593
rect 508604 323273 508646 323509
rect 508882 323273 508924 323509
rect 508604 323241 508924 323273
rect 524076 323829 524396 323861
rect 524076 323593 524118 323829
rect 524354 323593 524396 323829
rect 524076 323509 524396 323593
rect 524076 323273 524118 323509
rect 524354 323273 524396 323509
rect 524076 323241 524396 323273
rect 530340 323829 530660 323861
rect 530340 323593 530382 323829
rect 530618 323593 530660 323829
rect 530340 323509 530660 323593
rect 530340 323273 530382 323509
rect 530618 323273 530660 323509
rect 530340 323241 530660 323273
rect 536604 323829 536924 323861
rect 536604 323593 536646 323829
rect 536882 323593 536924 323829
rect 536604 323509 536924 323593
rect 536604 323273 536646 323509
rect 536882 323273 536924 323509
rect 536604 323241 536924 323273
rect 552076 323829 552396 323861
rect 552076 323593 552118 323829
rect 552354 323593 552396 323829
rect 552076 323509 552396 323593
rect 552076 323273 552118 323509
rect 552354 323273 552396 323509
rect 552076 323241 552396 323273
rect 558340 323829 558660 323861
rect 558340 323593 558382 323829
rect 558618 323593 558660 323829
rect 558340 323509 558660 323593
rect 558340 323273 558382 323509
rect 558618 323273 558660 323509
rect 558340 323241 558660 323273
rect 564604 323829 564924 323861
rect 564604 323593 564646 323829
rect 564882 323593 564924 323829
rect 564604 323509 564924 323593
rect 564604 323273 564646 323509
rect 564882 323273 564924 323509
rect 573494 323829 574114 350273
rect 573494 323593 573526 323829
rect 573762 323593 573846 323829
rect 574082 323593 574114 323829
rect 573494 323509 574114 323593
rect 568435 323372 568501 323373
rect 568435 323370 568436 323372
rect 564604 323241 564924 323273
rect 567334 323310 568436 323370
rect 456379 323236 456445 323237
rect 456379 323172 456380 323236
rect 456444 323172 456445 323236
rect 456379 323171 456445 323172
rect 393472 320454 393792 320486
rect 393472 320218 393514 320454
rect 393750 320218 393792 320454
rect 393472 320134 393792 320218
rect 393472 319898 393514 320134
rect 393750 319898 393792 320134
rect 393472 319866 393792 319898
rect 415208 320454 415528 320486
rect 415208 320218 415250 320454
rect 415486 320218 415528 320454
rect 415208 320134 415528 320218
rect 415208 319898 415250 320134
rect 415486 319898 415528 320134
rect 415208 319866 415528 319898
rect 421472 320454 421792 320486
rect 421472 320218 421514 320454
rect 421750 320218 421792 320454
rect 421472 320134 421792 320218
rect 421472 319898 421514 320134
rect 421750 319898 421792 320134
rect 421472 319866 421792 319898
rect 443208 320454 443528 320486
rect 443208 320218 443250 320454
rect 443486 320218 443528 320454
rect 443208 320134 443528 320218
rect 443208 319898 443250 320134
rect 443486 319898 443528 320134
rect 443208 319866 443528 319898
rect 449472 320454 449792 320486
rect 449472 320218 449514 320454
rect 449750 320218 449792 320454
rect 449472 320134 449792 320218
rect 449472 319898 449514 320134
rect 449750 319898 449792 320134
rect 449472 319866 449792 319898
rect 456382 316050 456442 323171
rect 471208 320454 471528 320486
rect 471208 320218 471250 320454
rect 471486 320218 471528 320454
rect 471208 320134 471528 320218
rect 471208 319898 471250 320134
rect 471486 319898 471528 320134
rect 471208 319866 471528 319898
rect 477472 320454 477792 320486
rect 477472 320218 477514 320454
rect 477750 320218 477792 320454
rect 477472 320134 477792 320218
rect 477472 319898 477514 320134
rect 477750 319898 477792 320134
rect 477472 319866 477792 319898
rect 499208 320454 499528 320486
rect 499208 320218 499250 320454
rect 499486 320218 499528 320454
rect 499208 320134 499528 320218
rect 499208 319898 499250 320134
rect 499486 319898 499528 320134
rect 499208 319866 499528 319898
rect 505472 320454 505792 320486
rect 505472 320218 505514 320454
rect 505750 320218 505792 320454
rect 505472 320134 505792 320218
rect 505472 319898 505514 320134
rect 505750 319898 505792 320134
rect 505472 319866 505792 319898
rect 527208 320454 527528 320486
rect 527208 320218 527250 320454
rect 527486 320218 527528 320454
rect 527208 320134 527528 320218
rect 527208 319898 527250 320134
rect 527486 319898 527528 320134
rect 527208 319866 527528 319898
rect 533472 320454 533792 320486
rect 533472 320218 533514 320454
rect 533750 320218 533792 320454
rect 533472 320134 533792 320218
rect 533472 319898 533514 320134
rect 533750 319898 533792 320134
rect 533472 319866 533792 319898
rect 555208 320454 555528 320486
rect 555208 320218 555250 320454
rect 555486 320218 555528 320454
rect 555208 320134 555528 320218
rect 555208 319898 555250 320134
rect 555486 319898 555528 320134
rect 555208 319866 555528 319898
rect 561472 320454 561792 320486
rect 561472 320218 561514 320454
rect 561750 320218 561792 320454
rect 561472 320134 561792 320218
rect 561472 319898 561514 320134
rect 561750 319898 561792 320134
rect 561472 319866 561792 319898
rect 567334 318810 567394 323310
rect 568435 323308 568436 323310
rect 568500 323308 568501 323372
rect 568435 323307 568501 323308
rect 455462 315990 456442 316050
rect 566966 318750 567394 318810
rect 573494 323273 573526 323509
rect 573762 323273 573846 323509
rect 574082 323273 574114 323509
rect 455462 315349 455522 315990
rect 566966 315349 567026 318750
rect 455459 315348 455525 315349
rect 455459 315284 455460 315348
rect 455524 315284 455525 315348
rect 455459 315283 455525 315284
rect 566963 315348 567029 315349
rect 566963 315284 566964 315348
rect 567028 315284 567029 315348
rect 566963 315283 567029 315284
rect 128307 311812 128373 311813
rect 128307 311748 128308 311812
rect 128372 311748 128373 311812
rect 128307 311747 128373 311748
rect 194731 311812 194797 311813
rect 194731 311748 194732 311812
rect 194796 311748 194797 311812
rect 194731 311747 194797 311748
rect 390875 311812 390941 311813
rect 390875 311748 390876 311812
rect 390940 311748 390941 311812
rect 390875 311747 390941 311748
rect 165659 306508 165725 306509
rect 165659 306444 165660 306508
rect 165724 306444 165725 306508
rect 165659 306443 165725 306444
rect 259499 306508 259565 306509
rect 259499 306444 259500 306508
rect 259564 306444 259565 306508
rect 259499 306443 259565 306444
rect 361619 306508 361685 306509
rect 361619 306444 361620 306508
rect 361684 306444 361685 306508
rect 361619 306443 361685 306444
rect 445707 306508 445773 306509
rect 445707 306444 445708 306508
rect 445772 306444 445773 306508
rect 445707 306443 445773 306444
rect 557579 306508 557645 306509
rect 557579 306444 557580 306508
rect 557644 306444 557645 306508
rect 557579 306443 557645 306444
rect -2006 296593 -1974 296829
rect -1738 296593 -1654 296829
rect -1418 296593 -1386 296829
rect -2006 296509 -1386 296593
rect -2006 296273 -1974 296509
rect -1738 296273 -1654 296509
rect -1418 296273 -1386 296509
rect -2006 269829 -1386 296273
rect 20076 296829 20396 296861
rect 20076 296593 20118 296829
rect 20354 296593 20396 296829
rect 20076 296509 20396 296593
rect 20076 296273 20118 296509
rect 20354 296273 20396 296509
rect 20076 296241 20396 296273
rect 26340 296829 26660 296861
rect 26340 296593 26382 296829
rect 26618 296593 26660 296829
rect 26340 296509 26660 296593
rect 26340 296273 26382 296509
rect 26618 296273 26660 296509
rect 26340 296241 26660 296273
rect 32604 296829 32924 296861
rect 32604 296593 32646 296829
rect 32882 296593 32924 296829
rect 32604 296509 32924 296593
rect 32604 296273 32646 296509
rect 32882 296273 32924 296509
rect 32604 296241 32924 296273
rect 48076 296829 48396 296861
rect 48076 296593 48118 296829
rect 48354 296593 48396 296829
rect 48076 296509 48396 296593
rect 48076 296273 48118 296509
rect 48354 296273 48396 296509
rect 48076 296241 48396 296273
rect 54340 296829 54660 296861
rect 54340 296593 54382 296829
rect 54618 296593 54660 296829
rect 54340 296509 54660 296593
rect 54340 296273 54382 296509
rect 54618 296273 54660 296509
rect 54340 296241 54660 296273
rect 60604 296829 60924 296861
rect 60604 296593 60646 296829
rect 60882 296593 60924 296829
rect 60604 296509 60924 296593
rect 60604 296273 60646 296509
rect 60882 296273 60924 296509
rect 60604 296241 60924 296273
rect 76076 296829 76396 296861
rect 76076 296593 76118 296829
rect 76354 296593 76396 296829
rect 76076 296509 76396 296593
rect 76076 296273 76118 296509
rect 76354 296273 76396 296509
rect 76076 296241 76396 296273
rect 82340 296829 82660 296861
rect 82340 296593 82382 296829
rect 82618 296593 82660 296829
rect 82340 296509 82660 296593
rect 82340 296273 82382 296509
rect 82618 296273 82660 296509
rect 82340 296241 82660 296273
rect 88604 296829 88924 296861
rect 88604 296593 88646 296829
rect 88882 296593 88924 296829
rect 88604 296509 88924 296593
rect 88604 296273 88646 296509
rect 88882 296273 88924 296509
rect 88604 296241 88924 296273
rect 104076 296829 104396 296861
rect 104076 296593 104118 296829
rect 104354 296593 104396 296829
rect 104076 296509 104396 296593
rect 104076 296273 104118 296509
rect 104354 296273 104396 296509
rect 104076 296241 104396 296273
rect 110340 296829 110660 296861
rect 110340 296593 110382 296829
rect 110618 296593 110660 296829
rect 110340 296509 110660 296593
rect 110340 296273 110382 296509
rect 110618 296273 110660 296509
rect 110340 296241 110660 296273
rect 116604 296829 116924 296861
rect 116604 296593 116646 296829
rect 116882 296593 116924 296829
rect 116604 296509 116924 296593
rect 116604 296273 116646 296509
rect 116882 296273 116924 296509
rect 116604 296241 116924 296273
rect 132076 296829 132396 296861
rect 132076 296593 132118 296829
rect 132354 296593 132396 296829
rect 132076 296509 132396 296593
rect 132076 296273 132118 296509
rect 132354 296273 132396 296509
rect 132076 296241 132396 296273
rect 138340 296829 138660 296861
rect 138340 296593 138382 296829
rect 138618 296593 138660 296829
rect 138340 296509 138660 296593
rect 138340 296273 138382 296509
rect 138618 296273 138660 296509
rect 138340 296241 138660 296273
rect 144604 296829 144924 296861
rect 144604 296593 144646 296829
rect 144882 296593 144924 296829
rect 144604 296509 144924 296593
rect 144604 296273 144646 296509
rect 144882 296273 144924 296509
rect 144604 296241 144924 296273
rect 160076 296829 160396 296861
rect 160076 296593 160118 296829
rect 160354 296593 160396 296829
rect 160076 296509 160396 296593
rect 160076 296273 160118 296509
rect 160354 296273 160396 296509
rect 160076 296241 160396 296273
rect 44587 295764 44653 295765
rect 44587 295700 44588 295764
rect 44652 295700 44653 295764
rect 44587 295699 44653 295700
rect 23208 293454 23528 293486
rect 23208 293218 23250 293454
rect 23486 293218 23528 293454
rect 23208 293134 23528 293218
rect 23208 292898 23250 293134
rect 23486 292898 23528 293134
rect 23208 292866 23528 292898
rect 29472 293454 29792 293486
rect 29472 293218 29514 293454
rect 29750 293218 29792 293454
rect 29472 293134 29792 293218
rect 29472 292898 29514 293134
rect 29750 292898 29792 293134
rect 29472 292866 29792 292898
rect 44590 287877 44650 295699
rect 51208 293454 51528 293486
rect 51208 293218 51250 293454
rect 51486 293218 51528 293454
rect 51208 293134 51528 293218
rect 51208 292898 51250 293134
rect 51486 292898 51528 293134
rect 51208 292866 51528 292898
rect 57472 293454 57792 293486
rect 57472 293218 57514 293454
rect 57750 293218 57792 293454
rect 57472 293134 57792 293218
rect 57472 292898 57514 293134
rect 57750 292898 57792 293134
rect 57472 292866 57792 292898
rect 79208 293454 79528 293486
rect 79208 293218 79250 293454
rect 79486 293218 79528 293454
rect 79208 293134 79528 293218
rect 79208 292898 79250 293134
rect 79486 292898 79528 293134
rect 79208 292866 79528 292898
rect 85472 293454 85792 293486
rect 85472 293218 85514 293454
rect 85750 293218 85792 293454
rect 85472 293134 85792 293218
rect 85472 292898 85514 293134
rect 85750 292898 85792 293134
rect 85472 292866 85792 292898
rect 107208 293454 107528 293486
rect 107208 293218 107250 293454
rect 107486 293218 107528 293454
rect 107208 293134 107528 293218
rect 107208 292898 107250 293134
rect 107486 292898 107528 293134
rect 107208 292866 107528 292898
rect 113472 293454 113792 293486
rect 113472 293218 113514 293454
rect 113750 293218 113792 293454
rect 113472 293134 113792 293218
rect 113472 292898 113514 293134
rect 113750 292898 113792 293134
rect 113472 292866 113792 292898
rect 135208 293454 135528 293486
rect 135208 293218 135250 293454
rect 135486 293218 135528 293454
rect 135208 293134 135528 293218
rect 135208 292898 135250 293134
rect 135486 292898 135528 293134
rect 135208 292866 135528 292898
rect 141472 293454 141792 293486
rect 141472 293218 141514 293454
rect 141750 293218 141792 293454
rect 141472 293134 141792 293218
rect 141472 292898 141514 293134
rect 141750 292898 141792 293134
rect 141472 292866 141792 292898
rect 163208 293454 163528 293486
rect 163208 293218 163250 293454
rect 163486 293218 163528 293454
rect 163208 293134 163528 293218
rect 163208 292898 163250 293134
rect 163486 292898 163528 293134
rect 163208 292866 163528 292898
rect 44587 287876 44653 287877
rect 44587 287812 44588 287876
rect 44652 287812 44653 287876
rect 44587 287811 44653 287812
rect 165662 284205 165722 306443
rect 166340 296829 166660 296861
rect 166340 296593 166382 296829
rect 166618 296593 166660 296829
rect 166340 296509 166660 296593
rect 166340 296273 166382 296509
rect 166618 296273 166660 296509
rect 166340 296241 166660 296273
rect 172604 296829 172924 296861
rect 172604 296593 172646 296829
rect 172882 296593 172924 296829
rect 172604 296509 172924 296593
rect 172604 296273 172646 296509
rect 172882 296273 172924 296509
rect 172604 296241 172924 296273
rect 188076 296829 188396 296861
rect 188076 296593 188118 296829
rect 188354 296593 188396 296829
rect 188076 296509 188396 296593
rect 188076 296273 188118 296509
rect 188354 296273 188396 296509
rect 188076 296241 188396 296273
rect 194340 296829 194660 296861
rect 194340 296593 194382 296829
rect 194618 296593 194660 296829
rect 194340 296509 194660 296593
rect 194340 296273 194382 296509
rect 194618 296273 194660 296509
rect 194340 296241 194660 296273
rect 200604 296829 200924 296861
rect 200604 296593 200646 296829
rect 200882 296593 200924 296829
rect 200604 296509 200924 296593
rect 200604 296273 200646 296509
rect 200882 296273 200924 296509
rect 200604 296241 200924 296273
rect 216076 296829 216396 296861
rect 216076 296593 216118 296829
rect 216354 296593 216396 296829
rect 216076 296509 216396 296593
rect 216076 296273 216118 296509
rect 216354 296273 216396 296509
rect 216076 296241 216396 296273
rect 222340 296829 222660 296861
rect 222340 296593 222382 296829
rect 222618 296593 222660 296829
rect 222340 296509 222660 296593
rect 222340 296273 222382 296509
rect 222618 296273 222660 296509
rect 222340 296241 222660 296273
rect 228604 296829 228924 296861
rect 228604 296593 228646 296829
rect 228882 296593 228924 296829
rect 228604 296509 228924 296593
rect 228604 296273 228646 296509
rect 228882 296273 228924 296509
rect 228604 296241 228924 296273
rect 244076 296829 244396 296861
rect 244076 296593 244118 296829
rect 244354 296593 244396 296829
rect 244076 296509 244396 296593
rect 244076 296273 244118 296509
rect 244354 296273 244396 296509
rect 244076 296241 244396 296273
rect 250340 296829 250660 296861
rect 250340 296593 250382 296829
rect 250618 296593 250660 296829
rect 250340 296509 250660 296593
rect 250340 296273 250382 296509
rect 250618 296273 250660 296509
rect 250340 296241 250660 296273
rect 256604 296829 256924 296861
rect 256604 296593 256646 296829
rect 256882 296593 256924 296829
rect 256604 296509 256924 296593
rect 256604 296273 256646 296509
rect 256882 296273 256924 296509
rect 256604 296241 256924 296273
rect 176331 295764 176397 295765
rect 176331 295700 176332 295764
rect 176396 295700 176397 295764
rect 176331 295699 176397 295700
rect 212579 295764 212645 295765
rect 212579 295700 212580 295764
rect 212644 295700 212645 295764
rect 212579 295699 212645 295700
rect 169472 293454 169792 293486
rect 169472 293218 169514 293454
rect 169750 293218 169792 293454
rect 169472 293134 169792 293218
rect 169472 292898 169514 293134
rect 169750 292898 169792 293134
rect 169472 292866 169792 292898
rect 176334 288013 176394 295699
rect 191208 293454 191528 293486
rect 191208 293218 191250 293454
rect 191486 293218 191528 293454
rect 191208 293134 191528 293218
rect 191208 292898 191250 293134
rect 191486 292898 191528 293134
rect 191208 292866 191528 292898
rect 197472 293454 197792 293486
rect 197472 293218 197514 293454
rect 197750 293218 197792 293454
rect 197472 293134 197792 293218
rect 197472 292898 197514 293134
rect 197750 292898 197792 293134
rect 197472 292866 197792 292898
rect 176331 288012 176397 288013
rect 176331 287948 176332 288012
rect 176396 287948 176397 288012
rect 176331 287947 176397 287948
rect 212582 287877 212642 295699
rect 219208 293454 219528 293486
rect 219208 293218 219250 293454
rect 219486 293218 219528 293454
rect 219208 293134 219528 293218
rect 219208 292898 219250 293134
rect 219486 292898 219528 293134
rect 219208 292866 219528 292898
rect 225472 293454 225792 293486
rect 225472 293218 225514 293454
rect 225750 293218 225792 293454
rect 225472 293134 225792 293218
rect 225472 292898 225514 293134
rect 225750 292898 225792 293134
rect 225472 292866 225792 292898
rect 247208 293454 247528 293486
rect 247208 293218 247250 293454
rect 247486 293218 247528 293454
rect 247208 293134 247528 293218
rect 247208 292898 247250 293134
rect 247486 292898 247528 293134
rect 247208 292866 247528 292898
rect 253472 293454 253792 293486
rect 253472 293218 253514 293454
rect 253750 293218 253792 293454
rect 253472 293134 253792 293218
rect 253472 292898 253514 293134
rect 253750 292898 253792 293134
rect 253472 292866 253792 292898
rect 212579 287876 212645 287877
rect 212579 287812 212580 287876
rect 212644 287812 212645 287876
rect 212579 287811 212645 287812
rect 259502 284205 259562 306443
rect 272076 296829 272396 296861
rect 272076 296593 272118 296829
rect 272354 296593 272396 296829
rect 272076 296509 272396 296593
rect 272076 296273 272118 296509
rect 272354 296273 272396 296509
rect 272076 296241 272396 296273
rect 278340 296829 278660 296861
rect 278340 296593 278382 296829
rect 278618 296593 278660 296829
rect 278340 296509 278660 296593
rect 278340 296273 278382 296509
rect 278618 296273 278660 296509
rect 278340 296241 278660 296273
rect 284604 296829 284924 296861
rect 284604 296593 284646 296829
rect 284882 296593 284924 296829
rect 284604 296509 284924 296593
rect 284604 296273 284646 296509
rect 284882 296273 284924 296509
rect 284604 296241 284924 296273
rect 300076 296829 300396 296861
rect 300076 296593 300118 296829
rect 300354 296593 300396 296829
rect 300076 296509 300396 296593
rect 300076 296273 300118 296509
rect 300354 296273 300396 296509
rect 300076 296241 300396 296273
rect 306340 296829 306660 296861
rect 306340 296593 306382 296829
rect 306618 296593 306660 296829
rect 306340 296509 306660 296593
rect 306340 296273 306382 296509
rect 306618 296273 306660 296509
rect 306340 296241 306660 296273
rect 312604 296829 312924 296861
rect 312604 296593 312646 296829
rect 312882 296593 312924 296829
rect 312604 296509 312924 296593
rect 312604 296273 312646 296509
rect 312882 296273 312924 296509
rect 312604 296241 312924 296273
rect 328076 296829 328396 296861
rect 328076 296593 328118 296829
rect 328354 296593 328396 296829
rect 328076 296509 328396 296593
rect 328076 296273 328118 296509
rect 328354 296273 328396 296509
rect 328076 296241 328396 296273
rect 334340 296829 334660 296861
rect 334340 296593 334382 296829
rect 334618 296593 334660 296829
rect 334340 296509 334660 296593
rect 334340 296273 334382 296509
rect 334618 296273 334660 296509
rect 334340 296241 334660 296273
rect 340604 296829 340924 296861
rect 340604 296593 340646 296829
rect 340882 296593 340924 296829
rect 340604 296509 340924 296593
rect 340604 296273 340646 296509
rect 340882 296273 340924 296509
rect 340604 296241 340924 296273
rect 356076 296829 356396 296861
rect 356076 296593 356118 296829
rect 356354 296593 356396 296829
rect 356076 296509 356396 296593
rect 356076 296273 356118 296509
rect 356354 296273 356396 296509
rect 356076 296241 356396 296273
rect 288387 295764 288453 295765
rect 288387 295700 288388 295764
rect 288452 295700 288453 295764
rect 288387 295699 288453 295700
rect 296483 295764 296549 295765
rect 296483 295700 296484 295764
rect 296548 295700 296549 295764
rect 296483 295699 296549 295700
rect 275208 293454 275528 293486
rect 275208 293218 275250 293454
rect 275486 293218 275528 293454
rect 275208 293134 275528 293218
rect 275208 292898 275250 293134
rect 275486 292898 275528 293134
rect 275208 292866 275528 292898
rect 281472 293454 281792 293486
rect 281472 293218 281514 293454
rect 281750 293218 281792 293454
rect 281472 293134 281792 293218
rect 281472 292898 281514 293134
rect 281750 292898 281792 293134
rect 281472 292866 281792 292898
rect 288390 287741 288450 295699
rect 296486 289830 296546 295699
rect 303208 293454 303528 293486
rect 303208 293218 303250 293454
rect 303486 293218 303528 293454
rect 303208 293134 303528 293218
rect 303208 292898 303250 293134
rect 303486 292898 303528 293134
rect 303208 292866 303528 292898
rect 309472 293454 309792 293486
rect 309472 293218 309514 293454
rect 309750 293218 309792 293454
rect 309472 293134 309792 293218
rect 309472 292898 309514 293134
rect 309750 292898 309792 293134
rect 309472 292866 309792 292898
rect 331208 293454 331528 293486
rect 331208 293218 331250 293454
rect 331486 293218 331528 293454
rect 331208 293134 331528 293218
rect 331208 292898 331250 293134
rect 331486 292898 331528 293134
rect 331208 292866 331528 292898
rect 337472 293454 337792 293486
rect 337472 293218 337514 293454
rect 337750 293218 337792 293454
rect 337472 293134 337792 293218
rect 337472 292898 337514 293134
rect 337750 292898 337792 293134
rect 337472 292866 337792 292898
rect 359208 293454 359528 293486
rect 359208 293218 359250 293454
rect 359486 293218 359528 293454
rect 359208 293134 359528 293218
rect 359208 292898 359250 293134
rect 359486 292898 359528 293134
rect 359208 292866 359528 292898
rect 296486 289770 296914 289830
rect 296854 287877 296914 289770
rect 296851 287876 296917 287877
rect 296851 287812 296852 287876
rect 296916 287812 296917 287876
rect 296851 287811 296917 287812
rect 288387 287740 288453 287741
rect 288387 287676 288388 287740
rect 288452 287676 288453 287740
rect 288387 287675 288453 287676
rect 361622 284205 361682 306443
rect 362340 296829 362660 296861
rect 362340 296593 362382 296829
rect 362618 296593 362660 296829
rect 362340 296509 362660 296593
rect 362340 296273 362382 296509
rect 362618 296273 362660 296509
rect 362340 296241 362660 296273
rect 368604 296829 368924 296861
rect 368604 296593 368646 296829
rect 368882 296593 368924 296829
rect 368604 296509 368924 296593
rect 368604 296273 368646 296509
rect 368882 296273 368924 296509
rect 368604 296241 368924 296273
rect 384076 296829 384396 296861
rect 384076 296593 384118 296829
rect 384354 296593 384396 296829
rect 384076 296509 384396 296593
rect 384076 296273 384118 296509
rect 384354 296273 384396 296509
rect 384076 296241 384396 296273
rect 390340 296829 390660 296861
rect 390340 296593 390382 296829
rect 390618 296593 390660 296829
rect 390340 296509 390660 296593
rect 390340 296273 390382 296509
rect 390618 296273 390660 296509
rect 390340 296241 390660 296273
rect 396604 296829 396924 296861
rect 396604 296593 396646 296829
rect 396882 296593 396924 296829
rect 396604 296509 396924 296593
rect 396604 296273 396646 296509
rect 396882 296273 396924 296509
rect 396604 296241 396924 296273
rect 412076 296829 412396 296861
rect 412076 296593 412118 296829
rect 412354 296593 412396 296829
rect 412076 296509 412396 296593
rect 412076 296273 412118 296509
rect 412354 296273 412396 296509
rect 412076 296241 412396 296273
rect 418340 296829 418660 296861
rect 418340 296593 418382 296829
rect 418618 296593 418660 296829
rect 418340 296509 418660 296593
rect 418340 296273 418382 296509
rect 418618 296273 418660 296509
rect 418340 296241 418660 296273
rect 424604 296829 424924 296861
rect 424604 296593 424646 296829
rect 424882 296593 424924 296829
rect 424604 296509 424924 296593
rect 424604 296273 424646 296509
rect 424882 296273 424924 296509
rect 424604 296241 424924 296273
rect 440076 296829 440396 296861
rect 440076 296593 440118 296829
rect 440354 296593 440396 296829
rect 440076 296509 440396 296593
rect 440076 296273 440118 296509
rect 440354 296273 440396 296509
rect 440076 296241 440396 296273
rect 372291 295764 372357 295765
rect 372291 295700 372292 295764
rect 372356 295700 372357 295764
rect 372291 295699 372357 295700
rect 408539 295764 408605 295765
rect 408539 295700 408540 295764
rect 408604 295700 408605 295764
rect 408539 295699 408605 295700
rect 365472 293454 365792 293486
rect 365472 293218 365514 293454
rect 365750 293218 365792 293454
rect 365472 293134 365792 293218
rect 365472 292898 365514 293134
rect 365750 292898 365792 293134
rect 365472 292866 365792 292898
rect 372294 288013 372354 295699
rect 387208 293454 387528 293486
rect 387208 293218 387250 293454
rect 387486 293218 387528 293454
rect 387208 293134 387528 293218
rect 387208 292898 387250 293134
rect 387486 292898 387528 293134
rect 387208 292866 387528 292898
rect 393472 293454 393792 293486
rect 393472 293218 393514 293454
rect 393750 293218 393792 293454
rect 393472 293134 393792 293218
rect 393472 292898 393514 293134
rect 393750 292898 393792 293134
rect 393472 292866 393792 292898
rect 372291 288012 372357 288013
rect 372291 287948 372292 288012
rect 372356 287948 372357 288012
rect 372291 287947 372357 287948
rect 408542 287877 408602 295699
rect 415208 293454 415528 293486
rect 415208 293218 415250 293454
rect 415486 293218 415528 293454
rect 415208 293134 415528 293218
rect 415208 292898 415250 293134
rect 415486 292898 415528 293134
rect 415208 292866 415528 292898
rect 421472 293454 421792 293486
rect 421472 293218 421514 293454
rect 421750 293218 421792 293454
rect 421472 293134 421792 293218
rect 421472 292898 421514 293134
rect 421750 292898 421792 293134
rect 421472 292866 421792 292898
rect 443208 293454 443528 293486
rect 443208 293218 443250 293454
rect 443486 293218 443528 293454
rect 443208 293134 443528 293218
rect 443208 292898 443250 293134
rect 443486 292898 443528 293134
rect 443208 292866 443528 292898
rect 408539 287876 408605 287877
rect 408539 287812 408540 287876
rect 408604 287812 408605 287876
rect 408539 287811 408605 287812
rect 445710 284205 445770 306443
rect 446340 296829 446660 296861
rect 446340 296593 446382 296829
rect 446618 296593 446660 296829
rect 446340 296509 446660 296593
rect 446340 296273 446382 296509
rect 446618 296273 446660 296509
rect 446340 296241 446660 296273
rect 452604 296829 452924 296861
rect 452604 296593 452646 296829
rect 452882 296593 452924 296829
rect 452604 296509 452924 296593
rect 452604 296273 452646 296509
rect 452882 296273 452924 296509
rect 452604 296241 452924 296273
rect 468076 296829 468396 296861
rect 468076 296593 468118 296829
rect 468354 296593 468396 296829
rect 468076 296509 468396 296593
rect 468076 296273 468118 296509
rect 468354 296273 468396 296509
rect 468076 296241 468396 296273
rect 474340 296829 474660 296861
rect 474340 296593 474382 296829
rect 474618 296593 474660 296829
rect 474340 296509 474660 296593
rect 474340 296273 474382 296509
rect 474618 296273 474660 296509
rect 474340 296241 474660 296273
rect 480604 296829 480924 296861
rect 480604 296593 480646 296829
rect 480882 296593 480924 296829
rect 480604 296509 480924 296593
rect 480604 296273 480646 296509
rect 480882 296273 480924 296509
rect 480604 296241 480924 296273
rect 496076 296829 496396 296861
rect 496076 296593 496118 296829
rect 496354 296593 496396 296829
rect 496076 296509 496396 296593
rect 496076 296273 496118 296509
rect 496354 296273 496396 296509
rect 496076 296241 496396 296273
rect 502340 296829 502660 296861
rect 502340 296593 502382 296829
rect 502618 296593 502660 296829
rect 502340 296509 502660 296593
rect 502340 296273 502382 296509
rect 502618 296273 502660 296509
rect 502340 296241 502660 296273
rect 508604 296829 508924 296861
rect 508604 296593 508646 296829
rect 508882 296593 508924 296829
rect 508604 296509 508924 296593
rect 508604 296273 508646 296509
rect 508882 296273 508924 296509
rect 508604 296241 508924 296273
rect 524076 296829 524396 296861
rect 524076 296593 524118 296829
rect 524354 296593 524396 296829
rect 524076 296509 524396 296593
rect 524076 296273 524118 296509
rect 524354 296273 524396 296509
rect 524076 296241 524396 296273
rect 530340 296829 530660 296861
rect 530340 296593 530382 296829
rect 530618 296593 530660 296829
rect 530340 296509 530660 296593
rect 530340 296273 530382 296509
rect 530618 296273 530660 296509
rect 530340 296241 530660 296273
rect 536604 296829 536924 296861
rect 536604 296593 536646 296829
rect 536882 296593 536924 296829
rect 536604 296509 536924 296593
rect 536604 296273 536646 296509
rect 536882 296273 536924 296509
rect 536604 296241 536924 296273
rect 552076 296829 552396 296861
rect 552076 296593 552118 296829
rect 552354 296593 552396 296829
rect 552076 296509 552396 296593
rect 552076 296273 552118 296509
rect 552354 296273 552396 296509
rect 552076 296241 552396 296273
rect 484347 295764 484413 295765
rect 484347 295700 484348 295764
rect 484412 295700 484413 295764
rect 484347 295699 484413 295700
rect 492627 295764 492693 295765
rect 492627 295700 492628 295764
rect 492692 295700 492693 295764
rect 492627 295699 492693 295700
rect 520595 295764 520661 295765
rect 520595 295700 520596 295764
rect 520660 295700 520661 295764
rect 520595 295699 520661 295700
rect 449472 293454 449792 293486
rect 449472 293218 449514 293454
rect 449750 293218 449792 293454
rect 449472 293134 449792 293218
rect 449472 292898 449514 293134
rect 449750 292898 449792 293134
rect 449472 292866 449792 292898
rect 471208 293454 471528 293486
rect 471208 293218 471250 293454
rect 471486 293218 471528 293454
rect 471208 293134 471528 293218
rect 471208 292898 471250 293134
rect 471486 292898 471528 293134
rect 471208 292866 471528 292898
rect 477472 293454 477792 293486
rect 477472 293218 477514 293454
rect 477750 293218 477792 293454
rect 477472 293134 477792 293218
rect 477472 292898 477514 293134
rect 477750 292898 477792 293134
rect 477472 292866 477792 292898
rect 484350 287741 484410 295699
rect 492630 287877 492690 295699
rect 499208 293454 499528 293486
rect 499208 293218 499250 293454
rect 499486 293218 499528 293454
rect 499208 293134 499528 293218
rect 499208 292898 499250 293134
rect 499486 292898 499528 293134
rect 499208 292866 499528 292898
rect 505472 293454 505792 293486
rect 505472 293218 505514 293454
rect 505750 293218 505792 293454
rect 505472 293134 505792 293218
rect 505472 292898 505514 293134
rect 505750 292898 505792 293134
rect 505472 292866 505792 292898
rect 520598 288013 520658 295699
rect 527208 293454 527528 293486
rect 527208 293218 527250 293454
rect 527486 293218 527528 293454
rect 527208 293134 527528 293218
rect 527208 292898 527250 293134
rect 527486 292898 527528 293134
rect 527208 292866 527528 292898
rect 533472 293454 533792 293486
rect 533472 293218 533514 293454
rect 533750 293218 533792 293454
rect 533472 293134 533792 293218
rect 533472 292898 533514 293134
rect 533750 292898 533792 293134
rect 533472 292866 533792 292898
rect 555208 293454 555528 293486
rect 555208 293218 555250 293454
rect 555486 293218 555528 293454
rect 555208 293134 555528 293218
rect 555208 292898 555250 293134
rect 555486 292898 555528 293134
rect 555208 292866 555528 292898
rect 520595 288012 520661 288013
rect 520595 287948 520596 288012
rect 520660 287948 520661 288012
rect 520595 287947 520661 287948
rect 492627 287876 492693 287877
rect 492627 287812 492628 287876
rect 492692 287812 492693 287876
rect 492627 287811 492693 287812
rect 484347 287740 484413 287741
rect 484347 287676 484348 287740
rect 484412 287676 484413 287740
rect 484347 287675 484413 287676
rect 557582 284205 557642 306443
rect 558340 296829 558660 296861
rect 558340 296593 558382 296829
rect 558618 296593 558660 296829
rect 558340 296509 558660 296593
rect 558340 296273 558382 296509
rect 558618 296273 558660 296509
rect 558340 296241 558660 296273
rect 564604 296829 564924 296861
rect 564604 296593 564646 296829
rect 564882 296593 564924 296829
rect 564604 296509 564924 296593
rect 564604 296273 564646 296509
rect 564882 296273 564924 296509
rect 564604 296241 564924 296273
rect 573494 296829 574114 323273
rect 573494 296593 573526 296829
rect 573762 296593 573846 296829
rect 574082 296593 574114 296829
rect 573494 296509 574114 296593
rect 573494 296273 573526 296509
rect 573762 296273 573846 296509
rect 574082 296273 574114 296509
rect 561472 293454 561792 293486
rect 561472 293218 561514 293454
rect 561750 293218 561792 293454
rect 561472 293134 561792 293218
rect 561472 292898 561514 293134
rect 561750 292898 561792 293134
rect 561472 292866 561792 292898
rect 165659 284204 165725 284205
rect 165659 284140 165660 284204
rect 165724 284140 165725 284204
rect 165659 284139 165725 284140
rect 259499 284204 259565 284205
rect 259499 284140 259500 284204
rect 259564 284140 259565 284204
rect 259499 284139 259565 284140
rect 361619 284204 361685 284205
rect 361619 284140 361620 284204
rect 361684 284140 361685 284204
rect 361619 284139 361685 284140
rect 445707 284204 445773 284205
rect 445707 284140 445708 284204
rect 445772 284140 445773 284204
rect 445707 284139 445773 284140
rect 557579 284204 557645 284205
rect 557579 284140 557580 284204
rect 557644 284140 557645 284204
rect 557579 284139 557645 284140
rect 277347 279852 277413 279853
rect 277347 279850 277348 279852
rect 277166 279790 277348 279850
rect 81387 279308 81453 279309
rect 81387 279244 81388 279308
rect 81452 279244 81453 279308
rect 81387 279243 81453 279244
rect 128307 279308 128373 279309
rect 128307 279244 128308 279308
rect 128372 279244 128373 279308
rect 128307 279243 128373 279244
rect 194731 279308 194797 279309
rect 194731 279244 194732 279308
rect 194796 279244 194797 279308
rect 194731 279243 194797 279244
rect -2006 269593 -1974 269829
rect -1738 269593 -1654 269829
rect -1418 269593 -1386 269829
rect -2006 269509 -1386 269593
rect -2006 269273 -1974 269509
rect -1738 269273 -1654 269509
rect -1418 269273 -1386 269509
rect -2006 242829 -1386 269273
rect 20076 269829 20396 269861
rect 20076 269593 20118 269829
rect 20354 269593 20396 269829
rect 20076 269509 20396 269593
rect 20076 269273 20118 269509
rect 20354 269273 20396 269509
rect 20076 269241 20396 269273
rect 26340 269829 26660 269861
rect 26340 269593 26382 269829
rect 26618 269593 26660 269829
rect 26340 269509 26660 269593
rect 26340 269273 26382 269509
rect 26618 269273 26660 269509
rect 26340 269241 26660 269273
rect 32604 269829 32924 269861
rect 32604 269593 32646 269829
rect 32882 269593 32924 269829
rect 32604 269509 32924 269593
rect 32604 269273 32646 269509
rect 32882 269273 32924 269509
rect 32604 269241 32924 269273
rect 48076 269829 48396 269861
rect 48076 269593 48118 269829
rect 48354 269593 48396 269829
rect 48076 269509 48396 269593
rect 48076 269273 48118 269509
rect 48354 269273 48396 269509
rect 48076 269241 48396 269273
rect 54340 269829 54660 269861
rect 54340 269593 54382 269829
rect 54618 269593 54660 269829
rect 54340 269509 54660 269593
rect 54340 269273 54382 269509
rect 54618 269273 54660 269509
rect 54340 269241 54660 269273
rect 60604 269829 60924 269861
rect 60604 269593 60646 269829
rect 60882 269593 60924 269829
rect 60604 269509 60924 269593
rect 60604 269273 60646 269509
rect 60882 269273 60924 269509
rect 60604 269241 60924 269273
rect 76076 269829 76396 269861
rect 76076 269593 76118 269829
rect 76354 269593 76396 269829
rect 76076 269509 76396 269593
rect 76076 269273 76118 269509
rect 76354 269273 76396 269509
rect 76076 269241 76396 269273
rect 23208 266454 23528 266486
rect 23208 266218 23250 266454
rect 23486 266218 23528 266454
rect 23208 266134 23528 266218
rect 23208 265898 23250 266134
rect 23486 265898 23528 266134
rect 23208 265866 23528 265898
rect 29472 266454 29792 266486
rect 29472 266218 29514 266454
rect 29750 266218 29792 266454
rect 29472 266134 29792 266218
rect 29472 265898 29514 266134
rect 29750 265898 29792 266134
rect 29472 265866 29792 265898
rect 51208 266454 51528 266486
rect 51208 266218 51250 266454
rect 51486 266218 51528 266454
rect 51208 266134 51528 266218
rect 51208 265898 51250 266134
rect 51486 265898 51528 266134
rect 51208 265866 51528 265898
rect 57472 266454 57792 266486
rect 57472 266218 57514 266454
rect 57750 266218 57792 266454
rect 57472 266134 57792 266218
rect 57472 265898 57514 266134
rect 57750 265898 57792 266134
rect 57472 265866 57792 265898
rect 79208 266454 79528 266486
rect 79208 266218 79250 266454
rect 79486 266218 79528 266454
rect 79208 266134 79528 266218
rect 79208 265898 79250 266134
rect 79486 265898 79528 266134
rect 79208 265866 79528 265898
rect 81390 256597 81450 279243
rect 82340 269829 82660 269861
rect 82340 269593 82382 269829
rect 82618 269593 82660 269829
rect 82340 269509 82660 269593
rect 82340 269273 82382 269509
rect 82618 269273 82660 269509
rect 82340 269241 82660 269273
rect 88604 269829 88924 269861
rect 88604 269593 88646 269829
rect 88882 269593 88924 269829
rect 88604 269509 88924 269593
rect 88604 269273 88646 269509
rect 88882 269273 88924 269509
rect 88604 269241 88924 269273
rect 104076 269829 104396 269861
rect 104076 269593 104118 269829
rect 104354 269593 104396 269829
rect 104076 269509 104396 269593
rect 104076 269273 104118 269509
rect 104354 269273 104396 269509
rect 104076 269241 104396 269273
rect 110340 269829 110660 269861
rect 110340 269593 110382 269829
rect 110618 269593 110660 269829
rect 110340 269509 110660 269593
rect 110340 269273 110382 269509
rect 110618 269273 110660 269509
rect 110340 269241 110660 269273
rect 116604 269829 116924 269861
rect 116604 269593 116646 269829
rect 116882 269593 116924 269829
rect 116604 269509 116924 269593
rect 116604 269273 116646 269509
rect 116882 269273 116924 269509
rect 116604 269241 116924 269273
rect 85472 266454 85792 266486
rect 85472 266218 85514 266454
rect 85750 266218 85792 266454
rect 85472 266134 85792 266218
rect 85472 265898 85514 266134
rect 85750 265898 85792 266134
rect 85472 265866 85792 265898
rect 107208 266454 107528 266486
rect 107208 266218 107250 266454
rect 107486 266218 107528 266454
rect 107208 266134 107528 266218
rect 107208 265898 107250 266134
rect 107486 265898 107528 266134
rect 107208 265866 107528 265898
rect 113472 266454 113792 266486
rect 113472 266218 113514 266454
rect 113750 266218 113792 266454
rect 113472 266134 113792 266218
rect 113472 265898 113514 266134
rect 113750 265898 113792 266134
rect 113472 265866 113792 265898
rect 128310 256597 128370 279243
rect 176331 278084 176397 278085
rect 176331 278020 176332 278084
rect 176396 278020 176397 278084
rect 176331 278019 176397 278020
rect 176334 270333 176394 278019
rect 176331 270332 176397 270333
rect 176331 270268 176332 270332
rect 176396 270268 176397 270332
rect 176331 270267 176397 270268
rect 132076 269829 132396 269861
rect 132076 269593 132118 269829
rect 132354 269593 132396 269829
rect 132076 269509 132396 269593
rect 132076 269273 132118 269509
rect 132354 269273 132396 269509
rect 132076 269241 132396 269273
rect 138340 269829 138660 269861
rect 138340 269593 138382 269829
rect 138618 269593 138660 269829
rect 138340 269509 138660 269593
rect 138340 269273 138382 269509
rect 138618 269273 138660 269509
rect 138340 269241 138660 269273
rect 144604 269829 144924 269861
rect 144604 269593 144646 269829
rect 144882 269593 144924 269829
rect 144604 269509 144924 269593
rect 144604 269273 144646 269509
rect 144882 269273 144924 269509
rect 144604 269241 144924 269273
rect 160076 269829 160396 269861
rect 160076 269593 160118 269829
rect 160354 269593 160396 269829
rect 160076 269509 160396 269593
rect 160076 269273 160118 269509
rect 160354 269273 160396 269509
rect 160076 269241 160396 269273
rect 166340 269829 166660 269861
rect 166340 269593 166382 269829
rect 166618 269593 166660 269829
rect 166340 269509 166660 269593
rect 166340 269273 166382 269509
rect 166618 269273 166660 269509
rect 166340 269241 166660 269273
rect 172604 269829 172924 269861
rect 172604 269593 172646 269829
rect 172882 269593 172924 269829
rect 172604 269509 172924 269593
rect 172604 269273 172646 269509
rect 172882 269273 172924 269509
rect 172604 269241 172924 269273
rect 188076 269829 188396 269861
rect 188076 269593 188118 269829
rect 188354 269593 188396 269829
rect 188076 269509 188396 269593
rect 188076 269273 188118 269509
rect 188354 269273 188396 269509
rect 188076 269241 188396 269273
rect 194340 269829 194660 269861
rect 194340 269593 194382 269829
rect 194618 269593 194660 269829
rect 194340 269509 194660 269593
rect 194340 269273 194382 269509
rect 194618 269273 194660 269509
rect 194340 269241 194660 269273
rect 135208 266454 135528 266486
rect 135208 266218 135250 266454
rect 135486 266218 135528 266454
rect 135208 266134 135528 266218
rect 135208 265898 135250 266134
rect 135486 265898 135528 266134
rect 135208 265866 135528 265898
rect 141472 266454 141792 266486
rect 141472 266218 141514 266454
rect 141750 266218 141792 266454
rect 141472 266134 141792 266218
rect 141472 265898 141514 266134
rect 141750 265898 141792 266134
rect 141472 265866 141792 265898
rect 163208 266454 163528 266486
rect 163208 266218 163250 266454
rect 163486 266218 163528 266454
rect 163208 266134 163528 266218
rect 163208 265898 163250 266134
rect 163486 265898 163528 266134
rect 163208 265866 163528 265898
rect 169472 266454 169792 266486
rect 169472 266218 169514 266454
rect 169750 266218 169792 266454
rect 169472 266134 169792 266218
rect 169472 265898 169514 266134
rect 169750 265898 169792 266134
rect 169472 265866 169792 265898
rect 191208 266454 191528 266486
rect 191208 266218 191250 266454
rect 191486 266218 191528 266454
rect 191208 266134 191528 266218
rect 191208 265898 191250 266134
rect 191486 265898 191528 266134
rect 191208 265866 191528 265898
rect 194734 256597 194794 279243
rect 200604 269829 200924 269861
rect 200604 269593 200646 269829
rect 200882 269593 200924 269829
rect 200604 269509 200924 269593
rect 200604 269273 200646 269509
rect 200882 269273 200924 269509
rect 200604 269241 200924 269273
rect 216076 269829 216396 269861
rect 216076 269593 216118 269829
rect 216354 269593 216396 269829
rect 216076 269509 216396 269593
rect 216076 269273 216118 269509
rect 216354 269273 216396 269509
rect 216076 269241 216396 269273
rect 222340 269829 222660 269861
rect 222340 269593 222382 269829
rect 222618 269593 222660 269829
rect 222340 269509 222660 269593
rect 222340 269273 222382 269509
rect 222618 269273 222660 269509
rect 222340 269241 222660 269273
rect 228604 269829 228924 269861
rect 228604 269593 228646 269829
rect 228882 269593 228924 269829
rect 228604 269509 228924 269593
rect 228604 269273 228646 269509
rect 228882 269273 228924 269509
rect 228604 269241 228924 269273
rect 244076 269829 244396 269861
rect 244076 269593 244118 269829
rect 244354 269593 244396 269829
rect 244076 269509 244396 269593
rect 244076 269273 244118 269509
rect 244354 269273 244396 269509
rect 244076 269241 244396 269273
rect 250340 269829 250660 269861
rect 250340 269593 250382 269829
rect 250618 269593 250660 269829
rect 250340 269509 250660 269593
rect 250340 269273 250382 269509
rect 250618 269273 250660 269509
rect 250340 269241 250660 269273
rect 256604 269829 256924 269861
rect 256604 269593 256646 269829
rect 256882 269593 256924 269829
rect 256604 269509 256924 269593
rect 256604 269273 256646 269509
rect 256882 269273 256924 269509
rect 256604 269241 256924 269273
rect 272076 269829 272396 269861
rect 272076 269593 272118 269829
rect 272354 269593 272396 269829
rect 272076 269509 272396 269593
rect 272076 269273 272118 269509
rect 272354 269273 272396 269509
rect 272076 269241 272396 269273
rect 197472 266454 197792 266486
rect 197472 266218 197514 266454
rect 197750 266218 197792 266454
rect 197472 266134 197792 266218
rect 197472 265898 197514 266134
rect 197750 265898 197792 266134
rect 197472 265866 197792 265898
rect 219208 266454 219528 266486
rect 219208 266218 219250 266454
rect 219486 266218 219528 266454
rect 219208 266134 219528 266218
rect 219208 265898 219250 266134
rect 219486 265898 219528 266134
rect 219208 265866 219528 265898
rect 225472 266454 225792 266486
rect 225472 266218 225514 266454
rect 225750 266218 225792 266454
rect 225472 266134 225792 266218
rect 225472 265898 225514 266134
rect 225750 265898 225792 266134
rect 225472 265866 225792 265898
rect 247208 266454 247528 266486
rect 247208 266218 247250 266454
rect 247486 266218 247528 266454
rect 247208 266134 247528 266218
rect 247208 265898 247250 266134
rect 247486 265898 247528 266134
rect 247208 265866 247528 265898
rect 253472 266454 253792 266486
rect 253472 266218 253514 266454
rect 253750 266218 253792 266454
rect 253472 266134 253792 266218
rect 253472 265898 253514 266134
rect 253750 265898 253792 266134
rect 253472 265866 253792 265898
rect 275208 266454 275528 266486
rect 275208 266218 275250 266454
rect 275486 266218 275528 266454
rect 275208 266134 275528 266218
rect 275208 265898 275250 266134
rect 275486 265898 275528 266134
rect 275208 265866 275528 265898
rect 277166 256597 277226 279790
rect 277347 279788 277348 279790
rect 277412 279788 277413 279852
rect 277347 279787 277413 279788
rect 390875 279308 390941 279309
rect 390875 279244 390876 279308
rect 390940 279244 390941 279308
rect 390875 279243 390941 279244
rect 473491 279308 473557 279309
rect 473491 279244 473492 279308
rect 473556 279244 473557 279308
rect 473491 279243 473557 279244
rect 520227 279308 520293 279309
rect 520227 279244 520228 279308
rect 520292 279244 520293 279308
rect 520227 279243 520293 279244
rect 278340 269829 278660 269861
rect 278340 269593 278382 269829
rect 278618 269593 278660 269829
rect 278340 269509 278660 269593
rect 278340 269273 278382 269509
rect 278618 269273 278660 269509
rect 278340 269241 278660 269273
rect 284604 269829 284924 269861
rect 284604 269593 284646 269829
rect 284882 269593 284924 269829
rect 284604 269509 284924 269593
rect 284604 269273 284646 269509
rect 284882 269273 284924 269509
rect 284604 269241 284924 269273
rect 300076 269829 300396 269861
rect 300076 269593 300118 269829
rect 300354 269593 300396 269829
rect 300076 269509 300396 269593
rect 300076 269273 300118 269509
rect 300354 269273 300396 269509
rect 300076 269241 300396 269273
rect 306340 269829 306660 269861
rect 306340 269593 306382 269829
rect 306618 269593 306660 269829
rect 306340 269509 306660 269593
rect 306340 269273 306382 269509
rect 306618 269273 306660 269509
rect 306340 269241 306660 269273
rect 312604 269829 312924 269861
rect 312604 269593 312646 269829
rect 312882 269593 312924 269829
rect 312604 269509 312924 269593
rect 312604 269273 312646 269509
rect 312882 269273 312924 269509
rect 312604 269241 312924 269273
rect 328076 269829 328396 269861
rect 328076 269593 328118 269829
rect 328354 269593 328396 269829
rect 328076 269509 328396 269593
rect 328076 269273 328118 269509
rect 328354 269273 328396 269509
rect 328076 269241 328396 269273
rect 334340 269829 334660 269861
rect 334340 269593 334382 269829
rect 334618 269593 334660 269829
rect 334340 269509 334660 269593
rect 334340 269273 334382 269509
rect 334618 269273 334660 269509
rect 334340 269241 334660 269273
rect 340604 269829 340924 269861
rect 340604 269593 340646 269829
rect 340882 269593 340924 269829
rect 340604 269509 340924 269593
rect 340604 269273 340646 269509
rect 340882 269273 340924 269509
rect 340604 269241 340924 269273
rect 356076 269829 356396 269861
rect 356076 269593 356118 269829
rect 356354 269593 356396 269829
rect 356076 269509 356396 269593
rect 356076 269273 356118 269509
rect 356354 269273 356396 269509
rect 356076 269241 356396 269273
rect 362340 269829 362660 269861
rect 362340 269593 362382 269829
rect 362618 269593 362660 269829
rect 362340 269509 362660 269593
rect 362340 269273 362382 269509
rect 362618 269273 362660 269509
rect 362340 269241 362660 269273
rect 368604 269829 368924 269861
rect 368604 269593 368646 269829
rect 368882 269593 368924 269829
rect 368604 269509 368924 269593
rect 368604 269273 368646 269509
rect 368882 269273 368924 269509
rect 368604 269241 368924 269273
rect 384076 269829 384396 269861
rect 384076 269593 384118 269829
rect 384354 269593 384396 269829
rect 384076 269509 384396 269593
rect 384076 269273 384118 269509
rect 384354 269273 384396 269509
rect 384076 269241 384396 269273
rect 390340 269829 390660 269861
rect 390340 269593 390382 269829
rect 390618 269593 390660 269829
rect 390340 269509 390660 269593
rect 390340 269273 390382 269509
rect 390618 269273 390660 269509
rect 390340 269241 390660 269273
rect 281472 266454 281792 266486
rect 281472 266218 281514 266454
rect 281750 266218 281792 266454
rect 281472 266134 281792 266218
rect 281472 265898 281514 266134
rect 281750 265898 281792 266134
rect 281472 265866 281792 265898
rect 303208 266454 303528 266486
rect 303208 266218 303250 266454
rect 303486 266218 303528 266454
rect 303208 266134 303528 266218
rect 303208 265898 303250 266134
rect 303486 265898 303528 266134
rect 303208 265866 303528 265898
rect 309472 266454 309792 266486
rect 309472 266218 309514 266454
rect 309750 266218 309792 266454
rect 309472 266134 309792 266218
rect 309472 265898 309514 266134
rect 309750 265898 309792 266134
rect 309472 265866 309792 265898
rect 331208 266454 331528 266486
rect 331208 266218 331250 266454
rect 331486 266218 331528 266454
rect 331208 266134 331528 266218
rect 331208 265898 331250 266134
rect 331486 265898 331528 266134
rect 331208 265866 331528 265898
rect 337472 266454 337792 266486
rect 337472 266218 337514 266454
rect 337750 266218 337792 266454
rect 337472 266134 337792 266218
rect 337472 265898 337514 266134
rect 337750 265898 337792 266134
rect 337472 265866 337792 265898
rect 359208 266454 359528 266486
rect 359208 266218 359250 266454
rect 359486 266218 359528 266454
rect 359208 266134 359528 266218
rect 359208 265898 359250 266134
rect 359486 265898 359528 266134
rect 359208 265866 359528 265898
rect 365472 266454 365792 266486
rect 365472 266218 365514 266454
rect 365750 266218 365792 266454
rect 365472 266134 365792 266218
rect 365472 265898 365514 266134
rect 365750 265898 365792 266134
rect 365472 265866 365792 265898
rect 387208 266454 387528 266486
rect 387208 266218 387250 266454
rect 387486 266218 387528 266454
rect 387208 266134 387528 266218
rect 387208 265898 387250 266134
rect 387486 265898 387528 266134
rect 387208 265866 387528 265898
rect 390878 256597 390938 279243
rect 456379 278084 456445 278085
rect 456379 278020 456380 278084
rect 456444 278020 456445 278084
rect 456379 278019 456445 278020
rect 456382 270333 456442 278019
rect 456379 270332 456445 270333
rect 456379 270268 456380 270332
rect 456444 270268 456445 270332
rect 456379 270267 456445 270268
rect 396604 269829 396924 269861
rect 396604 269593 396646 269829
rect 396882 269593 396924 269829
rect 396604 269509 396924 269593
rect 396604 269273 396646 269509
rect 396882 269273 396924 269509
rect 396604 269241 396924 269273
rect 412076 269829 412396 269861
rect 412076 269593 412118 269829
rect 412354 269593 412396 269829
rect 412076 269509 412396 269593
rect 412076 269273 412118 269509
rect 412354 269273 412396 269509
rect 412076 269241 412396 269273
rect 418340 269829 418660 269861
rect 418340 269593 418382 269829
rect 418618 269593 418660 269829
rect 418340 269509 418660 269593
rect 418340 269273 418382 269509
rect 418618 269273 418660 269509
rect 418340 269241 418660 269273
rect 424604 269829 424924 269861
rect 424604 269593 424646 269829
rect 424882 269593 424924 269829
rect 424604 269509 424924 269593
rect 424604 269273 424646 269509
rect 424882 269273 424924 269509
rect 424604 269241 424924 269273
rect 440076 269829 440396 269861
rect 440076 269593 440118 269829
rect 440354 269593 440396 269829
rect 440076 269509 440396 269593
rect 440076 269273 440118 269509
rect 440354 269273 440396 269509
rect 440076 269241 440396 269273
rect 446340 269829 446660 269861
rect 446340 269593 446382 269829
rect 446618 269593 446660 269829
rect 446340 269509 446660 269593
rect 446340 269273 446382 269509
rect 446618 269273 446660 269509
rect 446340 269241 446660 269273
rect 452604 269829 452924 269861
rect 452604 269593 452646 269829
rect 452882 269593 452924 269829
rect 452604 269509 452924 269593
rect 452604 269273 452646 269509
rect 452882 269273 452924 269509
rect 452604 269241 452924 269273
rect 468076 269829 468396 269861
rect 468076 269593 468118 269829
rect 468354 269593 468396 269829
rect 468076 269509 468396 269593
rect 468076 269273 468118 269509
rect 468354 269273 468396 269509
rect 468076 269241 468396 269273
rect 393472 266454 393792 266486
rect 393472 266218 393514 266454
rect 393750 266218 393792 266454
rect 393472 266134 393792 266218
rect 393472 265898 393514 266134
rect 393750 265898 393792 266134
rect 393472 265866 393792 265898
rect 415208 266454 415528 266486
rect 415208 266218 415250 266454
rect 415486 266218 415528 266454
rect 415208 266134 415528 266218
rect 415208 265898 415250 266134
rect 415486 265898 415528 266134
rect 415208 265866 415528 265898
rect 421472 266454 421792 266486
rect 421472 266218 421514 266454
rect 421750 266218 421792 266454
rect 421472 266134 421792 266218
rect 421472 265898 421514 266134
rect 421750 265898 421792 266134
rect 421472 265866 421792 265898
rect 443208 266454 443528 266486
rect 443208 266218 443250 266454
rect 443486 266218 443528 266454
rect 443208 266134 443528 266218
rect 443208 265898 443250 266134
rect 443486 265898 443528 266134
rect 443208 265866 443528 265898
rect 449472 266454 449792 266486
rect 449472 266218 449514 266454
rect 449750 266218 449792 266454
rect 449472 266134 449792 266218
rect 449472 265898 449514 266134
rect 449750 265898 449792 266134
rect 449472 265866 449792 265898
rect 471208 266454 471528 266486
rect 471208 266218 471250 266454
rect 471486 266218 471528 266454
rect 471208 266134 471528 266218
rect 471208 265898 471250 266134
rect 471486 265898 471528 266134
rect 471208 265866 471528 265898
rect 473494 256597 473554 279243
rect 474340 269829 474660 269861
rect 474340 269593 474382 269829
rect 474618 269593 474660 269829
rect 474340 269509 474660 269593
rect 474340 269273 474382 269509
rect 474618 269273 474660 269509
rect 474340 269241 474660 269273
rect 480604 269829 480924 269861
rect 480604 269593 480646 269829
rect 480882 269593 480924 269829
rect 480604 269509 480924 269593
rect 480604 269273 480646 269509
rect 480882 269273 480924 269509
rect 480604 269241 480924 269273
rect 496076 269829 496396 269861
rect 496076 269593 496118 269829
rect 496354 269593 496396 269829
rect 496076 269509 496396 269593
rect 496076 269273 496118 269509
rect 496354 269273 496396 269509
rect 496076 269241 496396 269273
rect 502340 269829 502660 269861
rect 502340 269593 502382 269829
rect 502618 269593 502660 269829
rect 502340 269509 502660 269593
rect 502340 269273 502382 269509
rect 502618 269273 502660 269509
rect 502340 269241 502660 269273
rect 508604 269829 508924 269861
rect 508604 269593 508646 269829
rect 508882 269593 508924 269829
rect 508604 269509 508924 269593
rect 508604 269273 508646 269509
rect 508882 269273 508924 269509
rect 508604 269241 508924 269273
rect 477472 266454 477792 266486
rect 477472 266218 477514 266454
rect 477750 266218 477792 266454
rect 477472 266134 477792 266218
rect 477472 265898 477514 266134
rect 477750 265898 477792 266134
rect 477472 265866 477792 265898
rect 499208 266454 499528 266486
rect 499208 266218 499250 266454
rect 499486 266218 499528 266454
rect 499208 266134 499528 266218
rect 499208 265898 499250 266134
rect 499486 265898 499528 266134
rect 499208 265866 499528 265898
rect 505472 266454 505792 266486
rect 505472 266218 505514 266454
rect 505750 266218 505792 266454
rect 505472 266134 505792 266218
rect 505472 265898 505514 266134
rect 505750 265898 505792 266134
rect 505472 265866 505792 265898
rect 520230 256597 520290 279243
rect 566963 278084 567029 278085
rect 566963 278020 566964 278084
rect 567028 278020 567029 278084
rect 566963 278019 567029 278020
rect 566966 270510 567026 278019
rect 566966 270450 568498 270510
rect 568438 270197 568498 270450
rect 568435 270196 568501 270197
rect 568435 270132 568436 270196
rect 568500 270132 568501 270196
rect 568435 270131 568501 270132
rect 524076 269829 524396 269861
rect 524076 269593 524118 269829
rect 524354 269593 524396 269829
rect 524076 269509 524396 269593
rect 524076 269273 524118 269509
rect 524354 269273 524396 269509
rect 524076 269241 524396 269273
rect 530340 269829 530660 269861
rect 530340 269593 530382 269829
rect 530618 269593 530660 269829
rect 530340 269509 530660 269593
rect 530340 269273 530382 269509
rect 530618 269273 530660 269509
rect 530340 269241 530660 269273
rect 536604 269829 536924 269861
rect 536604 269593 536646 269829
rect 536882 269593 536924 269829
rect 536604 269509 536924 269593
rect 536604 269273 536646 269509
rect 536882 269273 536924 269509
rect 536604 269241 536924 269273
rect 552076 269829 552396 269861
rect 552076 269593 552118 269829
rect 552354 269593 552396 269829
rect 552076 269509 552396 269593
rect 552076 269273 552118 269509
rect 552354 269273 552396 269509
rect 552076 269241 552396 269273
rect 558340 269829 558660 269861
rect 558340 269593 558382 269829
rect 558618 269593 558660 269829
rect 558340 269509 558660 269593
rect 558340 269273 558382 269509
rect 558618 269273 558660 269509
rect 558340 269241 558660 269273
rect 564604 269829 564924 269861
rect 564604 269593 564646 269829
rect 564882 269593 564924 269829
rect 564604 269509 564924 269593
rect 564604 269273 564646 269509
rect 564882 269273 564924 269509
rect 564604 269241 564924 269273
rect 573494 269829 574114 296273
rect 573494 269593 573526 269829
rect 573762 269593 573846 269829
rect 574082 269593 574114 269829
rect 573494 269509 574114 269593
rect 573494 269273 573526 269509
rect 573762 269273 573846 269509
rect 574082 269273 574114 269509
rect 527208 266454 527528 266486
rect 527208 266218 527250 266454
rect 527486 266218 527528 266454
rect 527208 266134 527528 266218
rect 527208 265898 527250 266134
rect 527486 265898 527528 266134
rect 527208 265866 527528 265898
rect 533472 266454 533792 266486
rect 533472 266218 533514 266454
rect 533750 266218 533792 266454
rect 533472 266134 533792 266218
rect 533472 265898 533514 266134
rect 533750 265898 533792 266134
rect 533472 265866 533792 265898
rect 555208 266454 555528 266486
rect 555208 266218 555250 266454
rect 555486 266218 555528 266454
rect 555208 266134 555528 266218
rect 555208 265898 555250 266134
rect 555486 265898 555528 266134
rect 555208 265866 555528 265898
rect 561472 266454 561792 266486
rect 561472 266218 561514 266454
rect 561750 266218 561792 266454
rect 561472 266134 561792 266218
rect 561472 265898 561514 266134
rect 561750 265898 561792 266134
rect 561472 265866 561792 265898
rect 81387 256596 81453 256597
rect 81387 256532 81388 256596
rect 81452 256532 81453 256596
rect 81387 256531 81453 256532
rect 128307 256596 128373 256597
rect 128307 256532 128308 256596
rect 128372 256532 128373 256596
rect 128307 256531 128373 256532
rect 194731 256596 194797 256597
rect 194731 256532 194732 256596
rect 194796 256532 194797 256596
rect 194731 256531 194797 256532
rect 277163 256596 277229 256597
rect 277163 256532 277164 256596
rect 277228 256532 277229 256596
rect 277163 256531 277229 256532
rect 390875 256596 390941 256597
rect 390875 256532 390876 256596
rect 390940 256532 390941 256596
rect 390875 256531 390941 256532
rect 473491 256596 473557 256597
rect 473491 256532 473492 256596
rect 473556 256532 473557 256596
rect 473491 256531 473557 256532
rect 520227 256596 520293 256597
rect 520227 256532 520228 256596
rect 520292 256532 520293 256596
rect 520227 256531 520293 256532
rect 165659 252652 165725 252653
rect 165659 252588 165660 252652
rect 165724 252588 165725 252652
rect 165659 252587 165725 252588
rect 259499 252652 259565 252653
rect 259499 252588 259500 252652
rect 259564 252588 259565 252652
rect 259499 252587 259565 252588
rect 361619 252652 361685 252653
rect 361619 252588 361620 252652
rect 361684 252588 361685 252652
rect 361619 252587 361685 252588
rect 445707 252652 445773 252653
rect 445707 252588 445708 252652
rect 445772 252588 445773 252652
rect 445707 252587 445773 252588
rect 557579 252652 557645 252653
rect 557579 252588 557580 252652
rect 557644 252588 557645 252652
rect 557579 252587 557645 252588
rect -2006 242593 -1974 242829
rect -1738 242593 -1654 242829
rect -1418 242593 -1386 242829
rect -2006 242509 -1386 242593
rect -2006 242273 -1974 242509
rect -1738 242273 -1654 242509
rect -1418 242273 -1386 242509
rect -2006 215829 -1386 242273
rect 20076 242829 20396 242861
rect 20076 242593 20118 242829
rect 20354 242593 20396 242829
rect 20076 242509 20396 242593
rect 20076 242273 20118 242509
rect 20354 242273 20396 242509
rect 20076 242241 20396 242273
rect 26340 242829 26660 242861
rect 26340 242593 26382 242829
rect 26618 242593 26660 242829
rect 26340 242509 26660 242593
rect 26340 242273 26382 242509
rect 26618 242273 26660 242509
rect 26340 242241 26660 242273
rect 32604 242829 32924 242861
rect 32604 242593 32646 242829
rect 32882 242593 32924 242829
rect 32604 242509 32924 242593
rect 32604 242273 32646 242509
rect 32882 242273 32924 242509
rect 32604 242241 32924 242273
rect 48076 242829 48396 242861
rect 48076 242593 48118 242829
rect 48354 242593 48396 242829
rect 48076 242509 48396 242593
rect 48076 242273 48118 242509
rect 48354 242273 48396 242509
rect 48076 242241 48396 242273
rect 54340 242829 54660 242861
rect 54340 242593 54382 242829
rect 54618 242593 54660 242829
rect 54340 242509 54660 242593
rect 54340 242273 54382 242509
rect 54618 242273 54660 242509
rect 54340 242241 54660 242273
rect 60604 242829 60924 242861
rect 60604 242593 60646 242829
rect 60882 242593 60924 242829
rect 60604 242509 60924 242593
rect 60604 242273 60646 242509
rect 60882 242273 60924 242509
rect 60604 242241 60924 242273
rect 76076 242829 76396 242861
rect 76076 242593 76118 242829
rect 76354 242593 76396 242829
rect 76076 242509 76396 242593
rect 76076 242273 76118 242509
rect 76354 242273 76396 242509
rect 76076 242241 76396 242273
rect 82340 242829 82660 242861
rect 82340 242593 82382 242829
rect 82618 242593 82660 242829
rect 82340 242509 82660 242593
rect 82340 242273 82382 242509
rect 82618 242273 82660 242509
rect 82340 242241 82660 242273
rect 88604 242829 88924 242861
rect 88604 242593 88646 242829
rect 88882 242593 88924 242829
rect 88604 242509 88924 242593
rect 88604 242273 88646 242509
rect 88882 242273 88924 242509
rect 88604 242241 88924 242273
rect 104076 242829 104396 242861
rect 104076 242593 104118 242829
rect 104354 242593 104396 242829
rect 104076 242509 104396 242593
rect 104076 242273 104118 242509
rect 104354 242273 104396 242509
rect 104076 242241 104396 242273
rect 110340 242829 110660 242861
rect 110340 242593 110382 242829
rect 110618 242593 110660 242829
rect 110340 242509 110660 242593
rect 110340 242273 110382 242509
rect 110618 242273 110660 242509
rect 110340 242241 110660 242273
rect 116604 242829 116924 242861
rect 116604 242593 116646 242829
rect 116882 242593 116924 242829
rect 116604 242509 116924 242593
rect 116604 242273 116646 242509
rect 116882 242273 116924 242509
rect 116604 242241 116924 242273
rect 132076 242829 132396 242861
rect 132076 242593 132118 242829
rect 132354 242593 132396 242829
rect 132076 242509 132396 242593
rect 132076 242273 132118 242509
rect 132354 242273 132396 242509
rect 132076 242241 132396 242273
rect 138340 242829 138660 242861
rect 138340 242593 138382 242829
rect 138618 242593 138660 242829
rect 138340 242509 138660 242593
rect 138340 242273 138382 242509
rect 138618 242273 138660 242509
rect 138340 242241 138660 242273
rect 144604 242829 144924 242861
rect 144604 242593 144646 242829
rect 144882 242593 144924 242829
rect 144604 242509 144924 242593
rect 144604 242273 144646 242509
rect 144882 242273 144924 242509
rect 144604 242241 144924 242273
rect 160076 242829 160396 242861
rect 160076 242593 160118 242829
rect 160354 242593 160396 242829
rect 160076 242509 160396 242593
rect 160076 242273 160118 242509
rect 160354 242273 160396 242509
rect 160076 242241 160396 242273
rect 23208 239454 23528 239486
rect 23208 239218 23250 239454
rect 23486 239218 23528 239454
rect 23208 239134 23528 239218
rect 23208 238898 23250 239134
rect 23486 238898 23528 239134
rect 23208 238866 23528 238898
rect 29472 239454 29792 239486
rect 29472 239218 29514 239454
rect 29750 239218 29792 239454
rect 29472 239134 29792 239218
rect 29472 238898 29514 239134
rect 29750 238898 29792 239134
rect 29472 238866 29792 238898
rect 51208 239454 51528 239486
rect 51208 239218 51250 239454
rect 51486 239218 51528 239454
rect 51208 239134 51528 239218
rect 51208 238898 51250 239134
rect 51486 238898 51528 239134
rect 51208 238866 51528 238898
rect 57472 239454 57792 239486
rect 57472 239218 57514 239454
rect 57750 239218 57792 239454
rect 57472 239134 57792 239218
rect 57472 238898 57514 239134
rect 57750 238898 57792 239134
rect 57472 238866 57792 238898
rect 79208 239454 79528 239486
rect 79208 239218 79250 239454
rect 79486 239218 79528 239454
rect 79208 239134 79528 239218
rect 79208 238898 79250 239134
rect 79486 238898 79528 239134
rect 79208 238866 79528 238898
rect 85472 239454 85792 239486
rect 85472 239218 85514 239454
rect 85750 239218 85792 239454
rect 85472 239134 85792 239218
rect 85472 238898 85514 239134
rect 85750 238898 85792 239134
rect 85472 238866 85792 238898
rect 107208 239454 107528 239486
rect 107208 239218 107250 239454
rect 107486 239218 107528 239454
rect 107208 239134 107528 239218
rect 107208 238898 107250 239134
rect 107486 238898 107528 239134
rect 107208 238866 107528 238898
rect 113472 239454 113792 239486
rect 113472 239218 113514 239454
rect 113750 239218 113792 239454
rect 113472 239134 113792 239218
rect 113472 238898 113514 239134
rect 113750 238898 113792 239134
rect 113472 238866 113792 238898
rect 135208 239454 135528 239486
rect 135208 239218 135250 239454
rect 135486 239218 135528 239454
rect 135208 239134 135528 239218
rect 135208 238898 135250 239134
rect 135486 238898 135528 239134
rect 135208 238866 135528 238898
rect 141472 239454 141792 239486
rect 141472 239218 141514 239454
rect 141750 239218 141792 239454
rect 141472 239134 141792 239218
rect 141472 238898 141514 239134
rect 141750 238898 141792 239134
rect 141472 238866 141792 238898
rect 163208 239454 163528 239486
rect 163208 239218 163250 239454
rect 163486 239218 163528 239454
rect 163208 239134 163528 239218
rect 163208 238898 163250 239134
rect 163486 238898 163528 239134
rect 163208 238866 163528 238898
rect 165662 230485 165722 252587
rect 166340 242829 166660 242861
rect 166340 242593 166382 242829
rect 166618 242593 166660 242829
rect 166340 242509 166660 242593
rect 166340 242273 166382 242509
rect 166618 242273 166660 242509
rect 166340 242241 166660 242273
rect 172604 242829 172924 242861
rect 172604 242593 172646 242829
rect 172882 242593 172924 242829
rect 172604 242509 172924 242593
rect 172604 242273 172646 242509
rect 172882 242273 172924 242509
rect 172604 242241 172924 242273
rect 188076 242829 188396 242861
rect 188076 242593 188118 242829
rect 188354 242593 188396 242829
rect 188076 242509 188396 242593
rect 188076 242273 188118 242509
rect 188354 242273 188396 242509
rect 188076 242241 188396 242273
rect 194340 242829 194660 242861
rect 194340 242593 194382 242829
rect 194618 242593 194660 242829
rect 194340 242509 194660 242593
rect 194340 242273 194382 242509
rect 194618 242273 194660 242509
rect 194340 242241 194660 242273
rect 200604 242829 200924 242861
rect 200604 242593 200646 242829
rect 200882 242593 200924 242829
rect 200604 242509 200924 242593
rect 200604 242273 200646 242509
rect 200882 242273 200924 242509
rect 200604 242241 200924 242273
rect 216076 242829 216396 242861
rect 216076 242593 216118 242829
rect 216354 242593 216396 242829
rect 216076 242509 216396 242593
rect 216076 242273 216118 242509
rect 216354 242273 216396 242509
rect 216076 242241 216396 242273
rect 222340 242829 222660 242861
rect 222340 242593 222382 242829
rect 222618 242593 222660 242829
rect 222340 242509 222660 242593
rect 222340 242273 222382 242509
rect 222618 242273 222660 242509
rect 222340 242241 222660 242273
rect 228604 242829 228924 242861
rect 228604 242593 228646 242829
rect 228882 242593 228924 242829
rect 228604 242509 228924 242593
rect 228604 242273 228646 242509
rect 228882 242273 228924 242509
rect 228604 242241 228924 242273
rect 244076 242829 244396 242861
rect 244076 242593 244118 242829
rect 244354 242593 244396 242829
rect 244076 242509 244396 242593
rect 244076 242273 244118 242509
rect 244354 242273 244396 242509
rect 244076 242241 244396 242273
rect 250340 242829 250660 242861
rect 250340 242593 250382 242829
rect 250618 242593 250660 242829
rect 250340 242509 250660 242593
rect 250340 242273 250382 242509
rect 250618 242273 250660 242509
rect 250340 242241 250660 242273
rect 256604 242829 256924 242861
rect 256604 242593 256646 242829
rect 256882 242593 256924 242829
rect 256604 242509 256924 242593
rect 256604 242273 256646 242509
rect 256882 242273 256924 242509
rect 256604 242241 256924 242273
rect 169472 239454 169792 239486
rect 169472 239218 169514 239454
rect 169750 239218 169792 239454
rect 169472 239134 169792 239218
rect 169472 238898 169514 239134
rect 169750 238898 169792 239134
rect 169472 238866 169792 238898
rect 191208 239454 191528 239486
rect 191208 239218 191250 239454
rect 191486 239218 191528 239454
rect 191208 239134 191528 239218
rect 191208 238898 191250 239134
rect 191486 238898 191528 239134
rect 191208 238866 191528 238898
rect 197472 239454 197792 239486
rect 197472 239218 197514 239454
rect 197750 239218 197792 239454
rect 197472 239134 197792 239218
rect 197472 238898 197514 239134
rect 197750 238898 197792 239134
rect 197472 238866 197792 238898
rect 219208 239454 219528 239486
rect 219208 239218 219250 239454
rect 219486 239218 219528 239454
rect 219208 239134 219528 239218
rect 219208 238898 219250 239134
rect 219486 238898 219528 239134
rect 219208 238866 219528 238898
rect 225472 239454 225792 239486
rect 225472 239218 225514 239454
rect 225750 239218 225792 239454
rect 225472 239134 225792 239218
rect 225472 238898 225514 239134
rect 225750 238898 225792 239134
rect 225472 238866 225792 238898
rect 247208 239454 247528 239486
rect 247208 239218 247250 239454
rect 247486 239218 247528 239454
rect 247208 239134 247528 239218
rect 247208 238898 247250 239134
rect 247486 238898 247528 239134
rect 247208 238866 247528 238898
rect 253472 239454 253792 239486
rect 253472 239218 253514 239454
rect 253750 239218 253792 239454
rect 253472 239134 253792 239218
rect 253472 238898 253514 239134
rect 253750 238898 253792 239134
rect 253472 238866 253792 238898
rect 259502 230485 259562 252587
rect 272076 242829 272396 242861
rect 272076 242593 272118 242829
rect 272354 242593 272396 242829
rect 272076 242509 272396 242593
rect 272076 242273 272118 242509
rect 272354 242273 272396 242509
rect 272076 242241 272396 242273
rect 278340 242829 278660 242861
rect 278340 242593 278382 242829
rect 278618 242593 278660 242829
rect 278340 242509 278660 242593
rect 278340 242273 278382 242509
rect 278618 242273 278660 242509
rect 278340 242241 278660 242273
rect 284604 242829 284924 242861
rect 284604 242593 284646 242829
rect 284882 242593 284924 242829
rect 284604 242509 284924 242593
rect 284604 242273 284646 242509
rect 284882 242273 284924 242509
rect 284604 242241 284924 242273
rect 300076 242829 300396 242861
rect 300076 242593 300118 242829
rect 300354 242593 300396 242829
rect 300076 242509 300396 242593
rect 300076 242273 300118 242509
rect 300354 242273 300396 242509
rect 300076 242241 300396 242273
rect 306340 242829 306660 242861
rect 306340 242593 306382 242829
rect 306618 242593 306660 242829
rect 306340 242509 306660 242593
rect 306340 242273 306382 242509
rect 306618 242273 306660 242509
rect 306340 242241 306660 242273
rect 312604 242829 312924 242861
rect 312604 242593 312646 242829
rect 312882 242593 312924 242829
rect 312604 242509 312924 242593
rect 312604 242273 312646 242509
rect 312882 242273 312924 242509
rect 312604 242241 312924 242273
rect 328076 242829 328396 242861
rect 328076 242593 328118 242829
rect 328354 242593 328396 242829
rect 328076 242509 328396 242593
rect 328076 242273 328118 242509
rect 328354 242273 328396 242509
rect 328076 242241 328396 242273
rect 334340 242829 334660 242861
rect 334340 242593 334382 242829
rect 334618 242593 334660 242829
rect 334340 242509 334660 242593
rect 334340 242273 334382 242509
rect 334618 242273 334660 242509
rect 334340 242241 334660 242273
rect 340604 242829 340924 242861
rect 340604 242593 340646 242829
rect 340882 242593 340924 242829
rect 340604 242509 340924 242593
rect 340604 242273 340646 242509
rect 340882 242273 340924 242509
rect 340604 242241 340924 242273
rect 356076 242829 356396 242861
rect 356076 242593 356118 242829
rect 356354 242593 356396 242829
rect 356076 242509 356396 242593
rect 356076 242273 356118 242509
rect 356354 242273 356396 242509
rect 356076 242241 356396 242273
rect 275208 239454 275528 239486
rect 275208 239218 275250 239454
rect 275486 239218 275528 239454
rect 275208 239134 275528 239218
rect 275208 238898 275250 239134
rect 275486 238898 275528 239134
rect 275208 238866 275528 238898
rect 281472 239454 281792 239486
rect 281472 239218 281514 239454
rect 281750 239218 281792 239454
rect 281472 239134 281792 239218
rect 281472 238898 281514 239134
rect 281750 238898 281792 239134
rect 281472 238866 281792 238898
rect 303208 239454 303528 239486
rect 303208 239218 303250 239454
rect 303486 239218 303528 239454
rect 303208 239134 303528 239218
rect 303208 238898 303250 239134
rect 303486 238898 303528 239134
rect 303208 238866 303528 238898
rect 309472 239454 309792 239486
rect 309472 239218 309514 239454
rect 309750 239218 309792 239454
rect 309472 239134 309792 239218
rect 309472 238898 309514 239134
rect 309750 238898 309792 239134
rect 309472 238866 309792 238898
rect 331208 239454 331528 239486
rect 331208 239218 331250 239454
rect 331486 239218 331528 239454
rect 331208 239134 331528 239218
rect 331208 238898 331250 239134
rect 331486 238898 331528 239134
rect 331208 238866 331528 238898
rect 337472 239454 337792 239486
rect 337472 239218 337514 239454
rect 337750 239218 337792 239454
rect 337472 239134 337792 239218
rect 337472 238898 337514 239134
rect 337750 238898 337792 239134
rect 337472 238866 337792 238898
rect 359208 239454 359528 239486
rect 359208 239218 359250 239454
rect 359486 239218 359528 239454
rect 359208 239134 359528 239218
rect 359208 238898 359250 239134
rect 359486 238898 359528 239134
rect 359208 238866 359528 238898
rect 361622 230485 361682 252587
rect 362340 242829 362660 242861
rect 362340 242593 362382 242829
rect 362618 242593 362660 242829
rect 362340 242509 362660 242593
rect 362340 242273 362382 242509
rect 362618 242273 362660 242509
rect 362340 242241 362660 242273
rect 368604 242829 368924 242861
rect 368604 242593 368646 242829
rect 368882 242593 368924 242829
rect 368604 242509 368924 242593
rect 368604 242273 368646 242509
rect 368882 242273 368924 242509
rect 368604 242241 368924 242273
rect 384076 242829 384396 242861
rect 384076 242593 384118 242829
rect 384354 242593 384396 242829
rect 384076 242509 384396 242593
rect 384076 242273 384118 242509
rect 384354 242273 384396 242509
rect 384076 242241 384396 242273
rect 390340 242829 390660 242861
rect 390340 242593 390382 242829
rect 390618 242593 390660 242829
rect 390340 242509 390660 242593
rect 390340 242273 390382 242509
rect 390618 242273 390660 242509
rect 390340 242241 390660 242273
rect 396604 242829 396924 242861
rect 396604 242593 396646 242829
rect 396882 242593 396924 242829
rect 396604 242509 396924 242593
rect 396604 242273 396646 242509
rect 396882 242273 396924 242509
rect 396604 242241 396924 242273
rect 412076 242829 412396 242861
rect 412076 242593 412118 242829
rect 412354 242593 412396 242829
rect 412076 242509 412396 242593
rect 412076 242273 412118 242509
rect 412354 242273 412396 242509
rect 412076 242241 412396 242273
rect 418340 242829 418660 242861
rect 418340 242593 418382 242829
rect 418618 242593 418660 242829
rect 418340 242509 418660 242593
rect 418340 242273 418382 242509
rect 418618 242273 418660 242509
rect 418340 242241 418660 242273
rect 424604 242829 424924 242861
rect 424604 242593 424646 242829
rect 424882 242593 424924 242829
rect 424604 242509 424924 242593
rect 424604 242273 424646 242509
rect 424882 242273 424924 242509
rect 424604 242241 424924 242273
rect 440076 242829 440396 242861
rect 440076 242593 440118 242829
rect 440354 242593 440396 242829
rect 440076 242509 440396 242593
rect 440076 242273 440118 242509
rect 440354 242273 440396 242509
rect 440076 242241 440396 242273
rect 365472 239454 365792 239486
rect 365472 239218 365514 239454
rect 365750 239218 365792 239454
rect 365472 239134 365792 239218
rect 365472 238898 365514 239134
rect 365750 238898 365792 239134
rect 365472 238866 365792 238898
rect 387208 239454 387528 239486
rect 387208 239218 387250 239454
rect 387486 239218 387528 239454
rect 387208 239134 387528 239218
rect 387208 238898 387250 239134
rect 387486 238898 387528 239134
rect 387208 238866 387528 238898
rect 393472 239454 393792 239486
rect 393472 239218 393514 239454
rect 393750 239218 393792 239454
rect 393472 239134 393792 239218
rect 393472 238898 393514 239134
rect 393750 238898 393792 239134
rect 393472 238866 393792 238898
rect 415208 239454 415528 239486
rect 415208 239218 415250 239454
rect 415486 239218 415528 239454
rect 415208 239134 415528 239218
rect 415208 238898 415250 239134
rect 415486 238898 415528 239134
rect 415208 238866 415528 238898
rect 421472 239454 421792 239486
rect 421472 239218 421514 239454
rect 421750 239218 421792 239454
rect 421472 239134 421792 239218
rect 421472 238898 421514 239134
rect 421750 238898 421792 239134
rect 421472 238866 421792 238898
rect 443208 239454 443528 239486
rect 443208 239218 443250 239454
rect 443486 239218 443528 239454
rect 443208 239134 443528 239218
rect 443208 238898 443250 239134
rect 443486 238898 443528 239134
rect 443208 238866 443528 238898
rect 445710 230485 445770 252587
rect 446340 242829 446660 242861
rect 446340 242593 446382 242829
rect 446618 242593 446660 242829
rect 446340 242509 446660 242593
rect 446340 242273 446382 242509
rect 446618 242273 446660 242509
rect 446340 242241 446660 242273
rect 452604 242829 452924 242861
rect 452604 242593 452646 242829
rect 452882 242593 452924 242829
rect 452604 242509 452924 242593
rect 452604 242273 452646 242509
rect 452882 242273 452924 242509
rect 452604 242241 452924 242273
rect 468076 242829 468396 242861
rect 468076 242593 468118 242829
rect 468354 242593 468396 242829
rect 468076 242509 468396 242593
rect 468076 242273 468118 242509
rect 468354 242273 468396 242509
rect 468076 242241 468396 242273
rect 474340 242829 474660 242861
rect 474340 242593 474382 242829
rect 474618 242593 474660 242829
rect 474340 242509 474660 242593
rect 474340 242273 474382 242509
rect 474618 242273 474660 242509
rect 474340 242241 474660 242273
rect 480604 242829 480924 242861
rect 480604 242593 480646 242829
rect 480882 242593 480924 242829
rect 480604 242509 480924 242593
rect 480604 242273 480646 242509
rect 480882 242273 480924 242509
rect 480604 242241 480924 242273
rect 496076 242829 496396 242861
rect 496076 242593 496118 242829
rect 496354 242593 496396 242829
rect 496076 242509 496396 242593
rect 496076 242273 496118 242509
rect 496354 242273 496396 242509
rect 496076 242241 496396 242273
rect 502340 242829 502660 242861
rect 502340 242593 502382 242829
rect 502618 242593 502660 242829
rect 502340 242509 502660 242593
rect 502340 242273 502382 242509
rect 502618 242273 502660 242509
rect 502340 242241 502660 242273
rect 508604 242829 508924 242861
rect 508604 242593 508646 242829
rect 508882 242593 508924 242829
rect 508604 242509 508924 242593
rect 508604 242273 508646 242509
rect 508882 242273 508924 242509
rect 508604 242241 508924 242273
rect 524076 242829 524396 242861
rect 524076 242593 524118 242829
rect 524354 242593 524396 242829
rect 524076 242509 524396 242593
rect 524076 242273 524118 242509
rect 524354 242273 524396 242509
rect 524076 242241 524396 242273
rect 530340 242829 530660 242861
rect 530340 242593 530382 242829
rect 530618 242593 530660 242829
rect 530340 242509 530660 242593
rect 530340 242273 530382 242509
rect 530618 242273 530660 242509
rect 530340 242241 530660 242273
rect 536604 242829 536924 242861
rect 536604 242593 536646 242829
rect 536882 242593 536924 242829
rect 536604 242509 536924 242593
rect 536604 242273 536646 242509
rect 536882 242273 536924 242509
rect 536604 242241 536924 242273
rect 552076 242829 552396 242861
rect 552076 242593 552118 242829
rect 552354 242593 552396 242829
rect 552076 242509 552396 242593
rect 552076 242273 552118 242509
rect 552354 242273 552396 242509
rect 552076 242241 552396 242273
rect 449472 239454 449792 239486
rect 449472 239218 449514 239454
rect 449750 239218 449792 239454
rect 449472 239134 449792 239218
rect 449472 238898 449514 239134
rect 449750 238898 449792 239134
rect 449472 238866 449792 238898
rect 471208 239454 471528 239486
rect 471208 239218 471250 239454
rect 471486 239218 471528 239454
rect 471208 239134 471528 239218
rect 471208 238898 471250 239134
rect 471486 238898 471528 239134
rect 471208 238866 471528 238898
rect 477472 239454 477792 239486
rect 477472 239218 477514 239454
rect 477750 239218 477792 239454
rect 477472 239134 477792 239218
rect 477472 238898 477514 239134
rect 477750 238898 477792 239134
rect 477472 238866 477792 238898
rect 499208 239454 499528 239486
rect 499208 239218 499250 239454
rect 499486 239218 499528 239454
rect 499208 239134 499528 239218
rect 499208 238898 499250 239134
rect 499486 238898 499528 239134
rect 499208 238866 499528 238898
rect 505472 239454 505792 239486
rect 505472 239218 505514 239454
rect 505750 239218 505792 239454
rect 505472 239134 505792 239218
rect 505472 238898 505514 239134
rect 505750 238898 505792 239134
rect 505472 238866 505792 238898
rect 527208 239454 527528 239486
rect 527208 239218 527250 239454
rect 527486 239218 527528 239454
rect 527208 239134 527528 239218
rect 527208 238898 527250 239134
rect 527486 238898 527528 239134
rect 527208 238866 527528 238898
rect 533472 239454 533792 239486
rect 533472 239218 533514 239454
rect 533750 239218 533792 239454
rect 533472 239134 533792 239218
rect 533472 238898 533514 239134
rect 533750 238898 533792 239134
rect 533472 238866 533792 238898
rect 555208 239454 555528 239486
rect 555208 239218 555250 239454
rect 555486 239218 555528 239454
rect 555208 239134 555528 239218
rect 555208 238898 555250 239134
rect 555486 238898 555528 239134
rect 555208 238866 555528 238898
rect 557582 230485 557642 252587
rect 558340 242829 558660 242861
rect 558340 242593 558382 242829
rect 558618 242593 558660 242829
rect 558340 242509 558660 242593
rect 558340 242273 558382 242509
rect 558618 242273 558660 242509
rect 558340 242241 558660 242273
rect 564604 242829 564924 242861
rect 564604 242593 564646 242829
rect 564882 242593 564924 242829
rect 564604 242509 564924 242593
rect 564604 242273 564646 242509
rect 564882 242273 564924 242509
rect 564604 242241 564924 242273
rect 573494 242829 574114 269273
rect 573494 242593 573526 242829
rect 573762 242593 573846 242829
rect 574082 242593 574114 242829
rect 573494 242509 574114 242593
rect 573494 242273 573526 242509
rect 573762 242273 573846 242509
rect 574082 242273 574114 242509
rect 561472 239454 561792 239486
rect 561472 239218 561514 239454
rect 561750 239218 561792 239454
rect 561472 239134 561792 239218
rect 561472 238898 561514 239134
rect 561750 238898 561792 239134
rect 561472 238866 561792 238898
rect 165659 230484 165725 230485
rect 165659 230420 165660 230484
rect 165724 230420 165725 230484
rect 165659 230419 165725 230420
rect 259499 230484 259565 230485
rect 259499 230420 259500 230484
rect 259564 230420 259565 230484
rect 259499 230419 259565 230420
rect 361619 230484 361685 230485
rect 361619 230420 361620 230484
rect 361684 230420 361685 230484
rect 361619 230419 361685 230420
rect 445707 230484 445773 230485
rect 445707 230420 445708 230484
rect 445772 230420 445773 230484
rect 445707 230419 445773 230420
rect 557579 230484 557645 230485
rect 557579 230420 557580 230484
rect 557644 230420 557645 230484
rect 557579 230419 557645 230420
rect 128307 225316 128373 225317
rect 128307 225252 128308 225316
rect 128372 225252 128373 225316
rect 128307 225251 128373 225252
rect 194731 225316 194797 225317
rect 194731 225252 194732 225316
rect 194796 225252 194797 225316
rect 194731 225251 194797 225252
rect 92427 224228 92493 224229
rect 92427 224164 92428 224228
rect 92492 224164 92493 224228
rect 92427 224163 92493 224164
rect 64459 224092 64525 224093
rect 64459 224028 64460 224092
rect 64524 224028 64525 224092
rect 64459 224027 64525 224028
rect 64462 216341 64522 224027
rect 92430 216341 92490 224163
rect 64459 216340 64525 216341
rect 64459 216276 64460 216340
rect 64524 216276 64525 216340
rect 64459 216275 64525 216276
rect 92427 216340 92493 216341
rect 92427 216276 92428 216340
rect 92492 216276 92493 216340
rect 92427 216275 92493 216276
rect -2006 215593 -1974 215829
rect -1738 215593 -1654 215829
rect -1418 215593 -1386 215829
rect -2006 215509 -1386 215593
rect -2006 215273 -1974 215509
rect -1738 215273 -1654 215509
rect -1418 215273 -1386 215509
rect -2006 188829 -1386 215273
rect 20076 215829 20396 215861
rect 20076 215593 20118 215829
rect 20354 215593 20396 215829
rect 20076 215509 20396 215593
rect 20076 215273 20118 215509
rect 20354 215273 20396 215509
rect 20076 215241 20396 215273
rect 26340 215829 26660 215861
rect 26340 215593 26382 215829
rect 26618 215593 26660 215829
rect 26340 215509 26660 215593
rect 26340 215273 26382 215509
rect 26618 215273 26660 215509
rect 26340 215241 26660 215273
rect 32604 215829 32924 215861
rect 32604 215593 32646 215829
rect 32882 215593 32924 215829
rect 32604 215509 32924 215593
rect 32604 215273 32646 215509
rect 32882 215273 32924 215509
rect 32604 215241 32924 215273
rect 48076 215829 48396 215861
rect 48076 215593 48118 215829
rect 48354 215593 48396 215829
rect 48076 215509 48396 215593
rect 48076 215273 48118 215509
rect 48354 215273 48396 215509
rect 48076 215241 48396 215273
rect 54340 215829 54660 215861
rect 54340 215593 54382 215829
rect 54618 215593 54660 215829
rect 54340 215509 54660 215593
rect 54340 215273 54382 215509
rect 54618 215273 54660 215509
rect 54340 215241 54660 215273
rect 60604 215829 60924 215861
rect 60604 215593 60646 215829
rect 60882 215593 60924 215829
rect 60604 215509 60924 215593
rect 60604 215273 60646 215509
rect 60882 215273 60924 215509
rect 60604 215241 60924 215273
rect 76076 215829 76396 215861
rect 76076 215593 76118 215829
rect 76354 215593 76396 215829
rect 76076 215509 76396 215593
rect 76076 215273 76118 215509
rect 76354 215273 76396 215509
rect 76076 215241 76396 215273
rect 82340 215829 82660 215861
rect 82340 215593 82382 215829
rect 82618 215593 82660 215829
rect 82340 215509 82660 215593
rect 82340 215273 82382 215509
rect 82618 215273 82660 215509
rect 82340 215241 82660 215273
rect 88604 215829 88924 215861
rect 88604 215593 88646 215829
rect 88882 215593 88924 215829
rect 88604 215509 88924 215593
rect 88604 215273 88646 215509
rect 88882 215273 88924 215509
rect 88604 215241 88924 215273
rect 104076 215829 104396 215861
rect 104076 215593 104118 215829
rect 104354 215593 104396 215829
rect 104076 215509 104396 215593
rect 104076 215273 104118 215509
rect 104354 215273 104396 215509
rect 104076 215241 104396 215273
rect 110340 215829 110660 215861
rect 110340 215593 110382 215829
rect 110618 215593 110660 215829
rect 110340 215509 110660 215593
rect 110340 215273 110382 215509
rect 110618 215273 110660 215509
rect 110340 215241 110660 215273
rect 116604 215829 116924 215861
rect 116604 215593 116646 215829
rect 116882 215593 116924 215829
rect 116604 215509 116924 215593
rect 116604 215273 116646 215509
rect 116882 215273 116924 215509
rect 116604 215241 116924 215273
rect 23208 212454 23528 212486
rect 23208 212218 23250 212454
rect 23486 212218 23528 212454
rect 23208 212134 23528 212218
rect 23208 211898 23250 212134
rect 23486 211898 23528 212134
rect 23208 211866 23528 211898
rect 29472 212454 29792 212486
rect 29472 212218 29514 212454
rect 29750 212218 29792 212454
rect 29472 212134 29792 212218
rect 29472 211898 29514 212134
rect 29750 211898 29792 212134
rect 29472 211866 29792 211898
rect 51208 212454 51528 212486
rect 51208 212218 51250 212454
rect 51486 212218 51528 212454
rect 51208 212134 51528 212218
rect 51208 211898 51250 212134
rect 51486 211898 51528 212134
rect 51208 211866 51528 211898
rect 57472 212454 57792 212486
rect 57472 212218 57514 212454
rect 57750 212218 57792 212454
rect 57472 212134 57792 212218
rect 57472 211898 57514 212134
rect 57750 211898 57792 212134
rect 57472 211866 57792 211898
rect 79208 212454 79528 212486
rect 79208 212218 79250 212454
rect 79486 212218 79528 212454
rect 79208 212134 79528 212218
rect 79208 211898 79250 212134
rect 79486 211898 79528 212134
rect 79208 211866 79528 211898
rect 85472 212454 85792 212486
rect 85472 212218 85514 212454
rect 85750 212218 85792 212454
rect 85472 212134 85792 212218
rect 85472 211898 85514 212134
rect 85750 211898 85792 212134
rect 85472 211866 85792 211898
rect 107208 212454 107528 212486
rect 107208 212218 107250 212454
rect 107486 212218 107528 212454
rect 107208 212134 107528 212218
rect 107208 211898 107250 212134
rect 107486 211898 107528 212134
rect 107208 211866 107528 211898
rect 113472 212454 113792 212486
rect 113472 212218 113514 212454
rect 113750 212218 113792 212454
rect 113472 212134 113792 212218
rect 113472 211898 113514 212134
rect 113750 211898 113792 212134
rect 113472 211866 113792 211898
rect 128310 202877 128370 225251
rect 148363 224228 148429 224229
rect 148363 224164 148364 224228
rect 148428 224164 148429 224228
rect 148363 224163 148429 224164
rect 148366 216341 148426 224163
rect 176331 224092 176397 224093
rect 176331 224028 176332 224092
rect 176396 224028 176397 224092
rect 176331 224027 176397 224028
rect 176334 216341 176394 224027
rect 148363 216340 148429 216341
rect 148363 216276 148364 216340
rect 148428 216276 148429 216340
rect 148363 216275 148429 216276
rect 176331 216340 176397 216341
rect 176331 216276 176332 216340
rect 176396 216276 176397 216340
rect 176331 216275 176397 216276
rect 132076 215829 132396 215861
rect 132076 215593 132118 215829
rect 132354 215593 132396 215829
rect 132076 215509 132396 215593
rect 132076 215273 132118 215509
rect 132354 215273 132396 215509
rect 132076 215241 132396 215273
rect 138340 215829 138660 215861
rect 138340 215593 138382 215829
rect 138618 215593 138660 215829
rect 138340 215509 138660 215593
rect 138340 215273 138382 215509
rect 138618 215273 138660 215509
rect 138340 215241 138660 215273
rect 144604 215829 144924 215861
rect 144604 215593 144646 215829
rect 144882 215593 144924 215829
rect 144604 215509 144924 215593
rect 144604 215273 144646 215509
rect 144882 215273 144924 215509
rect 144604 215241 144924 215273
rect 160076 215829 160396 215861
rect 160076 215593 160118 215829
rect 160354 215593 160396 215829
rect 160076 215509 160396 215593
rect 160076 215273 160118 215509
rect 160354 215273 160396 215509
rect 160076 215241 160396 215273
rect 166340 215829 166660 215861
rect 166340 215593 166382 215829
rect 166618 215593 166660 215829
rect 166340 215509 166660 215593
rect 166340 215273 166382 215509
rect 166618 215273 166660 215509
rect 166340 215241 166660 215273
rect 172604 215829 172924 215861
rect 172604 215593 172646 215829
rect 172882 215593 172924 215829
rect 172604 215509 172924 215593
rect 172604 215273 172646 215509
rect 172882 215273 172924 215509
rect 172604 215241 172924 215273
rect 187293 215829 187613 215861
rect 187293 215593 187335 215829
rect 187571 215593 187613 215829
rect 187293 215509 187613 215593
rect 187293 215273 187335 215509
rect 187571 215273 187613 215509
rect 187293 215241 187613 215273
rect 191991 215829 192311 215861
rect 191991 215593 192033 215829
rect 192269 215593 192311 215829
rect 191991 215509 192311 215593
rect 191991 215273 192033 215509
rect 192269 215273 192311 215509
rect 191991 215241 192311 215273
rect 135208 212454 135528 212486
rect 135208 212218 135250 212454
rect 135486 212218 135528 212454
rect 135208 212134 135528 212218
rect 135208 211898 135250 212134
rect 135486 211898 135528 212134
rect 135208 211866 135528 211898
rect 141472 212454 141792 212486
rect 141472 212218 141514 212454
rect 141750 212218 141792 212454
rect 141472 212134 141792 212218
rect 141472 211898 141514 212134
rect 141750 211898 141792 212134
rect 141472 211866 141792 211898
rect 163208 212454 163528 212486
rect 163208 212218 163250 212454
rect 163486 212218 163528 212454
rect 163208 212134 163528 212218
rect 163208 211898 163250 212134
rect 163486 211898 163528 212134
rect 163208 211866 163528 211898
rect 169472 212454 169792 212486
rect 169472 212218 169514 212454
rect 169750 212218 169792 212454
rect 169472 212134 169792 212218
rect 169472 211898 169514 212134
rect 169750 211898 169792 212134
rect 169472 211866 169792 211898
rect 189642 212454 189962 212486
rect 189642 212218 189684 212454
rect 189920 212218 189962 212454
rect 189642 212134 189962 212218
rect 189642 211898 189684 212134
rect 189920 211898 189962 212134
rect 189642 211866 189962 211898
rect 194340 212454 194660 212486
rect 194340 212218 194382 212454
rect 194618 212218 194660 212454
rect 194340 212134 194660 212218
rect 194340 211898 194382 212134
rect 194618 211898 194660 212134
rect 194340 211866 194660 211898
rect 194734 202877 194794 225251
rect 288387 224364 288453 224365
rect 288387 224300 288388 224364
rect 288452 224300 288453 224364
rect 288387 224299 288453 224300
rect 260419 224228 260485 224229
rect 260419 224164 260420 224228
rect 260484 224164 260485 224228
rect 260419 224163 260485 224164
rect 260422 216341 260482 224163
rect 288390 216341 288450 224299
rect 492627 224228 492693 224229
rect 492627 224164 492628 224228
rect 492692 224164 492693 224228
rect 492627 224163 492693 224164
rect 492630 216341 492690 224163
rect 520595 224092 520661 224093
rect 520595 224028 520596 224092
rect 520660 224028 520661 224092
rect 520595 224027 520661 224028
rect 520598 216341 520658 224027
rect 260419 216340 260485 216341
rect 260419 216276 260420 216340
rect 260484 216276 260485 216340
rect 260419 216275 260485 216276
rect 288387 216340 288453 216341
rect 288387 216276 288388 216340
rect 288452 216276 288453 216340
rect 288387 216275 288453 216276
rect 492627 216340 492693 216341
rect 492627 216276 492628 216340
rect 492692 216276 492693 216340
rect 492627 216275 492693 216276
rect 520595 216340 520661 216341
rect 520595 216276 520596 216340
rect 520660 216276 520661 216340
rect 520595 216275 520661 216276
rect 196689 215829 197009 215861
rect 196689 215593 196731 215829
rect 196967 215593 197009 215829
rect 196689 215509 197009 215593
rect 196689 215273 196731 215509
rect 196967 215273 197009 215509
rect 196689 215241 197009 215273
rect 201387 215829 201707 215861
rect 201387 215593 201429 215829
rect 201665 215593 201707 215829
rect 201387 215509 201707 215593
rect 201387 215273 201429 215509
rect 201665 215273 201707 215509
rect 201387 215241 201707 215273
rect 215293 215829 215613 215861
rect 215293 215593 215335 215829
rect 215571 215593 215613 215829
rect 215293 215509 215613 215593
rect 215293 215273 215335 215509
rect 215571 215273 215613 215509
rect 215293 215241 215613 215273
rect 219991 215829 220311 215861
rect 219991 215593 220033 215829
rect 220269 215593 220311 215829
rect 219991 215509 220311 215593
rect 219991 215273 220033 215509
rect 220269 215273 220311 215509
rect 219991 215241 220311 215273
rect 224689 215829 225009 215861
rect 224689 215593 224731 215829
rect 224967 215593 225009 215829
rect 224689 215509 225009 215593
rect 224689 215273 224731 215509
rect 224967 215273 225009 215509
rect 224689 215241 225009 215273
rect 229387 215829 229707 215861
rect 229387 215593 229429 215829
rect 229665 215593 229707 215829
rect 229387 215509 229707 215593
rect 229387 215273 229429 215509
rect 229665 215273 229707 215509
rect 229387 215241 229707 215273
rect 243293 215829 243613 215861
rect 243293 215593 243335 215829
rect 243571 215593 243613 215829
rect 243293 215509 243613 215593
rect 243293 215273 243335 215509
rect 243571 215273 243613 215509
rect 243293 215241 243613 215273
rect 247991 215829 248311 215861
rect 247991 215593 248033 215829
rect 248269 215593 248311 215829
rect 247991 215509 248311 215593
rect 247991 215273 248033 215509
rect 248269 215273 248311 215509
rect 247991 215241 248311 215273
rect 252689 215829 253009 215861
rect 252689 215593 252731 215829
rect 252967 215593 253009 215829
rect 252689 215509 253009 215593
rect 252689 215273 252731 215509
rect 252967 215273 253009 215509
rect 252689 215241 253009 215273
rect 257387 215829 257707 215861
rect 257387 215593 257429 215829
rect 257665 215593 257707 215829
rect 257387 215509 257707 215593
rect 257387 215273 257429 215509
rect 257665 215273 257707 215509
rect 257387 215241 257707 215273
rect 271293 215829 271613 215861
rect 271293 215593 271335 215829
rect 271571 215593 271613 215829
rect 271293 215509 271613 215593
rect 271293 215273 271335 215509
rect 271571 215273 271613 215509
rect 271293 215241 271613 215273
rect 275991 215829 276311 215861
rect 275991 215593 276033 215829
rect 276269 215593 276311 215829
rect 275991 215509 276311 215593
rect 275991 215273 276033 215509
rect 276269 215273 276311 215509
rect 275991 215241 276311 215273
rect 280689 215829 281009 215861
rect 280689 215593 280731 215829
rect 280967 215593 281009 215829
rect 280689 215509 281009 215593
rect 280689 215273 280731 215509
rect 280967 215273 281009 215509
rect 280689 215241 281009 215273
rect 285387 215829 285707 215861
rect 285387 215593 285429 215829
rect 285665 215593 285707 215829
rect 285387 215509 285707 215593
rect 285387 215273 285429 215509
rect 285665 215273 285707 215509
rect 285387 215241 285707 215273
rect 299293 215829 299613 215861
rect 299293 215593 299335 215829
rect 299571 215593 299613 215829
rect 299293 215509 299613 215593
rect 299293 215273 299335 215509
rect 299571 215273 299613 215509
rect 299293 215241 299613 215273
rect 303991 215829 304311 215861
rect 303991 215593 304033 215829
rect 304269 215593 304311 215829
rect 303991 215509 304311 215593
rect 303991 215273 304033 215509
rect 304269 215273 304311 215509
rect 303991 215241 304311 215273
rect 308689 215829 309009 215861
rect 308689 215593 308731 215829
rect 308967 215593 309009 215829
rect 308689 215509 309009 215593
rect 308689 215273 308731 215509
rect 308967 215273 309009 215509
rect 308689 215241 309009 215273
rect 313387 215829 313707 215861
rect 313387 215593 313429 215829
rect 313665 215593 313707 215829
rect 313387 215509 313707 215593
rect 313387 215273 313429 215509
rect 313665 215273 313707 215509
rect 313387 215241 313707 215273
rect 328076 215829 328396 215861
rect 328076 215593 328118 215829
rect 328354 215593 328396 215829
rect 328076 215509 328396 215593
rect 328076 215273 328118 215509
rect 328354 215273 328396 215509
rect 328076 215241 328396 215273
rect 334340 215829 334660 215861
rect 334340 215593 334382 215829
rect 334618 215593 334660 215829
rect 334340 215509 334660 215593
rect 334340 215273 334382 215509
rect 334618 215273 334660 215509
rect 334340 215241 334660 215273
rect 340604 215829 340924 215861
rect 340604 215593 340646 215829
rect 340882 215593 340924 215829
rect 340604 215509 340924 215593
rect 340604 215273 340646 215509
rect 340882 215273 340924 215509
rect 340604 215241 340924 215273
rect 355293 215829 355613 215861
rect 355293 215593 355335 215829
rect 355571 215593 355613 215829
rect 355293 215509 355613 215593
rect 355293 215273 355335 215509
rect 355571 215273 355613 215509
rect 355293 215241 355613 215273
rect 359991 215829 360311 215861
rect 359991 215593 360033 215829
rect 360269 215593 360311 215829
rect 359991 215509 360311 215593
rect 359991 215273 360033 215509
rect 360269 215273 360311 215509
rect 359991 215241 360311 215273
rect 364689 215829 365009 215861
rect 364689 215593 364731 215829
rect 364967 215593 365009 215829
rect 364689 215509 365009 215593
rect 364689 215273 364731 215509
rect 364967 215273 365009 215509
rect 364689 215241 365009 215273
rect 369387 215829 369707 215861
rect 369387 215593 369429 215829
rect 369665 215593 369707 215829
rect 369387 215509 369707 215593
rect 369387 215273 369429 215509
rect 369665 215273 369707 215509
rect 369387 215241 369707 215273
rect 383293 215829 383613 215861
rect 383293 215593 383335 215829
rect 383571 215593 383613 215829
rect 383293 215509 383613 215593
rect 383293 215273 383335 215509
rect 383571 215273 383613 215509
rect 383293 215241 383613 215273
rect 387991 215829 388311 215861
rect 387991 215593 388033 215829
rect 388269 215593 388311 215829
rect 387991 215509 388311 215593
rect 387991 215273 388033 215509
rect 388269 215273 388311 215509
rect 387991 215241 388311 215273
rect 392689 215829 393009 215861
rect 392689 215593 392731 215829
rect 392967 215593 393009 215829
rect 392689 215509 393009 215593
rect 392689 215273 392731 215509
rect 392967 215273 393009 215509
rect 392689 215241 393009 215273
rect 397387 215829 397707 215861
rect 397387 215593 397429 215829
rect 397665 215593 397707 215829
rect 397387 215509 397707 215593
rect 397387 215273 397429 215509
rect 397665 215273 397707 215509
rect 397387 215241 397707 215273
rect 411293 215829 411613 215861
rect 411293 215593 411335 215829
rect 411571 215593 411613 215829
rect 411293 215509 411613 215593
rect 411293 215273 411335 215509
rect 411571 215273 411613 215509
rect 411293 215241 411613 215273
rect 415991 215829 416311 215861
rect 415991 215593 416033 215829
rect 416269 215593 416311 215829
rect 415991 215509 416311 215593
rect 415991 215273 416033 215509
rect 416269 215273 416311 215509
rect 415991 215241 416311 215273
rect 420689 215829 421009 215861
rect 420689 215593 420731 215829
rect 420967 215593 421009 215829
rect 420689 215509 421009 215593
rect 420689 215273 420731 215509
rect 420967 215273 421009 215509
rect 420689 215241 421009 215273
rect 425387 215829 425707 215861
rect 425387 215593 425429 215829
rect 425665 215593 425707 215829
rect 425387 215509 425707 215593
rect 425387 215273 425429 215509
rect 425665 215273 425707 215509
rect 425387 215241 425707 215273
rect 439293 215829 439613 215861
rect 439293 215593 439335 215829
rect 439571 215593 439613 215829
rect 439293 215509 439613 215593
rect 439293 215273 439335 215509
rect 439571 215273 439613 215509
rect 439293 215241 439613 215273
rect 443991 215829 444311 215861
rect 443991 215593 444033 215829
rect 444269 215593 444311 215829
rect 443991 215509 444311 215593
rect 443991 215273 444033 215509
rect 444269 215273 444311 215509
rect 443991 215241 444311 215273
rect 448689 215829 449009 215861
rect 448689 215593 448731 215829
rect 448967 215593 449009 215829
rect 448689 215509 449009 215593
rect 448689 215273 448731 215509
rect 448967 215273 449009 215509
rect 448689 215241 449009 215273
rect 453387 215829 453707 215861
rect 453387 215593 453429 215829
rect 453665 215593 453707 215829
rect 453387 215509 453707 215593
rect 453387 215273 453429 215509
rect 453665 215273 453707 215509
rect 453387 215241 453707 215273
rect 467293 215829 467613 215861
rect 467293 215593 467335 215829
rect 467571 215593 467613 215829
rect 467293 215509 467613 215593
rect 467293 215273 467335 215509
rect 467571 215273 467613 215509
rect 467293 215241 467613 215273
rect 471991 215829 472311 215861
rect 471991 215593 472033 215829
rect 472269 215593 472311 215829
rect 471991 215509 472311 215593
rect 471991 215273 472033 215509
rect 472269 215273 472311 215509
rect 471991 215241 472311 215273
rect 476689 215829 477009 215861
rect 476689 215593 476731 215829
rect 476967 215593 477009 215829
rect 476689 215509 477009 215593
rect 476689 215273 476731 215509
rect 476967 215273 477009 215509
rect 476689 215241 477009 215273
rect 481387 215829 481707 215861
rect 481387 215593 481429 215829
rect 481665 215593 481707 215829
rect 481387 215509 481707 215593
rect 481387 215273 481429 215509
rect 481665 215273 481707 215509
rect 481387 215241 481707 215273
rect 495293 215829 495613 215861
rect 495293 215593 495335 215829
rect 495571 215593 495613 215829
rect 495293 215509 495613 215593
rect 495293 215273 495335 215509
rect 495571 215273 495613 215509
rect 495293 215241 495613 215273
rect 499991 215829 500311 215861
rect 499991 215593 500033 215829
rect 500269 215593 500311 215829
rect 499991 215509 500311 215593
rect 499991 215273 500033 215509
rect 500269 215273 500311 215509
rect 499991 215241 500311 215273
rect 504689 215829 505009 215861
rect 504689 215593 504731 215829
rect 504967 215593 505009 215829
rect 504689 215509 505009 215593
rect 504689 215273 504731 215509
rect 504967 215273 505009 215509
rect 504689 215241 505009 215273
rect 509387 215829 509707 215861
rect 509387 215593 509429 215829
rect 509665 215593 509707 215829
rect 509387 215509 509707 215593
rect 509387 215273 509429 215509
rect 509665 215273 509707 215509
rect 509387 215241 509707 215273
rect 523293 215829 523613 215861
rect 523293 215593 523335 215829
rect 523571 215593 523613 215829
rect 523293 215509 523613 215593
rect 523293 215273 523335 215509
rect 523571 215273 523613 215509
rect 523293 215241 523613 215273
rect 527991 215829 528311 215861
rect 527991 215593 528033 215829
rect 528269 215593 528311 215829
rect 527991 215509 528311 215593
rect 527991 215273 528033 215509
rect 528269 215273 528311 215509
rect 527991 215241 528311 215273
rect 532689 215829 533009 215861
rect 532689 215593 532731 215829
rect 532967 215593 533009 215829
rect 532689 215509 533009 215593
rect 532689 215273 532731 215509
rect 532967 215273 533009 215509
rect 532689 215241 533009 215273
rect 537387 215829 537707 215861
rect 537387 215593 537429 215829
rect 537665 215593 537707 215829
rect 537387 215509 537707 215593
rect 537387 215273 537429 215509
rect 537665 215273 537707 215509
rect 537387 215241 537707 215273
rect 551293 215829 551613 215861
rect 551293 215593 551335 215829
rect 551571 215593 551613 215829
rect 551293 215509 551613 215593
rect 551293 215273 551335 215509
rect 551571 215273 551613 215509
rect 551293 215241 551613 215273
rect 555991 215829 556311 215861
rect 555991 215593 556033 215829
rect 556269 215593 556311 215829
rect 555991 215509 556311 215593
rect 555991 215273 556033 215509
rect 556269 215273 556311 215509
rect 555991 215241 556311 215273
rect 560689 215829 561009 215861
rect 560689 215593 560731 215829
rect 560967 215593 561009 215829
rect 560689 215509 561009 215593
rect 560689 215273 560731 215509
rect 560967 215273 561009 215509
rect 560689 215241 561009 215273
rect 565387 215829 565707 215861
rect 565387 215593 565429 215829
rect 565665 215593 565707 215829
rect 565387 215509 565707 215593
rect 565387 215273 565429 215509
rect 565665 215273 565707 215509
rect 565387 215241 565707 215273
rect 573494 215829 574114 242273
rect 573494 215593 573526 215829
rect 573762 215593 573846 215829
rect 574082 215593 574114 215829
rect 573494 215509 574114 215593
rect 573494 215273 573526 215509
rect 573762 215273 573846 215509
rect 574082 215273 574114 215509
rect 199038 212454 199358 212486
rect 199038 212218 199080 212454
rect 199316 212218 199358 212454
rect 199038 212134 199358 212218
rect 199038 211898 199080 212134
rect 199316 211898 199358 212134
rect 199038 211866 199358 211898
rect 217642 212454 217962 212486
rect 217642 212218 217684 212454
rect 217920 212218 217962 212454
rect 217642 212134 217962 212218
rect 217642 211898 217684 212134
rect 217920 211898 217962 212134
rect 217642 211866 217962 211898
rect 222340 212454 222660 212486
rect 222340 212218 222382 212454
rect 222618 212218 222660 212454
rect 222340 212134 222660 212218
rect 222340 211898 222382 212134
rect 222618 211898 222660 212134
rect 222340 211866 222660 211898
rect 227038 212454 227358 212486
rect 227038 212218 227080 212454
rect 227316 212218 227358 212454
rect 227038 212134 227358 212218
rect 227038 211898 227080 212134
rect 227316 211898 227358 212134
rect 227038 211866 227358 211898
rect 245642 212454 245962 212486
rect 245642 212218 245684 212454
rect 245920 212218 245962 212454
rect 245642 212134 245962 212218
rect 245642 211898 245684 212134
rect 245920 211898 245962 212134
rect 245642 211866 245962 211898
rect 250340 212454 250660 212486
rect 250340 212218 250382 212454
rect 250618 212218 250660 212454
rect 250340 212134 250660 212218
rect 250340 211898 250382 212134
rect 250618 211898 250660 212134
rect 250340 211866 250660 211898
rect 255038 212454 255358 212486
rect 255038 212218 255080 212454
rect 255316 212218 255358 212454
rect 255038 212134 255358 212218
rect 255038 211898 255080 212134
rect 255316 211898 255358 212134
rect 255038 211866 255358 211898
rect 273642 212454 273962 212486
rect 273642 212218 273684 212454
rect 273920 212218 273962 212454
rect 273642 212134 273962 212218
rect 273642 211898 273684 212134
rect 273920 211898 273962 212134
rect 273642 211866 273962 211898
rect 278340 212454 278660 212486
rect 278340 212218 278382 212454
rect 278618 212218 278660 212454
rect 278340 212134 278660 212218
rect 278340 211898 278382 212134
rect 278618 211898 278660 212134
rect 278340 211866 278660 211898
rect 283038 212454 283358 212486
rect 283038 212218 283080 212454
rect 283316 212218 283358 212454
rect 283038 212134 283358 212218
rect 283038 211898 283080 212134
rect 283316 211898 283358 212134
rect 283038 211866 283358 211898
rect 301642 212454 301962 212486
rect 301642 212218 301684 212454
rect 301920 212218 301962 212454
rect 301642 212134 301962 212218
rect 301642 211898 301684 212134
rect 301920 211898 301962 212134
rect 301642 211866 301962 211898
rect 306340 212454 306660 212486
rect 306340 212218 306382 212454
rect 306618 212218 306660 212454
rect 306340 212134 306660 212218
rect 306340 211898 306382 212134
rect 306618 211898 306660 212134
rect 306340 211866 306660 211898
rect 311038 212454 311358 212486
rect 311038 212218 311080 212454
rect 311316 212218 311358 212454
rect 311038 212134 311358 212218
rect 311038 211898 311080 212134
rect 311316 211898 311358 212134
rect 311038 211866 311358 211898
rect 331208 212454 331528 212486
rect 331208 212218 331250 212454
rect 331486 212218 331528 212454
rect 331208 212134 331528 212218
rect 331208 211898 331250 212134
rect 331486 211898 331528 212134
rect 331208 211866 331528 211898
rect 337472 212454 337792 212486
rect 337472 212218 337514 212454
rect 337750 212218 337792 212454
rect 337472 212134 337792 212218
rect 337472 211898 337514 212134
rect 337750 211898 337792 212134
rect 337472 211866 337792 211898
rect 357642 212454 357962 212486
rect 357642 212218 357684 212454
rect 357920 212218 357962 212454
rect 357642 212134 357962 212218
rect 357642 211898 357684 212134
rect 357920 211898 357962 212134
rect 357642 211866 357962 211898
rect 362340 212454 362660 212486
rect 362340 212218 362382 212454
rect 362618 212218 362660 212454
rect 362340 212134 362660 212218
rect 362340 211898 362382 212134
rect 362618 211898 362660 212134
rect 362340 211866 362660 211898
rect 367038 212454 367358 212486
rect 367038 212218 367080 212454
rect 367316 212218 367358 212454
rect 367038 212134 367358 212218
rect 367038 211898 367080 212134
rect 367316 211898 367358 212134
rect 367038 211866 367358 211898
rect 385642 212454 385962 212486
rect 385642 212218 385684 212454
rect 385920 212218 385962 212454
rect 385642 212134 385962 212218
rect 385642 211898 385684 212134
rect 385920 211898 385962 212134
rect 385642 211866 385962 211898
rect 390340 212454 390660 212486
rect 390340 212218 390382 212454
rect 390618 212218 390660 212454
rect 390340 212134 390660 212218
rect 390340 211898 390382 212134
rect 390618 211898 390660 212134
rect 390340 211866 390660 211898
rect 395038 212454 395358 212486
rect 395038 212218 395080 212454
rect 395316 212218 395358 212454
rect 395038 212134 395358 212218
rect 395038 211898 395080 212134
rect 395316 211898 395358 212134
rect 395038 211866 395358 211898
rect 413642 212454 413962 212486
rect 413642 212218 413684 212454
rect 413920 212218 413962 212454
rect 413642 212134 413962 212218
rect 413642 211898 413684 212134
rect 413920 211898 413962 212134
rect 413642 211866 413962 211898
rect 418340 212454 418660 212486
rect 418340 212218 418382 212454
rect 418618 212218 418660 212454
rect 418340 212134 418660 212218
rect 418340 211898 418382 212134
rect 418618 211898 418660 212134
rect 418340 211866 418660 211898
rect 423038 212454 423358 212486
rect 423038 212218 423080 212454
rect 423316 212218 423358 212454
rect 423038 212134 423358 212218
rect 423038 211898 423080 212134
rect 423316 211898 423358 212134
rect 423038 211866 423358 211898
rect 441642 212454 441962 212486
rect 441642 212218 441684 212454
rect 441920 212218 441962 212454
rect 441642 212134 441962 212218
rect 441642 211898 441684 212134
rect 441920 211898 441962 212134
rect 441642 211866 441962 211898
rect 446340 212454 446660 212486
rect 446340 212218 446382 212454
rect 446618 212218 446660 212454
rect 446340 212134 446660 212218
rect 446340 211898 446382 212134
rect 446618 211898 446660 212134
rect 446340 211866 446660 211898
rect 451038 212454 451358 212486
rect 451038 212218 451080 212454
rect 451316 212218 451358 212454
rect 451038 212134 451358 212218
rect 451038 211898 451080 212134
rect 451316 211898 451358 212134
rect 451038 211866 451358 211898
rect 469642 212454 469962 212486
rect 469642 212218 469684 212454
rect 469920 212218 469962 212454
rect 469642 212134 469962 212218
rect 469642 211898 469684 212134
rect 469920 211898 469962 212134
rect 469642 211866 469962 211898
rect 474340 212454 474660 212486
rect 474340 212218 474382 212454
rect 474618 212218 474660 212454
rect 474340 212134 474660 212218
rect 474340 211898 474382 212134
rect 474618 211898 474660 212134
rect 474340 211866 474660 211898
rect 479038 212454 479358 212486
rect 479038 212218 479080 212454
rect 479316 212218 479358 212454
rect 479038 212134 479358 212218
rect 479038 211898 479080 212134
rect 479316 211898 479358 212134
rect 479038 211866 479358 211898
rect 497642 212454 497962 212486
rect 497642 212218 497684 212454
rect 497920 212218 497962 212454
rect 497642 212134 497962 212218
rect 497642 211898 497684 212134
rect 497920 211898 497962 212134
rect 497642 211866 497962 211898
rect 502340 212454 502660 212486
rect 502340 212218 502382 212454
rect 502618 212218 502660 212454
rect 502340 212134 502660 212218
rect 502340 211898 502382 212134
rect 502618 211898 502660 212134
rect 502340 211866 502660 211898
rect 507038 212454 507358 212486
rect 507038 212218 507080 212454
rect 507316 212218 507358 212454
rect 507038 212134 507358 212218
rect 507038 211898 507080 212134
rect 507316 211898 507358 212134
rect 507038 211866 507358 211898
rect 525642 212454 525962 212486
rect 525642 212218 525684 212454
rect 525920 212218 525962 212454
rect 525642 212134 525962 212218
rect 525642 211898 525684 212134
rect 525920 211898 525962 212134
rect 525642 211866 525962 211898
rect 530340 212454 530660 212486
rect 530340 212218 530382 212454
rect 530618 212218 530660 212454
rect 530340 212134 530660 212218
rect 530340 211898 530382 212134
rect 530618 211898 530660 212134
rect 530340 211866 530660 211898
rect 535038 212454 535358 212486
rect 535038 212218 535080 212454
rect 535316 212218 535358 212454
rect 535038 212134 535358 212218
rect 535038 211898 535080 212134
rect 535316 211898 535358 212134
rect 535038 211866 535358 211898
rect 553642 212454 553962 212486
rect 553642 212218 553684 212454
rect 553920 212218 553962 212454
rect 553642 212134 553962 212218
rect 553642 211898 553684 212134
rect 553920 211898 553962 212134
rect 553642 211866 553962 211898
rect 558340 212454 558660 212486
rect 558340 212218 558382 212454
rect 558618 212218 558660 212454
rect 558340 212134 558660 212218
rect 558340 211898 558382 212134
rect 558618 211898 558660 212134
rect 558340 211866 558660 211898
rect 563038 212454 563358 212486
rect 563038 212218 563080 212454
rect 563316 212218 563358 212454
rect 563038 212134 563358 212218
rect 563038 211898 563080 212134
rect 563316 211898 563358 212134
rect 563038 211866 563358 211898
rect 128307 202876 128373 202877
rect 128307 202812 128308 202876
rect 128372 202812 128373 202876
rect 128307 202811 128373 202812
rect 194731 202876 194797 202877
rect 194731 202812 194732 202876
rect 194796 202812 194797 202876
rect 194731 202811 194797 202812
rect 63723 201516 63789 201517
rect 63723 201452 63724 201516
rect 63788 201452 63789 201516
rect 63723 201451 63789 201452
rect -2006 188593 -1974 188829
rect -1738 188593 -1654 188829
rect -1418 188593 -1386 188829
rect -2006 188509 -1386 188593
rect -2006 188273 -1974 188509
rect -1738 188273 -1654 188509
rect -1418 188273 -1386 188509
rect -2006 161829 -1386 188273
rect 19293 188829 19613 188861
rect 19293 188593 19335 188829
rect 19571 188593 19613 188829
rect 19293 188509 19613 188593
rect 19293 188273 19335 188509
rect 19571 188273 19613 188509
rect 19293 188241 19613 188273
rect 23991 188829 24311 188861
rect 23991 188593 24033 188829
rect 24269 188593 24311 188829
rect 23991 188509 24311 188593
rect 23991 188273 24033 188509
rect 24269 188273 24311 188509
rect 23991 188241 24311 188273
rect 28689 188829 29009 188861
rect 28689 188593 28731 188829
rect 28967 188593 29009 188829
rect 28689 188509 29009 188593
rect 28689 188273 28731 188509
rect 28967 188273 29009 188509
rect 28689 188241 29009 188273
rect 33387 188829 33707 188861
rect 33387 188593 33429 188829
rect 33665 188593 33707 188829
rect 33387 188509 33707 188593
rect 33387 188273 33429 188509
rect 33665 188273 33707 188509
rect 33387 188241 33707 188273
rect 47293 188829 47613 188861
rect 47293 188593 47335 188829
rect 47571 188593 47613 188829
rect 47293 188509 47613 188593
rect 47293 188273 47335 188509
rect 47571 188273 47613 188509
rect 47293 188241 47613 188273
rect 51991 188829 52311 188861
rect 51991 188593 52033 188829
rect 52269 188593 52311 188829
rect 51991 188509 52311 188593
rect 51991 188273 52033 188509
rect 52269 188273 52311 188509
rect 51991 188241 52311 188273
rect 56689 188829 57009 188861
rect 56689 188593 56731 188829
rect 56967 188593 57009 188829
rect 56689 188509 57009 188593
rect 56689 188273 56731 188509
rect 56967 188273 57009 188509
rect 56689 188241 57009 188273
rect 61387 188829 61707 188861
rect 61387 188593 61429 188829
rect 61665 188593 61707 188829
rect 61387 188509 61707 188593
rect 61387 188273 61429 188509
rect 61665 188273 61707 188509
rect 61387 188241 61707 188273
rect 21642 185454 21962 185486
rect 21642 185218 21684 185454
rect 21920 185218 21962 185454
rect 21642 185134 21962 185218
rect 21642 184898 21684 185134
rect 21920 184898 21962 185134
rect 21642 184866 21962 184898
rect 26340 185454 26660 185486
rect 26340 185218 26382 185454
rect 26618 185218 26660 185454
rect 26340 185134 26660 185218
rect 26340 184898 26382 185134
rect 26618 184898 26660 185134
rect 26340 184866 26660 184898
rect 31038 185454 31358 185486
rect 31038 185218 31080 185454
rect 31316 185218 31358 185454
rect 31038 185134 31358 185218
rect 31038 184898 31080 185134
rect 31316 184898 31358 185134
rect 31038 184866 31358 184898
rect 49642 185454 49962 185486
rect 49642 185218 49684 185454
rect 49920 185218 49962 185454
rect 49642 185134 49962 185218
rect 49642 184898 49684 185134
rect 49920 184898 49962 185134
rect 49642 184866 49962 184898
rect 54340 185454 54660 185486
rect 54340 185218 54382 185454
rect 54618 185218 54660 185454
rect 54340 185134 54660 185218
rect 54340 184898 54382 185134
rect 54618 184898 54660 185134
rect 54340 184866 54660 184898
rect 59038 185454 59358 185486
rect 59038 185218 59080 185454
rect 59316 185218 59358 185454
rect 59038 185134 59358 185218
rect 59038 184898 59080 185134
rect 59316 184898 59358 185134
rect 59038 184866 59358 184898
rect -2006 161593 -1974 161829
rect -1738 161593 -1654 161829
rect -1418 161593 -1386 161829
rect -2006 161509 -1386 161593
rect -2006 161273 -1974 161509
rect -1738 161273 -1654 161509
rect -1418 161273 -1386 161509
rect -2006 134829 -1386 161273
rect 19293 161829 19613 161861
rect 19293 161593 19335 161829
rect 19571 161593 19613 161829
rect 19293 161509 19613 161593
rect 19293 161273 19335 161509
rect 19571 161273 19613 161509
rect 19293 161241 19613 161273
rect 23991 161829 24311 161861
rect 23991 161593 24033 161829
rect 24269 161593 24311 161829
rect 23991 161509 24311 161593
rect 23991 161273 24033 161509
rect 24269 161273 24311 161509
rect 23991 161241 24311 161273
rect 28689 161829 29009 161861
rect 28689 161593 28731 161829
rect 28967 161593 29009 161829
rect 28689 161509 29009 161593
rect 28689 161273 28731 161509
rect 28967 161273 29009 161509
rect 28689 161241 29009 161273
rect 33387 161829 33707 161861
rect 33387 161593 33429 161829
rect 33665 161593 33707 161829
rect 33387 161509 33707 161593
rect 33387 161273 33429 161509
rect 33665 161273 33707 161509
rect 33387 161241 33707 161273
rect 47293 161829 47613 161861
rect 47293 161593 47335 161829
rect 47571 161593 47613 161829
rect 47293 161509 47613 161593
rect 47293 161273 47335 161509
rect 47571 161273 47613 161509
rect 47293 161241 47613 161273
rect 51991 161829 52311 161861
rect 51991 161593 52033 161829
rect 52269 161593 52311 161829
rect 51991 161509 52311 161593
rect 51991 161273 52033 161509
rect 52269 161273 52311 161509
rect 51991 161241 52311 161273
rect 56689 161829 57009 161861
rect 56689 161593 56731 161829
rect 56967 161593 57009 161829
rect 56689 161509 57009 161593
rect 56689 161273 56731 161509
rect 56967 161273 57009 161509
rect 56689 161241 57009 161273
rect 61387 161829 61707 161861
rect 61387 161593 61429 161829
rect 61665 161593 61707 161829
rect 61387 161509 61707 161593
rect 61387 161273 61429 161509
rect 61665 161273 61707 161509
rect 61387 161241 61707 161273
rect 21642 158454 21962 158486
rect 21642 158218 21684 158454
rect 21920 158218 21962 158454
rect 21642 158134 21962 158218
rect 21642 157898 21684 158134
rect 21920 157898 21962 158134
rect 21642 157866 21962 157898
rect 26340 158454 26660 158486
rect 26340 158218 26382 158454
rect 26618 158218 26660 158454
rect 26340 158134 26660 158218
rect 26340 157898 26382 158134
rect 26618 157898 26660 158134
rect 26340 157866 26660 157898
rect 31038 158454 31358 158486
rect 31038 158218 31080 158454
rect 31316 158218 31358 158454
rect 31038 158134 31358 158218
rect 31038 157898 31080 158134
rect 31316 157898 31358 158134
rect 31038 157866 31358 157898
rect 49642 158454 49962 158486
rect 49642 158218 49684 158454
rect 49920 158218 49962 158454
rect 49642 158134 49962 158218
rect 49642 157898 49684 158134
rect 49920 157898 49962 158134
rect 49642 157866 49962 157898
rect 54340 158454 54660 158486
rect 54340 158218 54382 158454
rect 54618 158218 54660 158454
rect 54340 158134 54660 158218
rect 54340 157898 54382 158134
rect 54618 157898 54660 158134
rect 54340 157866 54660 157898
rect 59038 158454 59358 158486
rect 59038 158218 59080 158454
rect 59316 158218 59358 158454
rect 59038 158134 59358 158218
rect 59038 157898 59080 158134
rect 59316 157898 59358 158134
rect 59038 157866 59358 157898
rect -2006 134593 -1974 134829
rect -1738 134593 -1654 134829
rect -1418 134593 -1386 134829
rect -2006 134509 -1386 134593
rect -2006 134273 -1974 134509
rect -1738 134273 -1654 134509
rect -1418 134273 -1386 134509
rect -2006 107829 -1386 134273
rect 19293 134829 19613 134861
rect 19293 134593 19335 134829
rect 19571 134593 19613 134829
rect 19293 134509 19613 134593
rect 19293 134273 19335 134509
rect 19571 134273 19613 134509
rect 19293 134241 19613 134273
rect 23991 134829 24311 134861
rect 23991 134593 24033 134829
rect 24269 134593 24311 134829
rect 23991 134509 24311 134593
rect 23991 134273 24033 134509
rect 24269 134273 24311 134509
rect 23991 134241 24311 134273
rect 28689 134829 29009 134861
rect 28689 134593 28731 134829
rect 28967 134593 29009 134829
rect 28689 134509 29009 134593
rect 28689 134273 28731 134509
rect 28967 134273 29009 134509
rect 28689 134241 29009 134273
rect 33387 134829 33707 134861
rect 33387 134593 33429 134829
rect 33665 134593 33707 134829
rect 33387 134509 33707 134593
rect 33387 134273 33429 134509
rect 33665 134273 33707 134509
rect 33387 134241 33707 134273
rect 47293 134829 47613 134861
rect 47293 134593 47335 134829
rect 47571 134593 47613 134829
rect 47293 134509 47613 134593
rect 47293 134273 47335 134509
rect 47571 134273 47613 134509
rect 47293 134241 47613 134273
rect 51991 134829 52311 134861
rect 51991 134593 52033 134829
rect 52269 134593 52311 134829
rect 51991 134509 52311 134593
rect 51991 134273 52033 134509
rect 52269 134273 52311 134509
rect 51991 134241 52311 134273
rect 56689 134829 57009 134861
rect 56689 134593 56731 134829
rect 56967 134593 57009 134829
rect 56689 134509 57009 134593
rect 56689 134273 56731 134509
rect 56967 134273 57009 134509
rect 56689 134241 57009 134273
rect 61387 134829 61707 134861
rect 61387 134593 61429 134829
rect 61665 134593 61707 134829
rect 61387 134509 61707 134593
rect 61387 134273 61429 134509
rect 61665 134273 61707 134509
rect 61387 134241 61707 134273
rect 21642 131454 21962 131486
rect 21642 131218 21684 131454
rect 21920 131218 21962 131454
rect 21642 131134 21962 131218
rect 21642 130898 21684 131134
rect 21920 130898 21962 131134
rect 21642 130866 21962 130898
rect 26340 131454 26660 131486
rect 26340 131218 26382 131454
rect 26618 131218 26660 131454
rect 26340 131134 26660 131218
rect 26340 130898 26382 131134
rect 26618 130898 26660 131134
rect 26340 130866 26660 130898
rect 31038 131454 31358 131486
rect 31038 131218 31080 131454
rect 31316 131218 31358 131454
rect 31038 131134 31358 131218
rect 31038 130898 31080 131134
rect 31316 130898 31358 131134
rect 31038 130866 31358 130898
rect 49642 131454 49962 131486
rect 49642 131218 49684 131454
rect 49920 131218 49962 131454
rect 49642 131134 49962 131218
rect 49642 130898 49684 131134
rect 49920 130898 49962 131134
rect 49642 130866 49962 130898
rect 54340 131454 54660 131486
rect 54340 131218 54382 131454
rect 54618 131218 54660 131454
rect 54340 131134 54660 131218
rect 54340 130898 54382 131134
rect 54618 130898 54660 131134
rect 54340 130866 54660 130898
rect 59038 131454 59358 131486
rect 59038 131218 59080 131454
rect 59316 131218 59358 131454
rect 59038 131134 59358 131218
rect 59038 130898 59080 131134
rect 59316 130898 59358 131134
rect 59038 130866 59358 130898
rect -2006 107593 -1974 107829
rect -1738 107593 -1654 107829
rect -1418 107593 -1386 107829
rect -2006 107509 -1386 107593
rect -2006 107273 -1974 107509
rect -1738 107273 -1654 107509
rect -1418 107273 -1386 107509
rect -2006 80829 -1386 107273
rect 19293 107829 19613 107861
rect 19293 107593 19335 107829
rect 19571 107593 19613 107829
rect 19293 107509 19613 107593
rect 19293 107273 19335 107509
rect 19571 107273 19613 107509
rect 19293 107241 19613 107273
rect 23991 107829 24311 107861
rect 23991 107593 24033 107829
rect 24269 107593 24311 107829
rect 23991 107509 24311 107593
rect 23991 107273 24033 107509
rect 24269 107273 24311 107509
rect 23991 107241 24311 107273
rect 28689 107829 29009 107861
rect 28689 107593 28731 107829
rect 28967 107593 29009 107829
rect 28689 107509 29009 107593
rect 28689 107273 28731 107509
rect 28967 107273 29009 107509
rect 28689 107241 29009 107273
rect 33387 107829 33707 107861
rect 33387 107593 33429 107829
rect 33665 107593 33707 107829
rect 33387 107509 33707 107593
rect 33387 107273 33429 107509
rect 33665 107273 33707 107509
rect 33387 107241 33707 107273
rect 47293 107829 47613 107861
rect 47293 107593 47335 107829
rect 47571 107593 47613 107829
rect 47293 107509 47613 107593
rect 47293 107273 47335 107509
rect 47571 107273 47613 107509
rect 47293 107241 47613 107273
rect 51991 107829 52311 107861
rect 51991 107593 52033 107829
rect 52269 107593 52311 107829
rect 51991 107509 52311 107593
rect 51991 107273 52033 107509
rect 52269 107273 52311 107509
rect 51991 107241 52311 107273
rect 56689 107829 57009 107861
rect 56689 107593 56731 107829
rect 56967 107593 57009 107829
rect 56689 107509 57009 107593
rect 56689 107273 56731 107509
rect 56967 107273 57009 107509
rect 56689 107241 57009 107273
rect 61387 107829 61707 107861
rect 61387 107593 61429 107829
rect 61665 107593 61707 107829
rect 61387 107509 61707 107593
rect 61387 107273 61429 107509
rect 61665 107273 61707 107509
rect 61387 107241 61707 107273
rect 21642 104454 21962 104486
rect 21642 104218 21684 104454
rect 21920 104218 21962 104454
rect 21642 104134 21962 104218
rect 21642 103898 21684 104134
rect 21920 103898 21962 104134
rect 21642 103866 21962 103898
rect 26340 104454 26660 104486
rect 26340 104218 26382 104454
rect 26618 104218 26660 104454
rect 26340 104134 26660 104218
rect 26340 103898 26382 104134
rect 26618 103898 26660 104134
rect 26340 103866 26660 103898
rect 31038 104454 31358 104486
rect 31038 104218 31080 104454
rect 31316 104218 31358 104454
rect 31038 104134 31358 104218
rect 31038 103898 31080 104134
rect 31316 103898 31358 104134
rect 31038 103866 31358 103898
rect 49642 104454 49962 104486
rect 49642 104218 49684 104454
rect 49920 104218 49962 104454
rect 49642 104134 49962 104218
rect 49642 103898 49684 104134
rect 49920 103898 49962 104134
rect 49642 103866 49962 103898
rect 54340 104454 54660 104486
rect 54340 104218 54382 104454
rect 54618 104218 54660 104454
rect 54340 104134 54660 104218
rect 54340 103898 54382 104134
rect 54618 103898 54660 104134
rect 54340 103866 54660 103898
rect 59038 104454 59358 104486
rect 59038 104218 59080 104454
rect 59316 104218 59358 104454
rect 59038 104134 59358 104218
rect 59038 103898 59080 104134
rect 59316 103898 59358 104134
rect 59038 103866 59358 103898
rect 44587 88908 44653 88909
rect 44587 88844 44588 88908
rect 44652 88844 44653 88908
rect 44587 88843 44653 88844
rect 44590 80885 44650 88843
rect 44587 80884 44653 80885
rect -2006 80593 -1974 80829
rect -1738 80593 -1654 80829
rect -1418 80593 -1386 80829
rect -2006 80509 -1386 80593
rect -2006 80273 -1974 80509
rect -1738 80273 -1654 80509
rect -1418 80273 -1386 80509
rect -2006 53829 -1386 80273
rect 20076 80829 20396 80861
rect 20076 80593 20118 80829
rect 20354 80593 20396 80829
rect 20076 80509 20396 80593
rect 20076 80273 20118 80509
rect 20354 80273 20396 80509
rect 20076 80241 20396 80273
rect 26340 80829 26660 80861
rect 26340 80593 26382 80829
rect 26618 80593 26660 80829
rect 26340 80509 26660 80593
rect 26340 80273 26382 80509
rect 26618 80273 26660 80509
rect 26340 80241 26660 80273
rect 32604 80829 32924 80861
rect 32604 80593 32646 80829
rect 32882 80593 32924 80829
rect 44587 80820 44588 80884
rect 44652 80820 44653 80884
rect 44587 80819 44653 80820
rect 48076 80829 48396 80861
rect 32604 80509 32924 80593
rect 32604 80273 32646 80509
rect 32882 80273 32924 80509
rect 32604 80241 32924 80273
rect 48076 80593 48118 80829
rect 48354 80593 48396 80829
rect 48076 80509 48396 80593
rect 48076 80273 48118 80509
rect 48354 80273 48396 80509
rect 48076 80241 48396 80273
rect 54340 80829 54660 80861
rect 54340 80593 54382 80829
rect 54618 80593 54660 80829
rect 54340 80509 54660 80593
rect 54340 80273 54382 80509
rect 54618 80273 54660 80509
rect 54340 80241 54660 80273
rect 60604 80829 60924 80861
rect 60604 80593 60646 80829
rect 60882 80593 60924 80829
rect 60604 80509 60924 80593
rect 60604 80273 60646 80509
rect 60882 80273 60924 80509
rect 60604 80241 60924 80273
rect 23208 77454 23528 77486
rect 23208 77218 23250 77454
rect 23486 77218 23528 77454
rect 23208 77134 23528 77218
rect 23208 76898 23250 77134
rect 23486 76898 23528 77134
rect 23208 76866 23528 76898
rect 29472 77454 29792 77486
rect 29472 77218 29514 77454
rect 29750 77218 29792 77454
rect 29472 77134 29792 77218
rect 29472 76898 29514 77134
rect 29750 76898 29792 77134
rect 29472 76866 29792 76898
rect 51208 77454 51528 77486
rect 51208 77218 51250 77454
rect 51486 77218 51528 77454
rect 51208 77134 51528 77218
rect 51208 76898 51250 77134
rect 51486 76898 51528 77134
rect 51208 76866 51528 76898
rect 57472 77454 57792 77486
rect 57472 77218 57514 77454
rect 57750 77218 57792 77454
rect 57472 77134 57792 77218
rect 57472 76898 57514 77134
rect 57750 76898 57792 77134
rect 57472 76866 57792 76898
rect -2006 53593 -1974 53829
rect -1738 53593 -1654 53829
rect -1418 53593 -1386 53829
rect -2006 53509 -1386 53593
rect -2006 53273 -1974 53509
rect -1738 53273 -1654 53509
rect -1418 53273 -1386 53509
rect -2006 26829 -1386 53273
rect 20076 53829 20396 53861
rect 20076 53593 20118 53829
rect 20354 53593 20396 53829
rect 20076 53509 20396 53593
rect 20076 53273 20118 53509
rect 20354 53273 20396 53509
rect 20076 53241 20396 53273
rect 26340 53829 26660 53861
rect 26340 53593 26382 53829
rect 26618 53593 26660 53829
rect 26340 53509 26660 53593
rect 26340 53273 26382 53509
rect 26618 53273 26660 53509
rect 26340 53241 26660 53273
rect 32604 53829 32924 53861
rect 32604 53593 32646 53829
rect 32882 53593 32924 53829
rect 32604 53509 32924 53593
rect 32604 53273 32646 53509
rect 32882 53273 32924 53509
rect 32604 53241 32924 53273
rect 48076 53829 48396 53861
rect 48076 53593 48118 53829
rect 48354 53593 48396 53829
rect 48076 53509 48396 53593
rect 48076 53273 48118 53509
rect 48354 53273 48396 53509
rect 48076 53241 48396 53273
rect 54340 53829 54660 53861
rect 54340 53593 54382 53829
rect 54618 53593 54660 53829
rect 54340 53509 54660 53593
rect 54340 53273 54382 53509
rect 54618 53273 54660 53509
rect 54340 53241 54660 53273
rect 60604 53829 60924 53861
rect 60604 53593 60646 53829
rect 60882 53593 60924 53829
rect 60604 53509 60924 53593
rect 60604 53273 60646 53509
rect 60882 53273 60924 53509
rect 60604 53241 60924 53273
rect 23208 50454 23528 50486
rect 23208 50218 23250 50454
rect 23486 50218 23528 50454
rect 23208 50134 23528 50218
rect 23208 49898 23250 50134
rect 23486 49898 23528 50134
rect 23208 49866 23528 49898
rect 29472 50454 29792 50486
rect 29472 50218 29514 50454
rect 29750 50218 29792 50454
rect 29472 50134 29792 50218
rect 29472 49898 29514 50134
rect 29750 49898 29792 50134
rect 29472 49866 29792 49898
rect 51208 50454 51528 50486
rect 51208 50218 51250 50454
rect 51486 50218 51528 50454
rect 51208 50134 51528 50218
rect 51208 49898 51250 50134
rect 51486 49898 51528 50134
rect 51208 49866 51528 49898
rect 57472 50454 57792 50486
rect 57472 50218 57514 50454
rect 57750 50218 57792 50454
rect 57472 50134 57792 50218
rect 57472 49898 57514 50134
rect 57750 49898 57792 50134
rect 57472 49866 57792 49898
rect -2006 26593 -1974 26829
rect -1738 26593 -1654 26829
rect -1418 26593 -1386 26829
rect -2006 26509 -1386 26593
rect -2006 26273 -1974 26509
rect -1738 26273 -1654 26509
rect -1418 26273 -1386 26509
rect -2006 -346 -1386 26273
rect 22418 26829 22738 26861
rect 22418 26593 22460 26829
rect 22696 26593 22738 26829
rect 22418 26509 22738 26593
rect 22418 26273 22460 26509
rect 22696 26273 22738 26509
rect 22418 26241 22738 26273
rect 33366 26829 33686 26861
rect 33366 26593 33408 26829
rect 33644 26593 33686 26829
rect 33366 26509 33686 26593
rect 33366 26273 33408 26509
rect 33644 26273 33686 26509
rect 33366 26241 33686 26273
rect 44314 26829 44634 26861
rect 44314 26593 44356 26829
rect 44592 26593 44634 26829
rect 44314 26509 44634 26593
rect 44314 26273 44356 26509
rect 44592 26273 44634 26509
rect 44314 26241 44634 26273
rect 55262 26829 55582 26861
rect 55262 26593 55304 26829
rect 55540 26593 55582 26829
rect 55262 26509 55582 26593
rect 55262 26273 55304 26509
rect 55540 26273 55582 26509
rect 55262 26241 55582 26273
rect 27892 23454 28212 23486
rect 27892 23218 27934 23454
rect 28170 23218 28212 23454
rect 27892 23134 28212 23218
rect 27892 22898 27934 23134
rect 28170 22898 28212 23134
rect 27892 22866 28212 22898
rect 38840 23454 39160 23486
rect 38840 23218 38882 23454
rect 39118 23218 39160 23454
rect 38840 23134 39160 23218
rect 38840 22898 38882 23134
rect 39118 22898 39160 23134
rect 38840 22866 39160 22898
rect 49788 23454 50108 23486
rect 49788 23218 49830 23454
rect 50066 23218 50108 23454
rect 49788 23134 50108 23218
rect 49788 22898 49830 23134
rect 50066 22898 50108 23134
rect 49788 22866 50108 22898
rect 60736 23454 61056 23486
rect 60736 23218 60778 23454
rect 61014 23218 61056 23454
rect 60736 23134 61056 23218
rect 60736 22898 60778 23134
rect 61014 22898 61056 23134
rect 60736 22866 61056 22898
rect 63726 20229 63786 201451
rect 259499 198524 259565 198525
rect 259499 198460 259500 198524
rect 259564 198460 259565 198524
rect 259499 198459 259565 198460
rect 361619 198524 361685 198525
rect 361619 198460 361620 198524
rect 361684 198460 361685 198524
rect 361619 198459 361685 198460
rect 445707 198524 445773 198525
rect 445707 198460 445708 198524
rect 445772 198460 445773 198524
rect 445707 198459 445773 198460
rect 75293 188829 75613 188861
rect 75293 188593 75335 188829
rect 75571 188593 75613 188829
rect 75293 188509 75613 188593
rect 75293 188273 75335 188509
rect 75571 188273 75613 188509
rect 75293 188241 75613 188273
rect 79991 188829 80311 188861
rect 79991 188593 80033 188829
rect 80269 188593 80311 188829
rect 79991 188509 80311 188593
rect 79991 188273 80033 188509
rect 80269 188273 80311 188509
rect 79991 188241 80311 188273
rect 84689 188829 85009 188861
rect 84689 188593 84731 188829
rect 84967 188593 85009 188829
rect 84689 188509 85009 188593
rect 84689 188273 84731 188509
rect 84967 188273 85009 188509
rect 84689 188241 85009 188273
rect 89387 188829 89707 188861
rect 89387 188593 89429 188829
rect 89665 188593 89707 188829
rect 89387 188509 89707 188593
rect 89387 188273 89429 188509
rect 89665 188273 89707 188509
rect 89387 188241 89707 188273
rect 103293 188829 103613 188861
rect 103293 188593 103335 188829
rect 103571 188593 103613 188829
rect 103293 188509 103613 188593
rect 103293 188273 103335 188509
rect 103571 188273 103613 188509
rect 103293 188241 103613 188273
rect 107991 188829 108311 188861
rect 107991 188593 108033 188829
rect 108269 188593 108311 188829
rect 107991 188509 108311 188593
rect 107991 188273 108033 188509
rect 108269 188273 108311 188509
rect 107991 188241 108311 188273
rect 112689 188829 113009 188861
rect 112689 188593 112731 188829
rect 112967 188593 113009 188829
rect 112689 188509 113009 188593
rect 112689 188273 112731 188509
rect 112967 188273 113009 188509
rect 112689 188241 113009 188273
rect 117387 188829 117707 188861
rect 117387 188593 117429 188829
rect 117665 188593 117707 188829
rect 117387 188509 117707 188593
rect 117387 188273 117429 188509
rect 117665 188273 117707 188509
rect 117387 188241 117707 188273
rect 131293 188829 131613 188861
rect 131293 188593 131335 188829
rect 131571 188593 131613 188829
rect 131293 188509 131613 188593
rect 131293 188273 131335 188509
rect 131571 188273 131613 188509
rect 131293 188241 131613 188273
rect 135991 188829 136311 188861
rect 135991 188593 136033 188829
rect 136269 188593 136311 188829
rect 135991 188509 136311 188593
rect 135991 188273 136033 188509
rect 136269 188273 136311 188509
rect 135991 188241 136311 188273
rect 140689 188829 141009 188861
rect 140689 188593 140731 188829
rect 140967 188593 141009 188829
rect 140689 188509 141009 188593
rect 140689 188273 140731 188509
rect 140967 188273 141009 188509
rect 140689 188241 141009 188273
rect 145387 188829 145707 188861
rect 145387 188593 145429 188829
rect 145665 188593 145707 188829
rect 145387 188509 145707 188593
rect 145387 188273 145429 188509
rect 145665 188273 145707 188509
rect 145387 188241 145707 188273
rect 159293 188829 159613 188861
rect 159293 188593 159335 188829
rect 159571 188593 159613 188829
rect 159293 188509 159613 188593
rect 159293 188273 159335 188509
rect 159571 188273 159613 188509
rect 159293 188241 159613 188273
rect 163991 188829 164311 188861
rect 163991 188593 164033 188829
rect 164269 188593 164311 188829
rect 163991 188509 164311 188593
rect 163991 188273 164033 188509
rect 164269 188273 164311 188509
rect 163991 188241 164311 188273
rect 168689 188829 169009 188861
rect 168689 188593 168731 188829
rect 168967 188593 169009 188829
rect 168689 188509 169009 188593
rect 168689 188273 168731 188509
rect 168967 188273 169009 188509
rect 168689 188241 169009 188273
rect 173387 188829 173707 188861
rect 173387 188593 173429 188829
rect 173665 188593 173707 188829
rect 173387 188509 173707 188593
rect 173387 188273 173429 188509
rect 173665 188273 173707 188509
rect 173387 188241 173707 188273
rect 187293 188829 187613 188861
rect 187293 188593 187335 188829
rect 187571 188593 187613 188829
rect 187293 188509 187613 188593
rect 187293 188273 187335 188509
rect 187571 188273 187613 188509
rect 187293 188241 187613 188273
rect 191991 188829 192311 188861
rect 191991 188593 192033 188829
rect 192269 188593 192311 188829
rect 191991 188509 192311 188593
rect 191991 188273 192033 188509
rect 192269 188273 192311 188509
rect 191991 188241 192311 188273
rect 196689 188829 197009 188861
rect 196689 188593 196731 188829
rect 196967 188593 197009 188829
rect 196689 188509 197009 188593
rect 196689 188273 196731 188509
rect 196967 188273 197009 188509
rect 196689 188241 197009 188273
rect 201387 188829 201707 188861
rect 201387 188593 201429 188829
rect 201665 188593 201707 188829
rect 201387 188509 201707 188593
rect 201387 188273 201429 188509
rect 201665 188273 201707 188509
rect 201387 188241 201707 188273
rect 215293 188829 215613 188861
rect 215293 188593 215335 188829
rect 215571 188593 215613 188829
rect 215293 188509 215613 188593
rect 215293 188273 215335 188509
rect 215571 188273 215613 188509
rect 215293 188241 215613 188273
rect 219991 188829 220311 188861
rect 219991 188593 220033 188829
rect 220269 188593 220311 188829
rect 219991 188509 220311 188593
rect 219991 188273 220033 188509
rect 220269 188273 220311 188509
rect 219991 188241 220311 188273
rect 224689 188829 225009 188861
rect 224689 188593 224731 188829
rect 224967 188593 225009 188829
rect 224689 188509 225009 188593
rect 224689 188273 224731 188509
rect 224967 188273 225009 188509
rect 224689 188241 225009 188273
rect 229387 188829 229707 188861
rect 229387 188593 229429 188829
rect 229665 188593 229707 188829
rect 229387 188509 229707 188593
rect 229387 188273 229429 188509
rect 229665 188273 229707 188509
rect 229387 188241 229707 188273
rect 243293 188829 243613 188861
rect 243293 188593 243335 188829
rect 243571 188593 243613 188829
rect 243293 188509 243613 188593
rect 243293 188273 243335 188509
rect 243571 188273 243613 188509
rect 243293 188241 243613 188273
rect 247991 188829 248311 188861
rect 247991 188593 248033 188829
rect 248269 188593 248311 188829
rect 247991 188509 248311 188593
rect 247991 188273 248033 188509
rect 248269 188273 248311 188509
rect 247991 188241 248311 188273
rect 252689 188829 253009 188861
rect 252689 188593 252731 188829
rect 252967 188593 253009 188829
rect 252689 188509 253009 188593
rect 252689 188273 252731 188509
rect 252967 188273 253009 188509
rect 252689 188241 253009 188273
rect 257387 188829 257707 188861
rect 257387 188593 257429 188829
rect 257665 188593 257707 188829
rect 257387 188509 257707 188593
rect 257387 188273 257429 188509
rect 257665 188273 257707 188509
rect 257387 188241 257707 188273
rect 77642 185454 77962 185486
rect 77642 185218 77684 185454
rect 77920 185218 77962 185454
rect 77642 185134 77962 185218
rect 77642 184898 77684 185134
rect 77920 184898 77962 185134
rect 77642 184866 77962 184898
rect 82340 185454 82660 185486
rect 82340 185218 82382 185454
rect 82618 185218 82660 185454
rect 82340 185134 82660 185218
rect 82340 184898 82382 185134
rect 82618 184898 82660 185134
rect 82340 184866 82660 184898
rect 87038 185454 87358 185486
rect 87038 185218 87080 185454
rect 87316 185218 87358 185454
rect 87038 185134 87358 185218
rect 87038 184898 87080 185134
rect 87316 184898 87358 185134
rect 87038 184866 87358 184898
rect 105642 185454 105962 185486
rect 105642 185218 105684 185454
rect 105920 185218 105962 185454
rect 105642 185134 105962 185218
rect 105642 184898 105684 185134
rect 105920 184898 105962 185134
rect 105642 184866 105962 184898
rect 110340 185454 110660 185486
rect 110340 185218 110382 185454
rect 110618 185218 110660 185454
rect 110340 185134 110660 185218
rect 110340 184898 110382 185134
rect 110618 184898 110660 185134
rect 110340 184866 110660 184898
rect 115038 185454 115358 185486
rect 115038 185218 115080 185454
rect 115316 185218 115358 185454
rect 115038 185134 115358 185218
rect 115038 184898 115080 185134
rect 115316 184898 115358 185134
rect 115038 184866 115358 184898
rect 133642 185454 133962 185486
rect 133642 185218 133684 185454
rect 133920 185218 133962 185454
rect 133642 185134 133962 185218
rect 133642 184898 133684 185134
rect 133920 184898 133962 185134
rect 133642 184866 133962 184898
rect 138340 185454 138660 185486
rect 138340 185218 138382 185454
rect 138618 185218 138660 185454
rect 138340 185134 138660 185218
rect 138340 184898 138382 185134
rect 138618 184898 138660 185134
rect 138340 184866 138660 184898
rect 143038 185454 143358 185486
rect 143038 185218 143080 185454
rect 143316 185218 143358 185454
rect 143038 185134 143358 185218
rect 143038 184898 143080 185134
rect 143316 184898 143358 185134
rect 143038 184866 143358 184898
rect 161642 185454 161962 185486
rect 161642 185218 161684 185454
rect 161920 185218 161962 185454
rect 161642 185134 161962 185218
rect 161642 184898 161684 185134
rect 161920 184898 161962 185134
rect 161642 184866 161962 184898
rect 166340 185454 166660 185486
rect 166340 185218 166382 185454
rect 166618 185218 166660 185454
rect 166340 185134 166660 185218
rect 166340 184898 166382 185134
rect 166618 184898 166660 185134
rect 166340 184866 166660 184898
rect 171038 185454 171358 185486
rect 171038 185218 171080 185454
rect 171316 185218 171358 185454
rect 171038 185134 171358 185218
rect 171038 184898 171080 185134
rect 171316 184898 171358 185134
rect 171038 184866 171358 184898
rect 189642 185454 189962 185486
rect 189642 185218 189684 185454
rect 189920 185218 189962 185454
rect 189642 185134 189962 185218
rect 189642 184898 189684 185134
rect 189920 184898 189962 185134
rect 189642 184866 189962 184898
rect 194340 185454 194660 185486
rect 194340 185218 194382 185454
rect 194618 185218 194660 185454
rect 194340 185134 194660 185218
rect 194340 184898 194382 185134
rect 194618 184898 194660 185134
rect 194340 184866 194660 184898
rect 199038 185454 199358 185486
rect 199038 185218 199080 185454
rect 199316 185218 199358 185454
rect 199038 185134 199358 185218
rect 199038 184898 199080 185134
rect 199316 184898 199358 185134
rect 199038 184866 199358 184898
rect 217642 185454 217962 185486
rect 217642 185218 217684 185454
rect 217920 185218 217962 185454
rect 217642 185134 217962 185218
rect 217642 184898 217684 185134
rect 217920 184898 217962 185134
rect 217642 184866 217962 184898
rect 222340 185454 222660 185486
rect 222340 185218 222382 185454
rect 222618 185218 222660 185454
rect 222340 185134 222660 185218
rect 222340 184898 222382 185134
rect 222618 184898 222660 185134
rect 222340 184866 222660 184898
rect 227038 185454 227358 185486
rect 227038 185218 227080 185454
rect 227316 185218 227358 185454
rect 227038 185134 227358 185218
rect 227038 184898 227080 185134
rect 227316 184898 227358 185134
rect 227038 184866 227358 184898
rect 245642 185454 245962 185486
rect 245642 185218 245684 185454
rect 245920 185218 245962 185454
rect 245642 185134 245962 185218
rect 245642 184898 245684 185134
rect 245920 184898 245962 185134
rect 245642 184866 245962 184898
rect 250340 185454 250660 185486
rect 250340 185218 250382 185454
rect 250618 185218 250660 185454
rect 250340 185134 250660 185218
rect 250340 184898 250382 185134
rect 250618 184898 250660 185134
rect 250340 184866 250660 184898
rect 255038 185454 255358 185486
rect 255038 185218 255080 185454
rect 255316 185218 255358 185454
rect 255038 185134 255358 185218
rect 255038 184898 255080 185134
rect 255316 184898 255358 185134
rect 255038 184866 255358 184898
rect 259502 176629 259562 198459
rect 271293 188829 271613 188861
rect 271293 188593 271335 188829
rect 271571 188593 271613 188829
rect 271293 188509 271613 188593
rect 271293 188273 271335 188509
rect 271571 188273 271613 188509
rect 271293 188241 271613 188273
rect 275991 188829 276311 188861
rect 275991 188593 276033 188829
rect 276269 188593 276311 188829
rect 275991 188509 276311 188593
rect 275991 188273 276033 188509
rect 276269 188273 276311 188509
rect 275991 188241 276311 188273
rect 280689 188829 281009 188861
rect 280689 188593 280731 188829
rect 280967 188593 281009 188829
rect 280689 188509 281009 188593
rect 280689 188273 280731 188509
rect 280967 188273 281009 188509
rect 280689 188241 281009 188273
rect 285387 188829 285707 188861
rect 285387 188593 285429 188829
rect 285665 188593 285707 188829
rect 285387 188509 285707 188593
rect 285387 188273 285429 188509
rect 285665 188273 285707 188509
rect 285387 188241 285707 188273
rect 299293 188829 299613 188861
rect 299293 188593 299335 188829
rect 299571 188593 299613 188829
rect 299293 188509 299613 188593
rect 299293 188273 299335 188509
rect 299571 188273 299613 188509
rect 299293 188241 299613 188273
rect 303991 188829 304311 188861
rect 303991 188593 304033 188829
rect 304269 188593 304311 188829
rect 303991 188509 304311 188593
rect 303991 188273 304033 188509
rect 304269 188273 304311 188509
rect 303991 188241 304311 188273
rect 308689 188829 309009 188861
rect 308689 188593 308731 188829
rect 308967 188593 309009 188829
rect 308689 188509 309009 188593
rect 308689 188273 308731 188509
rect 308967 188273 309009 188509
rect 308689 188241 309009 188273
rect 313387 188829 313707 188861
rect 313387 188593 313429 188829
rect 313665 188593 313707 188829
rect 313387 188509 313707 188593
rect 313387 188273 313429 188509
rect 313665 188273 313707 188509
rect 313387 188241 313707 188273
rect 327293 188829 327613 188861
rect 327293 188593 327335 188829
rect 327571 188593 327613 188829
rect 327293 188509 327613 188593
rect 327293 188273 327335 188509
rect 327571 188273 327613 188509
rect 327293 188241 327613 188273
rect 331991 188829 332311 188861
rect 331991 188593 332033 188829
rect 332269 188593 332311 188829
rect 331991 188509 332311 188593
rect 331991 188273 332033 188509
rect 332269 188273 332311 188509
rect 331991 188241 332311 188273
rect 336689 188829 337009 188861
rect 336689 188593 336731 188829
rect 336967 188593 337009 188829
rect 336689 188509 337009 188593
rect 336689 188273 336731 188509
rect 336967 188273 337009 188509
rect 336689 188241 337009 188273
rect 341387 188829 341707 188861
rect 341387 188593 341429 188829
rect 341665 188593 341707 188829
rect 341387 188509 341707 188593
rect 341387 188273 341429 188509
rect 341665 188273 341707 188509
rect 341387 188241 341707 188273
rect 355293 188829 355613 188861
rect 355293 188593 355335 188829
rect 355571 188593 355613 188829
rect 355293 188509 355613 188593
rect 355293 188273 355335 188509
rect 355571 188273 355613 188509
rect 355293 188241 355613 188273
rect 359991 188829 360311 188861
rect 359991 188593 360033 188829
rect 360269 188593 360311 188829
rect 359991 188509 360311 188593
rect 359991 188273 360033 188509
rect 360269 188273 360311 188509
rect 359991 188241 360311 188273
rect 273642 185454 273962 185486
rect 273642 185218 273684 185454
rect 273920 185218 273962 185454
rect 273642 185134 273962 185218
rect 273642 184898 273684 185134
rect 273920 184898 273962 185134
rect 273642 184866 273962 184898
rect 278340 185454 278660 185486
rect 278340 185218 278382 185454
rect 278618 185218 278660 185454
rect 278340 185134 278660 185218
rect 278340 184898 278382 185134
rect 278618 184898 278660 185134
rect 278340 184866 278660 184898
rect 283038 185454 283358 185486
rect 283038 185218 283080 185454
rect 283316 185218 283358 185454
rect 283038 185134 283358 185218
rect 283038 184898 283080 185134
rect 283316 184898 283358 185134
rect 283038 184866 283358 184898
rect 301642 185454 301962 185486
rect 301642 185218 301684 185454
rect 301920 185218 301962 185454
rect 301642 185134 301962 185218
rect 301642 184898 301684 185134
rect 301920 184898 301962 185134
rect 301642 184866 301962 184898
rect 306340 185454 306660 185486
rect 306340 185218 306382 185454
rect 306618 185218 306660 185454
rect 306340 185134 306660 185218
rect 306340 184898 306382 185134
rect 306618 184898 306660 185134
rect 306340 184866 306660 184898
rect 311038 185454 311358 185486
rect 311038 185218 311080 185454
rect 311316 185218 311358 185454
rect 311038 185134 311358 185218
rect 311038 184898 311080 185134
rect 311316 184898 311358 185134
rect 311038 184866 311358 184898
rect 329642 185454 329962 185486
rect 329642 185218 329684 185454
rect 329920 185218 329962 185454
rect 329642 185134 329962 185218
rect 329642 184898 329684 185134
rect 329920 184898 329962 185134
rect 329642 184866 329962 184898
rect 334340 185454 334660 185486
rect 334340 185218 334382 185454
rect 334618 185218 334660 185454
rect 334340 185134 334660 185218
rect 334340 184898 334382 185134
rect 334618 184898 334660 185134
rect 334340 184866 334660 184898
rect 339038 185454 339358 185486
rect 339038 185218 339080 185454
rect 339316 185218 339358 185454
rect 339038 185134 339358 185218
rect 339038 184898 339080 185134
rect 339316 184898 339358 185134
rect 339038 184866 339358 184898
rect 357642 185454 357962 185486
rect 357642 185218 357684 185454
rect 357920 185218 357962 185454
rect 357642 185134 357962 185218
rect 357642 184898 357684 185134
rect 357920 184898 357962 185134
rect 357642 184866 357962 184898
rect 361622 176629 361682 198459
rect 364689 188829 365009 188861
rect 364689 188593 364731 188829
rect 364967 188593 365009 188829
rect 364689 188509 365009 188593
rect 364689 188273 364731 188509
rect 364967 188273 365009 188509
rect 364689 188241 365009 188273
rect 369387 188829 369707 188861
rect 369387 188593 369429 188829
rect 369665 188593 369707 188829
rect 369387 188509 369707 188593
rect 369387 188273 369429 188509
rect 369665 188273 369707 188509
rect 369387 188241 369707 188273
rect 383293 188829 383613 188861
rect 383293 188593 383335 188829
rect 383571 188593 383613 188829
rect 383293 188509 383613 188593
rect 383293 188273 383335 188509
rect 383571 188273 383613 188509
rect 383293 188241 383613 188273
rect 387991 188829 388311 188861
rect 387991 188593 388033 188829
rect 388269 188593 388311 188829
rect 387991 188509 388311 188593
rect 387991 188273 388033 188509
rect 388269 188273 388311 188509
rect 387991 188241 388311 188273
rect 392689 188829 393009 188861
rect 392689 188593 392731 188829
rect 392967 188593 393009 188829
rect 392689 188509 393009 188593
rect 392689 188273 392731 188509
rect 392967 188273 393009 188509
rect 392689 188241 393009 188273
rect 397387 188829 397707 188861
rect 397387 188593 397429 188829
rect 397665 188593 397707 188829
rect 397387 188509 397707 188593
rect 397387 188273 397429 188509
rect 397665 188273 397707 188509
rect 397387 188241 397707 188273
rect 411293 188829 411613 188861
rect 411293 188593 411335 188829
rect 411571 188593 411613 188829
rect 411293 188509 411613 188593
rect 411293 188273 411335 188509
rect 411571 188273 411613 188509
rect 411293 188241 411613 188273
rect 415991 188829 416311 188861
rect 415991 188593 416033 188829
rect 416269 188593 416311 188829
rect 415991 188509 416311 188593
rect 415991 188273 416033 188509
rect 416269 188273 416311 188509
rect 415991 188241 416311 188273
rect 420689 188829 421009 188861
rect 420689 188593 420731 188829
rect 420967 188593 421009 188829
rect 420689 188509 421009 188593
rect 420689 188273 420731 188509
rect 420967 188273 421009 188509
rect 420689 188241 421009 188273
rect 425387 188829 425707 188861
rect 425387 188593 425429 188829
rect 425665 188593 425707 188829
rect 425387 188509 425707 188593
rect 425387 188273 425429 188509
rect 425665 188273 425707 188509
rect 425387 188241 425707 188273
rect 439293 188829 439613 188861
rect 439293 188593 439335 188829
rect 439571 188593 439613 188829
rect 439293 188509 439613 188593
rect 439293 188273 439335 188509
rect 439571 188273 439613 188509
rect 439293 188241 439613 188273
rect 443991 188829 444311 188861
rect 443991 188593 444033 188829
rect 444269 188593 444311 188829
rect 443991 188509 444311 188593
rect 443991 188273 444033 188509
rect 444269 188273 444311 188509
rect 443991 188241 444311 188273
rect 362340 185454 362660 185486
rect 362340 185218 362382 185454
rect 362618 185218 362660 185454
rect 362340 185134 362660 185218
rect 362340 184898 362382 185134
rect 362618 184898 362660 185134
rect 362340 184866 362660 184898
rect 367038 185454 367358 185486
rect 367038 185218 367080 185454
rect 367316 185218 367358 185454
rect 367038 185134 367358 185218
rect 367038 184898 367080 185134
rect 367316 184898 367358 185134
rect 367038 184866 367358 184898
rect 385642 185454 385962 185486
rect 385642 185218 385684 185454
rect 385920 185218 385962 185454
rect 385642 185134 385962 185218
rect 385642 184898 385684 185134
rect 385920 184898 385962 185134
rect 385642 184866 385962 184898
rect 390340 185454 390660 185486
rect 390340 185218 390382 185454
rect 390618 185218 390660 185454
rect 390340 185134 390660 185218
rect 390340 184898 390382 185134
rect 390618 184898 390660 185134
rect 390340 184866 390660 184898
rect 395038 185454 395358 185486
rect 395038 185218 395080 185454
rect 395316 185218 395358 185454
rect 395038 185134 395358 185218
rect 395038 184898 395080 185134
rect 395316 184898 395358 185134
rect 395038 184866 395358 184898
rect 413642 185454 413962 185486
rect 413642 185218 413684 185454
rect 413920 185218 413962 185454
rect 413642 185134 413962 185218
rect 413642 184898 413684 185134
rect 413920 184898 413962 185134
rect 413642 184866 413962 184898
rect 418340 185454 418660 185486
rect 418340 185218 418382 185454
rect 418618 185218 418660 185454
rect 418340 185134 418660 185218
rect 418340 184898 418382 185134
rect 418618 184898 418660 185134
rect 418340 184866 418660 184898
rect 423038 185454 423358 185486
rect 423038 185218 423080 185454
rect 423316 185218 423358 185454
rect 423038 185134 423358 185218
rect 423038 184898 423080 185134
rect 423316 184898 423358 185134
rect 423038 184866 423358 184898
rect 441642 185454 441962 185486
rect 441642 185218 441684 185454
rect 441920 185218 441962 185454
rect 441642 185134 441962 185218
rect 441642 184898 441684 185134
rect 441920 184898 441962 185134
rect 441642 184866 441962 184898
rect 445710 176629 445770 198459
rect 448689 188829 449009 188861
rect 448689 188593 448731 188829
rect 448967 188593 449009 188829
rect 448689 188509 449009 188593
rect 448689 188273 448731 188509
rect 448967 188273 449009 188509
rect 448689 188241 449009 188273
rect 453387 188829 453707 188861
rect 453387 188593 453429 188829
rect 453665 188593 453707 188829
rect 453387 188509 453707 188593
rect 453387 188273 453429 188509
rect 453665 188273 453707 188509
rect 453387 188241 453707 188273
rect 467293 188829 467613 188861
rect 467293 188593 467335 188829
rect 467571 188593 467613 188829
rect 467293 188509 467613 188593
rect 467293 188273 467335 188509
rect 467571 188273 467613 188509
rect 467293 188241 467613 188273
rect 471991 188829 472311 188861
rect 471991 188593 472033 188829
rect 472269 188593 472311 188829
rect 471991 188509 472311 188593
rect 471991 188273 472033 188509
rect 472269 188273 472311 188509
rect 471991 188241 472311 188273
rect 476689 188829 477009 188861
rect 476689 188593 476731 188829
rect 476967 188593 477009 188829
rect 476689 188509 477009 188593
rect 476689 188273 476731 188509
rect 476967 188273 477009 188509
rect 476689 188241 477009 188273
rect 481387 188829 481707 188861
rect 481387 188593 481429 188829
rect 481665 188593 481707 188829
rect 481387 188509 481707 188593
rect 481387 188273 481429 188509
rect 481665 188273 481707 188509
rect 481387 188241 481707 188273
rect 495293 188829 495613 188861
rect 495293 188593 495335 188829
rect 495571 188593 495613 188829
rect 495293 188509 495613 188593
rect 495293 188273 495335 188509
rect 495571 188273 495613 188509
rect 495293 188241 495613 188273
rect 499991 188829 500311 188861
rect 499991 188593 500033 188829
rect 500269 188593 500311 188829
rect 499991 188509 500311 188593
rect 499991 188273 500033 188509
rect 500269 188273 500311 188509
rect 499991 188241 500311 188273
rect 504689 188829 505009 188861
rect 504689 188593 504731 188829
rect 504967 188593 505009 188829
rect 504689 188509 505009 188593
rect 504689 188273 504731 188509
rect 504967 188273 505009 188509
rect 504689 188241 505009 188273
rect 509387 188829 509707 188861
rect 509387 188593 509429 188829
rect 509665 188593 509707 188829
rect 509387 188509 509707 188593
rect 509387 188273 509429 188509
rect 509665 188273 509707 188509
rect 509387 188241 509707 188273
rect 523293 188829 523613 188861
rect 523293 188593 523335 188829
rect 523571 188593 523613 188829
rect 523293 188509 523613 188593
rect 523293 188273 523335 188509
rect 523571 188273 523613 188509
rect 523293 188241 523613 188273
rect 527991 188829 528311 188861
rect 527991 188593 528033 188829
rect 528269 188593 528311 188829
rect 527991 188509 528311 188593
rect 527991 188273 528033 188509
rect 528269 188273 528311 188509
rect 527991 188241 528311 188273
rect 532689 188829 533009 188861
rect 532689 188593 532731 188829
rect 532967 188593 533009 188829
rect 532689 188509 533009 188593
rect 532689 188273 532731 188509
rect 532967 188273 533009 188509
rect 532689 188241 533009 188273
rect 537387 188829 537707 188861
rect 537387 188593 537429 188829
rect 537665 188593 537707 188829
rect 537387 188509 537707 188593
rect 537387 188273 537429 188509
rect 537665 188273 537707 188509
rect 537387 188241 537707 188273
rect 551293 188829 551613 188861
rect 551293 188593 551335 188829
rect 551571 188593 551613 188829
rect 551293 188509 551613 188593
rect 551293 188273 551335 188509
rect 551571 188273 551613 188509
rect 551293 188241 551613 188273
rect 555991 188829 556311 188861
rect 555991 188593 556033 188829
rect 556269 188593 556311 188829
rect 555991 188509 556311 188593
rect 555991 188273 556033 188509
rect 556269 188273 556311 188509
rect 555991 188241 556311 188273
rect 560689 188829 561009 188861
rect 560689 188593 560731 188829
rect 560967 188593 561009 188829
rect 560689 188509 561009 188593
rect 560689 188273 560731 188509
rect 560967 188273 561009 188509
rect 560689 188241 561009 188273
rect 565387 188829 565707 188861
rect 565387 188593 565429 188829
rect 565665 188593 565707 188829
rect 565387 188509 565707 188593
rect 565387 188273 565429 188509
rect 565665 188273 565707 188509
rect 565387 188241 565707 188273
rect 573494 188829 574114 215273
rect 573494 188593 573526 188829
rect 573762 188593 573846 188829
rect 574082 188593 574114 188829
rect 573494 188509 574114 188593
rect 573494 188273 573526 188509
rect 573762 188273 573846 188509
rect 574082 188273 574114 188509
rect 446340 185454 446660 185486
rect 446340 185218 446382 185454
rect 446618 185218 446660 185454
rect 446340 185134 446660 185218
rect 446340 184898 446382 185134
rect 446618 184898 446660 185134
rect 446340 184866 446660 184898
rect 451038 185454 451358 185486
rect 451038 185218 451080 185454
rect 451316 185218 451358 185454
rect 451038 185134 451358 185218
rect 451038 184898 451080 185134
rect 451316 184898 451358 185134
rect 451038 184866 451358 184898
rect 469642 185454 469962 185486
rect 469642 185218 469684 185454
rect 469920 185218 469962 185454
rect 469642 185134 469962 185218
rect 469642 184898 469684 185134
rect 469920 184898 469962 185134
rect 469642 184866 469962 184898
rect 474340 185454 474660 185486
rect 474340 185218 474382 185454
rect 474618 185218 474660 185454
rect 474340 185134 474660 185218
rect 474340 184898 474382 185134
rect 474618 184898 474660 185134
rect 474340 184866 474660 184898
rect 479038 185454 479358 185486
rect 479038 185218 479080 185454
rect 479316 185218 479358 185454
rect 479038 185134 479358 185218
rect 479038 184898 479080 185134
rect 479316 184898 479358 185134
rect 479038 184866 479358 184898
rect 497642 185454 497962 185486
rect 497642 185218 497684 185454
rect 497920 185218 497962 185454
rect 497642 185134 497962 185218
rect 497642 184898 497684 185134
rect 497920 184898 497962 185134
rect 497642 184866 497962 184898
rect 502340 185454 502660 185486
rect 502340 185218 502382 185454
rect 502618 185218 502660 185454
rect 502340 185134 502660 185218
rect 502340 184898 502382 185134
rect 502618 184898 502660 185134
rect 502340 184866 502660 184898
rect 507038 185454 507358 185486
rect 507038 185218 507080 185454
rect 507316 185218 507358 185454
rect 507038 185134 507358 185218
rect 507038 184898 507080 185134
rect 507316 184898 507358 185134
rect 507038 184866 507358 184898
rect 525642 185454 525962 185486
rect 525642 185218 525684 185454
rect 525920 185218 525962 185454
rect 525642 185134 525962 185218
rect 525642 184898 525684 185134
rect 525920 184898 525962 185134
rect 525642 184866 525962 184898
rect 530340 185454 530660 185486
rect 530340 185218 530382 185454
rect 530618 185218 530660 185454
rect 530340 185134 530660 185218
rect 530340 184898 530382 185134
rect 530618 184898 530660 185134
rect 530340 184866 530660 184898
rect 535038 185454 535358 185486
rect 535038 185218 535080 185454
rect 535316 185218 535358 185454
rect 535038 185134 535358 185218
rect 535038 184898 535080 185134
rect 535316 184898 535358 185134
rect 535038 184866 535358 184898
rect 553642 185454 553962 185486
rect 553642 185218 553684 185454
rect 553920 185218 553962 185454
rect 553642 185134 553962 185218
rect 553642 184898 553684 185134
rect 553920 184898 553962 185134
rect 553642 184866 553962 184898
rect 558340 185454 558660 185486
rect 558340 185218 558382 185454
rect 558618 185218 558660 185454
rect 558340 185134 558660 185218
rect 558340 184898 558382 185134
rect 558618 184898 558660 185134
rect 558340 184866 558660 184898
rect 563038 185454 563358 185486
rect 563038 185218 563080 185454
rect 563316 185218 563358 185454
rect 563038 185134 563358 185218
rect 563038 184898 563080 185134
rect 563316 184898 563358 185134
rect 563038 184866 563358 184898
rect 259499 176628 259565 176629
rect 259499 176564 259500 176628
rect 259564 176564 259565 176628
rect 259499 176563 259565 176564
rect 361619 176628 361685 176629
rect 361619 176564 361620 176628
rect 361684 176564 361685 176628
rect 361619 176563 361685 176564
rect 445707 176628 445773 176629
rect 445707 176564 445708 176628
rect 445772 176564 445773 176628
rect 445707 176563 445773 176564
rect 148363 170644 148429 170645
rect 148363 170580 148364 170644
rect 148428 170580 148429 170644
rect 148363 170579 148429 170580
rect 128491 170372 128557 170373
rect 128491 170308 128492 170372
rect 128556 170308 128557 170372
rect 128491 170307 128557 170308
rect 128494 162349 128554 170307
rect 148366 162349 148426 170579
rect 372291 170372 372357 170373
rect 372291 170308 372292 170372
rect 372356 170308 372357 170372
rect 372291 170307 372357 170308
rect 344323 170236 344389 170237
rect 344323 170172 344324 170236
rect 344388 170172 344389 170236
rect 344323 170171 344389 170172
rect 344326 162349 344386 170171
rect 372294 162349 372354 170307
rect 540467 170236 540533 170237
rect 540467 170172 540468 170236
rect 540532 170172 540533 170236
rect 540467 170171 540533 170172
rect 408539 170100 408605 170101
rect 408539 170036 408540 170100
rect 408604 170036 408605 170100
rect 408539 170035 408605 170036
rect 520595 170100 520661 170101
rect 520595 170036 520596 170100
rect 520660 170036 520661 170100
rect 520595 170035 520661 170036
rect 408542 162349 408602 170035
rect 520598 162349 520658 170035
rect 540470 162349 540530 170171
rect 128491 162348 128557 162349
rect 128491 162284 128492 162348
rect 128556 162284 128557 162348
rect 128491 162283 128557 162284
rect 148363 162348 148429 162349
rect 148363 162284 148364 162348
rect 148428 162284 148429 162348
rect 148363 162283 148429 162284
rect 344323 162348 344389 162349
rect 344323 162284 344324 162348
rect 344388 162284 344389 162348
rect 344323 162283 344389 162284
rect 372291 162348 372357 162349
rect 372291 162284 372292 162348
rect 372356 162284 372357 162348
rect 372291 162283 372357 162284
rect 408539 162348 408605 162349
rect 408539 162284 408540 162348
rect 408604 162284 408605 162348
rect 408539 162283 408605 162284
rect 520595 162348 520661 162349
rect 520595 162284 520596 162348
rect 520660 162284 520661 162348
rect 520595 162283 520661 162284
rect 540467 162348 540533 162349
rect 540467 162284 540468 162348
rect 540532 162284 540533 162348
rect 540467 162283 540533 162284
rect 75293 161829 75613 161861
rect 75293 161593 75335 161829
rect 75571 161593 75613 161829
rect 75293 161509 75613 161593
rect 75293 161273 75335 161509
rect 75571 161273 75613 161509
rect 75293 161241 75613 161273
rect 79991 161829 80311 161861
rect 79991 161593 80033 161829
rect 80269 161593 80311 161829
rect 79991 161509 80311 161593
rect 79991 161273 80033 161509
rect 80269 161273 80311 161509
rect 79991 161241 80311 161273
rect 84689 161829 85009 161861
rect 84689 161593 84731 161829
rect 84967 161593 85009 161829
rect 84689 161509 85009 161593
rect 84689 161273 84731 161509
rect 84967 161273 85009 161509
rect 84689 161241 85009 161273
rect 89387 161829 89707 161861
rect 89387 161593 89429 161829
rect 89665 161593 89707 161829
rect 89387 161509 89707 161593
rect 89387 161273 89429 161509
rect 89665 161273 89707 161509
rect 89387 161241 89707 161273
rect 103293 161829 103613 161861
rect 103293 161593 103335 161829
rect 103571 161593 103613 161829
rect 103293 161509 103613 161593
rect 103293 161273 103335 161509
rect 103571 161273 103613 161509
rect 103293 161241 103613 161273
rect 107991 161829 108311 161861
rect 107991 161593 108033 161829
rect 108269 161593 108311 161829
rect 107991 161509 108311 161593
rect 107991 161273 108033 161509
rect 108269 161273 108311 161509
rect 107991 161241 108311 161273
rect 112689 161829 113009 161861
rect 112689 161593 112731 161829
rect 112967 161593 113009 161829
rect 112689 161509 113009 161593
rect 112689 161273 112731 161509
rect 112967 161273 113009 161509
rect 112689 161241 113009 161273
rect 117387 161829 117707 161861
rect 117387 161593 117429 161829
rect 117665 161593 117707 161829
rect 117387 161509 117707 161593
rect 117387 161273 117429 161509
rect 117665 161273 117707 161509
rect 117387 161241 117707 161273
rect 131293 161829 131613 161861
rect 131293 161593 131335 161829
rect 131571 161593 131613 161829
rect 131293 161509 131613 161593
rect 131293 161273 131335 161509
rect 131571 161273 131613 161509
rect 131293 161241 131613 161273
rect 135991 161829 136311 161861
rect 135991 161593 136033 161829
rect 136269 161593 136311 161829
rect 135991 161509 136311 161593
rect 135991 161273 136033 161509
rect 136269 161273 136311 161509
rect 135991 161241 136311 161273
rect 140689 161829 141009 161861
rect 140689 161593 140731 161829
rect 140967 161593 141009 161829
rect 140689 161509 141009 161593
rect 140689 161273 140731 161509
rect 140967 161273 141009 161509
rect 140689 161241 141009 161273
rect 145387 161829 145707 161861
rect 145387 161593 145429 161829
rect 145665 161593 145707 161829
rect 145387 161509 145707 161593
rect 145387 161273 145429 161509
rect 145665 161273 145707 161509
rect 145387 161241 145707 161273
rect 159293 161829 159613 161861
rect 159293 161593 159335 161829
rect 159571 161593 159613 161829
rect 159293 161509 159613 161593
rect 159293 161273 159335 161509
rect 159571 161273 159613 161509
rect 159293 161241 159613 161273
rect 163991 161829 164311 161861
rect 163991 161593 164033 161829
rect 164269 161593 164311 161829
rect 163991 161509 164311 161593
rect 163991 161273 164033 161509
rect 164269 161273 164311 161509
rect 163991 161241 164311 161273
rect 168689 161829 169009 161861
rect 168689 161593 168731 161829
rect 168967 161593 169009 161829
rect 168689 161509 169009 161593
rect 168689 161273 168731 161509
rect 168967 161273 169009 161509
rect 168689 161241 169009 161273
rect 173387 161829 173707 161861
rect 173387 161593 173429 161829
rect 173665 161593 173707 161829
rect 173387 161509 173707 161593
rect 173387 161273 173429 161509
rect 173665 161273 173707 161509
rect 173387 161241 173707 161273
rect 187293 161829 187613 161861
rect 187293 161593 187335 161829
rect 187571 161593 187613 161829
rect 187293 161509 187613 161593
rect 187293 161273 187335 161509
rect 187571 161273 187613 161509
rect 187293 161241 187613 161273
rect 191991 161829 192311 161861
rect 191991 161593 192033 161829
rect 192269 161593 192311 161829
rect 191991 161509 192311 161593
rect 191991 161273 192033 161509
rect 192269 161273 192311 161509
rect 191991 161241 192311 161273
rect 196689 161829 197009 161861
rect 196689 161593 196731 161829
rect 196967 161593 197009 161829
rect 196689 161509 197009 161593
rect 196689 161273 196731 161509
rect 196967 161273 197009 161509
rect 196689 161241 197009 161273
rect 201387 161829 201707 161861
rect 201387 161593 201429 161829
rect 201665 161593 201707 161829
rect 201387 161509 201707 161593
rect 201387 161273 201429 161509
rect 201665 161273 201707 161509
rect 201387 161241 201707 161273
rect 215293 161829 215613 161861
rect 215293 161593 215335 161829
rect 215571 161593 215613 161829
rect 215293 161509 215613 161593
rect 215293 161273 215335 161509
rect 215571 161273 215613 161509
rect 215293 161241 215613 161273
rect 219991 161829 220311 161861
rect 219991 161593 220033 161829
rect 220269 161593 220311 161829
rect 219991 161509 220311 161593
rect 219991 161273 220033 161509
rect 220269 161273 220311 161509
rect 219991 161241 220311 161273
rect 224689 161829 225009 161861
rect 224689 161593 224731 161829
rect 224967 161593 225009 161829
rect 224689 161509 225009 161593
rect 224689 161273 224731 161509
rect 224967 161273 225009 161509
rect 224689 161241 225009 161273
rect 229387 161829 229707 161861
rect 229387 161593 229429 161829
rect 229665 161593 229707 161829
rect 229387 161509 229707 161593
rect 229387 161273 229429 161509
rect 229665 161273 229707 161509
rect 229387 161241 229707 161273
rect 243293 161829 243613 161861
rect 243293 161593 243335 161829
rect 243571 161593 243613 161829
rect 243293 161509 243613 161593
rect 243293 161273 243335 161509
rect 243571 161273 243613 161509
rect 243293 161241 243613 161273
rect 247991 161829 248311 161861
rect 247991 161593 248033 161829
rect 248269 161593 248311 161829
rect 247991 161509 248311 161593
rect 247991 161273 248033 161509
rect 248269 161273 248311 161509
rect 247991 161241 248311 161273
rect 252689 161829 253009 161861
rect 252689 161593 252731 161829
rect 252967 161593 253009 161829
rect 252689 161509 253009 161593
rect 252689 161273 252731 161509
rect 252967 161273 253009 161509
rect 252689 161241 253009 161273
rect 257387 161829 257707 161861
rect 257387 161593 257429 161829
rect 257665 161593 257707 161829
rect 257387 161509 257707 161593
rect 257387 161273 257429 161509
rect 257665 161273 257707 161509
rect 257387 161241 257707 161273
rect 271293 161829 271613 161861
rect 271293 161593 271335 161829
rect 271571 161593 271613 161829
rect 271293 161509 271613 161593
rect 271293 161273 271335 161509
rect 271571 161273 271613 161509
rect 271293 161241 271613 161273
rect 275991 161829 276311 161861
rect 275991 161593 276033 161829
rect 276269 161593 276311 161829
rect 275991 161509 276311 161593
rect 275991 161273 276033 161509
rect 276269 161273 276311 161509
rect 275991 161241 276311 161273
rect 280689 161829 281009 161861
rect 280689 161593 280731 161829
rect 280967 161593 281009 161829
rect 280689 161509 281009 161593
rect 280689 161273 280731 161509
rect 280967 161273 281009 161509
rect 280689 161241 281009 161273
rect 285387 161829 285707 161861
rect 285387 161593 285429 161829
rect 285665 161593 285707 161829
rect 285387 161509 285707 161593
rect 285387 161273 285429 161509
rect 285665 161273 285707 161509
rect 285387 161241 285707 161273
rect 299293 161829 299613 161861
rect 299293 161593 299335 161829
rect 299571 161593 299613 161829
rect 299293 161509 299613 161593
rect 299293 161273 299335 161509
rect 299571 161273 299613 161509
rect 299293 161241 299613 161273
rect 303991 161829 304311 161861
rect 303991 161593 304033 161829
rect 304269 161593 304311 161829
rect 303991 161509 304311 161593
rect 303991 161273 304033 161509
rect 304269 161273 304311 161509
rect 303991 161241 304311 161273
rect 308689 161829 309009 161861
rect 308689 161593 308731 161829
rect 308967 161593 309009 161829
rect 308689 161509 309009 161593
rect 308689 161273 308731 161509
rect 308967 161273 309009 161509
rect 308689 161241 309009 161273
rect 313387 161829 313707 161861
rect 313387 161593 313429 161829
rect 313665 161593 313707 161829
rect 313387 161509 313707 161593
rect 313387 161273 313429 161509
rect 313665 161273 313707 161509
rect 313387 161241 313707 161273
rect 327293 161829 327613 161861
rect 327293 161593 327335 161829
rect 327571 161593 327613 161829
rect 327293 161509 327613 161593
rect 327293 161273 327335 161509
rect 327571 161273 327613 161509
rect 327293 161241 327613 161273
rect 331991 161829 332311 161861
rect 331991 161593 332033 161829
rect 332269 161593 332311 161829
rect 331991 161509 332311 161593
rect 331991 161273 332033 161509
rect 332269 161273 332311 161509
rect 331991 161241 332311 161273
rect 336689 161829 337009 161861
rect 336689 161593 336731 161829
rect 336967 161593 337009 161829
rect 336689 161509 337009 161593
rect 336689 161273 336731 161509
rect 336967 161273 337009 161509
rect 336689 161241 337009 161273
rect 341387 161829 341707 161861
rect 341387 161593 341429 161829
rect 341665 161593 341707 161829
rect 341387 161509 341707 161593
rect 341387 161273 341429 161509
rect 341665 161273 341707 161509
rect 341387 161241 341707 161273
rect 355293 161829 355613 161861
rect 355293 161593 355335 161829
rect 355571 161593 355613 161829
rect 355293 161509 355613 161593
rect 355293 161273 355335 161509
rect 355571 161273 355613 161509
rect 355293 161241 355613 161273
rect 359991 161829 360311 161861
rect 359991 161593 360033 161829
rect 360269 161593 360311 161829
rect 359991 161509 360311 161593
rect 359991 161273 360033 161509
rect 360269 161273 360311 161509
rect 359991 161241 360311 161273
rect 364689 161829 365009 161861
rect 364689 161593 364731 161829
rect 364967 161593 365009 161829
rect 364689 161509 365009 161593
rect 364689 161273 364731 161509
rect 364967 161273 365009 161509
rect 364689 161241 365009 161273
rect 369387 161829 369707 161861
rect 369387 161593 369429 161829
rect 369665 161593 369707 161829
rect 369387 161509 369707 161593
rect 369387 161273 369429 161509
rect 369665 161273 369707 161509
rect 369387 161241 369707 161273
rect 383293 161829 383613 161861
rect 383293 161593 383335 161829
rect 383571 161593 383613 161829
rect 383293 161509 383613 161593
rect 383293 161273 383335 161509
rect 383571 161273 383613 161509
rect 383293 161241 383613 161273
rect 387991 161829 388311 161861
rect 387991 161593 388033 161829
rect 388269 161593 388311 161829
rect 387991 161509 388311 161593
rect 387991 161273 388033 161509
rect 388269 161273 388311 161509
rect 387991 161241 388311 161273
rect 392689 161829 393009 161861
rect 392689 161593 392731 161829
rect 392967 161593 393009 161829
rect 392689 161509 393009 161593
rect 392689 161273 392731 161509
rect 392967 161273 393009 161509
rect 392689 161241 393009 161273
rect 397387 161829 397707 161861
rect 397387 161593 397429 161829
rect 397665 161593 397707 161829
rect 397387 161509 397707 161593
rect 397387 161273 397429 161509
rect 397665 161273 397707 161509
rect 397387 161241 397707 161273
rect 411293 161829 411613 161861
rect 411293 161593 411335 161829
rect 411571 161593 411613 161829
rect 411293 161509 411613 161593
rect 411293 161273 411335 161509
rect 411571 161273 411613 161509
rect 411293 161241 411613 161273
rect 415991 161829 416311 161861
rect 415991 161593 416033 161829
rect 416269 161593 416311 161829
rect 415991 161509 416311 161593
rect 415991 161273 416033 161509
rect 416269 161273 416311 161509
rect 415991 161241 416311 161273
rect 420689 161829 421009 161861
rect 420689 161593 420731 161829
rect 420967 161593 421009 161829
rect 420689 161509 421009 161593
rect 420689 161273 420731 161509
rect 420967 161273 421009 161509
rect 420689 161241 421009 161273
rect 425387 161829 425707 161861
rect 425387 161593 425429 161829
rect 425665 161593 425707 161829
rect 425387 161509 425707 161593
rect 425387 161273 425429 161509
rect 425665 161273 425707 161509
rect 425387 161241 425707 161273
rect 439293 161829 439613 161861
rect 439293 161593 439335 161829
rect 439571 161593 439613 161829
rect 439293 161509 439613 161593
rect 439293 161273 439335 161509
rect 439571 161273 439613 161509
rect 439293 161241 439613 161273
rect 443991 161829 444311 161861
rect 443991 161593 444033 161829
rect 444269 161593 444311 161829
rect 443991 161509 444311 161593
rect 443991 161273 444033 161509
rect 444269 161273 444311 161509
rect 443991 161241 444311 161273
rect 448689 161829 449009 161861
rect 448689 161593 448731 161829
rect 448967 161593 449009 161829
rect 448689 161509 449009 161593
rect 448689 161273 448731 161509
rect 448967 161273 449009 161509
rect 448689 161241 449009 161273
rect 453387 161829 453707 161861
rect 453387 161593 453429 161829
rect 453665 161593 453707 161829
rect 453387 161509 453707 161593
rect 453387 161273 453429 161509
rect 453665 161273 453707 161509
rect 453387 161241 453707 161273
rect 467293 161829 467613 161861
rect 467293 161593 467335 161829
rect 467571 161593 467613 161829
rect 467293 161509 467613 161593
rect 467293 161273 467335 161509
rect 467571 161273 467613 161509
rect 467293 161241 467613 161273
rect 471991 161829 472311 161861
rect 471991 161593 472033 161829
rect 472269 161593 472311 161829
rect 471991 161509 472311 161593
rect 471991 161273 472033 161509
rect 472269 161273 472311 161509
rect 471991 161241 472311 161273
rect 476689 161829 477009 161861
rect 476689 161593 476731 161829
rect 476967 161593 477009 161829
rect 476689 161509 477009 161593
rect 476689 161273 476731 161509
rect 476967 161273 477009 161509
rect 476689 161241 477009 161273
rect 481387 161829 481707 161861
rect 481387 161593 481429 161829
rect 481665 161593 481707 161829
rect 481387 161509 481707 161593
rect 481387 161273 481429 161509
rect 481665 161273 481707 161509
rect 481387 161241 481707 161273
rect 495293 161829 495613 161861
rect 495293 161593 495335 161829
rect 495571 161593 495613 161829
rect 495293 161509 495613 161593
rect 495293 161273 495335 161509
rect 495571 161273 495613 161509
rect 495293 161241 495613 161273
rect 499991 161829 500311 161861
rect 499991 161593 500033 161829
rect 500269 161593 500311 161829
rect 499991 161509 500311 161593
rect 499991 161273 500033 161509
rect 500269 161273 500311 161509
rect 499991 161241 500311 161273
rect 504689 161829 505009 161861
rect 504689 161593 504731 161829
rect 504967 161593 505009 161829
rect 504689 161509 505009 161593
rect 504689 161273 504731 161509
rect 504967 161273 505009 161509
rect 504689 161241 505009 161273
rect 509387 161829 509707 161861
rect 509387 161593 509429 161829
rect 509665 161593 509707 161829
rect 509387 161509 509707 161593
rect 509387 161273 509429 161509
rect 509665 161273 509707 161509
rect 509387 161241 509707 161273
rect 523293 161829 523613 161861
rect 523293 161593 523335 161829
rect 523571 161593 523613 161829
rect 523293 161509 523613 161593
rect 523293 161273 523335 161509
rect 523571 161273 523613 161509
rect 523293 161241 523613 161273
rect 527991 161829 528311 161861
rect 527991 161593 528033 161829
rect 528269 161593 528311 161829
rect 527991 161509 528311 161593
rect 527991 161273 528033 161509
rect 528269 161273 528311 161509
rect 527991 161241 528311 161273
rect 532689 161829 533009 161861
rect 532689 161593 532731 161829
rect 532967 161593 533009 161829
rect 532689 161509 533009 161593
rect 532689 161273 532731 161509
rect 532967 161273 533009 161509
rect 532689 161241 533009 161273
rect 537387 161829 537707 161861
rect 537387 161593 537429 161829
rect 537665 161593 537707 161829
rect 537387 161509 537707 161593
rect 537387 161273 537429 161509
rect 537665 161273 537707 161509
rect 537387 161241 537707 161273
rect 551293 161829 551613 161861
rect 551293 161593 551335 161829
rect 551571 161593 551613 161829
rect 551293 161509 551613 161593
rect 551293 161273 551335 161509
rect 551571 161273 551613 161509
rect 551293 161241 551613 161273
rect 555991 161829 556311 161861
rect 555991 161593 556033 161829
rect 556269 161593 556311 161829
rect 555991 161509 556311 161593
rect 555991 161273 556033 161509
rect 556269 161273 556311 161509
rect 555991 161241 556311 161273
rect 560689 161829 561009 161861
rect 560689 161593 560731 161829
rect 560967 161593 561009 161829
rect 560689 161509 561009 161593
rect 560689 161273 560731 161509
rect 560967 161273 561009 161509
rect 560689 161241 561009 161273
rect 565387 161829 565707 161861
rect 565387 161593 565429 161829
rect 565665 161593 565707 161829
rect 565387 161509 565707 161593
rect 565387 161273 565429 161509
rect 565665 161273 565707 161509
rect 565387 161241 565707 161273
rect 573494 161829 574114 188273
rect 573494 161593 573526 161829
rect 573762 161593 573846 161829
rect 574082 161593 574114 161829
rect 573494 161509 574114 161593
rect 573494 161273 573526 161509
rect 573762 161273 573846 161509
rect 574082 161273 574114 161509
rect 77642 158454 77962 158486
rect 77642 158218 77684 158454
rect 77920 158218 77962 158454
rect 77642 158134 77962 158218
rect 77642 157898 77684 158134
rect 77920 157898 77962 158134
rect 77642 157866 77962 157898
rect 82340 158454 82660 158486
rect 82340 158218 82382 158454
rect 82618 158218 82660 158454
rect 82340 158134 82660 158218
rect 82340 157898 82382 158134
rect 82618 157898 82660 158134
rect 82340 157866 82660 157898
rect 87038 158454 87358 158486
rect 87038 158218 87080 158454
rect 87316 158218 87358 158454
rect 87038 158134 87358 158218
rect 87038 157898 87080 158134
rect 87316 157898 87358 158134
rect 87038 157866 87358 157898
rect 105642 158454 105962 158486
rect 105642 158218 105684 158454
rect 105920 158218 105962 158454
rect 105642 158134 105962 158218
rect 105642 157898 105684 158134
rect 105920 157898 105962 158134
rect 105642 157866 105962 157898
rect 110340 158454 110660 158486
rect 110340 158218 110382 158454
rect 110618 158218 110660 158454
rect 110340 158134 110660 158218
rect 110340 157898 110382 158134
rect 110618 157898 110660 158134
rect 110340 157866 110660 157898
rect 115038 158454 115358 158486
rect 115038 158218 115080 158454
rect 115316 158218 115358 158454
rect 115038 158134 115358 158218
rect 115038 157898 115080 158134
rect 115316 157898 115358 158134
rect 115038 157866 115358 157898
rect 133642 158454 133962 158486
rect 133642 158218 133684 158454
rect 133920 158218 133962 158454
rect 133642 158134 133962 158218
rect 133642 157898 133684 158134
rect 133920 157898 133962 158134
rect 133642 157866 133962 157898
rect 138340 158454 138660 158486
rect 138340 158218 138382 158454
rect 138618 158218 138660 158454
rect 138340 158134 138660 158218
rect 138340 157898 138382 158134
rect 138618 157898 138660 158134
rect 138340 157866 138660 157898
rect 143038 158454 143358 158486
rect 143038 158218 143080 158454
rect 143316 158218 143358 158454
rect 143038 158134 143358 158218
rect 143038 157898 143080 158134
rect 143316 157898 143358 158134
rect 143038 157866 143358 157898
rect 161642 158454 161962 158486
rect 161642 158218 161684 158454
rect 161920 158218 161962 158454
rect 161642 158134 161962 158218
rect 161642 157898 161684 158134
rect 161920 157898 161962 158134
rect 161642 157866 161962 157898
rect 166340 158454 166660 158486
rect 166340 158218 166382 158454
rect 166618 158218 166660 158454
rect 166340 158134 166660 158218
rect 166340 157898 166382 158134
rect 166618 157898 166660 158134
rect 166340 157866 166660 157898
rect 171038 158454 171358 158486
rect 171038 158218 171080 158454
rect 171316 158218 171358 158454
rect 171038 158134 171358 158218
rect 171038 157898 171080 158134
rect 171316 157898 171358 158134
rect 171038 157866 171358 157898
rect 189642 158454 189962 158486
rect 189642 158218 189684 158454
rect 189920 158218 189962 158454
rect 189642 158134 189962 158218
rect 189642 157898 189684 158134
rect 189920 157898 189962 158134
rect 189642 157866 189962 157898
rect 194340 158454 194660 158486
rect 194340 158218 194382 158454
rect 194618 158218 194660 158454
rect 194340 158134 194660 158218
rect 194340 157898 194382 158134
rect 194618 157898 194660 158134
rect 194340 157866 194660 157898
rect 199038 158454 199358 158486
rect 199038 158218 199080 158454
rect 199316 158218 199358 158454
rect 199038 158134 199358 158218
rect 199038 157898 199080 158134
rect 199316 157898 199358 158134
rect 199038 157866 199358 157898
rect 217642 158454 217962 158486
rect 217642 158218 217684 158454
rect 217920 158218 217962 158454
rect 217642 158134 217962 158218
rect 217642 157898 217684 158134
rect 217920 157898 217962 158134
rect 217642 157866 217962 157898
rect 222340 158454 222660 158486
rect 222340 158218 222382 158454
rect 222618 158218 222660 158454
rect 222340 158134 222660 158218
rect 222340 157898 222382 158134
rect 222618 157898 222660 158134
rect 222340 157866 222660 157898
rect 227038 158454 227358 158486
rect 227038 158218 227080 158454
rect 227316 158218 227358 158454
rect 227038 158134 227358 158218
rect 227038 157898 227080 158134
rect 227316 157898 227358 158134
rect 227038 157866 227358 157898
rect 245642 158454 245962 158486
rect 245642 158218 245684 158454
rect 245920 158218 245962 158454
rect 245642 158134 245962 158218
rect 245642 157898 245684 158134
rect 245920 157898 245962 158134
rect 245642 157866 245962 157898
rect 250340 158454 250660 158486
rect 250340 158218 250382 158454
rect 250618 158218 250660 158454
rect 250340 158134 250660 158218
rect 250340 157898 250382 158134
rect 250618 157898 250660 158134
rect 250340 157866 250660 157898
rect 255038 158454 255358 158486
rect 255038 158218 255080 158454
rect 255316 158218 255358 158454
rect 255038 158134 255358 158218
rect 255038 157898 255080 158134
rect 255316 157898 255358 158134
rect 255038 157866 255358 157898
rect 273642 158454 273962 158486
rect 273642 158218 273684 158454
rect 273920 158218 273962 158454
rect 273642 158134 273962 158218
rect 273642 157898 273684 158134
rect 273920 157898 273962 158134
rect 273642 157866 273962 157898
rect 278340 158454 278660 158486
rect 278340 158218 278382 158454
rect 278618 158218 278660 158454
rect 278340 158134 278660 158218
rect 278340 157898 278382 158134
rect 278618 157898 278660 158134
rect 278340 157866 278660 157898
rect 283038 158454 283358 158486
rect 283038 158218 283080 158454
rect 283316 158218 283358 158454
rect 283038 158134 283358 158218
rect 283038 157898 283080 158134
rect 283316 157898 283358 158134
rect 283038 157866 283358 157898
rect 301642 158454 301962 158486
rect 301642 158218 301684 158454
rect 301920 158218 301962 158454
rect 301642 158134 301962 158218
rect 301642 157898 301684 158134
rect 301920 157898 301962 158134
rect 301642 157866 301962 157898
rect 306340 158454 306660 158486
rect 306340 158218 306382 158454
rect 306618 158218 306660 158454
rect 306340 158134 306660 158218
rect 306340 157898 306382 158134
rect 306618 157898 306660 158134
rect 306340 157866 306660 157898
rect 311038 158454 311358 158486
rect 311038 158218 311080 158454
rect 311316 158218 311358 158454
rect 311038 158134 311358 158218
rect 311038 157898 311080 158134
rect 311316 157898 311358 158134
rect 311038 157866 311358 157898
rect 329642 158454 329962 158486
rect 329642 158218 329684 158454
rect 329920 158218 329962 158454
rect 329642 158134 329962 158218
rect 329642 157898 329684 158134
rect 329920 157898 329962 158134
rect 329642 157866 329962 157898
rect 334340 158454 334660 158486
rect 334340 158218 334382 158454
rect 334618 158218 334660 158454
rect 334340 158134 334660 158218
rect 334340 157898 334382 158134
rect 334618 157898 334660 158134
rect 334340 157866 334660 157898
rect 339038 158454 339358 158486
rect 339038 158218 339080 158454
rect 339316 158218 339358 158454
rect 339038 158134 339358 158218
rect 339038 157898 339080 158134
rect 339316 157898 339358 158134
rect 339038 157866 339358 157898
rect 357642 158454 357962 158486
rect 357642 158218 357684 158454
rect 357920 158218 357962 158454
rect 357642 158134 357962 158218
rect 357642 157898 357684 158134
rect 357920 157898 357962 158134
rect 357642 157866 357962 157898
rect 362340 158454 362660 158486
rect 362340 158218 362382 158454
rect 362618 158218 362660 158454
rect 362340 158134 362660 158218
rect 362340 157898 362382 158134
rect 362618 157898 362660 158134
rect 362340 157866 362660 157898
rect 367038 158454 367358 158486
rect 367038 158218 367080 158454
rect 367316 158218 367358 158454
rect 367038 158134 367358 158218
rect 367038 157898 367080 158134
rect 367316 157898 367358 158134
rect 367038 157866 367358 157898
rect 385642 158454 385962 158486
rect 385642 158218 385684 158454
rect 385920 158218 385962 158454
rect 385642 158134 385962 158218
rect 385642 157898 385684 158134
rect 385920 157898 385962 158134
rect 385642 157866 385962 157898
rect 390340 158454 390660 158486
rect 390340 158218 390382 158454
rect 390618 158218 390660 158454
rect 390340 158134 390660 158218
rect 390340 157898 390382 158134
rect 390618 157898 390660 158134
rect 390340 157866 390660 157898
rect 395038 158454 395358 158486
rect 395038 158218 395080 158454
rect 395316 158218 395358 158454
rect 395038 158134 395358 158218
rect 395038 157898 395080 158134
rect 395316 157898 395358 158134
rect 395038 157866 395358 157898
rect 413642 158454 413962 158486
rect 413642 158218 413684 158454
rect 413920 158218 413962 158454
rect 413642 158134 413962 158218
rect 413642 157898 413684 158134
rect 413920 157898 413962 158134
rect 413642 157866 413962 157898
rect 418340 158454 418660 158486
rect 418340 158218 418382 158454
rect 418618 158218 418660 158454
rect 418340 158134 418660 158218
rect 418340 157898 418382 158134
rect 418618 157898 418660 158134
rect 418340 157866 418660 157898
rect 423038 158454 423358 158486
rect 423038 158218 423080 158454
rect 423316 158218 423358 158454
rect 423038 158134 423358 158218
rect 423038 157898 423080 158134
rect 423316 157898 423358 158134
rect 423038 157866 423358 157898
rect 441642 158454 441962 158486
rect 441642 158218 441684 158454
rect 441920 158218 441962 158454
rect 441642 158134 441962 158218
rect 441642 157898 441684 158134
rect 441920 157898 441962 158134
rect 441642 157866 441962 157898
rect 446340 158454 446660 158486
rect 446340 158218 446382 158454
rect 446618 158218 446660 158454
rect 446340 158134 446660 158218
rect 446340 157898 446382 158134
rect 446618 157898 446660 158134
rect 446340 157866 446660 157898
rect 451038 158454 451358 158486
rect 451038 158218 451080 158454
rect 451316 158218 451358 158454
rect 451038 158134 451358 158218
rect 451038 157898 451080 158134
rect 451316 157898 451358 158134
rect 451038 157866 451358 157898
rect 469642 158454 469962 158486
rect 469642 158218 469684 158454
rect 469920 158218 469962 158454
rect 469642 158134 469962 158218
rect 469642 157898 469684 158134
rect 469920 157898 469962 158134
rect 469642 157866 469962 157898
rect 474340 158454 474660 158486
rect 474340 158218 474382 158454
rect 474618 158218 474660 158454
rect 474340 158134 474660 158218
rect 474340 157898 474382 158134
rect 474618 157898 474660 158134
rect 474340 157866 474660 157898
rect 479038 158454 479358 158486
rect 479038 158218 479080 158454
rect 479316 158218 479358 158454
rect 479038 158134 479358 158218
rect 479038 157898 479080 158134
rect 479316 157898 479358 158134
rect 479038 157866 479358 157898
rect 497642 158454 497962 158486
rect 497642 158218 497684 158454
rect 497920 158218 497962 158454
rect 497642 158134 497962 158218
rect 497642 157898 497684 158134
rect 497920 157898 497962 158134
rect 497642 157866 497962 157898
rect 502340 158454 502660 158486
rect 502340 158218 502382 158454
rect 502618 158218 502660 158454
rect 502340 158134 502660 158218
rect 502340 157898 502382 158134
rect 502618 157898 502660 158134
rect 502340 157866 502660 157898
rect 507038 158454 507358 158486
rect 507038 158218 507080 158454
rect 507316 158218 507358 158454
rect 507038 158134 507358 158218
rect 507038 157898 507080 158134
rect 507316 157898 507358 158134
rect 507038 157866 507358 157898
rect 525642 158454 525962 158486
rect 525642 158218 525684 158454
rect 525920 158218 525962 158454
rect 525642 158134 525962 158218
rect 525642 157898 525684 158134
rect 525920 157898 525962 158134
rect 525642 157866 525962 157898
rect 530340 158454 530660 158486
rect 530340 158218 530382 158454
rect 530618 158218 530660 158454
rect 530340 158134 530660 158218
rect 530340 157898 530382 158134
rect 530618 157898 530660 158134
rect 530340 157866 530660 157898
rect 535038 158454 535358 158486
rect 535038 158218 535080 158454
rect 535316 158218 535358 158454
rect 535038 158134 535358 158218
rect 535038 157898 535080 158134
rect 535316 157898 535358 158134
rect 535038 157866 535358 157898
rect 553642 158454 553962 158486
rect 553642 158218 553684 158454
rect 553920 158218 553962 158454
rect 553642 158134 553962 158218
rect 553642 157898 553684 158134
rect 553920 157898 553962 158134
rect 553642 157866 553962 157898
rect 558340 158454 558660 158486
rect 558340 158218 558382 158454
rect 558618 158218 558660 158454
rect 558340 158134 558660 158218
rect 558340 157898 558382 158134
rect 558618 157898 558660 158134
rect 558340 157866 558660 157898
rect 563038 158454 563358 158486
rect 563038 158218 563080 158454
rect 563316 158218 563358 158454
rect 563038 158134 563358 158218
rect 563038 157898 563080 158134
rect 563316 157898 563358 158134
rect 563038 157866 563358 157898
rect 361619 144532 361685 144533
rect 361619 144468 361620 144532
rect 361684 144468 361685 144532
rect 361619 144467 361685 144468
rect 445707 144532 445773 144533
rect 445707 144468 445708 144532
rect 445772 144468 445773 144532
rect 445707 144467 445773 144468
rect 75293 134829 75613 134861
rect 75293 134593 75335 134829
rect 75571 134593 75613 134829
rect 75293 134509 75613 134593
rect 75293 134273 75335 134509
rect 75571 134273 75613 134509
rect 75293 134241 75613 134273
rect 79991 134829 80311 134861
rect 79991 134593 80033 134829
rect 80269 134593 80311 134829
rect 79991 134509 80311 134593
rect 79991 134273 80033 134509
rect 80269 134273 80311 134509
rect 79991 134241 80311 134273
rect 84689 134829 85009 134861
rect 84689 134593 84731 134829
rect 84967 134593 85009 134829
rect 84689 134509 85009 134593
rect 84689 134273 84731 134509
rect 84967 134273 85009 134509
rect 84689 134241 85009 134273
rect 89387 134829 89707 134861
rect 89387 134593 89429 134829
rect 89665 134593 89707 134829
rect 89387 134509 89707 134593
rect 89387 134273 89429 134509
rect 89665 134273 89707 134509
rect 89387 134241 89707 134273
rect 103293 134829 103613 134861
rect 103293 134593 103335 134829
rect 103571 134593 103613 134829
rect 103293 134509 103613 134593
rect 103293 134273 103335 134509
rect 103571 134273 103613 134509
rect 103293 134241 103613 134273
rect 107991 134829 108311 134861
rect 107991 134593 108033 134829
rect 108269 134593 108311 134829
rect 107991 134509 108311 134593
rect 107991 134273 108033 134509
rect 108269 134273 108311 134509
rect 107991 134241 108311 134273
rect 112689 134829 113009 134861
rect 112689 134593 112731 134829
rect 112967 134593 113009 134829
rect 112689 134509 113009 134593
rect 112689 134273 112731 134509
rect 112967 134273 113009 134509
rect 112689 134241 113009 134273
rect 117387 134829 117707 134861
rect 117387 134593 117429 134829
rect 117665 134593 117707 134829
rect 117387 134509 117707 134593
rect 117387 134273 117429 134509
rect 117665 134273 117707 134509
rect 117387 134241 117707 134273
rect 131293 134829 131613 134861
rect 131293 134593 131335 134829
rect 131571 134593 131613 134829
rect 131293 134509 131613 134593
rect 131293 134273 131335 134509
rect 131571 134273 131613 134509
rect 131293 134241 131613 134273
rect 135991 134829 136311 134861
rect 135991 134593 136033 134829
rect 136269 134593 136311 134829
rect 135991 134509 136311 134593
rect 135991 134273 136033 134509
rect 136269 134273 136311 134509
rect 135991 134241 136311 134273
rect 140689 134829 141009 134861
rect 140689 134593 140731 134829
rect 140967 134593 141009 134829
rect 140689 134509 141009 134593
rect 140689 134273 140731 134509
rect 140967 134273 141009 134509
rect 140689 134241 141009 134273
rect 145387 134829 145707 134861
rect 145387 134593 145429 134829
rect 145665 134593 145707 134829
rect 145387 134509 145707 134593
rect 145387 134273 145429 134509
rect 145665 134273 145707 134509
rect 145387 134241 145707 134273
rect 159293 134829 159613 134861
rect 159293 134593 159335 134829
rect 159571 134593 159613 134829
rect 159293 134509 159613 134593
rect 159293 134273 159335 134509
rect 159571 134273 159613 134509
rect 159293 134241 159613 134273
rect 163991 134829 164311 134861
rect 163991 134593 164033 134829
rect 164269 134593 164311 134829
rect 163991 134509 164311 134593
rect 163991 134273 164033 134509
rect 164269 134273 164311 134509
rect 163991 134241 164311 134273
rect 168689 134829 169009 134861
rect 168689 134593 168731 134829
rect 168967 134593 169009 134829
rect 168689 134509 169009 134593
rect 168689 134273 168731 134509
rect 168967 134273 169009 134509
rect 168689 134241 169009 134273
rect 173387 134829 173707 134861
rect 173387 134593 173429 134829
rect 173665 134593 173707 134829
rect 173387 134509 173707 134593
rect 173387 134273 173429 134509
rect 173665 134273 173707 134509
rect 173387 134241 173707 134273
rect 187293 134829 187613 134861
rect 187293 134593 187335 134829
rect 187571 134593 187613 134829
rect 187293 134509 187613 134593
rect 187293 134273 187335 134509
rect 187571 134273 187613 134509
rect 187293 134241 187613 134273
rect 191991 134829 192311 134861
rect 191991 134593 192033 134829
rect 192269 134593 192311 134829
rect 191991 134509 192311 134593
rect 191991 134273 192033 134509
rect 192269 134273 192311 134509
rect 191991 134241 192311 134273
rect 196689 134829 197009 134861
rect 196689 134593 196731 134829
rect 196967 134593 197009 134829
rect 196689 134509 197009 134593
rect 196689 134273 196731 134509
rect 196967 134273 197009 134509
rect 196689 134241 197009 134273
rect 201387 134829 201707 134861
rect 201387 134593 201429 134829
rect 201665 134593 201707 134829
rect 201387 134509 201707 134593
rect 201387 134273 201429 134509
rect 201665 134273 201707 134509
rect 201387 134241 201707 134273
rect 215293 134829 215613 134861
rect 215293 134593 215335 134829
rect 215571 134593 215613 134829
rect 215293 134509 215613 134593
rect 215293 134273 215335 134509
rect 215571 134273 215613 134509
rect 215293 134241 215613 134273
rect 219991 134829 220311 134861
rect 219991 134593 220033 134829
rect 220269 134593 220311 134829
rect 219991 134509 220311 134593
rect 219991 134273 220033 134509
rect 220269 134273 220311 134509
rect 219991 134241 220311 134273
rect 224689 134829 225009 134861
rect 224689 134593 224731 134829
rect 224967 134593 225009 134829
rect 224689 134509 225009 134593
rect 224689 134273 224731 134509
rect 224967 134273 225009 134509
rect 224689 134241 225009 134273
rect 229387 134829 229707 134861
rect 229387 134593 229429 134829
rect 229665 134593 229707 134829
rect 229387 134509 229707 134593
rect 229387 134273 229429 134509
rect 229665 134273 229707 134509
rect 229387 134241 229707 134273
rect 243293 134829 243613 134861
rect 243293 134593 243335 134829
rect 243571 134593 243613 134829
rect 243293 134509 243613 134593
rect 243293 134273 243335 134509
rect 243571 134273 243613 134509
rect 243293 134241 243613 134273
rect 247991 134829 248311 134861
rect 247991 134593 248033 134829
rect 248269 134593 248311 134829
rect 247991 134509 248311 134593
rect 247991 134273 248033 134509
rect 248269 134273 248311 134509
rect 247991 134241 248311 134273
rect 252689 134829 253009 134861
rect 252689 134593 252731 134829
rect 252967 134593 253009 134829
rect 252689 134509 253009 134593
rect 252689 134273 252731 134509
rect 252967 134273 253009 134509
rect 252689 134241 253009 134273
rect 257387 134829 257707 134861
rect 257387 134593 257429 134829
rect 257665 134593 257707 134829
rect 257387 134509 257707 134593
rect 257387 134273 257429 134509
rect 257665 134273 257707 134509
rect 257387 134241 257707 134273
rect 271293 134829 271613 134861
rect 271293 134593 271335 134829
rect 271571 134593 271613 134829
rect 271293 134509 271613 134593
rect 271293 134273 271335 134509
rect 271571 134273 271613 134509
rect 271293 134241 271613 134273
rect 275991 134829 276311 134861
rect 275991 134593 276033 134829
rect 276269 134593 276311 134829
rect 275991 134509 276311 134593
rect 275991 134273 276033 134509
rect 276269 134273 276311 134509
rect 275991 134241 276311 134273
rect 280689 134829 281009 134861
rect 280689 134593 280731 134829
rect 280967 134593 281009 134829
rect 280689 134509 281009 134593
rect 280689 134273 280731 134509
rect 280967 134273 281009 134509
rect 280689 134241 281009 134273
rect 285387 134829 285707 134861
rect 285387 134593 285429 134829
rect 285665 134593 285707 134829
rect 285387 134509 285707 134593
rect 285387 134273 285429 134509
rect 285665 134273 285707 134509
rect 285387 134241 285707 134273
rect 299293 134829 299613 134861
rect 299293 134593 299335 134829
rect 299571 134593 299613 134829
rect 299293 134509 299613 134593
rect 299293 134273 299335 134509
rect 299571 134273 299613 134509
rect 299293 134241 299613 134273
rect 303991 134829 304311 134861
rect 303991 134593 304033 134829
rect 304269 134593 304311 134829
rect 303991 134509 304311 134593
rect 303991 134273 304033 134509
rect 304269 134273 304311 134509
rect 303991 134241 304311 134273
rect 308689 134829 309009 134861
rect 308689 134593 308731 134829
rect 308967 134593 309009 134829
rect 308689 134509 309009 134593
rect 308689 134273 308731 134509
rect 308967 134273 309009 134509
rect 308689 134241 309009 134273
rect 313387 134829 313707 134861
rect 313387 134593 313429 134829
rect 313665 134593 313707 134829
rect 313387 134509 313707 134593
rect 313387 134273 313429 134509
rect 313665 134273 313707 134509
rect 313387 134241 313707 134273
rect 327293 134829 327613 134861
rect 327293 134593 327335 134829
rect 327571 134593 327613 134829
rect 327293 134509 327613 134593
rect 327293 134273 327335 134509
rect 327571 134273 327613 134509
rect 327293 134241 327613 134273
rect 331991 134829 332311 134861
rect 331991 134593 332033 134829
rect 332269 134593 332311 134829
rect 331991 134509 332311 134593
rect 331991 134273 332033 134509
rect 332269 134273 332311 134509
rect 331991 134241 332311 134273
rect 336689 134829 337009 134861
rect 336689 134593 336731 134829
rect 336967 134593 337009 134829
rect 336689 134509 337009 134593
rect 336689 134273 336731 134509
rect 336967 134273 337009 134509
rect 336689 134241 337009 134273
rect 341387 134829 341707 134861
rect 341387 134593 341429 134829
rect 341665 134593 341707 134829
rect 341387 134509 341707 134593
rect 341387 134273 341429 134509
rect 341665 134273 341707 134509
rect 341387 134241 341707 134273
rect 355293 134829 355613 134861
rect 355293 134593 355335 134829
rect 355571 134593 355613 134829
rect 355293 134509 355613 134593
rect 355293 134273 355335 134509
rect 355571 134273 355613 134509
rect 355293 134241 355613 134273
rect 359991 134829 360311 134861
rect 359991 134593 360033 134829
rect 360269 134593 360311 134829
rect 359991 134509 360311 134593
rect 359991 134273 360033 134509
rect 360269 134273 360311 134509
rect 359991 134241 360311 134273
rect 77642 131454 77962 131486
rect 77642 131218 77684 131454
rect 77920 131218 77962 131454
rect 77642 131134 77962 131218
rect 77642 130898 77684 131134
rect 77920 130898 77962 131134
rect 77642 130866 77962 130898
rect 82340 131454 82660 131486
rect 82340 131218 82382 131454
rect 82618 131218 82660 131454
rect 82340 131134 82660 131218
rect 82340 130898 82382 131134
rect 82618 130898 82660 131134
rect 82340 130866 82660 130898
rect 87038 131454 87358 131486
rect 87038 131218 87080 131454
rect 87316 131218 87358 131454
rect 87038 131134 87358 131218
rect 87038 130898 87080 131134
rect 87316 130898 87358 131134
rect 87038 130866 87358 130898
rect 105642 131454 105962 131486
rect 105642 131218 105684 131454
rect 105920 131218 105962 131454
rect 105642 131134 105962 131218
rect 105642 130898 105684 131134
rect 105920 130898 105962 131134
rect 105642 130866 105962 130898
rect 110340 131454 110660 131486
rect 110340 131218 110382 131454
rect 110618 131218 110660 131454
rect 110340 131134 110660 131218
rect 110340 130898 110382 131134
rect 110618 130898 110660 131134
rect 110340 130866 110660 130898
rect 115038 131454 115358 131486
rect 115038 131218 115080 131454
rect 115316 131218 115358 131454
rect 115038 131134 115358 131218
rect 115038 130898 115080 131134
rect 115316 130898 115358 131134
rect 115038 130866 115358 130898
rect 133642 131454 133962 131486
rect 133642 131218 133684 131454
rect 133920 131218 133962 131454
rect 133642 131134 133962 131218
rect 133642 130898 133684 131134
rect 133920 130898 133962 131134
rect 133642 130866 133962 130898
rect 138340 131454 138660 131486
rect 138340 131218 138382 131454
rect 138618 131218 138660 131454
rect 138340 131134 138660 131218
rect 138340 130898 138382 131134
rect 138618 130898 138660 131134
rect 138340 130866 138660 130898
rect 143038 131454 143358 131486
rect 143038 131218 143080 131454
rect 143316 131218 143358 131454
rect 143038 131134 143358 131218
rect 143038 130898 143080 131134
rect 143316 130898 143358 131134
rect 143038 130866 143358 130898
rect 161642 131454 161962 131486
rect 161642 131218 161684 131454
rect 161920 131218 161962 131454
rect 161642 131134 161962 131218
rect 161642 130898 161684 131134
rect 161920 130898 161962 131134
rect 161642 130866 161962 130898
rect 166340 131454 166660 131486
rect 166340 131218 166382 131454
rect 166618 131218 166660 131454
rect 166340 131134 166660 131218
rect 166340 130898 166382 131134
rect 166618 130898 166660 131134
rect 166340 130866 166660 130898
rect 171038 131454 171358 131486
rect 171038 131218 171080 131454
rect 171316 131218 171358 131454
rect 171038 131134 171358 131218
rect 171038 130898 171080 131134
rect 171316 130898 171358 131134
rect 171038 130866 171358 130898
rect 189642 131454 189962 131486
rect 189642 131218 189684 131454
rect 189920 131218 189962 131454
rect 189642 131134 189962 131218
rect 189642 130898 189684 131134
rect 189920 130898 189962 131134
rect 189642 130866 189962 130898
rect 194340 131454 194660 131486
rect 194340 131218 194382 131454
rect 194618 131218 194660 131454
rect 194340 131134 194660 131218
rect 194340 130898 194382 131134
rect 194618 130898 194660 131134
rect 194340 130866 194660 130898
rect 199038 131454 199358 131486
rect 199038 131218 199080 131454
rect 199316 131218 199358 131454
rect 199038 131134 199358 131218
rect 199038 130898 199080 131134
rect 199316 130898 199358 131134
rect 199038 130866 199358 130898
rect 217642 131454 217962 131486
rect 217642 131218 217684 131454
rect 217920 131218 217962 131454
rect 217642 131134 217962 131218
rect 217642 130898 217684 131134
rect 217920 130898 217962 131134
rect 217642 130866 217962 130898
rect 222340 131454 222660 131486
rect 222340 131218 222382 131454
rect 222618 131218 222660 131454
rect 222340 131134 222660 131218
rect 222340 130898 222382 131134
rect 222618 130898 222660 131134
rect 222340 130866 222660 130898
rect 227038 131454 227358 131486
rect 227038 131218 227080 131454
rect 227316 131218 227358 131454
rect 227038 131134 227358 131218
rect 227038 130898 227080 131134
rect 227316 130898 227358 131134
rect 227038 130866 227358 130898
rect 245642 131454 245962 131486
rect 245642 131218 245684 131454
rect 245920 131218 245962 131454
rect 245642 131134 245962 131218
rect 245642 130898 245684 131134
rect 245920 130898 245962 131134
rect 245642 130866 245962 130898
rect 250340 131454 250660 131486
rect 250340 131218 250382 131454
rect 250618 131218 250660 131454
rect 250340 131134 250660 131218
rect 250340 130898 250382 131134
rect 250618 130898 250660 131134
rect 250340 130866 250660 130898
rect 255038 131454 255358 131486
rect 255038 131218 255080 131454
rect 255316 131218 255358 131454
rect 255038 131134 255358 131218
rect 255038 130898 255080 131134
rect 255316 130898 255358 131134
rect 255038 130866 255358 130898
rect 273642 131454 273962 131486
rect 273642 131218 273684 131454
rect 273920 131218 273962 131454
rect 273642 131134 273962 131218
rect 273642 130898 273684 131134
rect 273920 130898 273962 131134
rect 273642 130866 273962 130898
rect 278340 131454 278660 131486
rect 278340 131218 278382 131454
rect 278618 131218 278660 131454
rect 278340 131134 278660 131218
rect 278340 130898 278382 131134
rect 278618 130898 278660 131134
rect 278340 130866 278660 130898
rect 283038 131454 283358 131486
rect 283038 131218 283080 131454
rect 283316 131218 283358 131454
rect 283038 131134 283358 131218
rect 283038 130898 283080 131134
rect 283316 130898 283358 131134
rect 283038 130866 283358 130898
rect 301642 131454 301962 131486
rect 301642 131218 301684 131454
rect 301920 131218 301962 131454
rect 301642 131134 301962 131218
rect 301642 130898 301684 131134
rect 301920 130898 301962 131134
rect 301642 130866 301962 130898
rect 306340 131454 306660 131486
rect 306340 131218 306382 131454
rect 306618 131218 306660 131454
rect 306340 131134 306660 131218
rect 306340 130898 306382 131134
rect 306618 130898 306660 131134
rect 306340 130866 306660 130898
rect 311038 131454 311358 131486
rect 311038 131218 311080 131454
rect 311316 131218 311358 131454
rect 311038 131134 311358 131218
rect 311038 130898 311080 131134
rect 311316 130898 311358 131134
rect 311038 130866 311358 130898
rect 329642 131454 329962 131486
rect 329642 131218 329684 131454
rect 329920 131218 329962 131454
rect 329642 131134 329962 131218
rect 329642 130898 329684 131134
rect 329920 130898 329962 131134
rect 329642 130866 329962 130898
rect 334340 131454 334660 131486
rect 334340 131218 334382 131454
rect 334618 131218 334660 131454
rect 334340 131134 334660 131218
rect 334340 130898 334382 131134
rect 334618 130898 334660 131134
rect 334340 130866 334660 130898
rect 339038 131454 339358 131486
rect 339038 131218 339080 131454
rect 339316 131218 339358 131454
rect 339038 131134 339358 131218
rect 339038 130898 339080 131134
rect 339316 130898 339358 131134
rect 339038 130866 339358 130898
rect 357642 131454 357962 131486
rect 357642 131218 357684 131454
rect 357920 131218 357962 131454
rect 357642 131134 357962 131218
rect 357642 130898 357684 131134
rect 357920 130898 357962 131134
rect 357642 130866 357962 130898
rect 361622 122773 361682 144467
rect 364689 134829 365009 134861
rect 364689 134593 364731 134829
rect 364967 134593 365009 134829
rect 364689 134509 365009 134593
rect 364689 134273 364731 134509
rect 364967 134273 365009 134509
rect 364689 134241 365009 134273
rect 369387 134829 369707 134861
rect 369387 134593 369429 134829
rect 369665 134593 369707 134829
rect 369387 134509 369707 134593
rect 369387 134273 369429 134509
rect 369665 134273 369707 134509
rect 369387 134241 369707 134273
rect 383293 134829 383613 134861
rect 383293 134593 383335 134829
rect 383571 134593 383613 134829
rect 383293 134509 383613 134593
rect 383293 134273 383335 134509
rect 383571 134273 383613 134509
rect 383293 134241 383613 134273
rect 387991 134829 388311 134861
rect 387991 134593 388033 134829
rect 388269 134593 388311 134829
rect 387991 134509 388311 134593
rect 387991 134273 388033 134509
rect 388269 134273 388311 134509
rect 387991 134241 388311 134273
rect 392689 134829 393009 134861
rect 392689 134593 392731 134829
rect 392967 134593 393009 134829
rect 392689 134509 393009 134593
rect 392689 134273 392731 134509
rect 392967 134273 393009 134509
rect 392689 134241 393009 134273
rect 397387 134829 397707 134861
rect 397387 134593 397429 134829
rect 397665 134593 397707 134829
rect 397387 134509 397707 134593
rect 397387 134273 397429 134509
rect 397665 134273 397707 134509
rect 397387 134241 397707 134273
rect 411293 134829 411613 134861
rect 411293 134593 411335 134829
rect 411571 134593 411613 134829
rect 411293 134509 411613 134593
rect 411293 134273 411335 134509
rect 411571 134273 411613 134509
rect 411293 134241 411613 134273
rect 415991 134829 416311 134861
rect 415991 134593 416033 134829
rect 416269 134593 416311 134829
rect 415991 134509 416311 134593
rect 415991 134273 416033 134509
rect 416269 134273 416311 134509
rect 415991 134241 416311 134273
rect 420689 134829 421009 134861
rect 420689 134593 420731 134829
rect 420967 134593 421009 134829
rect 420689 134509 421009 134593
rect 420689 134273 420731 134509
rect 420967 134273 421009 134509
rect 420689 134241 421009 134273
rect 425387 134829 425707 134861
rect 425387 134593 425429 134829
rect 425665 134593 425707 134829
rect 425387 134509 425707 134593
rect 425387 134273 425429 134509
rect 425665 134273 425707 134509
rect 425387 134241 425707 134273
rect 439293 134829 439613 134861
rect 439293 134593 439335 134829
rect 439571 134593 439613 134829
rect 439293 134509 439613 134593
rect 439293 134273 439335 134509
rect 439571 134273 439613 134509
rect 439293 134241 439613 134273
rect 443991 134829 444311 134861
rect 443991 134593 444033 134829
rect 444269 134593 444311 134829
rect 443991 134509 444311 134593
rect 443991 134273 444033 134509
rect 444269 134273 444311 134509
rect 443991 134241 444311 134273
rect 362340 131454 362660 131486
rect 362340 131218 362382 131454
rect 362618 131218 362660 131454
rect 362340 131134 362660 131218
rect 362340 130898 362382 131134
rect 362618 130898 362660 131134
rect 362340 130866 362660 130898
rect 367038 131454 367358 131486
rect 367038 131218 367080 131454
rect 367316 131218 367358 131454
rect 367038 131134 367358 131218
rect 367038 130898 367080 131134
rect 367316 130898 367358 131134
rect 367038 130866 367358 130898
rect 385642 131454 385962 131486
rect 385642 131218 385684 131454
rect 385920 131218 385962 131454
rect 385642 131134 385962 131218
rect 385642 130898 385684 131134
rect 385920 130898 385962 131134
rect 385642 130866 385962 130898
rect 390340 131454 390660 131486
rect 390340 131218 390382 131454
rect 390618 131218 390660 131454
rect 390340 131134 390660 131218
rect 390340 130898 390382 131134
rect 390618 130898 390660 131134
rect 390340 130866 390660 130898
rect 395038 131454 395358 131486
rect 395038 131218 395080 131454
rect 395316 131218 395358 131454
rect 395038 131134 395358 131218
rect 395038 130898 395080 131134
rect 395316 130898 395358 131134
rect 395038 130866 395358 130898
rect 413642 131454 413962 131486
rect 413642 131218 413684 131454
rect 413920 131218 413962 131454
rect 413642 131134 413962 131218
rect 413642 130898 413684 131134
rect 413920 130898 413962 131134
rect 413642 130866 413962 130898
rect 418340 131454 418660 131486
rect 418340 131218 418382 131454
rect 418618 131218 418660 131454
rect 418340 131134 418660 131218
rect 418340 130898 418382 131134
rect 418618 130898 418660 131134
rect 418340 130866 418660 130898
rect 423038 131454 423358 131486
rect 423038 131218 423080 131454
rect 423316 131218 423358 131454
rect 423038 131134 423358 131218
rect 423038 130898 423080 131134
rect 423316 130898 423358 131134
rect 423038 130866 423358 130898
rect 441642 131454 441962 131486
rect 441642 131218 441684 131454
rect 441920 131218 441962 131454
rect 441642 131134 441962 131218
rect 441642 130898 441684 131134
rect 441920 130898 441962 131134
rect 441642 130866 441962 130898
rect 445710 122773 445770 144467
rect 448689 134829 449009 134861
rect 448689 134593 448731 134829
rect 448967 134593 449009 134829
rect 448689 134509 449009 134593
rect 448689 134273 448731 134509
rect 448967 134273 449009 134509
rect 448689 134241 449009 134273
rect 453387 134829 453707 134861
rect 453387 134593 453429 134829
rect 453665 134593 453707 134829
rect 453387 134509 453707 134593
rect 453387 134273 453429 134509
rect 453665 134273 453707 134509
rect 453387 134241 453707 134273
rect 467293 134829 467613 134861
rect 467293 134593 467335 134829
rect 467571 134593 467613 134829
rect 467293 134509 467613 134593
rect 467293 134273 467335 134509
rect 467571 134273 467613 134509
rect 467293 134241 467613 134273
rect 471991 134829 472311 134861
rect 471991 134593 472033 134829
rect 472269 134593 472311 134829
rect 471991 134509 472311 134593
rect 471991 134273 472033 134509
rect 472269 134273 472311 134509
rect 471991 134241 472311 134273
rect 476689 134829 477009 134861
rect 476689 134593 476731 134829
rect 476967 134593 477009 134829
rect 476689 134509 477009 134593
rect 476689 134273 476731 134509
rect 476967 134273 477009 134509
rect 476689 134241 477009 134273
rect 481387 134829 481707 134861
rect 481387 134593 481429 134829
rect 481665 134593 481707 134829
rect 481387 134509 481707 134593
rect 481387 134273 481429 134509
rect 481665 134273 481707 134509
rect 481387 134241 481707 134273
rect 495293 134829 495613 134861
rect 495293 134593 495335 134829
rect 495571 134593 495613 134829
rect 495293 134509 495613 134593
rect 495293 134273 495335 134509
rect 495571 134273 495613 134509
rect 495293 134241 495613 134273
rect 499991 134829 500311 134861
rect 499991 134593 500033 134829
rect 500269 134593 500311 134829
rect 499991 134509 500311 134593
rect 499991 134273 500033 134509
rect 500269 134273 500311 134509
rect 499991 134241 500311 134273
rect 504689 134829 505009 134861
rect 504689 134593 504731 134829
rect 504967 134593 505009 134829
rect 504689 134509 505009 134593
rect 504689 134273 504731 134509
rect 504967 134273 505009 134509
rect 504689 134241 505009 134273
rect 509387 134829 509707 134861
rect 509387 134593 509429 134829
rect 509665 134593 509707 134829
rect 509387 134509 509707 134593
rect 509387 134273 509429 134509
rect 509665 134273 509707 134509
rect 509387 134241 509707 134273
rect 523293 134829 523613 134861
rect 523293 134593 523335 134829
rect 523571 134593 523613 134829
rect 523293 134509 523613 134593
rect 523293 134273 523335 134509
rect 523571 134273 523613 134509
rect 523293 134241 523613 134273
rect 527991 134829 528311 134861
rect 527991 134593 528033 134829
rect 528269 134593 528311 134829
rect 527991 134509 528311 134593
rect 527991 134273 528033 134509
rect 528269 134273 528311 134509
rect 527991 134241 528311 134273
rect 532689 134829 533009 134861
rect 532689 134593 532731 134829
rect 532967 134593 533009 134829
rect 532689 134509 533009 134593
rect 532689 134273 532731 134509
rect 532967 134273 533009 134509
rect 532689 134241 533009 134273
rect 537387 134829 537707 134861
rect 537387 134593 537429 134829
rect 537665 134593 537707 134829
rect 537387 134509 537707 134593
rect 537387 134273 537429 134509
rect 537665 134273 537707 134509
rect 537387 134241 537707 134273
rect 551293 134829 551613 134861
rect 551293 134593 551335 134829
rect 551571 134593 551613 134829
rect 551293 134509 551613 134593
rect 551293 134273 551335 134509
rect 551571 134273 551613 134509
rect 551293 134241 551613 134273
rect 555991 134829 556311 134861
rect 555991 134593 556033 134829
rect 556269 134593 556311 134829
rect 555991 134509 556311 134593
rect 555991 134273 556033 134509
rect 556269 134273 556311 134509
rect 555991 134241 556311 134273
rect 560689 134829 561009 134861
rect 560689 134593 560731 134829
rect 560967 134593 561009 134829
rect 560689 134509 561009 134593
rect 560689 134273 560731 134509
rect 560967 134273 561009 134509
rect 560689 134241 561009 134273
rect 565387 134829 565707 134861
rect 565387 134593 565429 134829
rect 565665 134593 565707 134829
rect 565387 134509 565707 134593
rect 565387 134273 565429 134509
rect 565665 134273 565707 134509
rect 565387 134241 565707 134273
rect 573494 134829 574114 161273
rect 573494 134593 573526 134829
rect 573762 134593 573846 134829
rect 574082 134593 574114 134829
rect 573494 134509 574114 134593
rect 573494 134273 573526 134509
rect 573762 134273 573846 134509
rect 574082 134273 574114 134509
rect 446340 131454 446660 131486
rect 446340 131218 446382 131454
rect 446618 131218 446660 131454
rect 446340 131134 446660 131218
rect 446340 130898 446382 131134
rect 446618 130898 446660 131134
rect 446340 130866 446660 130898
rect 451038 131454 451358 131486
rect 451038 131218 451080 131454
rect 451316 131218 451358 131454
rect 451038 131134 451358 131218
rect 451038 130898 451080 131134
rect 451316 130898 451358 131134
rect 451038 130866 451358 130898
rect 469642 131454 469962 131486
rect 469642 131218 469684 131454
rect 469920 131218 469962 131454
rect 469642 131134 469962 131218
rect 469642 130898 469684 131134
rect 469920 130898 469962 131134
rect 469642 130866 469962 130898
rect 474340 131454 474660 131486
rect 474340 131218 474382 131454
rect 474618 131218 474660 131454
rect 474340 131134 474660 131218
rect 474340 130898 474382 131134
rect 474618 130898 474660 131134
rect 474340 130866 474660 130898
rect 479038 131454 479358 131486
rect 479038 131218 479080 131454
rect 479316 131218 479358 131454
rect 479038 131134 479358 131218
rect 479038 130898 479080 131134
rect 479316 130898 479358 131134
rect 479038 130866 479358 130898
rect 497642 131454 497962 131486
rect 497642 131218 497684 131454
rect 497920 131218 497962 131454
rect 497642 131134 497962 131218
rect 497642 130898 497684 131134
rect 497920 130898 497962 131134
rect 497642 130866 497962 130898
rect 502340 131454 502660 131486
rect 502340 131218 502382 131454
rect 502618 131218 502660 131454
rect 502340 131134 502660 131218
rect 502340 130898 502382 131134
rect 502618 130898 502660 131134
rect 502340 130866 502660 130898
rect 507038 131454 507358 131486
rect 507038 131218 507080 131454
rect 507316 131218 507358 131454
rect 507038 131134 507358 131218
rect 507038 130898 507080 131134
rect 507316 130898 507358 131134
rect 507038 130866 507358 130898
rect 525642 131454 525962 131486
rect 525642 131218 525684 131454
rect 525920 131218 525962 131454
rect 525642 131134 525962 131218
rect 525642 130898 525684 131134
rect 525920 130898 525962 131134
rect 525642 130866 525962 130898
rect 530340 131454 530660 131486
rect 530340 131218 530382 131454
rect 530618 131218 530660 131454
rect 530340 131134 530660 131218
rect 530340 130898 530382 131134
rect 530618 130898 530660 131134
rect 530340 130866 530660 130898
rect 535038 131454 535358 131486
rect 535038 131218 535080 131454
rect 535316 131218 535358 131454
rect 535038 131134 535358 131218
rect 535038 130898 535080 131134
rect 535316 130898 535358 131134
rect 535038 130866 535358 130898
rect 553642 131454 553962 131486
rect 553642 131218 553684 131454
rect 553920 131218 553962 131454
rect 553642 131134 553962 131218
rect 553642 130898 553684 131134
rect 553920 130898 553962 131134
rect 553642 130866 553962 130898
rect 558340 131454 558660 131486
rect 558340 131218 558382 131454
rect 558618 131218 558660 131454
rect 558340 131134 558660 131218
rect 558340 130898 558382 131134
rect 558618 130898 558660 131134
rect 558340 130866 558660 130898
rect 563038 131454 563358 131486
rect 563038 131218 563080 131454
rect 563316 131218 563358 131454
rect 563038 131134 563358 131218
rect 563038 130898 563080 131134
rect 563316 130898 563358 131134
rect 563038 130866 563358 130898
rect 361619 122772 361685 122773
rect 361619 122708 361620 122772
rect 361684 122708 361685 122772
rect 361619 122707 361685 122708
rect 445707 122772 445773 122773
rect 445707 122708 445708 122772
rect 445772 122708 445773 122772
rect 445707 122707 445773 122708
rect 194731 117332 194797 117333
rect 194731 117268 194732 117332
rect 194796 117268 194797 117332
rect 194731 117267 194797 117268
rect 324267 117332 324333 117333
rect 324267 117268 324268 117332
rect 324332 117268 324333 117332
rect 324267 117267 324333 117268
rect 176331 116380 176397 116381
rect 176331 116316 176332 116380
rect 176396 116316 176397 116380
rect 176331 116315 176397 116316
rect 92427 116244 92493 116245
rect 92427 116180 92428 116244
rect 92492 116180 92493 116244
rect 92427 116179 92493 116180
rect 148363 116244 148429 116245
rect 148363 116180 148364 116244
rect 148428 116180 148429 116244
rect 148363 116179 148429 116180
rect 64459 116108 64525 116109
rect 64459 116044 64460 116108
rect 64524 116044 64525 116108
rect 64459 116043 64525 116044
rect 64462 108357 64522 116043
rect 92430 108357 92490 116179
rect 148366 108357 148426 116179
rect 176334 108357 176394 116315
rect 64459 108356 64525 108357
rect 64459 108292 64460 108356
rect 64524 108292 64525 108356
rect 64459 108291 64525 108292
rect 92427 108356 92493 108357
rect 92427 108292 92428 108356
rect 92492 108292 92493 108356
rect 92427 108291 92493 108292
rect 148363 108356 148429 108357
rect 148363 108292 148364 108356
rect 148428 108292 148429 108356
rect 148363 108291 148429 108292
rect 176331 108356 176397 108357
rect 176331 108292 176332 108356
rect 176396 108292 176397 108356
rect 176331 108291 176397 108292
rect 75293 107829 75613 107861
rect 75293 107593 75335 107829
rect 75571 107593 75613 107829
rect 75293 107509 75613 107593
rect 75293 107273 75335 107509
rect 75571 107273 75613 107509
rect 75293 107241 75613 107273
rect 79991 107829 80311 107861
rect 79991 107593 80033 107829
rect 80269 107593 80311 107829
rect 79991 107509 80311 107593
rect 79991 107273 80033 107509
rect 80269 107273 80311 107509
rect 79991 107241 80311 107273
rect 84689 107829 85009 107861
rect 84689 107593 84731 107829
rect 84967 107593 85009 107829
rect 84689 107509 85009 107593
rect 84689 107273 84731 107509
rect 84967 107273 85009 107509
rect 84689 107241 85009 107273
rect 89387 107829 89707 107861
rect 89387 107593 89429 107829
rect 89665 107593 89707 107829
rect 89387 107509 89707 107593
rect 89387 107273 89429 107509
rect 89665 107273 89707 107509
rect 89387 107241 89707 107273
rect 103293 107829 103613 107861
rect 103293 107593 103335 107829
rect 103571 107593 103613 107829
rect 103293 107509 103613 107593
rect 103293 107273 103335 107509
rect 103571 107273 103613 107509
rect 103293 107241 103613 107273
rect 107991 107829 108311 107861
rect 107991 107593 108033 107829
rect 108269 107593 108311 107829
rect 107991 107509 108311 107593
rect 107991 107273 108033 107509
rect 108269 107273 108311 107509
rect 107991 107241 108311 107273
rect 112689 107829 113009 107861
rect 112689 107593 112731 107829
rect 112967 107593 113009 107829
rect 112689 107509 113009 107593
rect 112689 107273 112731 107509
rect 112967 107273 113009 107509
rect 112689 107241 113009 107273
rect 117387 107829 117707 107861
rect 117387 107593 117429 107829
rect 117665 107593 117707 107829
rect 117387 107509 117707 107593
rect 117387 107273 117429 107509
rect 117665 107273 117707 107509
rect 117387 107241 117707 107273
rect 131293 107829 131613 107861
rect 131293 107593 131335 107829
rect 131571 107593 131613 107829
rect 131293 107509 131613 107593
rect 131293 107273 131335 107509
rect 131571 107273 131613 107509
rect 131293 107241 131613 107273
rect 135991 107829 136311 107861
rect 135991 107593 136033 107829
rect 136269 107593 136311 107829
rect 135991 107509 136311 107593
rect 135991 107273 136033 107509
rect 136269 107273 136311 107509
rect 135991 107241 136311 107273
rect 140689 107829 141009 107861
rect 140689 107593 140731 107829
rect 140967 107593 141009 107829
rect 140689 107509 141009 107593
rect 140689 107273 140731 107509
rect 140967 107273 141009 107509
rect 140689 107241 141009 107273
rect 145387 107829 145707 107861
rect 145387 107593 145429 107829
rect 145665 107593 145707 107829
rect 145387 107509 145707 107593
rect 145387 107273 145429 107509
rect 145665 107273 145707 107509
rect 145387 107241 145707 107273
rect 159293 107829 159613 107861
rect 159293 107593 159335 107829
rect 159571 107593 159613 107829
rect 159293 107509 159613 107593
rect 159293 107273 159335 107509
rect 159571 107273 159613 107509
rect 159293 107241 159613 107273
rect 163991 107829 164311 107861
rect 163991 107593 164033 107829
rect 164269 107593 164311 107829
rect 163991 107509 164311 107593
rect 163991 107273 164033 107509
rect 164269 107273 164311 107509
rect 163991 107241 164311 107273
rect 168689 107829 169009 107861
rect 168689 107593 168731 107829
rect 168967 107593 169009 107829
rect 168689 107509 169009 107593
rect 168689 107273 168731 107509
rect 168967 107273 169009 107509
rect 168689 107241 169009 107273
rect 173387 107829 173707 107861
rect 173387 107593 173429 107829
rect 173665 107593 173707 107829
rect 173387 107509 173707 107593
rect 173387 107273 173429 107509
rect 173665 107273 173707 107509
rect 173387 107241 173707 107273
rect 187293 107829 187613 107861
rect 187293 107593 187335 107829
rect 187571 107593 187613 107829
rect 187293 107509 187613 107593
rect 187293 107273 187335 107509
rect 187571 107273 187613 107509
rect 187293 107241 187613 107273
rect 191991 107829 192311 107861
rect 191991 107593 192033 107829
rect 192269 107593 192311 107829
rect 191991 107509 192311 107593
rect 191991 107273 192033 107509
rect 192269 107273 192311 107509
rect 191991 107241 192311 107273
rect 77642 104454 77962 104486
rect 77642 104218 77684 104454
rect 77920 104218 77962 104454
rect 77642 104134 77962 104218
rect 77642 103898 77684 104134
rect 77920 103898 77962 104134
rect 77642 103866 77962 103898
rect 82340 104454 82660 104486
rect 82340 104218 82382 104454
rect 82618 104218 82660 104454
rect 82340 104134 82660 104218
rect 82340 103898 82382 104134
rect 82618 103898 82660 104134
rect 82340 103866 82660 103898
rect 87038 104454 87358 104486
rect 87038 104218 87080 104454
rect 87316 104218 87358 104454
rect 87038 104134 87358 104218
rect 87038 103898 87080 104134
rect 87316 103898 87358 104134
rect 87038 103866 87358 103898
rect 105642 104454 105962 104486
rect 105642 104218 105684 104454
rect 105920 104218 105962 104454
rect 105642 104134 105962 104218
rect 105642 103898 105684 104134
rect 105920 103898 105962 104134
rect 105642 103866 105962 103898
rect 110340 104454 110660 104486
rect 110340 104218 110382 104454
rect 110618 104218 110660 104454
rect 110340 104134 110660 104218
rect 110340 103898 110382 104134
rect 110618 103898 110660 104134
rect 110340 103866 110660 103898
rect 115038 104454 115358 104486
rect 115038 104218 115080 104454
rect 115316 104218 115358 104454
rect 115038 104134 115358 104218
rect 115038 103898 115080 104134
rect 115316 103898 115358 104134
rect 115038 103866 115358 103898
rect 133642 104454 133962 104486
rect 133642 104218 133684 104454
rect 133920 104218 133962 104454
rect 133642 104134 133962 104218
rect 133642 103898 133684 104134
rect 133920 103898 133962 104134
rect 133642 103866 133962 103898
rect 138340 104454 138660 104486
rect 138340 104218 138382 104454
rect 138618 104218 138660 104454
rect 138340 104134 138660 104218
rect 138340 103898 138382 104134
rect 138618 103898 138660 104134
rect 138340 103866 138660 103898
rect 143038 104454 143358 104486
rect 143038 104218 143080 104454
rect 143316 104218 143358 104454
rect 143038 104134 143358 104218
rect 143038 103898 143080 104134
rect 143316 103898 143358 104134
rect 143038 103866 143358 103898
rect 161642 104454 161962 104486
rect 161642 104218 161684 104454
rect 161920 104218 161962 104454
rect 161642 104134 161962 104218
rect 161642 103898 161684 104134
rect 161920 103898 161962 104134
rect 161642 103866 161962 103898
rect 166340 104454 166660 104486
rect 166340 104218 166382 104454
rect 166618 104218 166660 104454
rect 166340 104134 166660 104218
rect 166340 103898 166382 104134
rect 166618 103898 166660 104134
rect 166340 103866 166660 103898
rect 171038 104454 171358 104486
rect 171038 104218 171080 104454
rect 171316 104218 171358 104454
rect 171038 104134 171358 104218
rect 171038 103898 171080 104134
rect 171316 103898 171358 104134
rect 171038 103866 171358 103898
rect 189642 104454 189962 104486
rect 189642 104218 189684 104454
rect 189920 104218 189962 104454
rect 189642 104134 189962 104218
rect 189642 103898 189684 104134
rect 189920 103898 189962 104134
rect 189642 103866 189962 103898
rect 194340 104454 194660 104486
rect 194340 104218 194382 104454
rect 194618 104218 194660 104454
rect 194340 104134 194660 104218
rect 194340 103898 194382 104134
rect 194618 103898 194660 104134
rect 194340 103866 194660 103898
rect 194734 95165 194794 117267
rect 260419 116516 260485 116517
rect 260419 116452 260420 116516
rect 260484 116452 260485 116516
rect 260419 116451 260485 116452
rect 260422 108357 260482 116451
rect 260419 108356 260485 108357
rect 260419 108292 260420 108356
rect 260484 108292 260485 108356
rect 260419 108291 260485 108292
rect 196689 107829 197009 107861
rect 196689 107593 196731 107829
rect 196967 107593 197009 107829
rect 196689 107509 197009 107593
rect 196689 107273 196731 107509
rect 196967 107273 197009 107509
rect 196689 107241 197009 107273
rect 201387 107829 201707 107861
rect 201387 107593 201429 107829
rect 201665 107593 201707 107829
rect 201387 107509 201707 107593
rect 201387 107273 201429 107509
rect 201665 107273 201707 107509
rect 201387 107241 201707 107273
rect 215293 107829 215613 107861
rect 215293 107593 215335 107829
rect 215571 107593 215613 107829
rect 215293 107509 215613 107593
rect 215293 107273 215335 107509
rect 215571 107273 215613 107509
rect 215293 107241 215613 107273
rect 219991 107829 220311 107861
rect 219991 107593 220033 107829
rect 220269 107593 220311 107829
rect 219991 107509 220311 107593
rect 219991 107273 220033 107509
rect 220269 107273 220311 107509
rect 219991 107241 220311 107273
rect 224689 107829 225009 107861
rect 224689 107593 224731 107829
rect 224967 107593 225009 107829
rect 224689 107509 225009 107593
rect 224689 107273 224731 107509
rect 224967 107273 225009 107509
rect 224689 107241 225009 107273
rect 229387 107829 229707 107861
rect 229387 107593 229429 107829
rect 229665 107593 229707 107829
rect 229387 107509 229707 107593
rect 229387 107273 229429 107509
rect 229665 107273 229707 107509
rect 229387 107241 229707 107273
rect 244076 107829 244396 107861
rect 244076 107593 244118 107829
rect 244354 107593 244396 107829
rect 244076 107509 244396 107593
rect 244076 107273 244118 107509
rect 244354 107273 244396 107509
rect 244076 107241 244396 107273
rect 250340 107829 250660 107861
rect 250340 107593 250382 107829
rect 250618 107593 250660 107829
rect 250340 107509 250660 107593
rect 250340 107273 250382 107509
rect 250618 107273 250660 107509
rect 250340 107241 250660 107273
rect 256604 107829 256924 107861
rect 256604 107593 256646 107829
rect 256882 107593 256924 107829
rect 256604 107509 256924 107593
rect 256604 107273 256646 107509
rect 256882 107273 256924 107509
rect 256604 107241 256924 107273
rect 271293 107829 271613 107861
rect 271293 107593 271335 107829
rect 271571 107593 271613 107829
rect 271293 107509 271613 107593
rect 271293 107273 271335 107509
rect 271571 107273 271613 107509
rect 271293 107241 271613 107273
rect 275991 107829 276311 107861
rect 275991 107593 276033 107829
rect 276269 107593 276311 107829
rect 275991 107509 276311 107593
rect 275991 107273 276033 107509
rect 276269 107273 276311 107509
rect 275991 107241 276311 107273
rect 280689 107829 281009 107861
rect 280689 107593 280731 107829
rect 280967 107593 281009 107829
rect 280689 107509 281009 107593
rect 280689 107273 280731 107509
rect 280967 107273 281009 107509
rect 280689 107241 281009 107273
rect 285387 107829 285707 107861
rect 285387 107593 285429 107829
rect 285665 107593 285707 107829
rect 285387 107509 285707 107593
rect 285387 107273 285429 107509
rect 285665 107273 285707 107509
rect 285387 107241 285707 107273
rect 299293 107829 299613 107861
rect 299293 107593 299335 107829
rect 299571 107593 299613 107829
rect 299293 107509 299613 107593
rect 299293 107273 299335 107509
rect 299571 107273 299613 107509
rect 299293 107241 299613 107273
rect 303991 107829 304311 107861
rect 303991 107593 304033 107829
rect 304269 107593 304311 107829
rect 303991 107509 304311 107593
rect 303991 107273 304033 107509
rect 304269 107273 304311 107509
rect 303991 107241 304311 107273
rect 308689 107829 309009 107861
rect 308689 107593 308731 107829
rect 308967 107593 309009 107829
rect 308689 107509 309009 107593
rect 308689 107273 308731 107509
rect 308967 107273 309009 107509
rect 308689 107241 309009 107273
rect 313387 107829 313707 107861
rect 313387 107593 313429 107829
rect 313665 107593 313707 107829
rect 313387 107509 313707 107593
rect 313387 107273 313429 107509
rect 313665 107273 313707 107509
rect 313387 107241 313707 107273
rect 199038 104454 199358 104486
rect 199038 104218 199080 104454
rect 199316 104218 199358 104454
rect 199038 104134 199358 104218
rect 199038 103898 199080 104134
rect 199316 103898 199358 104134
rect 199038 103866 199358 103898
rect 217642 104454 217962 104486
rect 217642 104218 217684 104454
rect 217920 104218 217962 104454
rect 217642 104134 217962 104218
rect 217642 103898 217684 104134
rect 217920 103898 217962 104134
rect 217642 103866 217962 103898
rect 222340 104454 222660 104486
rect 222340 104218 222382 104454
rect 222618 104218 222660 104454
rect 222340 104134 222660 104218
rect 222340 103898 222382 104134
rect 222618 103898 222660 104134
rect 222340 103866 222660 103898
rect 227038 104454 227358 104486
rect 227038 104218 227080 104454
rect 227316 104218 227358 104454
rect 227038 104134 227358 104218
rect 227038 103898 227080 104134
rect 227316 103898 227358 104134
rect 227038 103866 227358 103898
rect 247208 104454 247528 104486
rect 247208 104218 247250 104454
rect 247486 104218 247528 104454
rect 247208 104134 247528 104218
rect 247208 103898 247250 104134
rect 247486 103898 247528 104134
rect 247208 103866 247528 103898
rect 253472 104454 253792 104486
rect 253472 104218 253514 104454
rect 253750 104218 253792 104454
rect 253472 104134 253792 104218
rect 253472 103898 253514 104134
rect 253750 103898 253792 104134
rect 253472 103866 253792 103898
rect 273642 104454 273962 104486
rect 273642 104218 273684 104454
rect 273920 104218 273962 104454
rect 273642 104134 273962 104218
rect 273642 103898 273684 104134
rect 273920 103898 273962 104134
rect 273642 103866 273962 103898
rect 278340 104454 278660 104486
rect 278340 104218 278382 104454
rect 278618 104218 278660 104454
rect 278340 104134 278660 104218
rect 278340 103898 278382 104134
rect 278618 103898 278660 104134
rect 278340 103866 278660 103898
rect 283038 104454 283358 104486
rect 283038 104218 283080 104454
rect 283316 104218 283358 104454
rect 283038 104134 283358 104218
rect 283038 103898 283080 104134
rect 283316 103898 283358 104134
rect 283038 103866 283358 103898
rect 301642 104454 301962 104486
rect 301642 104218 301684 104454
rect 301920 104218 301962 104454
rect 301642 104134 301962 104218
rect 301642 103898 301684 104134
rect 301920 103898 301962 104134
rect 301642 103866 301962 103898
rect 306340 104454 306660 104486
rect 306340 104218 306382 104454
rect 306618 104218 306660 104454
rect 306340 104134 306660 104218
rect 306340 103898 306382 104134
rect 306618 103898 306660 104134
rect 306340 103866 306660 103898
rect 311038 104454 311358 104486
rect 311038 104218 311080 104454
rect 311316 104218 311358 104454
rect 311038 104134 311358 104218
rect 311038 103898 311080 104134
rect 311316 103898 311358 104134
rect 311038 103866 311358 103898
rect 324270 95165 324330 117267
rect 540467 116244 540533 116245
rect 540467 116180 540468 116244
rect 540532 116180 540533 116244
rect 540467 116179 540533 116180
rect 408539 116108 408605 116109
rect 408539 116044 408540 116108
rect 408604 116044 408605 116108
rect 408539 116043 408605 116044
rect 520595 116108 520661 116109
rect 520595 116044 520596 116108
rect 520660 116044 520661 116108
rect 520595 116043 520661 116044
rect 408542 108357 408602 116043
rect 520598 108357 520658 116043
rect 540470 108357 540530 116179
rect 408539 108356 408605 108357
rect 408539 108292 408540 108356
rect 408604 108292 408605 108356
rect 408539 108291 408605 108292
rect 520595 108356 520661 108357
rect 520595 108292 520596 108356
rect 520660 108292 520661 108356
rect 520595 108291 520661 108292
rect 540467 108356 540533 108357
rect 540467 108292 540468 108356
rect 540532 108292 540533 108356
rect 540467 108291 540533 108292
rect 328076 107829 328396 107861
rect 328076 107593 328118 107829
rect 328354 107593 328396 107829
rect 328076 107509 328396 107593
rect 328076 107273 328118 107509
rect 328354 107273 328396 107509
rect 328076 107241 328396 107273
rect 334340 107829 334660 107861
rect 334340 107593 334382 107829
rect 334618 107593 334660 107829
rect 334340 107509 334660 107593
rect 334340 107273 334382 107509
rect 334618 107273 334660 107509
rect 334340 107241 334660 107273
rect 340604 107829 340924 107861
rect 340604 107593 340646 107829
rect 340882 107593 340924 107829
rect 340604 107509 340924 107593
rect 340604 107273 340646 107509
rect 340882 107273 340924 107509
rect 340604 107241 340924 107273
rect 355293 107829 355613 107861
rect 355293 107593 355335 107829
rect 355571 107593 355613 107829
rect 355293 107509 355613 107593
rect 355293 107273 355335 107509
rect 355571 107273 355613 107509
rect 355293 107241 355613 107273
rect 359991 107829 360311 107861
rect 359991 107593 360033 107829
rect 360269 107593 360311 107829
rect 359991 107509 360311 107593
rect 359991 107273 360033 107509
rect 360269 107273 360311 107509
rect 359991 107241 360311 107273
rect 364689 107829 365009 107861
rect 364689 107593 364731 107829
rect 364967 107593 365009 107829
rect 364689 107509 365009 107593
rect 364689 107273 364731 107509
rect 364967 107273 365009 107509
rect 364689 107241 365009 107273
rect 369387 107829 369707 107861
rect 369387 107593 369429 107829
rect 369665 107593 369707 107829
rect 369387 107509 369707 107593
rect 369387 107273 369429 107509
rect 369665 107273 369707 107509
rect 369387 107241 369707 107273
rect 383293 107829 383613 107861
rect 383293 107593 383335 107829
rect 383571 107593 383613 107829
rect 383293 107509 383613 107593
rect 383293 107273 383335 107509
rect 383571 107273 383613 107509
rect 383293 107241 383613 107273
rect 387991 107829 388311 107861
rect 387991 107593 388033 107829
rect 388269 107593 388311 107829
rect 387991 107509 388311 107593
rect 387991 107273 388033 107509
rect 388269 107273 388311 107509
rect 387991 107241 388311 107273
rect 392689 107829 393009 107861
rect 392689 107593 392731 107829
rect 392967 107593 393009 107829
rect 392689 107509 393009 107593
rect 392689 107273 392731 107509
rect 392967 107273 393009 107509
rect 392689 107241 393009 107273
rect 397387 107829 397707 107861
rect 397387 107593 397429 107829
rect 397665 107593 397707 107829
rect 397387 107509 397707 107593
rect 397387 107273 397429 107509
rect 397665 107273 397707 107509
rect 397387 107241 397707 107273
rect 411293 107829 411613 107861
rect 411293 107593 411335 107829
rect 411571 107593 411613 107829
rect 411293 107509 411613 107593
rect 411293 107273 411335 107509
rect 411571 107273 411613 107509
rect 411293 107241 411613 107273
rect 415991 107829 416311 107861
rect 415991 107593 416033 107829
rect 416269 107593 416311 107829
rect 415991 107509 416311 107593
rect 415991 107273 416033 107509
rect 416269 107273 416311 107509
rect 415991 107241 416311 107273
rect 420689 107829 421009 107861
rect 420689 107593 420731 107829
rect 420967 107593 421009 107829
rect 420689 107509 421009 107593
rect 420689 107273 420731 107509
rect 420967 107273 421009 107509
rect 420689 107241 421009 107273
rect 425387 107829 425707 107861
rect 425387 107593 425429 107829
rect 425665 107593 425707 107829
rect 425387 107509 425707 107593
rect 425387 107273 425429 107509
rect 425665 107273 425707 107509
rect 425387 107241 425707 107273
rect 439293 107829 439613 107861
rect 439293 107593 439335 107829
rect 439571 107593 439613 107829
rect 439293 107509 439613 107593
rect 439293 107273 439335 107509
rect 439571 107273 439613 107509
rect 439293 107241 439613 107273
rect 443991 107829 444311 107861
rect 443991 107593 444033 107829
rect 444269 107593 444311 107829
rect 443991 107509 444311 107593
rect 443991 107273 444033 107509
rect 444269 107273 444311 107509
rect 443991 107241 444311 107273
rect 448689 107829 449009 107861
rect 448689 107593 448731 107829
rect 448967 107593 449009 107829
rect 448689 107509 449009 107593
rect 448689 107273 448731 107509
rect 448967 107273 449009 107509
rect 448689 107241 449009 107273
rect 453387 107829 453707 107861
rect 453387 107593 453429 107829
rect 453665 107593 453707 107829
rect 453387 107509 453707 107593
rect 453387 107273 453429 107509
rect 453665 107273 453707 107509
rect 453387 107241 453707 107273
rect 467293 107829 467613 107861
rect 467293 107593 467335 107829
rect 467571 107593 467613 107829
rect 467293 107509 467613 107593
rect 467293 107273 467335 107509
rect 467571 107273 467613 107509
rect 467293 107241 467613 107273
rect 471991 107829 472311 107861
rect 471991 107593 472033 107829
rect 472269 107593 472311 107829
rect 471991 107509 472311 107593
rect 471991 107273 472033 107509
rect 472269 107273 472311 107509
rect 471991 107241 472311 107273
rect 476689 107829 477009 107861
rect 476689 107593 476731 107829
rect 476967 107593 477009 107829
rect 476689 107509 477009 107593
rect 476689 107273 476731 107509
rect 476967 107273 477009 107509
rect 476689 107241 477009 107273
rect 481387 107829 481707 107861
rect 481387 107593 481429 107829
rect 481665 107593 481707 107829
rect 481387 107509 481707 107593
rect 481387 107273 481429 107509
rect 481665 107273 481707 107509
rect 481387 107241 481707 107273
rect 495293 107829 495613 107861
rect 495293 107593 495335 107829
rect 495571 107593 495613 107829
rect 495293 107509 495613 107593
rect 495293 107273 495335 107509
rect 495571 107273 495613 107509
rect 495293 107241 495613 107273
rect 499991 107829 500311 107861
rect 499991 107593 500033 107829
rect 500269 107593 500311 107829
rect 499991 107509 500311 107593
rect 499991 107273 500033 107509
rect 500269 107273 500311 107509
rect 499991 107241 500311 107273
rect 504689 107829 505009 107861
rect 504689 107593 504731 107829
rect 504967 107593 505009 107829
rect 504689 107509 505009 107593
rect 504689 107273 504731 107509
rect 504967 107273 505009 107509
rect 504689 107241 505009 107273
rect 509387 107829 509707 107861
rect 509387 107593 509429 107829
rect 509665 107593 509707 107829
rect 509387 107509 509707 107593
rect 509387 107273 509429 107509
rect 509665 107273 509707 107509
rect 509387 107241 509707 107273
rect 523293 107829 523613 107861
rect 523293 107593 523335 107829
rect 523571 107593 523613 107829
rect 523293 107509 523613 107593
rect 523293 107273 523335 107509
rect 523571 107273 523613 107509
rect 523293 107241 523613 107273
rect 527991 107829 528311 107861
rect 527991 107593 528033 107829
rect 528269 107593 528311 107829
rect 527991 107509 528311 107593
rect 527991 107273 528033 107509
rect 528269 107273 528311 107509
rect 527991 107241 528311 107273
rect 532689 107829 533009 107861
rect 532689 107593 532731 107829
rect 532967 107593 533009 107829
rect 532689 107509 533009 107593
rect 532689 107273 532731 107509
rect 532967 107273 533009 107509
rect 532689 107241 533009 107273
rect 537387 107829 537707 107861
rect 537387 107593 537429 107829
rect 537665 107593 537707 107829
rect 537387 107509 537707 107593
rect 537387 107273 537429 107509
rect 537665 107273 537707 107509
rect 537387 107241 537707 107273
rect 551293 107829 551613 107861
rect 551293 107593 551335 107829
rect 551571 107593 551613 107829
rect 551293 107509 551613 107593
rect 551293 107273 551335 107509
rect 551571 107273 551613 107509
rect 551293 107241 551613 107273
rect 555991 107829 556311 107861
rect 555991 107593 556033 107829
rect 556269 107593 556311 107829
rect 555991 107509 556311 107593
rect 555991 107273 556033 107509
rect 556269 107273 556311 107509
rect 555991 107241 556311 107273
rect 560689 107829 561009 107861
rect 560689 107593 560731 107829
rect 560967 107593 561009 107829
rect 560689 107509 561009 107593
rect 560689 107273 560731 107509
rect 560967 107273 561009 107509
rect 560689 107241 561009 107273
rect 565387 107829 565707 107861
rect 565387 107593 565429 107829
rect 565665 107593 565707 107829
rect 565387 107509 565707 107593
rect 565387 107273 565429 107509
rect 565665 107273 565707 107509
rect 565387 107241 565707 107273
rect 573494 107829 574114 134273
rect 573494 107593 573526 107829
rect 573762 107593 573846 107829
rect 574082 107593 574114 107829
rect 573494 107509 574114 107593
rect 573494 107273 573526 107509
rect 573762 107273 573846 107509
rect 574082 107273 574114 107509
rect 331208 104454 331528 104486
rect 331208 104218 331250 104454
rect 331486 104218 331528 104454
rect 331208 104134 331528 104218
rect 331208 103898 331250 104134
rect 331486 103898 331528 104134
rect 331208 103866 331528 103898
rect 337472 104454 337792 104486
rect 337472 104218 337514 104454
rect 337750 104218 337792 104454
rect 337472 104134 337792 104218
rect 337472 103898 337514 104134
rect 337750 103898 337792 104134
rect 337472 103866 337792 103898
rect 357642 104454 357962 104486
rect 357642 104218 357684 104454
rect 357920 104218 357962 104454
rect 357642 104134 357962 104218
rect 357642 103898 357684 104134
rect 357920 103898 357962 104134
rect 357642 103866 357962 103898
rect 362340 104454 362660 104486
rect 362340 104218 362382 104454
rect 362618 104218 362660 104454
rect 362340 104134 362660 104218
rect 362340 103898 362382 104134
rect 362618 103898 362660 104134
rect 362340 103866 362660 103898
rect 367038 104454 367358 104486
rect 367038 104218 367080 104454
rect 367316 104218 367358 104454
rect 367038 104134 367358 104218
rect 367038 103898 367080 104134
rect 367316 103898 367358 104134
rect 367038 103866 367358 103898
rect 385642 104454 385962 104486
rect 385642 104218 385684 104454
rect 385920 104218 385962 104454
rect 385642 104134 385962 104218
rect 385642 103898 385684 104134
rect 385920 103898 385962 104134
rect 385642 103866 385962 103898
rect 390340 104454 390660 104486
rect 390340 104218 390382 104454
rect 390618 104218 390660 104454
rect 390340 104134 390660 104218
rect 390340 103898 390382 104134
rect 390618 103898 390660 104134
rect 390340 103866 390660 103898
rect 395038 104454 395358 104486
rect 395038 104218 395080 104454
rect 395316 104218 395358 104454
rect 395038 104134 395358 104218
rect 395038 103898 395080 104134
rect 395316 103898 395358 104134
rect 395038 103866 395358 103898
rect 413642 104454 413962 104486
rect 413642 104218 413684 104454
rect 413920 104218 413962 104454
rect 413642 104134 413962 104218
rect 413642 103898 413684 104134
rect 413920 103898 413962 104134
rect 413642 103866 413962 103898
rect 418340 104454 418660 104486
rect 418340 104218 418382 104454
rect 418618 104218 418660 104454
rect 418340 104134 418660 104218
rect 418340 103898 418382 104134
rect 418618 103898 418660 104134
rect 418340 103866 418660 103898
rect 423038 104454 423358 104486
rect 423038 104218 423080 104454
rect 423316 104218 423358 104454
rect 423038 104134 423358 104218
rect 423038 103898 423080 104134
rect 423316 103898 423358 104134
rect 423038 103866 423358 103898
rect 441642 104454 441962 104486
rect 441642 104218 441684 104454
rect 441920 104218 441962 104454
rect 441642 104134 441962 104218
rect 441642 103898 441684 104134
rect 441920 103898 441962 104134
rect 441642 103866 441962 103898
rect 446340 104454 446660 104486
rect 446340 104218 446382 104454
rect 446618 104218 446660 104454
rect 446340 104134 446660 104218
rect 446340 103898 446382 104134
rect 446618 103898 446660 104134
rect 446340 103866 446660 103898
rect 451038 104454 451358 104486
rect 451038 104218 451080 104454
rect 451316 104218 451358 104454
rect 451038 104134 451358 104218
rect 451038 103898 451080 104134
rect 451316 103898 451358 104134
rect 451038 103866 451358 103898
rect 469642 104454 469962 104486
rect 469642 104218 469684 104454
rect 469920 104218 469962 104454
rect 469642 104134 469962 104218
rect 469642 103898 469684 104134
rect 469920 103898 469962 104134
rect 469642 103866 469962 103898
rect 474340 104454 474660 104486
rect 474340 104218 474382 104454
rect 474618 104218 474660 104454
rect 474340 104134 474660 104218
rect 474340 103898 474382 104134
rect 474618 103898 474660 104134
rect 474340 103866 474660 103898
rect 479038 104454 479358 104486
rect 479038 104218 479080 104454
rect 479316 104218 479358 104454
rect 479038 104134 479358 104218
rect 479038 103898 479080 104134
rect 479316 103898 479358 104134
rect 479038 103866 479358 103898
rect 497642 104454 497962 104486
rect 497642 104218 497684 104454
rect 497920 104218 497962 104454
rect 497642 104134 497962 104218
rect 497642 103898 497684 104134
rect 497920 103898 497962 104134
rect 497642 103866 497962 103898
rect 502340 104454 502660 104486
rect 502340 104218 502382 104454
rect 502618 104218 502660 104454
rect 502340 104134 502660 104218
rect 502340 103898 502382 104134
rect 502618 103898 502660 104134
rect 502340 103866 502660 103898
rect 507038 104454 507358 104486
rect 507038 104218 507080 104454
rect 507316 104218 507358 104454
rect 507038 104134 507358 104218
rect 507038 103898 507080 104134
rect 507316 103898 507358 104134
rect 507038 103866 507358 103898
rect 525642 104454 525962 104486
rect 525642 104218 525684 104454
rect 525920 104218 525962 104454
rect 525642 104134 525962 104218
rect 525642 103898 525684 104134
rect 525920 103898 525962 104134
rect 525642 103866 525962 103898
rect 530340 104454 530660 104486
rect 530340 104218 530382 104454
rect 530618 104218 530660 104454
rect 530340 104134 530660 104218
rect 530340 103898 530382 104134
rect 530618 103898 530660 104134
rect 530340 103866 530660 103898
rect 535038 104454 535358 104486
rect 535038 104218 535080 104454
rect 535316 104218 535358 104454
rect 535038 104134 535358 104218
rect 535038 103898 535080 104134
rect 535316 103898 535358 104134
rect 535038 103866 535358 103898
rect 553642 104454 553962 104486
rect 553642 104218 553684 104454
rect 553920 104218 553962 104454
rect 553642 104134 553962 104218
rect 553642 103898 553684 104134
rect 553920 103898 553962 104134
rect 553642 103866 553962 103898
rect 558340 104454 558660 104486
rect 558340 104218 558382 104454
rect 558618 104218 558660 104454
rect 558340 104134 558660 104218
rect 558340 103898 558382 104134
rect 558618 103898 558660 104134
rect 558340 103866 558660 103898
rect 563038 104454 563358 104486
rect 563038 104218 563080 104454
rect 563316 104218 563358 104454
rect 563038 104134 563358 104218
rect 563038 103898 563080 104134
rect 563316 103898 563358 104134
rect 563038 103866 563358 103898
rect 194731 95164 194797 95165
rect 194731 95100 194732 95164
rect 194796 95100 194797 95164
rect 194731 95099 194797 95100
rect 324267 95164 324333 95165
rect 324267 95100 324268 95164
rect 324332 95100 324333 95164
rect 324267 95099 324333 95100
rect 372291 89044 372357 89045
rect 372291 88980 372292 89044
rect 372356 88980 372357 89044
rect 372291 88979 372357 88980
rect 288387 88908 288453 88909
rect 288387 88844 288388 88908
rect 288452 88844 288453 88908
rect 288387 88843 288453 88844
rect 296851 88908 296917 88909
rect 296851 88844 296852 88908
rect 296916 88844 296917 88908
rect 296851 88843 296917 88844
rect 176331 88772 176397 88773
rect 176331 88708 176332 88772
rect 176396 88708 176397 88772
rect 176331 88707 176397 88708
rect 176334 80885 176394 88707
rect 288390 80885 288450 88843
rect 296854 86970 296914 88843
rect 296486 86910 296914 86970
rect 296486 80885 296546 86910
rect 372294 80885 372354 88979
rect 484347 88908 484413 88909
rect 484347 88844 484348 88908
rect 484412 88844 484413 88908
rect 484347 88843 484413 88844
rect 484350 80885 484410 88843
rect 520595 88772 520661 88773
rect 520595 88708 520596 88772
rect 520660 88708 520661 88772
rect 520595 88707 520661 88708
rect 520598 80885 520658 88707
rect 176331 80884 176397 80885
rect 76076 80829 76396 80861
rect 76076 80593 76118 80829
rect 76354 80593 76396 80829
rect 76076 80509 76396 80593
rect 76076 80273 76118 80509
rect 76354 80273 76396 80509
rect 76076 80241 76396 80273
rect 82340 80829 82660 80861
rect 82340 80593 82382 80829
rect 82618 80593 82660 80829
rect 82340 80509 82660 80593
rect 82340 80273 82382 80509
rect 82618 80273 82660 80509
rect 82340 80241 82660 80273
rect 88604 80829 88924 80861
rect 88604 80593 88646 80829
rect 88882 80593 88924 80829
rect 88604 80509 88924 80593
rect 88604 80273 88646 80509
rect 88882 80273 88924 80509
rect 88604 80241 88924 80273
rect 103293 80829 103613 80861
rect 103293 80593 103335 80829
rect 103571 80593 103613 80829
rect 103293 80509 103613 80593
rect 103293 80273 103335 80509
rect 103571 80273 103613 80509
rect 103293 80241 103613 80273
rect 107991 80829 108311 80861
rect 107991 80593 108033 80829
rect 108269 80593 108311 80829
rect 107991 80509 108311 80593
rect 107991 80273 108033 80509
rect 108269 80273 108311 80509
rect 107991 80241 108311 80273
rect 112689 80829 113009 80861
rect 112689 80593 112731 80829
rect 112967 80593 113009 80829
rect 112689 80509 113009 80593
rect 112689 80273 112731 80509
rect 112967 80273 113009 80509
rect 112689 80241 113009 80273
rect 117387 80829 117707 80861
rect 117387 80593 117429 80829
rect 117665 80593 117707 80829
rect 117387 80509 117707 80593
rect 117387 80273 117429 80509
rect 117665 80273 117707 80509
rect 117387 80241 117707 80273
rect 131293 80829 131613 80861
rect 131293 80593 131335 80829
rect 131571 80593 131613 80829
rect 131293 80509 131613 80593
rect 131293 80273 131335 80509
rect 131571 80273 131613 80509
rect 131293 80241 131613 80273
rect 135991 80829 136311 80861
rect 135991 80593 136033 80829
rect 136269 80593 136311 80829
rect 135991 80509 136311 80593
rect 135991 80273 136033 80509
rect 136269 80273 136311 80509
rect 135991 80241 136311 80273
rect 140689 80829 141009 80861
rect 140689 80593 140731 80829
rect 140967 80593 141009 80829
rect 140689 80509 141009 80593
rect 140689 80273 140731 80509
rect 140967 80273 141009 80509
rect 140689 80241 141009 80273
rect 145387 80829 145707 80861
rect 145387 80593 145429 80829
rect 145665 80593 145707 80829
rect 145387 80509 145707 80593
rect 145387 80273 145429 80509
rect 145665 80273 145707 80509
rect 145387 80241 145707 80273
rect 159293 80829 159613 80861
rect 159293 80593 159335 80829
rect 159571 80593 159613 80829
rect 159293 80509 159613 80593
rect 159293 80273 159335 80509
rect 159571 80273 159613 80509
rect 159293 80241 159613 80273
rect 163991 80829 164311 80861
rect 163991 80593 164033 80829
rect 164269 80593 164311 80829
rect 163991 80509 164311 80593
rect 163991 80273 164033 80509
rect 164269 80273 164311 80509
rect 163991 80241 164311 80273
rect 168689 80829 169009 80861
rect 168689 80593 168731 80829
rect 168967 80593 169009 80829
rect 168689 80509 169009 80593
rect 168689 80273 168731 80509
rect 168967 80273 169009 80509
rect 168689 80241 169009 80273
rect 173387 80829 173707 80861
rect 173387 80593 173429 80829
rect 173665 80593 173707 80829
rect 176331 80820 176332 80884
rect 176396 80820 176397 80884
rect 288387 80884 288453 80885
rect 176331 80819 176397 80820
rect 188076 80829 188396 80861
rect 173387 80509 173707 80593
rect 173387 80273 173429 80509
rect 173665 80273 173707 80509
rect 173387 80241 173707 80273
rect 188076 80593 188118 80829
rect 188354 80593 188396 80829
rect 188076 80509 188396 80593
rect 188076 80273 188118 80509
rect 188354 80273 188396 80509
rect 188076 80241 188396 80273
rect 194340 80829 194660 80861
rect 194340 80593 194382 80829
rect 194618 80593 194660 80829
rect 194340 80509 194660 80593
rect 194340 80273 194382 80509
rect 194618 80273 194660 80509
rect 194340 80241 194660 80273
rect 200604 80829 200924 80861
rect 200604 80593 200646 80829
rect 200882 80593 200924 80829
rect 200604 80509 200924 80593
rect 200604 80273 200646 80509
rect 200882 80273 200924 80509
rect 200604 80241 200924 80273
rect 216076 80829 216396 80861
rect 216076 80593 216118 80829
rect 216354 80593 216396 80829
rect 216076 80509 216396 80593
rect 216076 80273 216118 80509
rect 216354 80273 216396 80509
rect 216076 80241 216396 80273
rect 222340 80829 222660 80861
rect 222340 80593 222382 80829
rect 222618 80593 222660 80829
rect 222340 80509 222660 80593
rect 222340 80273 222382 80509
rect 222618 80273 222660 80509
rect 222340 80241 222660 80273
rect 228604 80829 228924 80861
rect 228604 80593 228646 80829
rect 228882 80593 228924 80829
rect 228604 80509 228924 80593
rect 228604 80273 228646 80509
rect 228882 80273 228924 80509
rect 228604 80241 228924 80273
rect 244076 80829 244396 80861
rect 244076 80593 244118 80829
rect 244354 80593 244396 80829
rect 244076 80509 244396 80593
rect 244076 80273 244118 80509
rect 244354 80273 244396 80509
rect 244076 80241 244396 80273
rect 250340 80829 250660 80861
rect 250340 80593 250382 80829
rect 250618 80593 250660 80829
rect 250340 80509 250660 80593
rect 250340 80273 250382 80509
rect 250618 80273 250660 80509
rect 250340 80241 250660 80273
rect 256604 80829 256924 80861
rect 256604 80593 256646 80829
rect 256882 80593 256924 80829
rect 256604 80509 256924 80593
rect 256604 80273 256646 80509
rect 256882 80273 256924 80509
rect 256604 80241 256924 80273
rect 272076 80829 272396 80861
rect 272076 80593 272118 80829
rect 272354 80593 272396 80829
rect 272076 80509 272396 80593
rect 272076 80273 272118 80509
rect 272354 80273 272396 80509
rect 272076 80241 272396 80273
rect 278340 80829 278660 80861
rect 278340 80593 278382 80829
rect 278618 80593 278660 80829
rect 278340 80509 278660 80593
rect 278340 80273 278382 80509
rect 278618 80273 278660 80509
rect 278340 80241 278660 80273
rect 284604 80829 284924 80861
rect 284604 80593 284646 80829
rect 284882 80593 284924 80829
rect 288387 80820 288388 80884
rect 288452 80820 288453 80884
rect 288387 80819 288453 80820
rect 296483 80884 296549 80885
rect 296483 80820 296484 80884
rect 296548 80820 296549 80884
rect 372291 80884 372357 80885
rect 296483 80819 296549 80820
rect 300076 80829 300396 80861
rect 284604 80509 284924 80593
rect 284604 80273 284646 80509
rect 284882 80273 284924 80509
rect 284604 80241 284924 80273
rect 300076 80593 300118 80829
rect 300354 80593 300396 80829
rect 300076 80509 300396 80593
rect 300076 80273 300118 80509
rect 300354 80273 300396 80509
rect 300076 80241 300396 80273
rect 306340 80829 306660 80861
rect 306340 80593 306382 80829
rect 306618 80593 306660 80829
rect 306340 80509 306660 80593
rect 306340 80273 306382 80509
rect 306618 80273 306660 80509
rect 306340 80241 306660 80273
rect 312604 80829 312924 80861
rect 312604 80593 312646 80829
rect 312882 80593 312924 80829
rect 312604 80509 312924 80593
rect 312604 80273 312646 80509
rect 312882 80273 312924 80509
rect 312604 80241 312924 80273
rect 328076 80829 328396 80861
rect 328076 80593 328118 80829
rect 328354 80593 328396 80829
rect 328076 80509 328396 80593
rect 328076 80273 328118 80509
rect 328354 80273 328396 80509
rect 328076 80241 328396 80273
rect 334340 80829 334660 80861
rect 334340 80593 334382 80829
rect 334618 80593 334660 80829
rect 334340 80509 334660 80593
rect 334340 80273 334382 80509
rect 334618 80273 334660 80509
rect 334340 80241 334660 80273
rect 340604 80829 340924 80861
rect 340604 80593 340646 80829
rect 340882 80593 340924 80829
rect 340604 80509 340924 80593
rect 340604 80273 340646 80509
rect 340882 80273 340924 80509
rect 340604 80241 340924 80273
rect 355293 80829 355613 80861
rect 355293 80593 355335 80829
rect 355571 80593 355613 80829
rect 355293 80509 355613 80593
rect 355293 80273 355335 80509
rect 355571 80273 355613 80509
rect 355293 80241 355613 80273
rect 359991 80829 360311 80861
rect 359991 80593 360033 80829
rect 360269 80593 360311 80829
rect 359991 80509 360311 80593
rect 359991 80273 360033 80509
rect 360269 80273 360311 80509
rect 359991 80241 360311 80273
rect 364689 80829 365009 80861
rect 364689 80593 364731 80829
rect 364967 80593 365009 80829
rect 364689 80509 365009 80593
rect 364689 80273 364731 80509
rect 364967 80273 365009 80509
rect 364689 80241 365009 80273
rect 369387 80829 369707 80861
rect 369387 80593 369429 80829
rect 369665 80593 369707 80829
rect 372291 80820 372292 80884
rect 372356 80820 372357 80884
rect 484347 80884 484413 80885
rect 372291 80819 372357 80820
rect 383293 80829 383613 80861
rect 369387 80509 369707 80593
rect 369387 80273 369429 80509
rect 369665 80273 369707 80509
rect 369387 80241 369707 80273
rect 383293 80593 383335 80829
rect 383571 80593 383613 80829
rect 383293 80509 383613 80593
rect 383293 80273 383335 80509
rect 383571 80273 383613 80509
rect 383293 80241 383613 80273
rect 387991 80829 388311 80861
rect 387991 80593 388033 80829
rect 388269 80593 388311 80829
rect 387991 80509 388311 80593
rect 387991 80273 388033 80509
rect 388269 80273 388311 80509
rect 387991 80241 388311 80273
rect 392689 80829 393009 80861
rect 392689 80593 392731 80829
rect 392967 80593 393009 80829
rect 392689 80509 393009 80593
rect 392689 80273 392731 80509
rect 392967 80273 393009 80509
rect 392689 80241 393009 80273
rect 397387 80829 397707 80861
rect 397387 80593 397429 80829
rect 397665 80593 397707 80829
rect 397387 80509 397707 80593
rect 397387 80273 397429 80509
rect 397665 80273 397707 80509
rect 397387 80241 397707 80273
rect 411293 80829 411613 80861
rect 411293 80593 411335 80829
rect 411571 80593 411613 80829
rect 411293 80509 411613 80593
rect 411293 80273 411335 80509
rect 411571 80273 411613 80509
rect 411293 80241 411613 80273
rect 415991 80829 416311 80861
rect 415991 80593 416033 80829
rect 416269 80593 416311 80829
rect 415991 80509 416311 80593
rect 415991 80273 416033 80509
rect 416269 80273 416311 80509
rect 415991 80241 416311 80273
rect 420689 80829 421009 80861
rect 420689 80593 420731 80829
rect 420967 80593 421009 80829
rect 420689 80509 421009 80593
rect 420689 80273 420731 80509
rect 420967 80273 421009 80509
rect 420689 80241 421009 80273
rect 425387 80829 425707 80861
rect 425387 80593 425429 80829
rect 425665 80593 425707 80829
rect 425387 80509 425707 80593
rect 425387 80273 425429 80509
rect 425665 80273 425707 80509
rect 425387 80241 425707 80273
rect 439293 80829 439613 80861
rect 439293 80593 439335 80829
rect 439571 80593 439613 80829
rect 439293 80509 439613 80593
rect 439293 80273 439335 80509
rect 439571 80273 439613 80509
rect 439293 80241 439613 80273
rect 443991 80829 444311 80861
rect 443991 80593 444033 80829
rect 444269 80593 444311 80829
rect 443991 80509 444311 80593
rect 443991 80273 444033 80509
rect 444269 80273 444311 80509
rect 443991 80241 444311 80273
rect 448689 80829 449009 80861
rect 448689 80593 448731 80829
rect 448967 80593 449009 80829
rect 448689 80509 449009 80593
rect 448689 80273 448731 80509
rect 448967 80273 449009 80509
rect 448689 80241 449009 80273
rect 453387 80829 453707 80861
rect 453387 80593 453429 80829
rect 453665 80593 453707 80829
rect 453387 80509 453707 80593
rect 453387 80273 453429 80509
rect 453665 80273 453707 80509
rect 453387 80241 453707 80273
rect 467293 80829 467613 80861
rect 467293 80593 467335 80829
rect 467571 80593 467613 80829
rect 467293 80509 467613 80593
rect 467293 80273 467335 80509
rect 467571 80273 467613 80509
rect 467293 80241 467613 80273
rect 471991 80829 472311 80861
rect 471991 80593 472033 80829
rect 472269 80593 472311 80829
rect 471991 80509 472311 80593
rect 471991 80273 472033 80509
rect 472269 80273 472311 80509
rect 471991 80241 472311 80273
rect 476689 80829 477009 80861
rect 476689 80593 476731 80829
rect 476967 80593 477009 80829
rect 476689 80509 477009 80593
rect 476689 80273 476731 80509
rect 476967 80273 477009 80509
rect 476689 80241 477009 80273
rect 481387 80829 481707 80861
rect 481387 80593 481429 80829
rect 481665 80593 481707 80829
rect 484347 80820 484348 80884
rect 484412 80820 484413 80884
rect 520595 80884 520661 80885
rect 484347 80819 484413 80820
rect 495293 80829 495613 80861
rect 481387 80509 481707 80593
rect 481387 80273 481429 80509
rect 481665 80273 481707 80509
rect 481387 80241 481707 80273
rect 495293 80593 495335 80829
rect 495571 80593 495613 80829
rect 495293 80509 495613 80593
rect 495293 80273 495335 80509
rect 495571 80273 495613 80509
rect 495293 80241 495613 80273
rect 499991 80829 500311 80861
rect 499991 80593 500033 80829
rect 500269 80593 500311 80829
rect 499991 80509 500311 80593
rect 499991 80273 500033 80509
rect 500269 80273 500311 80509
rect 499991 80241 500311 80273
rect 504689 80829 505009 80861
rect 504689 80593 504731 80829
rect 504967 80593 505009 80829
rect 504689 80509 505009 80593
rect 504689 80273 504731 80509
rect 504967 80273 505009 80509
rect 504689 80241 505009 80273
rect 509387 80829 509707 80861
rect 509387 80593 509429 80829
rect 509665 80593 509707 80829
rect 520595 80820 520596 80884
rect 520660 80820 520661 80884
rect 520595 80819 520661 80820
rect 523293 80829 523613 80861
rect 509387 80509 509707 80593
rect 509387 80273 509429 80509
rect 509665 80273 509707 80509
rect 509387 80241 509707 80273
rect 523293 80593 523335 80829
rect 523571 80593 523613 80829
rect 523293 80509 523613 80593
rect 523293 80273 523335 80509
rect 523571 80273 523613 80509
rect 523293 80241 523613 80273
rect 527991 80829 528311 80861
rect 527991 80593 528033 80829
rect 528269 80593 528311 80829
rect 527991 80509 528311 80593
rect 527991 80273 528033 80509
rect 528269 80273 528311 80509
rect 527991 80241 528311 80273
rect 532689 80829 533009 80861
rect 532689 80593 532731 80829
rect 532967 80593 533009 80829
rect 532689 80509 533009 80593
rect 532689 80273 532731 80509
rect 532967 80273 533009 80509
rect 532689 80241 533009 80273
rect 537387 80829 537707 80861
rect 537387 80593 537429 80829
rect 537665 80593 537707 80829
rect 537387 80509 537707 80593
rect 537387 80273 537429 80509
rect 537665 80273 537707 80509
rect 537387 80241 537707 80273
rect 551293 80829 551613 80861
rect 551293 80593 551335 80829
rect 551571 80593 551613 80829
rect 551293 80509 551613 80593
rect 551293 80273 551335 80509
rect 551571 80273 551613 80509
rect 551293 80241 551613 80273
rect 555991 80829 556311 80861
rect 555991 80593 556033 80829
rect 556269 80593 556311 80829
rect 555991 80509 556311 80593
rect 555991 80273 556033 80509
rect 556269 80273 556311 80509
rect 555991 80241 556311 80273
rect 560689 80829 561009 80861
rect 560689 80593 560731 80829
rect 560967 80593 561009 80829
rect 560689 80509 561009 80593
rect 560689 80273 560731 80509
rect 560967 80273 561009 80509
rect 560689 80241 561009 80273
rect 565387 80829 565707 80861
rect 565387 80593 565429 80829
rect 565665 80593 565707 80829
rect 565387 80509 565707 80593
rect 565387 80273 565429 80509
rect 565665 80273 565707 80509
rect 565387 80241 565707 80273
rect 573494 80829 574114 107273
rect 573494 80593 573526 80829
rect 573762 80593 573846 80829
rect 574082 80593 574114 80829
rect 573494 80509 574114 80593
rect 573494 80273 573526 80509
rect 573762 80273 573846 80509
rect 574082 80273 574114 80509
rect 79208 77454 79528 77486
rect 79208 77218 79250 77454
rect 79486 77218 79528 77454
rect 79208 77134 79528 77218
rect 79208 76898 79250 77134
rect 79486 76898 79528 77134
rect 79208 76866 79528 76898
rect 85472 77454 85792 77486
rect 85472 77218 85514 77454
rect 85750 77218 85792 77454
rect 85472 77134 85792 77218
rect 85472 76898 85514 77134
rect 85750 76898 85792 77134
rect 85472 76866 85792 76898
rect 105642 77454 105962 77486
rect 105642 77218 105684 77454
rect 105920 77218 105962 77454
rect 105642 77134 105962 77218
rect 105642 76898 105684 77134
rect 105920 76898 105962 77134
rect 105642 76866 105962 76898
rect 110340 77454 110660 77486
rect 110340 77218 110382 77454
rect 110618 77218 110660 77454
rect 110340 77134 110660 77218
rect 110340 76898 110382 77134
rect 110618 76898 110660 77134
rect 110340 76866 110660 76898
rect 115038 77454 115358 77486
rect 115038 77218 115080 77454
rect 115316 77218 115358 77454
rect 115038 77134 115358 77218
rect 115038 76898 115080 77134
rect 115316 76898 115358 77134
rect 115038 76866 115358 76898
rect 133642 77454 133962 77486
rect 133642 77218 133684 77454
rect 133920 77218 133962 77454
rect 133642 77134 133962 77218
rect 133642 76898 133684 77134
rect 133920 76898 133962 77134
rect 133642 76866 133962 76898
rect 138340 77454 138660 77486
rect 138340 77218 138382 77454
rect 138618 77218 138660 77454
rect 138340 77134 138660 77218
rect 138340 76898 138382 77134
rect 138618 76898 138660 77134
rect 138340 76866 138660 76898
rect 143038 77454 143358 77486
rect 143038 77218 143080 77454
rect 143316 77218 143358 77454
rect 143038 77134 143358 77218
rect 143038 76898 143080 77134
rect 143316 76898 143358 77134
rect 143038 76866 143358 76898
rect 161642 77454 161962 77486
rect 161642 77218 161684 77454
rect 161920 77218 161962 77454
rect 161642 77134 161962 77218
rect 161642 76898 161684 77134
rect 161920 76898 161962 77134
rect 161642 76866 161962 76898
rect 166340 77454 166660 77486
rect 166340 77218 166382 77454
rect 166618 77218 166660 77454
rect 166340 77134 166660 77218
rect 166340 76898 166382 77134
rect 166618 76898 166660 77134
rect 166340 76866 166660 76898
rect 171038 77454 171358 77486
rect 171038 77218 171080 77454
rect 171316 77218 171358 77454
rect 171038 77134 171358 77218
rect 171038 76898 171080 77134
rect 171316 76898 171358 77134
rect 171038 76866 171358 76898
rect 191208 77454 191528 77486
rect 191208 77218 191250 77454
rect 191486 77218 191528 77454
rect 191208 77134 191528 77218
rect 191208 76898 191250 77134
rect 191486 76898 191528 77134
rect 191208 76866 191528 76898
rect 197472 77454 197792 77486
rect 197472 77218 197514 77454
rect 197750 77218 197792 77454
rect 197472 77134 197792 77218
rect 197472 76898 197514 77134
rect 197750 76898 197792 77134
rect 197472 76866 197792 76898
rect 219208 77454 219528 77486
rect 219208 77218 219250 77454
rect 219486 77218 219528 77454
rect 219208 77134 219528 77218
rect 219208 76898 219250 77134
rect 219486 76898 219528 77134
rect 219208 76866 219528 76898
rect 225472 77454 225792 77486
rect 225472 77218 225514 77454
rect 225750 77218 225792 77454
rect 225472 77134 225792 77218
rect 225472 76898 225514 77134
rect 225750 76898 225792 77134
rect 225472 76866 225792 76898
rect 247208 77454 247528 77486
rect 247208 77218 247250 77454
rect 247486 77218 247528 77454
rect 247208 77134 247528 77218
rect 247208 76898 247250 77134
rect 247486 76898 247528 77134
rect 247208 76866 247528 76898
rect 253472 77454 253792 77486
rect 253472 77218 253514 77454
rect 253750 77218 253792 77454
rect 253472 77134 253792 77218
rect 253472 76898 253514 77134
rect 253750 76898 253792 77134
rect 253472 76866 253792 76898
rect 275208 77454 275528 77486
rect 275208 77218 275250 77454
rect 275486 77218 275528 77454
rect 275208 77134 275528 77218
rect 275208 76898 275250 77134
rect 275486 76898 275528 77134
rect 275208 76866 275528 76898
rect 281472 77454 281792 77486
rect 281472 77218 281514 77454
rect 281750 77218 281792 77454
rect 281472 77134 281792 77218
rect 281472 76898 281514 77134
rect 281750 76898 281792 77134
rect 281472 76866 281792 76898
rect 303208 77454 303528 77486
rect 303208 77218 303250 77454
rect 303486 77218 303528 77454
rect 303208 77134 303528 77218
rect 303208 76898 303250 77134
rect 303486 76898 303528 77134
rect 303208 76866 303528 76898
rect 309472 77454 309792 77486
rect 309472 77218 309514 77454
rect 309750 77218 309792 77454
rect 309472 77134 309792 77218
rect 309472 76898 309514 77134
rect 309750 76898 309792 77134
rect 309472 76866 309792 76898
rect 331208 77454 331528 77486
rect 331208 77218 331250 77454
rect 331486 77218 331528 77454
rect 331208 77134 331528 77218
rect 331208 76898 331250 77134
rect 331486 76898 331528 77134
rect 331208 76866 331528 76898
rect 337472 77454 337792 77486
rect 337472 77218 337514 77454
rect 337750 77218 337792 77454
rect 337472 77134 337792 77218
rect 337472 76898 337514 77134
rect 337750 76898 337792 77134
rect 337472 76866 337792 76898
rect 357642 77454 357962 77486
rect 357642 77218 357684 77454
rect 357920 77218 357962 77454
rect 357642 77134 357962 77218
rect 357642 76898 357684 77134
rect 357920 76898 357962 77134
rect 357642 76866 357962 76898
rect 362340 77454 362660 77486
rect 362340 77218 362382 77454
rect 362618 77218 362660 77454
rect 362340 77134 362660 77218
rect 362340 76898 362382 77134
rect 362618 76898 362660 77134
rect 362340 76866 362660 76898
rect 367038 77454 367358 77486
rect 367038 77218 367080 77454
rect 367316 77218 367358 77454
rect 367038 77134 367358 77218
rect 367038 76898 367080 77134
rect 367316 76898 367358 77134
rect 367038 76866 367358 76898
rect 385642 77454 385962 77486
rect 385642 77218 385684 77454
rect 385920 77218 385962 77454
rect 385642 77134 385962 77218
rect 385642 76898 385684 77134
rect 385920 76898 385962 77134
rect 385642 76866 385962 76898
rect 390340 77454 390660 77486
rect 390340 77218 390382 77454
rect 390618 77218 390660 77454
rect 390340 77134 390660 77218
rect 390340 76898 390382 77134
rect 390618 76898 390660 77134
rect 390340 76866 390660 76898
rect 395038 77454 395358 77486
rect 395038 77218 395080 77454
rect 395316 77218 395358 77454
rect 395038 77134 395358 77218
rect 395038 76898 395080 77134
rect 395316 76898 395358 77134
rect 395038 76866 395358 76898
rect 413642 77454 413962 77486
rect 413642 77218 413684 77454
rect 413920 77218 413962 77454
rect 413642 77134 413962 77218
rect 413642 76898 413684 77134
rect 413920 76898 413962 77134
rect 413642 76866 413962 76898
rect 418340 77454 418660 77486
rect 418340 77218 418382 77454
rect 418618 77218 418660 77454
rect 418340 77134 418660 77218
rect 418340 76898 418382 77134
rect 418618 76898 418660 77134
rect 418340 76866 418660 76898
rect 423038 77454 423358 77486
rect 423038 77218 423080 77454
rect 423316 77218 423358 77454
rect 423038 77134 423358 77218
rect 423038 76898 423080 77134
rect 423316 76898 423358 77134
rect 423038 76866 423358 76898
rect 441642 77454 441962 77486
rect 441642 77218 441684 77454
rect 441920 77218 441962 77454
rect 441642 77134 441962 77218
rect 441642 76898 441684 77134
rect 441920 76898 441962 77134
rect 441642 76866 441962 76898
rect 446340 77454 446660 77486
rect 446340 77218 446382 77454
rect 446618 77218 446660 77454
rect 446340 77134 446660 77218
rect 446340 76898 446382 77134
rect 446618 76898 446660 77134
rect 446340 76866 446660 76898
rect 451038 77454 451358 77486
rect 451038 77218 451080 77454
rect 451316 77218 451358 77454
rect 451038 77134 451358 77218
rect 451038 76898 451080 77134
rect 451316 76898 451358 77134
rect 451038 76866 451358 76898
rect 469642 77454 469962 77486
rect 469642 77218 469684 77454
rect 469920 77218 469962 77454
rect 469642 77134 469962 77218
rect 469642 76898 469684 77134
rect 469920 76898 469962 77134
rect 469642 76866 469962 76898
rect 474340 77454 474660 77486
rect 474340 77218 474382 77454
rect 474618 77218 474660 77454
rect 474340 77134 474660 77218
rect 474340 76898 474382 77134
rect 474618 76898 474660 77134
rect 474340 76866 474660 76898
rect 479038 77454 479358 77486
rect 479038 77218 479080 77454
rect 479316 77218 479358 77454
rect 479038 77134 479358 77218
rect 479038 76898 479080 77134
rect 479316 76898 479358 77134
rect 479038 76866 479358 76898
rect 497642 77454 497962 77486
rect 497642 77218 497684 77454
rect 497920 77218 497962 77454
rect 497642 77134 497962 77218
rect 497642 76898 497684 77134
rect 497920 76898 497962 77134
rect 497642 76866 497962 76898
rect 502340 77454 502660 77486
rect 502340 77218 502382 77454
rect 502618 77218 502660 77454
rect 502340 77134 502660 77218
rect 502340 76898 502382 77134
rect 502618 76898 502660 77134
rect 502340 76866 502660 76898
rect 507038 77454 507358 77486
rect 507038 77218 507080 77454
rect 507316 77218 507358 77454
rect 507038 77134 507358 77218
rect 507038 76898 507080 77134
rect 507316 76898 507358 77134
rect 507038 76866 507358 76898
rect 525642 77454 525962 77486
rect 525642 77218 525684 77454
rect 525920 77218 525962 77454
rect 525642 77134 525962 77218
rect 525642 76898 525684 77134
rect 525920 76898 525962 77134
rect 525642 76866 525962 76898
rect 530340 77454 530660 77486
rect 530340 77218 530382 77454
rect 530618 77218 530660 77454
rect 530340 77134 530660 77218
rect 530340 76898 530382 77134
rect 530618 76898 530660 77134
rect 530340 76866 530660 76898
rect 535038 77454 535358 77486
rect 535038 77218 535080 77454
rect 535316 77218 535358 77454
rect 535038 77134 535358 77218
rect 535038 76898 535080 77134
rect 535316 76898 535358 77134
rect 535038 76866 535358 76898
rect 553642 77454 553962 77486
rect 553642 77218 553684 77454
rect 553920 77218 553962 77454
rect 553642 77134 553962 77218
rect 553642 76898 553684 77134
rect 553920 76898 553962 77134
rect 553642 76866 553962 76898
rect 558340 77454 558660 77486
rect 558340 77218 558382 77454
rect 558618 77218 558660 77454
rect 558340 77134 558660 77218
rect 558340 76898 558382 77134
rect 558618 76898 558660 77134
rect 558340 76866 558660 76898
rect 563038 77454 563358 77486
rect 563038 77218 563080 77454
rect 563316 77218 563358 77454
rect 563038 77134 563358 77218
rect 563038 76898 563080 77134
rect 563316 76898 563358 77134
rect 563038 76866 563358 76898
rect 76076 53829 76396 53861
rect 76076 53593 76118 53829
rect 76354 53593 76396 53829
rect 76076 53509 76396 53593
rect 64459 53412 64525 53413
rect 64459 53410 64460 53412
rect 63910 53350 64460 53410
rect 63910 45389 63970 53350
rect 64459 53348 64460 53350
rect 64524 53348 64525 53412
rect 64459 53347 64525 53348
rect 76076 53273 76118 53509
rect 76354 53273 76396 53509
rect 76076 53241 76396 53273
rect 82340 53829 82660 53861
rect 82340 53593 82382 53829
rect 82618 53593 82660 53829
rect 82340 53509 82660 53593
rect 82340 53273 82382 53509
rect 82618 53273 82660 53509
rect 82340 53241 82660 53273
rect 88604 53829 88924 53861
rect 88604 53593 88646 53829
rect 88882 53593 88924 53829
rect 88604 53509 88924 53593
rect 88604 53273 88646 53509
rect 88882 53273 88924 53509
rect 104076 53829 104396 53861
rect 104076 53593 104118 53829
rect 104354 53593 104396 53829
rect 104076 53509 104396 53593
rect 88604 53241 88924 53273
rect 92427 53276 92493 53277
rect 92427 53212 92428 53276
rect 92492 53212 92493 53276
rect 104076 53273 104118 53509
rect 104354 53273 104396 53509
rect 104076 53241 104396 53273
rect 110340 53829 110660 53861
rect 110340 53593 110382 53829
rect 110618 53593 110660 53829
rect 110340 53509 110660 53593
rect 110340 53273 110382 53509
rect 110618 53273 110660 53509
rect 110340 53241 110660 53273
rect 116604 53829 116924 53861
rect 116604 53593 116646 53829
rect 116882 53593 116924 53829
rect 116604 53509 116924 53593
rect 116604 53273 116646 53509
rect 116882 53273 116924 53509
rect 116604 53241 116924 53273
rect 132076 53829 132396 53861
rect 132076 53593 132118 53829
rect 132354 53593 132396 53829
rect 132076 53509 132396 53593
rect 132076 53273 132118 53509
rect 132354 53273 132396 53509
rect 132076 53241 132396 53273
rect 138340 53829 138660 53861
rect 138340 53593 138382 53829
rect 138618 53593 138660 53829
rect 138340 53509 138660 53593
rect 138340 53273 138382 53509
rect 138618 53273 138660 53509
rect 138340 53241 138660 53273
rect 144604 53829 144924 53861
rect 144604 53593 144646 53829
rect 144882 53593 144924 53829
rect 144604 53509 144924 53593
rect 144604 53273 144646 53509
rect 144882 53273 144924 53509
rect 160076 53829 160396 53861
rect 160076 53593 160118 53829
rect 160354 53593 160396 53829
rect 160076 53509 160396 53593
rect 144604 53241 144924 53273
rect 148363 53276 148429 53277
rect 92427 53211 92493 53212
rect 148363 53212 148364 53276
rect 148428 53212 148429 53276
rect 160076 53273 160118 53509
rect 160354 53273 160396 53509
rect 160076 53241 160396 53273
rect 166340 53829 166660 53861
rect 166340 53593 166382 53829
rect 166618 53593 166660 53829
rect 166340 53509 166660 53593
rect 166340 53273 166382 53509
rect 166618 53273 166660 53509
rect 166340 53241 166660 53273
rect 172604 53829 172924 53861
rect 172604 53593 172646 53829
rect 172882 53593 172924 53829
rect 172604 53509 172924 53593
rect 172604 53273 172646 53509
rect 172882 53273 172924 53509
rect 188076 53829 188396 53861
rect 188076 53593 188118 53829
rect 188354 53593 188396 53829
rect 188076 53509 188396 53593
rect 172604 53241 172924 53273
rect 176331 53276 176397 53277
rect 148363 53211 148429 53212
rect 176331 53212 176332 53276
rect 176396 53212 176397 53276
rect 188076 53273 188118 53509
rect 188354 53273 188396 53509
rect 188076 53241 188396 53273
rect 194340 53829 194660 53861
rect 194340 53593 194382 53829
rect 194618 53593 194660 53829
rect 194340 53509 194660 53593
rect 194340 53273 194382 53509
rect 194618 53273 194660 53509
rect 194340 53241 194660 53273
rect 200604 53829 200924 53861
rect 200604 53593 200646 53829
rect 200882 53593 200924 53829
rect 200604 53509 200924 53593
rect 200604 53273 200646 53509
rect 200882 53273 200924 53509
rect 200604 53241 200924 53273
rect 215293 53829 215613 53861
rect 215293 53593 215335 53829
rect 215571 53593 215613 53829
rect 215293 53509 215613 53593
rect 215293 53273 215335 53509
rect 215571 53273 215613 53509
rect 215293 53241 215613 53273
rect 219991 53829 220311 53861
rect 219991 53593 220033 53829
rect 220269 53593 220311 53829
rect 219991 53509 220311 53593
rect 219991 53273 220033 53509
rect 220269 53273 220311 53509
rect 219991 53241 220311 53273
rect 224689 53829 225009 53861
rect 224689 53593 224731 53829
rect 224967 53593 225009 53829
rect 224689 53509 225009 53593
rect 224689 53273 224731 53509
rect 224967 53273 225009 53509
rect 224689 53241 225009 53273
rect 229387 53829 229707 53861
rect 229387 53593 229429 53829
rect 229665 53593 229707 53829
rect 229387 53509 229707 53593
rect 229387 53273 229429 53509
rect 229665 53273 229707 53509
rect 229387 53241 229707 53273
rect 244076 53829 244396 53861
rect 244076 53593 244118 53829
rect 244354 53593 244396 53829
rect 244076 53509 244396 53593
rect 244076 53273 244118 53509
rect 244354 53273 244396 53509
rect 244076 53241 244396 53273
rect 250340 53829 250660 53861
rect 250340 53593 250382 53829
rect 250618 53593 250660 53829
rect 250340 53509 250660 53593
rect 250340 53273 250382 53509
rect 250618 53273 250660 53509
rect 250340 53241 250660 53273
rect 256604 53829 256924 53861
rect 256604 53593 256646 53829
rect 256882 53593 256924 53829
rect 256604 53509 256924 53593
rect 256604 53273 256646 53509
rect 256882 53273 256924 53509
rect 272076 53829 272396 53861
rect 272076 53593 272118 53829
rect 272354 53593 272396 53829
rect 272076 53509 272396 53593
rect 256604 53241 256924 53273
rect 260419 53276 260485 53277
rect 176331 53211 176397 53212
rect 260419 53212 260420 53276
rect 260484 53212 260485 53276
rect 272076 53273 272118 53509
rect 272354 53273 272396 53509
rect 272076 53241 272396 53273
rect 278340 53829 278660 53861
rect 278340 53593 278382 53829
rect 278618 53593 278660 53829
rect 278340 53509 278660 53593
rect 278340 53273 278382 53509
rect 278618 53273 278660 53509
rect 278340 53241 278660 53273
rect 284604 53829 284924 53861
rect 284604 53593 284646 53829
rect 284882 53593 284924 53829
rect 284604 53509 284924 53593
rect 284604 53273 284646 53509
rect 284882 53273 284924 53509
rect 300076 53829 300396 53861
rect 300076 53593 300118 53829
rect 300354 53593 300396 53829
rect 300076 53509 300396 53593
rect 284604 53241 284924 53273
rect 288387 53276 288453 53277
rect 260419 53211 260485 53212
rect 288387 53212 288388 53276
rect 288452 53212 288453 53276
rect 300076 53273 300118 53509
rect 300354 53273 300396 53509
rect 300076 53241 300396 53273
rect 306340 53829 306660 53861
rect 306340 53593 306382 53829
rect 306618 53593 306660 53829
rect 306340 53509 306660 53593
rect 306340 53273 306382 53509
rect 306618 53273 306660 53509
rect 306340 53241 306660 53273
rect 312604 53829 312924 53861
rect 312604 53593 312646 53829
rect 312882 53593 312924 53829
rect 312604 53509 312924 53593
rect 312604 53273 312646 53509
rect 312882 53273 312924 53509
rect 312604 53241 312924 53273
rect 327293 53829 327613 53861
rect 327293 53593 327335 53829
rect 327571 53593 327613 53829
rect 327293 53509 327613 53593
rect 327293 53273 327335 53509
rect 327571 53273 327613 53509
rect 327293 53241 327613 53273
rect 331991 53829 332311 53861
rect 331991 53593 332033 53829
rect 332269 53593 332311 53829
rect 331991 53509 332311 53593
rect 331991 53273 332033 53509
rect 332269 53273 332311 53509
rect 331991 53241 332311 53273
rect 336689 53829 337009 53861
rect 336689 53593 336731 53829
rect 336967 53593 337009 53829
rect 336689 53509 337009 53593
rect 336689 53273 336731 53509
rect 336967 53273 337009 53509
rect 336689 53241 337009 53273
rect 341387 53829 341707 53861
rect 341387 53593 341429 53829
rect 341665 53593 341707 53829
rect 341387 53509 341707 53593
rect 341387 53273 341429 53509
rect 341665 53273 341707 53509
rect 356076 53829 356396 53861
rect 356076 53593 356118 53829
rect 356354 53593 356396 53829
rect 356076 53509 356396 53593
rect 341387 53241 341707 53273
rect 344323 53276 344389 53277
rect 288387 53211 288453 53212
rect 344323 53212 344324 53276
rect 344388 53212 344389 53276
rect 356076 53273 356118 53509
rect 356354 53273 356396 53509
rect 356076 53241 356396 53273
rect 362340 53829 362660 53861
rect 362340 53593 362382 53829
rect 362618 53593 362660 53829
rect 362340 53509 362660 53593
rect 362340 53273 362382 53509
rect 362618 53273 362660 53509
rect 362340 53241 362660 53273
rect 368604 53829 368924 53861
rect 368604 53593 368646 53829
rect 368882 53593 368924 53829
rect 368604 53509 368924 53593
rect 368604 53273 368646 53509
rect 368882 53273 368924 53509
rect 384076 53829 384396 53861
rect 384076 53593 384118 53829
rect 384354 53593 384396 53829
rect 384076 53509 384396 53593
rect 368604 53241 368924 53273
rect 372291 53276 372357 53277
rect 344323 53211 344389 53212
rect 372291 53212 372292 53276
rect 372356 53212 372357 53276
rect 384076 53273 384118 53509
rect 384354 53273 384396 53509
rect 384076 53241 384396 53273
rect 390340 53829 390660 53861
rect 390340 53593 390382 53829
rect 390618 53593 390660 53829
rect 390340 53509 390660 53593
rect 390340 53273 390382 53509
rect 390618 53273 390660 53509
rect 390340 53241 390660 53273
rect 396604 53829 396924 53861
rect 396604 53593 396646 53829
rect 396882 53593 396924 53829
rect 396604 53509 396924 53593
rect 396604 53273 396646 53509
rect 396882 53273 396924 53509
rect 396604 53241 396924 53273
rect 412076 53829 412396 53861
rect 412076 53593 412118 53829
rect 412354 53593 412396 53829
rect 412076 53509 412396 53593
rect 412076 53273 412118 53509
rect 412354 53273 412396 53509
rect 412076 53241 412396 53273
rect 418340 53829 418660 53861
rect 418340 53593 418382 53829
rect 418618 53593 418660 53829
rect 418340 53509 418660 53593
rect 418340 53273 418382 53509
rect 418618 53273 418660 53509
rect 418340 53241 418660 53273
rect 424604 53829 424924 53861
rect 424604 53593 424646 53829
rect 424882 53593 424924 53829
rect 424604 53509 424924 53593
rect 424604 53273 424646 53509
rect 424882 53273 424924 53509
rect 424604 53241 424924 53273
rect 440076 53829 440396 53861
rect 440076 53593 440118 53829
rect 440354 53593 440396 53829
rect 440076 53509 440396 53593
rect 440076 53273 440118 53509
rect 440354 53273 440396 53509
rect 440076 53241 440396 53273
rect 446340 53829 446660 53861
rect 446340 53593 446382 53829
rect 446618 53593 446660 53829
rect 446340 53509 446660 53593
rect 446340 53273 446382 53509
rect 446618 53273 446660 53509
rect 446340 53241 446660 53273
rect 452604 53829 452924 53861
rect 452604 53593 452646 53829
rect 452882 53593 452924 53829
rect 452604 53509 452924 53593
rect 452604 53273 452646 53509
rect 452882 53273 452924 53509
rect 468076 53829 468396 53861
rect 468076 53593 468118 53829
rect 468354 53593 468396 53829
rect 468076 53509 468396 53593
rect 452604 53241 452924 53273
rect 456379 53276 456445 53277
rect 372291 53211 372357 53212
rect 456379 53212 456380 53276
rect 456444 53212 456445 53276
rect 468076 53273 468118 53509
rect 468354 53273 468396 53509
rect 468076 53241 468396 53273
rect 474340 53829 474660 53861
rect 474340 53593 474382 53829
rect 474618 53593 474660 53829
rect 474340 53509 474660 53593
rect 474340 53273 474382 53509
rect 474618 53273 474660 53509
rect 474340 53241 474660 53273
rect 480604 53829 480924 53861
rect 480604 53593 480646 53829
rect 480882 53593 480924 53829
rect 480604 53509 480924 53593
rect 480604 53273 480646 53509
rect 480882 53273 480924 53509
rect 495293 53829 495613 53861
rect 495293 53593 495335 53829
rect 495571 53593 495613 53829
rect 495293 53509 495613 53593
rect 480604 53241 480924 53273
rect 484347 53276 484413 53277
rect 456379 53211 456445 53212
rect 484347 53212 484348 53276
rect 484412 53212 484413 53276
rect 495293 53273 495335 53509
rect 495571 53273 495613 53509
rect 495293 53241 495613 53273
rect 499991 53829 500311 53861
rect 499991 53593 500033 53829
rect 500269 53593 500311 53829
rect 499991 53509 500311 53593
rect 499991 53273 500033 53509
rect 500269 53273 500311 53509
rect 499991 53241 500311 53273
rect 504689 53829 505009 53861
rect 504689 53593 504731 53829
rect 504967 53593 505009 53829
rect 504689 53509 505009 53593
rect 504689 53273 504731 53509
rect 504967 53273 505009 53509
rect 504689 53241 505009 53273
rect 509387 53829 509707 53861
rect 509387 53593 509429 53829
rect 509665 53593 509707 53829
rect 509387 53509 509707 53593
rect 509387 53273 509429 53509
rect 509665 53273 509707 53509
rect 524076 53829 524396 53861
rect 524076 53593 524118 53829
rect 524354 53593 524396 53829
rect 524076 53509 524396 53593
rect 509387 53241 509707 53273
rect 520595 53276 520661 53277
rect 484347 53211 484413 53212
rect 520595 53212 520596 53276
rect 520660 53212 520661 53276
rect 524076 53273 524118 53509
rect 524354 53273 524396 53509
rect 524076 53241 524396 53273
rect 530340 53829 530660 53861
rect 530340 53593 530382 53829
rect 530618 53593 530660 53829
rect 530340 53509 530660 53593
rect 530340 53273 530382 53509
rect 530618 53273 530660 53509
rect 530340 53241 530660 53273
rect 536604 53829 536924 53861
rect 536604 53593 536646 53829
rect 536882 53593 536924 53829
rect 536604 53509 536924 53593
rect 536604 53273 536646 53509
rect 536882 53273 536924 53509
rect 536604 53241 536924 53273
rect 552076 53829 552396 53861
rect 552076 53593 552118 53829
rect 552354 53593 552396 53829
rect 552076 53509 552396 53593
rect 552076 53273 552118 53509
rect 552354 53273 552396 53509
rect 552076 53241 552396 53273
rect 558340 53829 558660 53861
rect 558340 53593 558382 53829
rect 558618 53593 558660 53829
rect 558340 53509 558660 53593
rect 558340 53273 558382 53509
rect 558618 53273 558660 53509
rect 558340 53241 558660 53273
rect 564604 53829 564924 53861
rect 564604 53593 564646 53829
rect 564882 53593 564924 53829
rect 564604 53509 564924 53593
rect 564604 53273 564646 53509
rect 564882 53273 564924 53509
rect 564604 53241 564924 53273
rect 573494 53829 574114 80273
rect 573494 53593 573526 53829
rect 573762 53593 573846 53829
rect 574082 53593 574114 53829
rect 573494 53509 574114 53593
rect 573494 53273 573526 53509
rect 573762 53273 573846 53509
rect 574082 53273 574114 53509
rect 520595 53211 520661 53212
rect 79208 50454 79528 50486
rect 79208 50218 79250 50454
rect 79486 50218 79528 50454
rect 79208 50134 79528 50218
rect 79208 49898 79250 50134
rect 79486 49898 79528 50134
rect 79208 49866 79528 49898
rect 85472 50454 85792 50486
rect 85472 50218 85514 50454
rect 85750 50218 85792 50454
rect 85472 50134 85792 50218
rect 85472 49898 85514 50134
rect 85750 49898 85792 50134
rect 85472 49866 85792 49898
rect 92430 45570 92490 53211
rect 107208 50454 107528 50486
rect 107208 50218 107250 50454
rect 107486 50218 107528 50454
rect 107208 50134 107528 50218
rect 107208 49898 107250 50134
rect 107486 49898 107528 50134
rect 107208 49866 107528 49898
rect 113472 50454 113792 50486
rect 113472 50218 113514 50454
rect 113750 50218 113792 50454
rect 113472 50134 113792 50218
rect 113472 49898 113514 50134
rect 113750 49898 113792 50134
rect 113472 49866 113792 49898
rect 135208 50454 135528 50486
rect 135208 50218 135250 50454
rect 135486 50218 135528 50454
rect 135208 50134 135528 50218
rect 135208 49898 135250 50134
rect 135486 49898 135528 50134
rect 135208 49866 135528 49898
rect 141472 50454 141792 50486
rect 141472 50218 141514 50454
rect 141750 50218 141792 50454
rect 141472 50134 141792 50218
rect 141472 49898 141514 50134
rect 141750 49898 141792 50134
rect 141472 49866 141792 49898
rect 148366 45570 148426 53211
rect 163208 50454 163528 50486
rect 163208 50218 163250 50454
rect 163486 50218 163528 50454
rect 163208 50134 163528 50218
rect 163208 49898 163250 50134
rect 163486 49898 163528 50134
rect 163208 49866 163528 49898
rect 169472 50454 169792 50486
rect 169472 50218 169514 50454
rect 169750 50218 169792 50454
rect 169472 50134 169792 50218
rect 169472 49898 169514 50134
rect 169750 49898 169792 50134
rect 169472 49866 169792 49898
rect 176334 45570 176394 53211
rect 191208 50454 191528 50486
rect 191208 50218 191250 50454
rect 191486 50218 191528 50454
rect 191208 50134 191528 50218
rect 191208 49898 191250 50134
rect 191486 49898 191528 50134
rect 191208 49866 191528 49898
rect 197472 50454 197792 50486
rect 197472 50218 197514 50454
rect 197750 50218 197792 50454
rect 197472 50134 197792 50218
rect 197472 49898 197514 50134
rect 197750 49898 197792 50134
rect 197472 49866 197792 49898
rect 217642 50454 217962 50486
rect 217642 50218 217684 50454
rect 217920 50218 217962 50454
rect 217642 50134 217962 50218
rect 217642 49898 217684 50134
rect 217920 49898 217962 50134
rect 217642 49866 217962 49898
rect 222340 50454 222660 50486
rect 222340 50218 222382 50454
rect 222618 50218 222660 50454
rect 222340 50134 222660 50218
rect 222340 49898 222382 50134
rect 222618 49898 222660 50134
rect 222340 49866 222660 49898
rect 227038 50454 227358 50486
rect 227038 50218 227080 50454
rect 227316 50218 227358 50454
rect 227038 50134 227358 50218
rect 227038 49898 227080 50134
rect 227316 49898 227358 50134
rect 227038 49866 227358 49898
rect 247208 50454 247528 50486
rect 247208 50218 247250 50454
rect 247486 50218 247528 50454
rect 247208 50134 247528 50218
rect 247208 49898 247250 50134
rect 247486 49898 247528 50134
rect 247208 49866 247528 49898
rect 253472 50454 253792 50486
rect 253472 50218 253514 50454
rect 253750 50218 253792 50454
rect 253472 50134 253792 50218
rect 253472 49898 253514 50134
rect 253750 49898 253792 50134
rect 253472 49866 253792 49898
rect 260422 45570 260482 53211
rect 275208 50454 275528 50486
rect 275208 50218 275250 50454
rect 275486 50218 275528 50454
rect 275208 50134 275528 50218
rect 275208 49898 275250 50134
rect 275486 49898 275528 50134
rect 275208 49866 275528 49898
rect 281472 50454 281792 50486
rect 281472 50218 281514 50454
rect 281750 50218 281792 50454
rect 281472 50134 281792 50218
rect 281472 49898 281514 50134
rect 281750 49898 281792 50134
rect 281472 49866 281792 49898
rect 288390 45570 288450 53211
rect 303208 50454 303528 50486
rect 303208 50218 303250 50454
rect 303486 50218 303528 50454
rect 303208 50134 303528 50218
rect 303208 49898 303250 50134
rect 303486 49898 303528 50134
rect 303208 49866 303528 49898
rect 309472 50454 309792 50486
rect 309472 50218 309514 50454
rect 309750 50218 309792 50454
rect 309472 50134 309792 50218
rect 309472 49898 309514 50134
rect 309750 49898 309792 50134
rect 309472 49866 309792 49898
rect 329642 50454 329962 50486
rect 329642 50218 329684 50454
rect 329920 50218 329962 50454
rect 329642 50134 329962 50218
rect 329642 49898 329684 50134
rect 329920 49898 329962 50134
rect 329642 49866 329962 49898
rect 334340 50454 334660 50486
rect 334340 50218 334382 50454
rect 334618 50218 334660 50454
rect 334340 50134 334660 50218
rect 334340 49898 334382 50134
rect 334618 49898 334660 50134
rect 334340 49866 334660 49898
rect 339038 50454 339358 50486
rect 339038 50218 339080 50454
rect 339316 50218 339358 50454
rect 339038 50134 339358 50218
rect 339038 49898 339080 50134
rect 339316 49898 339358 50134
rect 339038 49866 339358 49898
rect 344326 45570 344386 53211
rect 359208 50454 359528 50486
rect 359208 50218 359250 50454
rect 359486 50218 359528 50454
rect 359208 50134 359528 50218
rect 359208 49898 359250 50134
rect 359486 49898 359528 50134
rect 359208 49866 359528 49898
rect 365472 50454 365792 50486
rect 365472 50218 365514 50454
rect 365750 50218 365792 50454
rect 365472 50134 365792 50218
rect 365472 49898 365514 50134
rect 365750 49898 365792 50134
rect 365472 49866 365792 49898
rect 372294 45570 372354 53211
rect 387208 50454 387528 50486
rect 387208 50218 387250 50454
rect 387486 50218 387528 50454
rect 387208 50134 387528 50218
rect 387208 49898 387250 50134
rect 387486 49898 387528 50134
rect 387208 49866 387528 49898
rect 393472 50454 393792 50486
rect 393472 50218 393514 50454
rect 393750 50218 393792 50454
rect 393472 50134 393792 50218
rect 393472 49898 393514 50134
rect 393750 49898 393792 50134
rect 393472 49866 393792 49898
rect 415208 50454 415528 50486
rect 415208 50218 415250 50454
rect 415486 50218 415528 50454
rect 415208 50134 415528 50218
rect 415208 49898 415250 50134
rect 415486 49898 415528 50134
rect 415208 49866 415528 49898
rect 421472 50454 421792 50486
rect 421472 50218 421514 50454
rect 421750 50218 421792 50454
rect 421472 50134 421792 50218
rect 421472 49898 421514 50134
rect 421750 49898 421792 50134
rect 421472 49866 421792 49898
rect 443208 50454 443528 50486
rect 443208 50218 443250 50454
rect 443486 50218 443528 50454
rect 443208 50134 443528 50218
rect 443208 49898 443250 50134
rect 443486 49898 443528 50134
rect 443208 49866 443528 49898
rect 449472 50454 449792 50486
rect 449472 50218 449514 50454
rect 449750 50218 449792 50454
rect 449472 50134 449792 50218
rect 449472 49898 449514 50134
rect 449750 49898 449792 50134
rect 449472 49866 449792 49898
rect 456382 45570 456442 53211
rect 471208 50454 471528 50486
rect 471208 50218 471250 50454
rect 471486 50218 471528 50454
rect 471208 50134 471528 50218
rect 471208 49898 471250 50134
rect 471486 49898 471528 50134
rect 471208 49866 471528 49898
rect 477472 50454 477792 50486
rect 477472 50218 477514 50454
rect 477750 50218 477792 50454
rect 477472 50134 477792 50218
rect 477472 49898 477514 50134
rect 477750 49898 477792 50134
rect 477472 49866 477792 49898
rect 484350 45570 484410 53211
rect 497642 50454 497962 50486
rect 497642 50218 497684 50454
rect 497920 50218 497962 50454
rect 497642 50134 497962 50218
rect 497642 49898 497684 50134
rect 497920 49898 497962 50134
rect 497642 49866 497962 49898
rect 502340 50454 502660 50486
rect 502340 50218 502382 50454
rect 502618 50218 502660 50454
rect 502340 50134 502660 50218
rect 502340 49898 502382 50134
rect 502618 49898 502660 50134
rect 502340 49866 502660 49898
rect 507038 50454 507358 50486
rect 507038 50218 507080 50454
rect 507316 50218 507358 50454
rect 507038 50134 507358 50218
rect 507038 49898 507080 50134
rect 507316 49898 507358 50134
rect 507038 49866 507358 49898
rect 91142 45510 92490 45570
rect 147630 45510 148426 45570
rect 175230 45510 176394 45570
rect 259502 45510 260482 45570
rect 287102 45510 288450 45570
rect 343590 45510 344386 45570
rect 371190 45510 372354 45570
rect 455462 45510 456442 45570
rect 483062 45510 484410 45570
rect 520598 45570 520658 53211
rect 527208 50454 527528 50486
rect 527208 50218 527250 50454
rect 527486 50218 527528 50454
rect 527208 50134 527528 50218
rect 527208 49898 527250 50134
rect 527486 49898 527528 50134
rect 527208 49866 527528 49898
rect 533472 50454 533792 50486
rect 533472 50218 533514 50454
rect 533750 50218 533792 50454
rect 533472 50134 533792 50218
rect 533472 49898 533514 50134
rect 533750 49898 533792 50134
rect 533472 49866 533792 49898
rect 555208 50454 555528 50486
rect 555208 50218 555250 50454
rect 555486 50218 555528 50454
rect 555208 50134 555528 50218
rect 555208 49898 555250 50134
rect 555486 49898 555528 50134
rect 555208 49866 555528 49898
rect 561472 50454 561792 50486
rect 561472 50218 561514 50454
rect 561750 50218 561792 50454
rect 561472 50134 561792 50218
rect 561472 49898 561514 50134
rect 561750 49898 561792 50134
rect 561472 49866 561792 49898
rect 520598 45510 520842 45570
rect 63907 45388 63973 45389
rect 63907 45324 63908 45388
rect 63972 45324 63973 45388
rect 63907 45323 63973 45324
rect 91142 45253 91202 45510
rect 147630 45253 147690 45510
rect 175230 45389 175290 45510
rect 175227 45388 175293 45389
rect 175227 45324 175228 45388
rect 175292 45324 175293 45388
rect 175227 45323 175293 45324
rect 259502 45253 259562 45510
rect 91139 45252 91205 45253
rect 91139 45188 91140 45252
rect 91204 45188 91205 45252
rect 91139 45187 91205 45188
rect 147627 45252 147693 45253
rect 147627 45188 147628 45252
rect 147692 45188 147693 45252
rect 147627 45187 147693 45188
rect 259499 45252 259565 45253
rect 259499 45188 259500 45252
rect 259564 45188 259565 45252
rect 259499 45187 259565 45188
rect 287102 45117 287162 45510
rect 343590 45253 343650 45510
rect 343587 45252 343653 45253
rect 343587 45188 343588 45252
rect 343652 45188 343653 45252
rect 343587 45187 343653 45188
rect 371190 45117 371250 45510
rect 455462 45389 455522 45510
rect 455459 45388 455525 45389
rect 455459 45324 455460 45388
rect 455524 45324 455525 45388
rect 455459 45323 455525 45324
rect 483062 45253 483122 45510
rect 520782 45389 520842 45510
rect 520779 45388 520845 45389
rect 520779 45324 520780 45388
rect 520844 45324 520845 45388
rect 520779 45323 520845 45324
rect 483059 45252 483125 45253
rect 483059 45188 483060 45252
rect 483124 45188 483125 45252
rect 483059 45187 483125 45188
rect 287099 45116 287165 45117
rect 287099 45052 287100 45116
rect 287164 45052 287165 45116
rect 287099 45051 287165 45052
rect 371187 45116 371253 45117
rect 371187 45052 371188 45116
rect 371252 45052 371253 45116
rect 371187 45051 371253 45052
rect 65994 23454 66614 41000
rect 249747 36548 249813 36549
rect 249747 36484 249748 36548
rect 249812 36484 249813 36548
rect 249747 36483 249813 36484
rect 455459 36548 455525 36549
rect 455459 36484 455460 36548
rect 455524 36484 455525 36548
rect 455459 36483 455525 36484
rect 557579 36548 557645 36549
rect 557579 36484 557580 36548
rect 557644 36484 557645 36548
rect 557579 36483 557645 36484
rect 128491 34916 128557 34917
rect 128491 34852 128492 34916
rect 128556 34852 128557 34916
rect 128491 34851 128557 34852
rect 240547 34916 240613 34917
rect 240547 34852 240548 34916
rect 240612 34852 240613 34916
rect 240547 34851 240613 34852
rect 128494 26893 128554 34851
rect 212579 34780 212645 34781
rect 212579 34716 212580 34780
rect 212644 34716 212645 34780
rect 212579 34715 212645 34716
rect 212582 26893 212642 34715
rect 240550 26893 240610 34851
rect 128491 26892 128557 26893
rect 76076 26829 76396 26861
rect 76076 26593 76118 26829
rect 76354 26593 76396 26829
rect 76076 26509 76396 26593
rect 76076 26273 76118 26509
rect 76354 26273 76396 26509
rect 76076 26241 76396 26273
rect 82340 26829 82660 26861
rect 82340 26593 82382 26829
rect 82618 26593 82660 26829
rect 82340 26509 82660 26593
rect 82340 26273 82382 26509
rect 82618 26273 82660 26509
rect 82340 26241 82660 26273
rect 88604 26829 88924 26861
rect 88604 26593 88646 26829
rect 88882 26593 88924 26829
rect 88604 26509 88924 26593
rect 88604 26273 88646 26509
rect 88882 26273 88924 26509
rect 88604 26241 88924 26273
rect 104076 26829 104396 26861
rect 104076 26593 104118 26829
rect 104354 26593 104396 26829
rect 104076 26509 104396 26593
rect 104076 26273 104118 26509
rect 104354 26273 104396 26509
rect 104076 26241 104396 26273
rect 110340 26829 110660 26861
rect 110340 26593 110382 26829
rect 110618 26593 110660 26829
rect 110340 26509 110660 26593
rect 110340 26273 110382 26509
rect 110618 26273 110660 26509
rect 110340 26241 110660 26273
rect 116604 26829 116924 26861
rect 116604 26593 116646 26829
rect 116882 26593 116924 26829
rect 128491 26828 128492 26892
rect 128556 26828 128557 26892
rect 212579 26892 212645 26893
rect 128491 26827 128557 26828
rect 132076 26829 132396 26861
rect 116604 26509 116924 26593
rect 116604 26273 116646 26509
rect 116882 26273 116924 26509
rect 116604 26241 116924 26273
rect 132076 26593 132118 26829
rect 132354 26593 132396 26829
rect 132076 26509 132396 26593
rect 132076 26273 132118 26509
rect 132354 26273 132396 26509
rect 132076 26241 132396 26273
rect 138340 26829 138660 26861
rect 138340 26593 138382 26829
rect 138618 26593 138660 26829
rect 138340 26509 138660 26593
rect 138340 26273 138382 26509
rect 138618 26273 138660 26509
rect 138340 26241 138660 26273
rect 144604 26829 144924 26861
rect 144604 26593 144646 26829
rect 144882 26593 144924 26829
rect 144604 26509 144924 26593
rect 144604 26273 144646 26509
rect 144882 26273 144924 26509
rect 144604 26241 144924 26273
rect 160076 26829 160396 26861
rect 160076 26593 160118 26829
rect 160354 26593 160396 26829
rect 160076 26509 160396 26593
rect 160076 26273 160118 26509
rect 160354 26273 160396 26509
rect 160076 26241 160396 26273
rect 166340 26829 166660 26861
rect 166340 26593 166382 26829
rect 166618 26593 166660 26829
rect 166340 26509 166660 26593
rect 166340 26273 166382 26509
rect 166618 26273 166660 26509
rect 166340 26241 166660 26273
rect 172604 26829 172924 26861
rect 172604 26593 172646 26829
rect 172882 26593 172924 26829
rect 172604 26509 172924 26593
rect 172604 26273 172646 26509
rect 172882 26273 172924 26509
rect 172604 26241 172924 26273
rect 188076 26829 188396 26861
rect 188076 26593 188118 26829
rect 188354 26593 188396 26829
rect 188076 26509 188396 26593
rect 188076 26273 188118 26509
rect 188354 26273 188396 26509
rect 188076 26241 188396 26273
rect 194340 26829 194660 26861
rect 194340 26593 194382 26829
rect 194618 26593 194660 26829
rect 194340 26509 194660 26593
rect 194340 26273 194382 26509
rect 194618 26273 194660 26509
rect 194340 26241 194660 26273
rect 200604 26829 200924 26861
rect 200604 26593 200646 26829
rect 200882 26593 200924 26829
rect 212579 26828 212580 26892
rect 212644 26828 212645 26892
rect 240547 26892 240613 26893
rect 212579 26827 212645 26828
rect 216076 26829 216396 26861
rect 200604 26509 200924 26593
rect 200604 26273 200646 26509
rect 200882 26273 200924 26509
rect 200604 26241 200924 26273
rect 216076 26593 216118 26829
rect 216354 26593 216396 26829
rect 216076 26509 216396 26593
rect 216076 26273 216118 26509
rect 216354 26273 216396 26509
rect 216076 26241 216396 26273
rect 222340 26829 222660 26861
rect 222340 26593 222382 26829
rect 222618 26593 222660 26829
rect 222340 26509 222660 26593
rect 222340 26273 222382 26509
rect 222618 26273 222660 26509
rect 222340 26241 222660 26273
rect 228604 26829 228924 26861
rect 228604 26593 228646 26829
rect 228882 26593 228924 26829
rect 240547 26828 240548 26892
rect 240612 26828 240613 26892
rect 240547 26827 240613 26828
rect 244076 26829 244396 26861
rect 228604 26509 228924 26593
rect 228604 26273 228646 26509
rect 228882 26273 228924 26509
rect 228604 26241 228924 26273
rect 244076 26593 244118 26829
rect 244354 26593 244396 26829
rect 244076 26509 244396 26593
rect 244076 26273 244118 26509
rect 244354 26273 244396 26509
rect 244076 26241 244396 26273
rect 65994 23218 66026 23454
rect 66262 23218 66346 23454
rect 66582 23218 66614 23454
rect 65994 23134 66614 23218
rect 65994 22898 66026 23134
rect 66262 22898 66346 23134
rect 66582 22898 66614 23134
rect 63723 20228 63789 20229
rect 63723 20164 63724 20228
rect 63788 20164 63789 20228
rect 63723 20163 63789 20164
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 65994 -1306 66614 22898
rect 79208 23454 79528 23486
rect 79208 23218 79250 23454
rect 79486 23218 79528 23454
rect 79208 23134 79528 23218
rect 79208 22898 79250 23134
rect 79486 22898 79528 23134
rect 79208 22866 79528 22898
rect 85472 23454 85792 23486
rect 85472 23218 85514 23454
rect 85750 23218 85792 23454
rect 85472 23134 85792 23218
rect 85472 22898 85514 23134
rect 85750 22898 85792 23134
rect 85472 22866 85792 22898
rect 107208 23454 107528 23486
rect 107208 23218 107250 23454
rect 107486 23218 107528 23454
rect 107208 23134 107528 23218
rect 107208 22898 107250 23134
rect 107486 22898 107528 23134
rect 107208 22866 107528 22898
rect 113472 23454 113792 23486
rect 113472 23218 113514 23454
rect 113750 23218 113792 23454
rect 113472 23134 113792 23218
rect 113472 22898 113514 23134
rect 113750 22898 113792 23134
rect 113472 22866 113792 22898
rect 135208 23454 135528 23486
rect 135208 23218 135250 23454
rect 135486 23218 135528 23454
rect 135208 23134 135528 23218
rect 135208 22898 135250 23134
rect 135486 22898 135528 23134
rect 135208 22866 135528 22898
rect 141472 23454 141792 23486
rect 141472 23218 141514 23454
rect 141750 23218 141792 23454
rect 141472 23134 141792 23218
rect 141472 22898 141514 23134
rect 141750 22898 141792 23134
rect 141472 22866 141792 22898
rect 163208 23454 163528 23486
rect 163208 23218 163250 23454
rect 163486 23218 163528 23454
rect 163208 23134 163528 23218
rect 163208 22898 163250 23134
rect 163486 22898 163528 23134
rect 163208 22866 163528 22898
rect 169472 23454 169792 23486
rect 169472 23218 169514 23454
rect 169750 23218 169792 23454
rect 169472 23134 169792 23218
rect 169472 22898 169514 23134
rect 169750 22898 169792 23134
rect 169472 22866 169792 22898
rect 191208 23454 191528 23486
rect 191208 23218 191250 23454
rect 191486 23218 191528 23454
rect 191208 23134 191528 23218
rect 191208 22898 191250 23134
rect 191486 22898 191528 23134
rect 191208 22866 191528 22898
rect 197472 23454 197792 23486
rect 197472 23218 197514 23454
rect 197750 23218 197792 23454
rect 197472 23134 197792 23218
rect 197472 22898 197514 23134
rect 197750 22898 197792 23134
rect 197472 22866 197792 22898
rect 219208 23454 219528 23486
rect 219208 23218 219250 23454
rect 219486 23218 219528 23454
rect 219208 23134 219528 23218
rect 219208 22898 219250 23134
rect 219486 22898 219528 23134
rect 219208 22866 219528 22898
rect 225472 23454 225792 23486
rect 225472 23218 225514 23454
rect 225750 23218 225792 23454
rect 225472 23134 225792 23218
rect 225472 22898 225514 23134
rect 225750 22898 225792 23134
rect 225472 22866 225792 22898
rect 247208 23454 247528 23486
rect 247208 23218 247250 23454
rect 247486 23218 247528 23454
rect 247208 23134 247528 23218
rect 247208 22898 247250 23134
rect 247486 22898 247528 23134
rect 247208 22866 247528 22898
rect 249750 13429 249810 36483
rect 296851 35052 296917 35053
rect 296851 34988 296852 35052
rect 296916 34988 296917 35052
rect 296851 34987 296917 34988
rect 296854 29010 296914 34987
rect 324635 34916 324701 34917
rect 324635 34852 324636 34916
rect 324700 34852 324701 34916
rect 324635 34851 324701 34852
rect 436507 34916 436573 34917
rect 436507 34852 436508 34916
rect 436572 34852 436573 34916
rect 436507 34851 436573 34852
rect 296486 28950 296914 29010
rect 296486 26893 296546 28950
rect 324638 26893 324698 34851
rect 408539 34780 408605 34781
rect 408539 34716 408540 34780
rect 408604 34716 408605 34780
rect 408539 34715 408605 34716
rect 408542 26893 408602 34715
rect 436510 26893 436570 34851
rect 296483 26892 296549 26893
rect 250340 26829 250660 26861
rect 250340 26593 250382 26829
rect 250618 26593 250660 26829
rect 250340 26509 250660 26593
rect 250340 26273 250382 26509
rect 250618 26273 250660 26509
rect 250340 26241 250660 26273
rect 256604 26829 256924 26861
rect 256604 26593 256646 26829
rect 256882 26593 256924 26829
rect 256604 26509 256924 26593
rect 256604 26273 256646 26509
rect 256882 26273 256924 26509
rect 256604 26241 256924 26273
rect 272076 26829 272396 26861
rect 272076 26593 272118 26829
rect 272354 26593 272396 26829
rect 272076 26509 272396 26593
rect 272076 26273 272118 26509
rect 272354 26273 272396 26509
rect 272076 26241 272396 26273
rect 278340 26829 278660 26861
rect 278340 26593 278382 26829
rect 278618 26593 278660 26829
rect 278340 26509 278660 26593
rect 278340 26273 278382 26509
rect 278618 26273 278660 26509
rect 278340 26241 278660 26273
rect 284604 26829 284924 26861
rect 284604 26593 284646 26829
rect 284882 26593 284924 26829
rect 296483 26828 296484 26892
rect 296548 26828 296549 26892
rect 324635 26892 324701 26893
rect 296483 26827 296549 26828
rect 300076 26829 300396 26861
rect 284604 26509 284924 26593
rect 284604 26273 284646 26509
rect 284882 26273 284924 26509
rect 284604 26241 284924 26273
rect 300076 26593 300118 26829
rect 300354 26593 300396 26829
rect 300076 26509 300396 26593
rect 300076 26273 300118 26509
rect 300354 26273 300396 26509
rect 300076 26241 300396 26273
rect 306340 26829 306660 26861
rect 306340 26593 306382 26829
rect 306618 26593 306660 26829
rect 306340 26509 306660 26593
rect 306340 26273 306382 26509
rect 306618 26273 306660 26509
rect 306340 26241 306660 26273
rect 312604 26829 312924 26861
rect 312604 26593 312646 26829
rect 312882 26593 312924 26829
rect 324635 26828 324636 26892
rect 324700 26828 324701 26892
rect 408539 26892 408605 26893
rect 324635 26827 324701 26828
rect 328076 26829 328396 26861
rect 312604 26509 312924 26593
rect 312604 26273 312646 26509
rect 312882 26273 312924 26509
rect 312604 26241 312924 26273
rect 328076 26593 328118 26829
rect 328354 26593 328396 26829
rect 328076 26509 328396 26593
rect 328076 26273 328118 26509
rect 328354 26273 328396 26509
rect 328076 26241 328396 26273
rect 334340 26829 334660 26861
rect 334340 26593 334382 26829
rect 334618 26593 334660 26829
rect 334340 26509 334660 26593
rect 334340 26273 334382 26509
rect 334618 26273 334660 26509
rect 334340 26241 334660 26273
rect 340604 26829 340924 26861
rect 340604 26593 340646 26829
rect 340882 26593 340924 26829
rect 340604 26509 340924 26593
rect 340604 26273 340646 26509
rect 340882 26273 340924 26509
rect 340604 26241 340924 26273
rect 355293 26829 355613 26861
rect 355293 26593 355335 26829
rect 355571 26593 355613 26829
rect 355293 26509 355613 26593
rect 355293 26273 355335 26509
rect 355571 26273 355613 26509
rect 355293 26241 355613 26273
rect 359991 26829 360311 26861
rect 359991 26593 360033 26829
rect 360269 26593 360311 26829
rect 359991 26509 360311 26593
rect 359991 26273 360033 26509
rect 360269 26273 360311 26509
rect 359991 26241 360311 26273
rect 364689 26829 365009 26861
rect 364689 26593 364731 26829
rect 364967 26593 365009 26829
rect 364689 26509 365009 26593
rect 364689 26273 364731 26509
rect 364967 26273 365009 26509
rect 364689 26241 365009 26273
rect 369387 26829 369707 26861
rect 369387 26593 369429 26829
rect 369665 26593 369707 26829
rect 369387 26509 369707 26593
rect 369387 26273 369429 26509
rect 369665 26273 369707 26509
rect 369387 26241 369707 26273
rect 384076 26829 384396 26861
rect 384076 26593 384118 26829
rect 384354 26593 384396 26829
rect 384076 26509 384396 26593
rect 384076 26273 384118 26509
rect 384354 26273 384396 26509
rect 384076 26241 384396 26273
rect 390340 26829 390660 26861
rect 390340 26593 390382 26829
rect 390618 26593 390660 26829
rect 390340 26509 390660 26593
rect 390340 26273 390382 26509
rect 390618 26273 390660 26509
rect 390340 26241 390660 26273
rect 396604 26829 396924 26861
rect 396604 26593 396646 26829
rect 396882 26593 396924 26829
rect 408539 26828 408540 26892
rect 408604 26828 408605 26892
rect 436507 26892 436573 26893
rect 408539 26827 408605 26828
rect 412076 26829 412396 26861
rect 396604 26509 396924 26593
rect 396604 26273 396646 26509
rect 396882 26273 396924 26509
rect 396604 26241 396924 26273
rect 412076 26593 412118 26829
rect 412354 26593 412396 26829
rect 412076 26509 412396 26593
rect 412076 26273 412118 26509
rect 412354 26273 412396 26509
rect 412076 26241 412396 26273
rect 418340 26829 418660 26861
rect 418340 26593 418382 26829
rect 418618 26593 418660 26829
rect 418340 26509 418660 26593
rect 418340 26273 418382 26509
rect 418618 26273 418660 26509
rect 418340 26241 418660 26273
rect 424604 26829 424924 26861
rect 424604 26593 424646 26829
rect 424882 26593 424924 26829
rect 436507 26828 436508 26892
rect 436572 26828 436573 26892
rect 436507 26827 436573 26828
rect 440076 26829 440396 26861
rect 424604 26509 424924 26593
rect 424604 26273 424646 26509
rect 424882 26273 424924 26509
rect 424604 26241 424924 26273
rect 440076 26593 440118 26829
rect 440354 26593 440396 26829
rect 440076 26509 440396 26593
rect 440076 26273 440118 26509
rect 440354 26273 440396 26509
rect 440076 26241 440396 26273
rect 446340 26829 446660 26861
rect 446340 26593 446382 26829
rect 446618 26593 446660 26829
rect 446340 26509 446660 26593
rect 446340 26273 446382 26509
rect 446618 26273 446660 26509
rect 446340 26241 446660 26273
rect 452604 26829 452924 26861
rect 452604 26593 452646 26829
rect 452882 26593 452924 26829
rect 452604 26509 452924 26593
rect 452604 26273 452646 26509
rect 452882 26273 452924 26509
rect 452604 26241 452924 26273
rect 253472 23454 253792 23486
rect 253472 23218 253514 23454
rect 253750 23218 253792 23454
rect 253472 23134 253792 23218
rect 253472 22898 253514 23134
rect 253750 22898 253792 23134
rect 253472 22866 253792 22898
rect 275208 23454 275528 23486
rect 275208 23218 275250 23454
rect 275486 23218 275528 23454
rect 275208 23134 275528 23218
rect 275208 22898 275250 23134
rect 275486 22898 275528 23134
rect 275208 22866 275528 22898
rect 281472 23454 281792 23486
rect 281472 23218 281514 23454
rect 281750 23218 281792 23454
rect 281472 23134 281792 23218
rect 281472 22898 281514 23134
rect 281750 22898 281792 23134
rect 281472 22866 281792 22898
rect 303208 23454 303528 23486
rect 303208 23218 303250 23454
rect 303486 23218 303528 23454
rect 303208 23134 303528 23218
rect 303208 22898 303250 23134
rect 303486 22898 303528 23134
rect 303208 22866 303528 22898
rect 309472 23454 309792 23486
rect 309472 23218 309514 23454
rect 309750 23218 309792 23454
rect 309472 23134 309792 23218
rect 309472 22898 309514 23134
rect 309750 22898 309792 23134
rect 309472 22866 309792 22898
rect 331208 23454 331528 23486
rect 331208 23218 331250 23454
rect 331486 23218 331528 23454
rect 331208 23134 331528 23218
rect 331208 22898 331250 23134
rect 331486 22898 331528 23134
rect 331208 22866 331528 22898
rect 337472 23454 337792 23486
rect 337472 23218 337514 23454
rect 337750 23218 337792 23454
rect 337472 23134 337792 23218
rect 337472 22898 337514 23134
rect 337750 22898 337792 23134
rect 337472 22866 337792 22898
rect 357642 23454 357962 23486
rect 357642 23218 357684 23454
rect 357920 23218 357962 23454
rect 357642 23134 357962 23218
rect 357642 22898 357684 23134
rect 357920 22898 357962 23134
rect 357642 22866 357962 22898
rect 362340 23454 362660 23486
rect 362340 23218 362382 23454
rect 362618 23218 362660 23454
rect 362340 23134 362660 23218
rect 362340 22898 362382 23134
rect 362618 22898 362660 23134
rect 362340 22866 362660 22898
rect 367038 23454 367358 23486
rect 367038 23218 367080 23454
rect 367316 23218 367358 23454
rect 367038 23134 367358 23218
rect 367038 22898 367080 23134
rect 367316 22898 367358 23134
rect 367038 22866 367358 22898
rect 387208 23454 387528 23486
rect 387208 23218 387250 23454
rect 387486 23218 387528 23454
rect 387208 23134 387528 23218
rect 387208 22898 387250 23134
rect 387486 22898 387528 23134
rect 387208 22866 387528 22898
rect 393472 23454 393792 23486
rect 393472 23218 393514 23454
rect 393750 23218 393792 23454
rect 393472 23134 393792 23218
rect 393472 22898 393514 23134
rect 393750 22898 393792 23134
rect 393472 22866 393792 22898
rect 415208 23454 415528 23486
rect 415208 23218 415250 23454
rect 415486 23218 415528 23454
rect 415208 23134 415528 23218
rect 415208 22898 415250 23134
rect 415486 22898 415528 23134
rect 415208 22866 415528 22898
rect 421472 23454 421792 23486
rect 421472 23218 421514 23454
rect 421750 23218 421792 23454
rect 421472 23134 421792 23218
rect 421472 22898 421514 23134
rect 421750 22898 421792 23134
rect 421472 22866 421792 22898
rect 443208 23454 443528 23486
rect 443208 23218 443250 23454
rect 443486 23218 443528 23454
rect 443208 23134 443528 23218
rect 443208 22898 443250 23134
rect 443486 22898 443528 23134
rect 443208 22866 443528 22898
rect 449472 23454 449792 23486
rect 449472 23218 449514 23454
rect 449750 23218 449792 23454
rect 449472 23134 449792 23218
rect 449472 22898 449514 23134
rect 449750 22898 449792 23134
rect 449472 22866 449792 22898
rect 455462 13429 455522 36483
rect 492627 34916 492693 34917
rect 492627 34852 492628 34916
rect 492692 34852 492693 34916
rect 492627 34851 492693 34852
rect 492630 26893 492690 34851
rect 520595 34780 520661 34781
rect 520595 34716 520596 34780
rect 520660 34716 520661 34780
rect 520595 34715 520661 34716
rect 520598 26893 520658 34715
rect 492627 26892 492693 26893
rect 468076 26829 468396 26861
rect 468076 26593 468118 26829
rect 468354 26593 468396 26829
rect 468076 26509 468396 26593
rect 468076 26273 468118 26509
rect 468354 26273 468396 26509
rect 468076 26241 468396 26273
rect 474340 26829 474660 26861
rect 474340 26593 474382 26829
rect 474618 26593 474660 26829
rect 474340 26509 474660 26593
rect 474340 26273 474382 26509
rect 474618 26273 474660 26509
rect 474340 26241 474660 26273
rect 480604 26829 480924 26861
rect 480604 26593 480646 26829
rect 480882 26593 480924 26829
rect 492627 26828 492628 26892
rect 492692 26828 492693 26892
rect 520595 26892 520661 26893
rect 492627 26827 492693 26828
rect 496076 26829 496396 26861
rect 480604 26509 480924 26593
rect 480604 26273 480646 26509
rect 480882 26273 480924 26509
rect 480604 26241 480924 26273
rect 496076 26593 496118 26829
rect 496354 26593 496396 26829
rect 496076 26509 496396 26593
rect 496076 26273 496118 26509
rect 496354 26273 496396 26509
rect 496076 26241 496396 26273
rect 502340 26829 502660 26861
rect 502340 26593 502382 26829
rect 502618 26593 502660 26829
rect 502340 26509 502660 26593
rect 502340 26273 502382 26509
rect 502618 26273 502660 26509
rect 502340 26241 502660 26273
rect 508604 26829 508924 26861
rect 508604 26593 508646 26829
rect 508882 26593 508924 26829
rect 520595 26828 520596 26892
rect 520660 26828 520661 26892
rect 520595 26827 520661 26828
rect 524076 26829 524396 26861
rect 508604 26509 508924 26593
rect 508604 26273 508646 26509
rect 508882 26273 508924 26509
rect 508604 26241 508924 26273
rect 524076 26593 524118 26829
rect 524354 26593 524396 26829
rect 524076 26509 524396 26593
rect 524076 26273 524118 26509
rect 524354 26273 524396 26509
rect 524076 26241 524396 26273
rect 530340 26829 530660 26861
rect 530340 26593 530382 26829
rect 530618 26593 530660 26829
rect 530340 26509 530660 26593
rect 530340 26273 530382 26509
rect 530618 26273 530660 26509
rect 530340 26241 530660 26273
rect 536604 26829 536924 26861
rect 536604 26593 536646 26829
rect 536882 26593 536924 26829
rect 536604 26509 536924 26593
rect 536604 26273 536646 26509
rect 536882 26273 536924 26509
rect 536604 26241 536924 26273
rect 552076 26829 552396 26861
rect 552076 26593 552118 26829
rect 552354 26593 552396 26829
rect 552076 26509 552396 26593
rect 552076 26273 552118 26509
rect 552354 26273 552396 26509
rect 552076 26241 552396 26273
rect 471208 23454 471528 23486
rect 471208 23218 471250 23454
rect 471486 23218 471528 23454
rect 471208 23134 471528 23218
rect 471208 22898 471250 23134
rect 471486 22898 471528 23134
rect 471208 22866 471528 22898
rect 477472 23454 477792 23486
rect 477472 23218 477514 23454
rect 477750 23218 477792 23454
rect 477472 23134 477792 23218
rect 477472 22898 477514 23134
rect 477750 22898 477792 23134
rect 477472 22866 477792 22898
rect 499208 23454 499528 23486
rect 499208 23218 499250 23454
rect 499486 23218 499528 23454
rect 499208 23134 499528 23218
rect 499208 22898 499250 23134
rect 499486 22898 499528 23134
rect 499208 22866 499528 22898
rect 505472 23454 505792 23486
rect 505472 23218 505514 23454
rect 505750 23218 505792 23454
rect 505472 23134 505792 23218
rect 505472 22898 505514 23134
rect 505750 22898 505792 23134
rect 505472 22866 505792 22898
rect 527208 23454 527528 23486
rect 527208 23218 527250 23454
rect 527486 23218 527528 23454
rect 527208 23134 527528 23218
rect 527208 22898 527250 23134
rect 527486 22898 527528 23134
rect 527208 22866 527528 22898
rect 533472 23454 533792 23486
rect 533472 23218 533514 23454
rect 533750 23218 533792 23454
rect 533472 23134 533792 23218
rect 533472 22898 533514 23134
rect 533750 22898 533792 23134
rect 533472 22866 533792 22898
rect 555208 23454 555528 23486
rect 555208 23218 555250 23454
rect 555486 23218 555528 23454
rect 555208 23134 555528 23218
rect 555208 22898 555250 23134
rect 555486 22898 555528 23134
rect 555208 22866 555528 22898
rect 557582 13429 557642 36483
rect 558340 26829 558660 26861
rect 558340 26593 558382 26829
rect 558618 26593 558660 26829
rect 558340 26509 558660 26593
rect 558340 26273 558382 26509
rect 558618 26273 558660 26509
rect 558340 26241 558660 26273
rect 564604 26829 564924 26861
rect 564604 26593 564646 26829
rect 564882 26593 564924 26829
rect 564604 26509 564924 26593
rect 564604 26273 564646 26509
rect 564882 26273 564924 26509
rect 564604 26241 564924 26273
rect 573494 26829 574114 53273
rect 580214 37909 580274 697171
rect 585310 674829 585930 701273
rect 585310 674593 585342 674829
rect 585578 674593 585662 674829
rect 585898 674593 585930 674829
rect 585310 674509 585930 674593
rect 585310 674273 585342 674509
rect 585578 674273 585662 674509
rect 585898 674273 585930 674509
rect 580395 670716 580461 670717
rect 580395 670652 580396 670716
rect 580460 670652 580461 670716
rect 580395 670651 580461 670652
rect 580211 37908 580277 37909
rect 580211 37844 580212 37908
rect 580276 37844 580277 37908
rect 580211 37843 580277 37844
rect 573494 26593 573526 26829
rect 573762 26593 573846 26829
rect 574082 26593 574114 26829
rect 573494 26509 574114 26593
rect 573494 26273 573526 26509
rect 573762 26273 573846 26509
rect 574082 26273 574114 26509
rect 561472 23454 561792 23486
rect 561472 23218 561514 23454
rect 561750 23218 561792 23454
rect 561472 23134 561792 23218
rect 561472 22898 561514 23134
rect 561750 22898 561792 23134
rect 561472 22866 561792 22898
rect 249747 13428 249813 13429
rect 249747 13364 249748 13428
rect 249812 13364 249813 13428
rect 249747 13363 249813 13364
rect 455459 13428 455525 13429
rect 455459 13364 455460 13428
rect 455524 13364 455525 13428
rect 455459 13363 455525 13364
rect 557579 13428 557645 13429
rect 557579 13364 557580 13428
rect 557644 13364 557645 13428
rect 557579 13363 557645 13364
rect 65994 -1542 66026 -1306
rect 66262 -1542 66346 -1306
rect 66582 -1542 66614 -1306
rect 65994 -1626 66614 -1542
rect 65994 -1862 66026 -1626
rect 66262 -1862 66346 -1626
rect 66582 -1862 66614 -1626
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 65994 -7654 66614 -1862
rect 573494 -346 574114 26273
rect 580398 13565 580458 670651
rect 585310 647829 585930 674273
rect 585310 647593 585342 647829
rect 585578 647593 585662 647829
rect 585898 647593 585930 647829
rect 585310 647509 585930 647593
rect 585310 647273 585342 647509
rect 585578 647273 585662 647509
rect 585898 647273 585930 647509
rect 580579 644060 580645 644061
rect 580579 643996 580580 644060
rect 580644 643996 580645 644060
rect 580579 643995 580645 643996
rect 580582 13701 580642 643995
rect 585310 620829 585930 647273
rect 585310 620593 585342 620829
rect 585578 620593 585662 620829
rect 585898 620593 585930 620829
rect 585310 620509 585930 620593
rect 585310 620273 585342 620509
rect 585578 620273 585662 620509
rect 585898 620273 585930 620509
rect 585310 593829 585930 620273
rect 585310 593593 585342 593829
rect 585578 593593 585662 593829
rect 585898 593593 585930 593829
rect 585310 593509 585930 593593
rect 585310 593273 585342 593509
rect 585578 593273 585662 593509
rect 585898 593273 585930 593509
rect 585310 566829 585930 593273
rect 585310 566593 585342 566829
rect 585578 566593 585662 566829
rect 585898 566593 585930 566829
rect 585310 566509 585930 566593
rect 585310 566273 585342 566509
rect 585578 566273 585662 566509
rect 585898 566273 585930 566509
rect 585310 539829 585930 566273
rect 585310 539593 585342 539829
rect 585578 539593 585662 539829
rect 585898 539593 585930 539829
rect 585310 539509 585930 539593
rect 585310 539273 585342 539509
rect 585578 539273 585662 539509
rect 585898 539273 585930 539509
rect 585310 512829 585930 539273
rect 585310 512593 585342 512829
rect 585578 512593 585662 512829
rect 585898 512593 585930 512829
rect 585310 512509 585930 512593
rect 585310 512273 585342 512509
rect 585578 512273 585662 512509
rect 585898 512273 585930 512509
rect 585310 485829 585930 512273
rect 585310 485593 585342 485829
rect 585578 485593 585662 485829
rect 585898 485593 585930 485829
rect 585310 485509 585930 485593
rect 585310 485273 585342 485509
rect 585578 485273 585662 485509
rect 585898 485273 585930 485509
rect 585310 458829 585930 485273
rect 585310 458593 585342 458829
rect 585578 458593 585662 458829
rect 585898 458593 585930 458829
rect 585310 458509 585930 458593
rect 585310 458273 585342 458509
rect 585578 458273 585662 458509
rect 585898 458273 585930 458509
rect 585310 431829 585930 458273
rect 585310 431593 585342 431829
rect 585578 431593 585662 431829
rect 585898 431593 585930 431829
rect 585310 431509 585930 431593
rect 585310 431273 585342 431509
rect 585578 431273 585662 431509
rect 585898 431273 585930 431509
rect 585310 404829 585930 431273
rect 585310 404593 585342 404829
rect 585578 404593 585662 404829
rect 585898 404593 585930 404829
rect 585310 404509 585930 404593
rect 585310 404273 585342 404509
rect 585578 404273 585662 404509
rect 585898 404273 585930 404509
rect 585310 377829 585930 404273
rect 585310 377593 585342 377829
rect 585578 377593 585662 377829
rect 585898 377593 585930 377829
rect 585310 377509 585930 377593
rect 585310 377273 585342 377509
rect 585578 377273 585662 377509
rect 585898 377273 585930 377509
rect 585310 350829 585930 377273
rect 585310 350593 585342 350829
rect 585578 350593 585662 350829
rect 585898 350593 585930 350829
rect 585310 350509 585930 350593
rect 585310 350273 585342 350509
rect 585578 350273 585662 350509
rect 585898 350273 585930 350509
rect 585310 323829 585930 350273
rect 585310 323593 585342 323829
rect 585578 323593 585662 323829
rect 585898 323593 585930 323829
rect 585310 323509 585930 323593
rect 585310 323273 585342 323509
rect 585578 323273 585662 323509
rect 585898 323273 585930 323509
rect 585310 296829 585930 323273
rect 585310 296593 585342 296829
rect 585578 296593 585662 296829
rect 585898 296593 585930 296829
rect 585310 296509 585930 296593
rect 585310 296273 585342 296509
rect 585578 296273 585662 296509
rect 585898 296273 585930 296509
rect 585310 269829 585930 296273
rect 585310 269593 585342 269829
rect 585578 269593 585662 269829
rect 585898 269593 585930 269829
rect 585310 269509 585930 269593
rect 585310 269273 585342 269509
rect 585578 269273 585662 269509
rect 585898 269273 585930 269509
rect 585310 242829 585930 269273
rect 585310 242593 585342 242829
rect 585578 242593 585662 242829
rect 585898 242593 585930 242829
rect 585310 242509 585930 242593
rect 585310 242273 585342 242509
rect 585578 242273 585662 242509
rect 585898 242273 585930 242509
rect 585310 215829 585930 242273
rect 585310 215593 585342 215829
rect 585578 215593 585662 215829
rect 585898 215593 585930 215829
rect 585310 215509 585930 215593
rect 585310 215273 585342 215509
rect 585578 215273 585662 215509
rect 585898 215273 585930 215509
rect 585310 188829 585930 215273
rect 585310 188593 585342 188829
rect 585578 188593 585662 188829
rect 585898 188593 585930 188829
rect 585310 188509 585930 188593
rect 585310 188273 585342 188509
rect 585578 188273 585662 188509
rect 585898 188273 585930 188509
rect 585310 161829 585930 188273
rect 585310 161593 585342 161829
rect 585578 161593 585662 161829
rect 585898 161593 585930 161829
rect 585310 161509 585930 161593
rect 585310 161273 585342 161509
rect 585578 161273 585662 161509
rect 585898 161273 585930 161509
rect 585310 134829 585930 161273
rect 585310 134593 585342 134829
rect 585578 134593 585662 134829
rect 585898 134593 585930 134829
rect 585310 134509 585930 134593
rect 585310 134273 585342 134509
rect 585578 134273 585662 134509
rect 585898 134273 585930 134509
rect 585310 107829 585930 134273
rect 585310 107593 585342 107829
rect 585578 107593 585662 107829
rect 585898 107593 585930 107829
rect 585310 107509 585930 107593
rect 585310 107273 585342 107509
rect 585578 107273 585662 107509
rect 585898 107273 585930 107509
rect 585310 80829 585930 107273
rect 585310 80593 585342 80829
rect 585578 80593 585662 80829
rect 585898 80593 585930 80829
rect 585310 80509 585930 80593
rect 585310 80273 585342 80509
rect 585578 80273 585662 80509
rect 585898 80273 585930 80509
rect 585310 53829 585930 80273
rect 585310 53593 585342 53829
rect 585578 53593 585662 53829
rect 585898 53593 585930 53829
rect 585310 53509 585930 53593
rect 585310 53273 585342 53509
rect 585578 53273 585662 53509
rect 585898 53273 585930 53509
rect 585310 26829 585930 53273
rect 585310 26593 585342 26829
rect 585578 26593 585662 26829
rect 585898 26593 585930 26829
rect 585310 26509 585930 26593
rect 585310 26273 585342 26509
rect 585578 26273 585662 26509
rect 585898 26273 585930 26509
rect 580579 13700 580645 13701
rect 580579 13636 580580 13700
rect 580644 13636 580645 13700
rect 580579 13635 580645 13636
rect 580395 13564 580461 13565
rect 580395 13500 580396 13564
rect 580460 13500 580461 13564
rect 580395 13499 580461 13500
rect 573494 -582 573526 -346
rect 573762 -582 573846 -346
rect 574082 -582 574114 -346
rect 573494 -666 574114 -582
rect 573494 -902 573526 -666
rect 573762 -902 573846 -666
rect 574082 -902 574114 -666
rect 573494 -7654 574114 -902
rect 585310 -346 585930 26273
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 698454 586890 705242
rect 586270 698218 586302 698454
rect 586538 698218 586622 698454
rect 586858 698218 586890 698454
rect 586270 698134 586890 698218
rect 586270 697898 586302 698134
rect 586538 697898 586622 698134
rect 586858 697898 586890 698134
rect 586270 671454 586890 697898
rect 586270 671218 586302 671454
rect 586538 671218 586622 671454
rect 586858 671218 586890 671454
rect 586270 671134 586890 671218
rect 586270 670898 586302 671134
rect 586538 670898 586622 671134
rect 586858 670898 586890 671134
rect 586270 644454 586890 670898
rect 586270 644218 586302 644454
rect 586538 644218 586622 644454
rect 586858 644218 586890 644454
rect 586270 644134 586890 644218
rect 586270 643898 586302 644134
rect 586538 643898 586622 644134
rect 586858 643898 586890 644134
rect 586270 617454 586890 643898
rect 586270 617218 586302 617454
rect 586538 617218 586622 617454
rect 586858 617218 586890 617454
rect 586270 617134 586890 617218
rect 586270 616898 586302 617134
rect 586538 616898 586622 617134
rect 586858 616898 586890 617134
rect 586270 590454 586890 616898
rect 586270 590218 586302 590454
rect 586538 590218 586622 590454
rect 586858 590218 586890 590454
rect 586270 590134 586890 590218
rect 586270 589898 586302 590134
rect 586538 589898 586622 590134
rect 586858 589898 586890 590134
rect 586270 563454 586890 589898
rect 586270 563218 586302 563454
rect 586538 563218 586622 563454
rect 586858 563218 586890 563454
rect 586270 563134 586890 563218
rect 586270 562898 586302 563134
rect 586538 562898 586622 563134
rect 586858 562898 586890 563134
rect 586270 536454 586890 562898
rect 586270 536218 586302 536454
rect 586538 536218 586622 536454
rect 586858 536218 586890 536454
rect 586270 536134 586890 536218
rect 586270 535898 586302 536134
rect 586538 535898 586622 536134
rect 586858 535898 586890 536134
rect 586270 509454 586890 535898
rect 586270 509218 586302 509454
rect 586538 509218 586622 509454
rect 586858 509218 586890 509454
rect 586270 509134 586890 509218
rect 586270 508898 586302 509134
rect 586538 508898 586622 509134
rect 586858 508898 586890 509134
rect 586270 482454 586890 508898
rect 586270 482218 586302 482454
rect 586538 482218 586622 482454
rect 586858 482218 586890 482454
rect 586270 482134 586890 482218
rect 586270 481898 586302 482134
rect 586538 481898 586622 482134
rect 586858 481898 586890 482134
rect 586270 455454 586890 481898
rect 586270 455218 586302 455454
rect 586538 455218 586622 455454
rect 586858 455218 586890 455454
rect 586270 455134 586890 455218
rect 586270 454898 586302 455134
rect 586538 454898 586622 455134
rect 586858 454898 586890 455134
rect 586270 428454 586890 454898
rect 586270 428218 586302 428454
rect 586538 428218 586622 428454
rect 586858 428218 586890 428454
rect 586270 428134 586890 428218
rect 586270 427898 586302 428134
rect 586538 427898 586622 428134
rect 586858 427898 586890 428134
rect 586270 401454 586890 427898
rect 586270 401218 586302 401454
rect 586538 401218 586622 401454
rect 586858 401218 586890 401454
rect 586270 401134 586890 401218
rect 586270 400898 586302 401134
rect 586538 400898 586622 401134
rect 586858 400898 586890 401134
rect 586270 374454 586890 400898
rect 586270 374218 586302 374454
rect 586538 374218 586622 374454
rect 586858 374218 586890 374454
rect 586270 374134 586890 374218
rect 586270 373898 586302 374134
rect 586538 373898 586622 374134
rect 586858 373898 586890 374134
rect 586270 347454 586890 373898
rect 586270 347218 586302 347454
rect 586538 347218 586622 347454
rect 586858 347218 586890 347454
rect 586270 347134 586890 347218
rect 586270 346898 586302 347134
rect 586538 346898 586622 347134
rect 586858 346898 586890 347134
rect 586270 320454 586890 346898
rect 586270 320218 586302 320454
rect 586538 320218 586622 320454
rect 586858 320218 586890 320454
rect 586270 320134 586890 320218
rect 586270 319898 586302 320134
rect 586538 319898 586622 320134
rect 586858 319898 586890 320134
rect 586270 293454 586890 319898
rect 586270 293218 586302 293454
rect 586538 293218 586622 293454
rect 586858 293218 586890 293454
rect 586270 293134 586890 293218
rect 586270 292898 586302 293134
rect 586538 292898 586622 293134
rect 586858 292898 586890 293134
rect 586270 266454 586890 292898
rect 586270 266218 586302 266454
rect 586538 266218 586622 266454
rect 586858 266218 586890 266454
rect 586270 266134 586890 266218
rect 586270 265898 586302 266134
rect 586538 265898 586622 266134
rect 586858 265898 586890 266134
rect 586270 239454 586890 265898
rect 586270 239218 586302 239454
rect 586538 239218 586622 239454
rect 586858 239218 586890 239454
rect 586270 239134 586890 239218
rect 586270 238898 586302 239134
rect 586538 238898 586622 239134
rect 586858 238898 586890 239134
rect 586270 212454 586890 238898
rect 586270 212218 586302 212454
rect 586538 212218 586622 212454
rect 586858 212218 586890 212454
rect 586270 212134 586890 212218
rect 586270 211898 586302 212134
rect 586538 211898 586622 212134
rect 586858 211898 586890 212134
rect 586270 185454 586890 211898
rect 586270 185218 586302 185454
rect 586538 185218 586622 185454
rect 586858 185218 586890 185454
rect 586270 185134 586890 185218
rect 586270 184898 586302 185134
rect 586538 184898 586622 185134
rect 586858 184898 586890 185134
rect 586270 158454 586890 184898
rect 586270 158218 586302 158454
rect 586538 158218 586622 158454
rect 586858 158218 586890 158454
rect 586270 158134 586890 158218
rect 586270 157898 586302 158134
rect 586538 157898 586622 158134
rect 586858 157898 586890 158134
rect 586270 131454 586890 157898
rect 586270 131218 586302 131454
rect 586538 131218 586622 131454
rect 586858 131218 586890 131454
rect 586270 131134 586890 131218
rect 586270 130898 586302 131134
rect 586538 130898 586622 131134
rect 586858 130898 586890 131134
rect 586270 104454 586890 130898
rect 586270 104218 586302 104454
rect 586538 104218 586622 104454
rect 586858 104218 586890 104454
rect 586270 104134 586890 104218
rect 586270 103898 586302 104134
rect 586538 103898 586622 104134
rect 586858 103898 586890 104134
rect 586270 77454 586890 103898
rect 586270 77218 586302 77454
rect 586538 77218 586622 77454
rect 586858 77218 586890 77454
rect 586270 77134 586890 77218
rect 586270 76898 586302 77134
rect 586538 76898 586622 77134
rect 586858 76898 586890 77134
rect 586270 50454 586890 76898
rect 586270 50218 586302 50454
rect 586538 50218 586622 50454
rect 586858 50218 586890 50454
rect 586270 50134 586890 50218
rect 586270 49898 586302 50134
rect 586538 49898 586622 50134
rect 586858 49898 586890 50134
rect 586270 23454 586890 49898
rect 586270 23218 586302 23454
rect 586538 23218 586622 23454
rect 586858 23218 586890 23454
rect 586270 23134 586890 23218
rect 586270 22898 586302 23134
rect 586538 22898 586622 23134
rect 586858 22898 586890 23134
rect 586270 -1306 586890 22898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 -2266 587850 706202
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 -3226 588810 707162
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 -4186 589770 708122
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 -5146 590730 709082
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 -6106 591690 710042
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 -7066 592650 711002
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect 38026 705562 38262 705798
rect 38346 705562 38582 705798
rect 38026 705242 38262 705478
rect 38346 705242 38582 705478
rect -2934 698218 -2698 698454
rect -2614 698218 -2378 698454
rect -2934 697898 -2698 698134
rect -2614 697898 -2378 698134
rect -2934 671218 -2698 671454
rect -2614 671218 -2378 671454
rect -2934 670898 -2698 671134
rect -2614 670898 -2378 671134
rect -2934 644218 -2698 644454
rect -2614 644218 -2378 644454
rect -2934 643898 -2698 644134
rect -2614 643898 -2378 644134
rect -2934 617218 -2698 617454
rect -2614 617218 -2378 617454
rect -2934 616898 -2698 617134
rect -2614 616898 -2378 617134
rect -2934 590218 -2698 590454
rect -2614 590218 -2378 590454
rect -2934 589898 -2698 590134
rect -2614 589898 -2378 590134
rect -2934 563218 -2698 563454
rect -2614 563218 -2378 563454
rect -2934 562898 -2698 563134
rect -2614 562898 -2378 563134
rect -2934 536218 -2698 536454
rect -2614 536218 -2378 536454
rect -2934 535898 -2698 536134
rect -2614 535898 -2378 536134
rect -2934 509218 -2698 509454
rect -2614 509218 -2378 509454
rect -2934 508898 -2698 509134
rect -2614 508898 -2378 509134
rect -2934 482218 -2698 482454
rect -2614 482218 -2378 482454
rect -2934 481898 -2698 482134
rect -2614 481898 -2378 482134
rect -2934 455218 -2698 455454
rect -2614 455218 -2378 455454
rect -2934 454898 -2698 455134
rect -2614 454898 -2378 455134
rect -2934 428218 -2698 428454
rect -2614 428218 -2378 428454
rect -2934 427898 -2698 428134
rect -2614 427898 -2378 428134
rect -2934 401218 -2698 401454
rect -2614 401218 -2378 401454
rect -2934 400898 -2698 401134
rect -2614 400898 -2378 401134
rect -2934 374218 -2698 374454
rect -2614 374218 -2378 374454
rect -2934 373898 -2698 374134
rect -2614 373898 -2378 374134
rect -2934 347218 -2698 347454
rect -2614 347218 -2378 347454
rect -2934 346898 -2698 347134
rect -2614 346898 -2378 347134
rect -2934 320218 -2698 320454
rect -2614 320218 -2378 320454
rect -2934 319898 -2698 320134
rect -2614 319898 -2378 320134
rect -2934 293218 -2698 293454
rect -2614 293218 -2378 293454
rect -2934 292898 -2698 293134
rect -2614 292898 -2378 293134
rect -2934 266218 -2698 266454
rect -2614 266218 -2378 266454
rect -2934 265898 -2698 266134
rect -2614 265898 -2378 266134
rect -2934 239218 -2698 239454
rect -2614 239218 -2378 239454
rect -2934 238898 -2698 239134
rect -2614 238898 -2378 239134
rect -2934 212218 -2698 212454
rect -2614 212218 -2378 212454
rect -2934 211898 -2698 212134
rect -2614 211898 -2378 212134
rect -2934 185218 -2698 185454
rect -2614 185218 -2378 185454
rect -2934 184898 -2698 185134
rect -2614 184898 -2378 185134
rect -2934 158218 -2698 158454
rect -2614 158218 -2378 158454
rect -2934 157898 -2698 158134
rect -2614 157898 -2378 158134
rect -2934 131218 -2698 131454
rect -2614 131218 -2378 131454
rect -2934 130898 -2698 131134
rect -2614 130898 -2378 131134
rect -2934 104218 -2698 104454
rect -2614 104218 -2378 104454
rect -2934 103898 -2698 104134
rect -2614 103898 -2378 104134
rect -2934 77218 -2698 77454
rect -2614 77218 -2378 77454
rect -2934 76898 -2698 77134
rect -2614 76898 -2378 77134
rect -2934 50218 -2698 50454
rect -2614 50218 -2378 50454
rect -2934 49898 -2698 50134
rect -2614 49898 -2378 50134
rect -2934 23218 -2698 23454
rect -2614 23218 -2378 23454
rect -2934 22898 -2698 23134
rect -2614 22898 -2378 23134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 701593 -1738 701829
rect -1654 701593 -1418 701829
rect -1974 701273 -1738 701509
rect -1654 701273 -1418 701509
rect 38026 698218 38262 698454
rect 38346 698218 38582 698454
rect 38026 697898 38262 698134
rect 38346 697898 38582 698134
rect 41526 704602 41762 704838
rect 41846 704602 42082 704838
rect 41526 704282 41762 704518
rect 41846 704282 42082 704518
rect 41526 701593 41762 701829
rect 41846 701593 42082 701829
rect 41526 701273 41762 701509
rect 41846 701273 42082 701509
rect 66026 705562 66262 705798
rect 66346 705562 66582 705798
rect 66026 705242 66262 705478
rect 66346 705242 66582 705478
rect 66026 698218 66262 698454
rect 66346 698218 66582 698454
rect 66026 697898 66262 698134
rect 66346 697898 66582 698134
rect 69526 704602 69762 704838
rect 69846 704602 70082 704838
rect 69526 704282 69762 704518
rect 69846 704282 70082 704518
rect 69526 701593 69762 701829
rect 69846 701593 70082 701829
rect 69526 701273 69762 701509
rect 69846 701273 70082 701509
rect 94026 705562 94262 705798
rect 94346 705562 94582 705798
rect 94026 705242 94262 705478
rect 94346 705242 94582 705478
rect 94026 698218 94262 698454
rect 94346 698218 94582 698454
rect 94026 697898 94262 698134
rect 94346 697898 94582 698134
rect 97526 704602 97762 704838
rect 97846 704602 98082 704838
rect 97526 704282 97762 704518
rect 97846 704282 98082 704518
rect 97526 701593 97762 701829
rect 97846 701593 98082 701829
rect 97526 701273 97762 701509
rect 97846 701273 98082 701509
rect 122026 705562 122262 705798
rect 122346 705562 122582 705798
rect 122026 705242 122262 705478
rect 122346 705242 122582 705478
rect 122026 698218 122262 698454
rect 122346 698218 122582 698454
rect 122026 697898 122262 698134
rect 122346 697898 122582 698134
rect 125526 704602 125762 704838
rect 125846 704602 126082 704838
rect 125526 704282 125762 704518
rect 125846 704282 126082 704518
rect 125526 701593 125762 701829
rect 125846 701593 126082 701829
rect 125526 701273 125762 701509
rect 125846 701273 126082 701509
rect 150026 705562 150262 705798
rect 150346 705562 150582 705798
rect 150026 705242 150262 705478
rect 150346 705242 150582 705478
rect 150026 698218 150262 698454
rect 150346 698218 150582 698454
rect 150026 697898 150262 698134
rect 150346 697898 150582 698134
rect 153526 704602 153762 704838
rect 153846 704602 154082 704838
rect 153526 704282 153762 704518
rect 153846 704282 154082 704518
rect 153526 701593 153762 701829
rect 153846 701593 154082 701829
rect 153526 701273 153762 701509
rect 153846 701273 154082 701509
rect 178026 705562 178262 705798
rect 178346 705562 178582 705798
rect 178026 705242 178262 705478
rect 178346 705242 178582 705478
rect 178026 698218 178262 698454
rect 178346 698218 178582 698454
rect 178026 697898 178262 698134
rect 178346 697898 178582 698134
rect 181526 704602 181762 704838
rect 181846 704602 182082 704838
rect 181526 704282 181762 704518
rect 181846 704282 182082 704518
rect 181526 701593 181762 701829
rect 181846 701593 182082 701829
rect 181526 701273 181762 701509
rect 181846 701273 182082 701509
rect 206026 705562 206262 705798
rect 206346 705562 206582 705798
rect 206026 705242 206262 705478
rect 206346 705242 206582 705478
rect 206026 698218 206262 698454
rect 206346 698218 206582 698454
rect 206026 697898 206262 698134
rect 206346 697898 206582 698134
rect 209526 704602 209762 704838
rect 209846 704602 210082 704838
rect 209526 704282 209762 704518
rect 209846 704282 210082 704518
rect 209526 701593 209762 701829
rect 209846 701593 210082 701829
rect 209526 701273 209762 701509
rect 209846 701273 210082 701509
rect 234026 705562 234262 705798
rect 234346 705562 234582 705798
rect 234026 705242 234262 705478
rect 234346 705242 234582 705478
rect 234026 698218 234262 698454
rect 234346 698218 234582 698454
rect 234026 697898 234262 698134
rect 234346 697898 234582 698134
rect 237526 704602 237762 704838
rect 237846 704602 238082 704838
rect 237526 704282 237762 704518
rect 237846 704282 238082 704518
rect 237526 701593 237762 701829
rect 237846 701593 238082 701829
rect 237526 701273 237762 701509
rect 237846 701273 238082 701509
rect 262026 705562 262262 705798
rect 262346 705562 262582 705798
rect 262026 705242 262262 705478
rect 262346 705242 262582 705478
rect 262026 698218 262262 698454
rect 262346 698218 262582 698454
rect 262026 697898 262262 698134
rect 262346 697898 262582 698134
rect 265526 704602 265762 704838
rect 265846 704602 266082 704838
rect 265526 704282 265762 704518
rect 265846 704282 266082 704518
rect 265526 701593 265762 701829
rect 265846 701593 266082 701829
rect 265526 701273 265762 701509
rect 265846 701273 266082 701509
rect 290026 705562 290262 705798
rect 290346 705562 290582 705798
rect 290026 705242 290262 705478
rect 290346 705242 290582 705478
rect 290026 698218 290262 698454
rect 290346 698218 290582 698454
rect 290026 697898 290262 698134
rect 290346 697898 290582 698134
rect 293526 704602 293762 704838
rect 293846 704602 294082 704838
rect 293526 704282 293762 704518
rect 293846 704282 294082 704518
rect 293526 701593 293762 701829
rect 293846 701593 294082 701829
rect 293526 701273 293762 701509
rect 293846 701273 294082 701509
rect 318026 705562 318262 705798
rect 318346 705562 318582 705798
rect 318026 705242 318262 705478
rect 318346 705242 318582 705478
rect 318026 698218 318262 698454
rect 318346 698218 318582 698454
rect 318026 697898 318262 698134
rect 318346 697898 318582 698134
rect 321526 704602 321762 704838
rect 321846 704602 322082 704838
rect 321526 704282 321762 704518
rect 321846 704282 322082 704518
rect 321526 701593 321762 701829
rect 321846 701593 322082 701829
rect 321526 701273 321762 701509
rect 321846 701273 322082 701509
rect 346026 705562 346262 705798
rect 346346 705562 346582 705798
rect 346026 705242 346262 705478
rect 346346 705242 346582 705478
rect 346026 698218 346262 698454
rect 346346 698218 346582 698454
rect 346026 697898 346262 698134
rect 346346 697898 346582 698134
rect 349526 704602 349762 704838
rect 349846 704602 350082 704838
rect 349526 704282 349762 704518
rect 349846 704282 350082 704518
rect 349526 701593 349762 701829
rect 349846 701593 350082 701829
rect 349526 701273 349762 701509
rect 349846 701273 350082 701509
rect 374026 705562 374262 705798
rect 374346 705562 374582 705798
rect 374026 705242 374262 705478
rect 374346 705242 374582 705478
rect 374026 698218 374262 698454
rect 374346 698218 374582 698454
rect 374026 697898 374262 698134
rect 374346 697898 374582 698134
rect 377526 704602 377762 704838
rect 377846 704602 378082 704838
rect 377526 704282 377762 704518
rect 377846 704282 378082 704518
rect 377526 701593 377762 701829
rect 377846 701593 378082 701829
rect 377526 701273 377762 701509
rect 377846 701273 378082 701509
rect 402026 705562 402262 705798
rect 402346 705562 402582 705798
rect 402026 705242 402262 705478
rect 402346 705242 402582 705478
rect 402026 698218 402262 698454
rect 402346 698218 402582 698454
rect 402026 697898 402262 698134
rect 402346 697898 402582 698134
rect 405526 704602 405762 704838
rect 405846 704602 406082 704838
rect 405526 704282 405762 704518
rect 405846 704282 406082 704518
rect 405526 701593 405762 701829
rect 405846 701593 406082 701829
rect 405526 701273 405762 701509
rect 405846 701273 406082 701509
rect 430026 705562 430262 705798
rect 430346 705562 430582 705798
rect 430026 705242 430262 705478
rect 430346 705242 430582 705478
rect 430026 698218 430262 698454
rect 430346 698218 430582 698454
rect 430026 697898 430262 698134
rect 430346 697898 430582 698134
rect 433526 704602 433762 704838
rect 433846 704602 434082 704838
rect 433526 704282 433762 704518
rect 433846 704282 434082 704518
rect 433526 701593 433762 701829
rect 433846 701593 434082 701829
rect 433526 701273 433762 701509
rect 433846 701273 434082 701509
rect 458026 705562 458262 705798
rect 458346 705562 458582 705798
rect 458026 705242 458262 705478
rect 458346 705242 458582 705478
rect 458026 698218 458262 698454
rect 458346 698218 458582 698454
rect 458026 697898 458262 698134
rect 458346 697898 458582 698134
rect 461526 704602 461762 704838
rect 461846 704602 462082 704838
rect 461526 704282 461762 704518
rect 461846 704282 462082 704518
rect 461526 701593 461762 701829
rect 461846 701593 462082 701829
rect 461526 701273 461762 701509
rect 461846 701273 462082 701509
rect 486026 705562 486262 705798
rect 486346 705562 486582 705798
rect 486026 705242 486262 705478
rect 486346 705242 486582 705478
rect 486026 698218 486262 698454
rect 486346 698218 486582 698454
rect 486026 697898 486262 698134
rect 486346 697898 486582 698134
rect 489526 704602 489762 704838
rect 489846 704602 490082 704838
rect 489526 704282 489762 704518
rect 489846 704282 490082 704518
rect 489526 701593 489762 701829
rect 489846 701593 490082 701829
rect 489526 701273 489762 701509
rect 489846 701273 490082 701509
rect 514026 705562 514262 705798
rect 514346 705562 514582 705798
rect 514026 705242 514262 705478
rect 514346 705242 514582 705478
rect 514026 698218 514262 698454
rect 514346 698218 514582 698454
rect 514026 697898 514262 698134
rect 514346 697898 514582 698134
rect 517526 704602 517762 704838
rect 517846 704602 518082 704838
rect 517526 704282 517762 704518
rect 517846 704282 518082 704518
rect 517526 701593 517762 701829
rect 517846 701593 518082 701829
rect 517526 701273 517762 701509
rect 517846 701273 518082 701509
rect 542026 705562 542262 705798
rect 542346 705562 542582 705798
rect 542026 705242 542262 705478
rect 542346 705242 542582 705478
rect 542026 698218 542262 698454
rect 542346 698218 542582 698454
rect 542026 697898 542262 698134
rect 542346 697898 542582 698134
rect 545526 704602 545762 704838
rect 545846 704602 546082 704838
rect 545526 704282 545762 704518
rect 545846 704282 546082 704518
rect 545526 701593 545762 701829
rect 545846 701593 546082 701829
rect 545526 701273 545762 701509
rect 545846 701273 546082 701509
rect 570026 705562 570262 705798
rect 570346 705562 570582 705798
rect 570026 705242 570262 705478
rect 570346 705242 570582 705478
rect 570026 698218 570262 698454
rect 570346 698218 570582 698454
rect 570026 697898 570262 698134
rect 570346 697898 570582 698134
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 573526 704602 573762 704838
rect 573846 704602 574082 704838
rect 573526 704282 573762 704518
rect 573846 704282 574082 704518
rect 573526 701593 573762 701829
rect 573846 701593 574082 701829
rect 573526 701273 573762 701509
rect 573846 701273 574082 701509
rect -1974 674593 -1738 674829
rect -1654 674593 -1418 674829
rect -1974 674273 -1738 674509
rect -1654 674273 -1418 674509
rect 20118 674593 20354 674829
rect 20118 674273 20354 674509
rect 26382 674593 26618 674829
rect 26382 674273 26618 674509
rect 32646 674593 32882 674829
rect 32646 674273 32882 674509
rect 48118 674593 48354 674829
rect 48118 674273 48354 674509
rect 54382 674593 54618 674829
rect 54382 674273 54618 674509
rect 60646 674593 60882 674829
rect 60646 674273 60882 674509
rect 76118 674593 76354 674829
rect 76118 674273 76354 674509
rect 82382 674593 82618 674829
rect 82382 674273 82618 674509
rect 88646 674593 88882 674829
rect 88646 674273 88882 674509
rect 104118 674593 104354 674829
rect 104118 674273 104354 674509
rect 110382 674593 110618 674829
rect 110382 674273 110618 674509
rect 116646 674593 116882 674829
rect 116646 674273 116882 674509
rect 132118 674593 132354 674829
rect 132118 674273 132354 674509
rect 138382 674593 138618 674829
rect 138382 674273 138618 674509
rect 144646 674593 144882 674829
rect 144646 674273 144882 674509
rect 160118 674593 160354 674829
rect 160118 674273 160354 674509
rect 23250 671218 23486 671454
rect 23250 670898 23486 671134
rect 29514 671218 29750 671454
rect 29514 670898 29750 671134
rect 51250 671218 51486 671454
rect 51250 670898 51486 671134
rect 57514 671218 57750 671454
rect 57514 670898 57750 671134
rect 79250 671218 79486 671454
rect 79250 670898 79486 671134
rect 85514 671218 85750 671454
rect 85514 670898 85750 671134
rect 107250 671218 107486 671454
rect 107250 670898 107486 671134
rect 113514 671218 113750 671454
rect 113514 670898 113750 671134
rect 135250 671218 135486 671454
rect 135250 670898 135486 671134
rect 141514 671218 141750 671454
rect 141514 670898 141750 671134
rect 163250 671218 163486 671454
rect 163250 670898 163486 671134
rect 166382 674593 166618 674829
rect 166382 674273 166618 674509
rect 172646 674593 172882 674829
rect 172646 674273 172882 674509
rect 188118 674593 188354 674829
rect 188118 674273 188354 674509
rect 194382 674593 194618 674829
rect 194382 674273 194618 674509
rect 200646 674593 200882 674829
rect 200646 674273 200882 674509
rect 216118 674593 216354 674829
rect 216118 674273 216354 674509
rect 222382 674593 222618 674829
rect 222382 674273 222618 674509
rect 228646 674593 228882 674829
rect 228646 674273 228882 674509
rect 244118 674593 244354 674829
rect 244118 674273 244354 674509
rect 250382 674593 250618 674829
rect 250382 674273 250618 674509
rect 256646 674593 256882 674829
rect 256646 674273 256882 674509
rect 169514 671218 169750 671454
rect 169514 670898 169750 671134
rect 191250 671218 191486 671454
rect 191250 670898 191486 671134
rect 197514 671218 197750 671454
rect 197514 670898 197750 671134
rect 219250 671218 219486 671454
rect 219250 670898 219486 671134
rect 225514 671218 225750 671454
rect 225514 670898 225750 671134
rect 247250 671218 247486 671454
rect 247250 670898 247486 671134
rect 253514 671218 253750 671454
rect 253514 670898 253750 671134
rect 272118 674593 272354 674829
rect 272118 674273 272354 674509
rect 278382 674593 278618 674829
rect 278382 674273 278618 674509
rect 284646 674593 284882 674829
rect 284646 674273 284882 674509
rect 300118 674593 300354 674829
rect 300118 674273 300354 674509
rect 306382 674593 306618 674829
rect 306382 674273 306618 674509
rect 312646 674593 312882 674829
rect 312646 674273 312882 674509
rect 328118 674593 328354 674829
rect 328118 674273 328354 674509
rect 334382 674593 334618 674829
rect 334382 674273 334618 674509
rect 340646 674593 340882 674829
rect 340646 674273 340882 674509
rect 356118 674593 356354 674829
rect 356118 674273 356354 674509
rect 275250 671218 275486 671454
rect 275250 670898 275486 671134
rect 281514 671218 281750 671454
rect 281514 670898 281750 671134
rect 303250 671218 303486 671454
rect 303250 670898 303486 671134
rect 309514 671218 309750 671454
rect 309514 670898 309750 671134
rect 331250 671218 331486 671454
rect 331250 670898 331486 671134
rect 337514 671218 337750 671454
rect 337514 670898 337750 671134
rect 359250 671218 359486 671454
rect 359250 670898 359486 671134
rect 362382 674593 362618 674829
rect 362382 674273 362618 674509
rect 368646 674593 368882 674829
rect 368646 674273 368882 674509
rect 384118 674593 384354 674829
rect 384118 674273 384354 674509
rect 390382 674593 390618 674829
rect 390382 674273 390618 674509
rect 396646 674593 396882 674829
rect 396646 674273 396882 674509
rect 412118 674593 412354 674829
rect 412118 674273 412354 674509
rect 418382 674593 418618 674829
rect 418382 674273 418618 674509
rect 424646 674593 424882 674829
rect 424646 674273 424882 674509
rect 440118 674593 440354 674829
rect 440118 674273 440354 674509
rect 365514 671218 365750 671454
rect 365514 670898 365750 671134
rect 387250 671218 387486 671454
rect 387250 670898 387486 671134
rect 393514 671218 393750 671454
rect 393514 670898 393750 671134
rect 415250 671218 415486 671454
rect 415250 670898 415486 671134
rect 421514 671218 421750 671454
rect 421514 670898 421750 671134
rect 443250 671218 443486 671454
rect 443250 670898 443486 671134
rect 446382 674593 446618 674829
rect 446382 674273 446618 674509
rect 452646 674593 452882 674829
rect 452646 674273 452882 674509
rect 468118 674593 468354 674829
rect 468118 674273 468354 674509
rect 474382 674593 474618 674829
rect 474382 674273 474618 674509
rect 480646 674593 480882 674829
rect 480646 674273 480882 674509
rect 496118 674593 496354 674829
rect 496118 674273 496354 674509
rect 502382 674593 502618 674829
rect 502382 674273 502618 674509
rect 508646 674593 508882 674829
rect 508646 674273 508882 674509
rect 524118 674593 524354 674829
rect 524118 674273 524354 674509
rect 530382 674593 530618 674829
rect 530382 674273 530618 674509
rect 536646 674593 536882 674829
rect 536646 674273 536882 674509
rect 552118 674593 552354 674829
rect 552118 674273 552354 674509
rect 449514 671218 449750 671454
rect 449514 670898 449750 671134
rect 471250 671218 471486 671454
rect 471250 670898 471486 671134
rect 477514 671218 477750 671454
rect 477514 670898 477750 671134
rect 499250 671218 499486 671454
rect 499250 670898 499486 671134
rect 505514 671218 505750 671454
rect 505514 670898 505750 671134
rect 527250 671218 527486 671454
rect 527250 670898 527486 671134
rect 533514 671218 533750 671454
rect 533514 670898 533750 671134
rect 555250 671218 555486 671454
rect 555250 670898 555486 671134
rect 558382 674593 558618 674829
rect 558382 674273 558618 674509
rect 564646 674593 564882 674829
rect 564646 674273 564882 674509
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 701593 585578 701829
rect 585662 701593 585898 701829
rect 585342 701273 585578 701509
rect 585662 701273 585898 701509
rect 573526 674593 573762 674829
rect 573846 674593 574082 674829
rect 573526 674273 573762 674509
rect 573846 674273 574082 674509
rect 561514 671218 561750 671454
rect 561514 670898 561750 671134
rect -1974 647593 -1738 647829
rect -1654 647593 -1418 647829
rect -1974 647273 -1738 647509
rect -1654 647273 -1418 647509
rect 20118 647593 20354 647829
rect 20118 647273 20354 647509
rect 26382 647593 26618 647829
rect 26382 647273 26618 647509
rect 32646 647593 32882 647829
rect 32646 647273 32882 647509
rect 48118 647593 48354 647829
rect 48118 647273 48354 647509
rect 54382 647593 54618 647829
rect 54382 647273 54618 647509
rect 60646 647593 60882 647829
rect 60646 647273 60882 647509
rect 76118 647593 76354 647829
rect 76118 647273 76354 647509
rect 23250 644218 23486 644454
rect 23250 643898 23486 644134
rect 29514 644218 29750 644454
rect 29514 643898 29750 644134
rect 51250 644218 51486 644454
rect 51250 643898 51486 644134
rect 57514 644218 57750 644454
rect 57514 643898 57750 644134
rect 79250 644218 79486 644454
rect 79250 643898 79486 644134
rect 82382 647593 82618 647829
rect 82382 647273 82618 647509
rect 88646 647593 88882 647829
rect 88646 647273 88882 647509
rect 104118 647593 104354 647829
rect 104118 647273 104354 647509
rect 110382 647593 110618 647829
rect 110382 647273 110618 647509
rect 116646 647593 116882 647829
rect 116646 647273 116882 647509
rect 85514 644218 85750 644454
rect 85514 643898 85750 644134
rect 107250 644218 107486 644454
rect 107250 643898 107486 644134
rect 113514 644218 113750 644454
rect 113514 643898 113750 644134
rect 132118 647593 132354 647829
rect 132118 647273 132354 647509
rect 138382 647593 138618 647829
rect 138382 647273 138618 647509
rect 144646 647593 144882 647829
rect 144646 647273 144882 647509
rect 160118 647593 160354 647829
rect 160118 647273 160354 647509
rect 166382 647593 166618 647829
rect 166382 647273 166618 647509
rect 172646 647593 172882 647829
rect 172646 647273 172882 647509
rect 188118 647593 188354 647829
rect 188118 647273 188354 647509
rect 194382 647593 194618 647829
rect 194382 647273 194618 647509
rect 135250 644218 135486 644454
rect 135250 643898 135486 644134
rect 141514 644218 141750 644454
rect 141514 643898 141750 644134
rect 163250 644218 163486 644454
rect 163250 643898 163486 644134
rect 169514 644218 169750 644454
rect 169514 643898 169750 644134
rect 191250 644218 191486 644454
rect 191250 643898 191486 644134
rect 200646 647593 200882 647829
rect 200646 647273 200882 647509
rect 216118 647593 216354 647829
rect 216118 647273 216354 647509
rect 222382 647593 222618 647829
rect 222382 647273 222618 647509
rect 228646 647593 228882 647829
rect 228646 647273 228882 647509
rect 244118 647593 244354 647829
rect 244118 647273 244354 647509
rect 250382 647593 250618 647829
rect 250382 647273 250618 647509
rect 256646 647593 256882 647829
rect 256646 647273 256882 647509
rect 272118 647593 272354 647829
rect 272118 647273 272354 647509
rect 197514 644218 197750 644454
rect 197514 643898 197750 644134
rect 219250 644218 219486 644454
rect 219250 643898 219486 644134
rect 225514 644218 225750 644454
rect 225514 643898 225750 644134
rect 247250 644218 247486 644454
rect 247250 643898 247486 644134
rect 253514 644218 253750 644454
rect 253514 643898 253750 644134
rect 275250 644218 275486 644454
rect 275250 643898 275486 644134
rect 278382 647593 278618 647829
rect 278382 647273 278618 647509
rect 284646 647593 284882 647829
rect 284646 647273 284882 647509
rect 300118 647593 300354 647829
rect 300118 647273 300354 647509
rect 306382 647593 306618 647829
rect 306382 647273 306618 647509
rect 312646 647593 312882 647829
rect 312646 647273 312882 647509
rect 328118 647593 328354 647829
rect 328118 647273 328354 647509
rect 334382 647593 334618 647829
rect 334382 647273 334618 647509
rect 340646 647593 340882 647829
rect 340646 647273 340882 647509
rect 356118 647593 356354 647829
rect 356118 647273 356354 647509
rect 362382 647593 362618 647829
rect 362382 647273 362618 647509
rect 368646 647593 368882 647829
rect 368646 647273 368882 647509
rect 384118 647593 384354 647829
rect 384118 647273 384354 647509
rect 390382 647593 390618 647829
rect 390382 647273 390618 647509
rect 281514 644218 281750 644454
rect 281514 643898 281750 644134
rect 303250 644218 303486 644454
rect 303250 643898 303486 644134
rect 309514 644218 309750 644454
rect 309514 643898 309750 644134
rect 331250 644218 331486 644454
rect 331250 643898 331486 644134
rect 337514 644218 337750 644454
rect 337514 643898 337750 644134
rect 359250 644218 359486 644454
rect 359250 643898 359486 644134
rect 365514 644218 365750 644454
rect 365514 643898 365750 644134
rect 387250 644218 387486 644454
rect 387250 643898 387486 644134
rect 396646 647593 396882 647829
rect 396646 647273 396882 647509
rect 412118 647593 412354 647829
rect 412118 647273 412354 647509
rect 418382 647593 418618 647829
rect 418382 647273 418618 647509
rect 424646 647593 424882 647829
rect 424646 647273 424882 647509
rect 440118 647593 440354 647829
rect 440118 647273 440354 647509
rect 446382 647593 446618 647829
rect 446382 647273 446618 647509
rect 452646 647593 452882 647829
rect 452646 647273 452882 647509
rect 468118 647593 468354 647829
rect 468118 647273 468354 647509
rect 393514 644218 393750 644454
rect 393514 643898 393750 644134
rect 415250 644218 415486 644454
rect 415250 643898 415486 644134
rect 421514 644218 421750 644454
rect 421514 643898 421750 644134
rect 443250 644218 443486 644454
rect 443250 643898 443486 644134
rect 449514 644218 449750 644454
rect 449514 643898 449750 644134
rect 471250 644218 471486 644454
rect 471250 643898 471486 644134
rect 474382 647593 474618 647829
rect 474382 647273 474618 647509
rect 480646 647593 480882 647829
rect 480646 647273 480882 647509
rect 496118 647593 496354 647829
rect 496118 647273 496354 647509
rect 502382 647593 502618 647829
rect 502382 647273 502618 647509
rect 508646 647593 508882 647829
rect 508646 647273 508882 647509
rect 477514 644218 477750 644454
rect 477514 643898 477750 644134
rect 499250 644218 499486 644454
rect 499250 643898 499486 644134
rect 505514 644218 505750 644454
rect 505514 643898 505750 644134
rect 524118 647593 524354 647829
rect 524118 647273 524354 647509
rect 530382 647593 530618 647829
rect 530382 647273 530618 647509
rect 536646 647593 536882 647829
rect 536646 647273 536882 647509
rect 552118 647593 552354 647829
rect 552118 647273 552354 647509
rect 558382 647593 558618 647829
rect 558382 647273 558618 647509
rect 564646 647593 564882 647829
rect 564646 647273 564882 647509
rect 573526 647593 573762 647829
rect 573846 647593 574082 647829
rect 573526 647273 573762 647509
rect 573846 647273 574082 647509
rect 527250 644218 527486 644454
rect 527250 643898 527486 644134
rect 533514 644218 533750 644454
rect 533514 643898 533750 644134
rect 555250 644218 555486 644454
rect 555250 643898 555486 644134
rect 561514 644218 561750 644454
rect 561514 643898 561750 644134
rect -1974 620593 -1738 620829
rect -1654 620593 -1418 620829
rect -1974 620273 -1738 620509
rect -1654 620273 -1418 620509
rect 20118 620593 20354 620829
rect 20118 620273 20354 620509
rect 26382 620593 26618 620829
rect 26382 620273 26618 620509
rect 32646 620593 32882 620829
rect 32646 620273 32882 620509
rect 48118 620593 48354 620829
rect 48118 620273 48354 620509
rect 54382 620593 54618 620829
rect 54382 620273 54618 620509
rect 60646 620593 60882 620829
rect 60646 620273 60882 620509
rect 76118 620593 76354 620829
rect 76118 620273 76354 620509
rect 82382 620593 82618 620829
rect 82382 620273 82618 620509
rect 88646 620593 88882 620829
rect 88646 620273 88882 620509
rect 104118 620593 104354 620829
rect 104118 620273 104354 620509
rect 110382 620593 110618 620829
rect 110382 620273 110618 620509
rect 116646 620593 116882 620829
rect 116646 620273 116882 620509
rect 132118 620593 132354 620829
rect 132118 620273 132354 620509
rect 138382 620593 138618 620829
rect 138382 620273 138618 620509
rect 144646 620593 144882 620829
rect 144646 620273 144882 620509
rect 160118 620593 160354 620829
rect 160118 620273 160354 620509
rect 23250 617218 23486 617454
rect 23250 616898 23486 617134
rect 29514 617218 29750 617454
rect 29514 616898 29750 617134
rect 51250 617218 51486 617454
rect 51250 616898 51486 617134
rect 57514 617218 57750 617454
rect 57514 616898 57750 617134
rect 79250 617218 79486 617454
rect 79250 616898 79486 617134
rect 85514 617218 85750 617454
rect 85514 616898 85750 617134
rect 107250 617218 107486 617454
rect 107250 616898 107486 617134
rect 113514 617218 113750 617454
rect 113514 616898 113750 617134
rect 135250 617218 135486 617454
rect 135250 616898 135486 617134
rect 141514 617218 141750 617454
rect 141514 616898 141750 617134
rect 163250 617218 163486 617454
rect 163250 616898 163486 617134
rect 166382 620593 166618 620829
rect 166382 620273 166618 620509
rect 172646 620593 172882 620829
rect 172646 620273 172882 620509
rect 188118 620593 188354 620829
rect 188118 620273 188354 620509
rect 194382 620593 194618 620829
rect 194382 620273 194618 620509
rect 200646 620593 200882 620829
rect 200646 620273 200882 620509
rect 216118 620593 216354 620829
rect 216118 620273 216354 620509
rect 222382 620593 222618 620829
rect 222382 620273 222618 620509
rect 228646 620593 228882 620829
rect 228646 620273 228882 620509
rect 244118 620593 244354 620829
rect 244118 620273 244354 620509
rect 250382 620593 250618 620829
rect 250382 620273 250618 620509
rect 256646 620593 256882 620829
rect 256646 620273 256882 620509
rect 169514 617218 169750 617454
rect 169514 616898 169750 617134
rect 191250 617218 191486 617454
rect 191250 616898 191486 617134
rect 197514 617218 197750 617454
rect 197514 616898 197750 617134
rect 219250 617218 219486 617454
rect 219250 616898 219486 617134
rect 225514 617218 225750 617454
rect 225514 616898 225750 617134
rect 247250 617218 247486 617454
rect 247250 616898 247486 617134
rect 253514 617218 253750 617454
rect 253514 616898 253750 617134
rect 272118 620593 272354 620829
rect 272118 620273 272354 620509
rect 278382 620593 278618 620829
rect 278382 620273 278618 620509
rect 284646 620593 284882 620829
rect 284646 620273 284882 620509
rect 300118 620593 300354 620829
rect 300118 620273 300354 620509
rect 306382 620593 306618 620829
rect 306382 620273 306618 620509
rect 312646 620593 312882 620829
rect 312646 620273 312882 620509
rect 328118 620593 328354 620829
rect 328118 620273 328354 620509
rect 334382 620593 334618 620829
rect 334382 620273 334618 620509
rect 340646 620593 340882 620829
rect 340646 620273 340882 620509
rect 356118 620593 356354 620829
rect 356118 620273 356354 620509
rect 275250 617218 275486 617454
rect 275250 616898 275486 617134
rect 281514 617218 281750 617454
rect 281514 616898 281750 617134
rect 303250 617218 303486 617454
rect 303250 616898 303486 617134
rect 309514 617218 309750 617454
rect 309514 616898 309750 617134
rect 331250 617218 331486 617454
rect 331250 616898 331486 617134
rect 337514 617218 337750 617454
rect 337514 616898 337750 617134
rect 359250 617218 359486 617454
rect 359250 616898 359486 617134
rect 362382 620593 362618 620829
rect 362382 620273 362618 620509
rect 368646 620593 368882 620829
rect 368646 620273 368882 620509
rect 384118 620593 384354 620829
rect 384118 620273 384354 620509
rect 390382 620593 390618 620829
rect 390382 620273 390618 620509
rect 396646 620593 396882 620829
rect 396646 620273 396882 620509
rect 412118 620593 412354 620829
rect 412118 620273 412354 620509
rect 418382 620593 418618 620829
rect 418382 620273 418618 620509
rect 424646 620593 424882 620829
rect 424646 620273 424882 620509
rect 440118 620593 440354 620829
rect 440118 620273 440354 620509
rect 365514 617218 365750 617454
rect 365514 616898 365750 617134
rect 387250 617218 387486 617454
rect 387250 616898 387486 617134
rect 393514 617218 393750 617454
rect 393514 616898 393750 617134
rect 415250 617218 415486 617454
rect 415250 616898 415486 617134
rect 421514 617218 421750 617454
rect 421514 616898 421750 617134
rect 443250 617218 443486 617454
rect 443250 616898 443486 617134
rect 446382 620593 446618 620829
rect 446382 620273 446618 620509
rect 452646 620593 452882 620829
rect 452646 620273 452882 620509
rect 468118 620593 468354 620829
rect 468118 620273 468354 620509
rect 474382 620593 474618 620829
rect 474382 620273 474618 620509
rect 480646 620593 480882 620829
rect 480646 620273 480882 620509
rect 496118 620593 496354 620829
rect 496118 620273 496354 620509
rect 502382 620593 502618 620829
rect 502382 620273 502618 620509
rect 508646 620593 508882 620829
rect 508646 620273 508882 620509
rect 524118 620593 524354 620829
rect 524118 620273 524354 620509
rect 530382 620593 530618 620829
rect 530382 620273 530618 620509
rect 536646 620593 536882 620829
rect 536646 620273 536882 620509
rect 552118 620593 552354 620829
rect 552118 620273 552354 620509
rect 449514 617218 449750 617454
rect 449514 616898 449750 617134
rect 471250 617218 471486 617454
rect 471250 616898 471486 617134
rect 477514 617218 477750 617454
rect 477514 616898 477750 617134
rect 499250 617218 499486 617454
rect 499250 616898 499486 617134
rect 505514 617218 505750 617454
rect 505514 616898 505750 617134
rect 527250 617218 527486 617454
rect 527250 616898 527486 617134
rect 533514 617218 533750 617454
rect 533514 616898 533750 617134
rect 555250 617218 555486 617454
rect 555250 616898 555486 617134
rect 558382 620593 558618 620829
rect 558382 620273 558618 620509
rect 564646 620593 564882 620829
rect 564646 620273 564882 620509
rect 573526 620593 573762 620829
rect 573846 620593 574082 620829
rect 573526 620273 573762 620509
rect 573846 620273 574082 620509
rect 561514 617218 561750 617454
rect 561514 616898 561750 617134
rect -1974 593593 -1738 593829
rect -1654 593593 -1418 593829
rect -1974 593273 -1738 593509
rect -1654 593273 -1418 593509
rect 20118 593593 20354 593829
rect 20118 593273 20354 593509
rect 26382 593593 26618 593829
rect 26382 593273 26618 593509
rect 32646 593593 32882 593829
rect 32646 593273 32882 593509
rect 48118 593593 48354 593829
rect 48118 593273 48354 593509
rect 54382 593593 54618 593829
rect 54382 593273 54618 593509
rect 60646 593593 60882 593829
rect 60646 593273 60882 593509
rect 76118 593593 76354 593829
rect 76118 593273 76354 593509
rect 82382 593593 82618 593829
rect 82382 593273 82618 593509
rect 88646 593593 88882 593829
rect 88646 593273 88882 593509
rect 104118 593593 104354 593829
rect 104118 593273 104354 593509
rect 110382 593593 110618 593829
rect 110382 593273 110618 593509
rect 116646 593593 116882 593829
rect 116646 593273 116882 593509
rect 23250 590218 23486 590454
rect 23250 589898 23486 590134
rect 29514 590218 29750 590454
rect 29514 589898 29750 590134
rect 51250 590218 51486 590454
rect 51250 589898 51486 590134
rect 57514 590218 57750 590454
rect 57514 589898 57750 590134
rect 79250 590218 79486 590454
rect 79250 589898 79486 590134
rect 85514 590218 85750 590454
rect 85514 589898 85750 590134
rect 107250 590218 107486 590454
rect 107250 589898 107486 590134
rect 113514 590218 113750 590454
rect 113514 589898 113750 590134
rect 132118 593593 132354 593829
rect 132118 593273 132354 593509
rect 138382 593593 138618 593829
rect 138382 593273 138618 593509
rect 144646 593593 144882 593829
rect 144646 593273 144882 593509
rect 160118 593593 160354 593829
rect 160118 593273 160354 593509
rect 166382 593593 166618 593829
rect 166382 593273 166618 593509
rect 172646 593593 172882 593829
rect 172646 593273 172882 593509
rect 188118 593593 188354 593829
rect 188118 593273 188354 593509
rect 194382 593593 194618 593829
rect 194382 593273 194618 593509
rect 135250 590218 135486 590454
rect 135250 589898 135486 590134
rect 141514 590218 141750 590454
rect 141514 589898 141750 590134
rect 163250 590218 163486 590454
rect 163250 589898 163486 590134
rect 169514 590218 169750 590454
rect 169514 589898 169750 590134
rect 191250 590218 191486 590454
rect 191250 589898 191486 590134
rect 200646 593593 200882 593829
rect 200646 593273 200882 593509
rect 216118 593593 216354 593829
rect 216118 593273 216354 593509
rect 222382 593593 222618 593829
rect 222382 593273 222618 593509
rect 228646 593593 228882 593829
rect 228646 593273 228882 593509
rect 244118 593593 244354 593829
rect 244118 593273 244354 593509
rect 250382 593593 250618 593829
rect 250382 593273 250618 593509
rect 256646 593593 256882 593829
rect 256646 593273 256882 593509
rect 272118 593593 272354 593829
rect 272118 593273 272354 593509
rect 278382 593593 278618 593829
rect 278382 593273 278618 593509
rect 284646 593593 284882 593829
rect 284646 593273 284882 593509
rect 300118 593593 300354 593829
rect 300118 593273 300354 593509
rect 306382 593593 306618 593829
rect 306382 593273 306618 593509
rect 312646 593593 312882 593829
rect 312646 593273 312882 593509
rect 328118 593593 328354 593829
rect 328118 593273 328354 593509
rect 334382 593593 334618 593829
rect 334382 593273 334618 593509
rect 340646 593593 340882 593829
rect 340646 593273 340882 593509
rect 356118 593593 356354 593829
rect 356118 593273 356354 593509
rect 362382 593593 362618 593829
rect 362382 593273 362618 593509
rect 368646 593593 368882 593829
rect 368646 593273 368882 593509
rect 384118 593593 384354 593829
rect 384118 593273 384354 593509
rect 390382 593593 390618 593829
rect 390382 593273 390618 593509
rect 197514 590218 197750 590454
rect 197514 589898 197750 590134
rect 219250 590218 219486 590454
rect 219250 589898 219486 590134
rect 225514 590218 225750 590454
rect 225514 589898 225750 590134
rect 247250 590218 247486 590454
rect 247250 589898 247486 590134
rect 253514 590218 253750 590454
rect 253514 589898 253750 590134
rect 275250 590218 275486 590454
rect 275250 589898 275486 590134
rect 281514 590218 281750 590454
rect 281514 589898 281750 590134
rect 303250 590218 303486 590454
rect 303250 589898 303486 590134
rect 309514 590218 309750 590454
rect 309514 589898 309750 590134
rect 331250 590218 331486 590454
rect 331250 589898 331486 590134
rect 337514 590218 337750 590454
rect 337514 589898 337750 590134
rect 359250 590218 359486 590454
rect 359250 589898 359486 590134
rect 365514 590218 365750 590454
rect 365514 589898 365750 590134
rect 387250 590218 387486 590454
rect 387250 589898 387486 590134
rect 396646 593593 396882 593829
rect 396646 593273 396882 593509
rect 412118 593593 412354 593829
rect 412118 593273 412354 593509
rect 418382 593593 418618 593829
rect 418382 593273 418618 593509
rect 424646 593593 424882 593829
rect 424646 593273 424882 593509
rect 440118 593593 440354 593829
rect 440118 593273 440354 593509
rect 446382 593593 446618 593829
rect 446382 593273 446618 593509
rect 452646 593593 452882 593829
rect 452646 593273 452882 593509
rect 468118 593593 468354 593829
rect 468118 593273 468354 593509
rect 474382 593593 474618 593829
rect 474382 593273 474618 593509
rect 480646 593593 480882 593829
rect 480646 593273 480882 593509
rect 496118 593593 496354 593829
rect 496118 593273 496354 593509
rect 502382 593593 502618 593829
rect 502382 593273 502618 593509
rect 508646 593593 508882 593829
rect 508646 593273 508882 593509
rect 524118 593593 524354 593829
rect 524118 593273 524354 593509
rect 530382 593593 530618 593829
rect 530382 593273 530618 593509
rect 536646 593593 536882 593829
rect 536646 593273 536882 593509
rect 552118 593593 552354 593829
rect 552118 593273 552354 593509
rect 558382 593593 558618 593829
rect 558382 593273 558618 593509
rect 564646 593593 564882 593829
rect 564646 593273 564882 593509
rect 573526 593593 573762 593829
rect 573846 593593 574082 593829
rect 573526 593273 573762 593509
rect 573846 593273 574082 593509
rect 393514 590218 393750 590454
rect 393514 589898 393750 590134
rect 415250 590218 415486 590454
rect 415250 589898 415486 590134
rect 421514 590218 421750 590454
rect 421514 589898 421750 590134
rect 443250 590218 443486 590454
rect 443250 589898 443486 590134
rect 449514 590218 449750 590454
rect 449514 589898 449750 590134
rect 471250 590218 471486 590454
rect 471250 589898 471486 590134
rect 477514 590218 477750 590454
rect 477514 589898 477750 590134
rect 499250 590218 499486 590454
rect 499250 589898 499486 590134
rect 505514 590218 505750 590454
rect 505514 589898 505750 590134
rect 527250 590218 527486 590454
rect 527250 589898 527486 590134
rect 533514 590218 533750 590454
rect 533514 589898 533750 590134
rect 555250 590218 555486 590454
rect 555250 589898 555486 590134
rect 561514 590218 561750 590454
rect 561514 589898 561750 590134
rect -1974 566593 -1738 566829
rect -1654 566593 -1418 566829
rect -1974 566273 -1738 566509
rect -1654 566273 -1418 566509
rect 20118 566593 20354 566829
rect 20118 566273 20354 566509
rect 26382 566593 26618 566829
rect 26382 566273 26618 566509
rect 32646 566593 32882 566829
rect 32646 566273 32882 566509
rect 48118 566593 48354 566829
rect 48118 566273 48354 566509
rect 54382 566593 54618 566829
rect 54382 566273 54618 566509
rect 60646 566593 60882 566829
rect 60646 566273 60882 566509
rect 76118 566593 76354 566829
rect 76118 566273 76354 566509
rect 82382 566593 82618 566829
rect 82382 566273 82618 566509
rect 88646 566593 88882 566829
rect 88646 566273 88882 566509
rect 104118 566593 104354 566829
rect 104118 566273 104354 566509
rect 110382 566593 110618 566829
rect 110382 566273 110618 566509
rect 116646 566593 116882 566829
rect 116646 566273 116882 566509
rect 132118 566593 132354 566829
rect 132118 566273 132354 566509
rect 138382 566593 138618 566829
rect 138382 566273 138618 566509
rect 144646 566593 144882 566829
rect 144646 566273 144882 566509
rect 160118 566593 160354 566829
rect 160118 566273 160354 566509
rect 23250 563218 23486 563454
rect 23250 562898 23486 563134
rect 29514 563218 29750 563454
rect 29514 562898 29750 563134
rect 51250 563218 51486 563454
rect 51250 562898 51486 563134
rect 57514 563218 57750 563454
rect 57514 562898 57750 563134
rect 79250 563218 79486 563454
rect 79250 562898 79486 563134
rect 85514 563218 85750 563454
rect 85514 562898 85750 563134
rect 107250 563218 107486 563454
rect 107250 562898 107486 563134
rect 113514 563218 113750 563454
rect 113514 562898 113750 563134
rect 135250 563218 135486 563454
rect 135250 562898 135486 563134
rect 141514 563218 141750 563454
rect 141514 562898 141750 563134
rect 163250 563218 163486 563454
rect 163250 562898 163486 563134
rect 166382 566593 166618 566829
rect 166382 566273 166618 566509
rect 172646 566593 172882 566829
rect 172646 566273 172882 566509
rect 188118 566593 188354 566829
rect 188118 566273 188354 566509
rect 194382 566593 194618 566829
rect 194382 566273 194618 566509
rect 200646 566593 200882 566829
rect 200646 566273 200882 566509
rect 216118 566593 216354 566829
rect 216118 566273 216354 566509
rect 222382 566593 222618 566829
rect 222382 566273 222618 566509
rect 228646 566593 228882 566829
rect 228646 566273 228882 566509
rect 244118 566593 244354 566829
rect 244118 566273 244354 566509
rect 250382 566593 250618 566829
rect 250382 566273 250618 566509
rect 256646 566593 256882 566829
rect 256646 566273 256882 566509
rect 169514 563218 169750 563454
rect 169514 562898 169750 563134
rect 191250 563218 191486 563454
rect 191250 562898 191486 563134
rect 197514 563218 197750 563454
rect 197514 562898 197750 563134
rect 219250 563218 219486 563454
rect 219250 562898 219486 563134
rect 225514 563218 225750 563454
rect 225514 562898 225750 563134
rect 247250 563218 247486 563454
rect 247250 562898 247486 563134
rect 253514 563218 253750 563454
rect 253514 562898 253750 563134
rect 272118 566593 272354 566829
rect 272118 566273 272354 566509
rect 278382 566593 278618 566829
rect 278382 566273 278618 566509
rect 284646 566593 284882 566829
rect 284646 566273 284882 566509
rect 300118 566593 300354 566829
rect 300118 566273 300354 566509
rect 306382 566593 306618 566829
rect 306382 566273 306618 566509
rect 312646 566593 312882 566829
rect 312646 566273 312882 566509
rect 328118 566593 328354 566829
rect 328118 566273 328354 566509
rect 334382 566593 334618 566829
rect 334382 566273 334618 566509
rect 340646 566593 340882 566829
rect 340646 566273 340882 566509
rect 356118 566593 356354 566829
rect 356118 566273 356354 566509
rect 275250 563218 275486 563454
rect 275250 562898 275486 563134
rect 281514 563218 281750 563454
rect 281514 562898 281750 563134
rect 303250 563218 303486 563454
rect 303250 562898 303486 563134
rect 309514 563218 309750 563454
rect 309514 562898 309750 563134
rect 331250 563218 331486 563454
rect 331250 562898 331486 563134
rect 337514 563218 337750 563454
rect 337514 562898 337750 563134
rect 359250 563218 359486 563454
rect 359250 562898 359486 563134
rect 362382 566593 362618 566829
rect 362382 566273 362618 566509
rect 368646 566593 368882 566829
rect 368646 566273 368882 566509
rect 384118 566593 384354 566829
rect 384118 566273 384354 566509
rect 390382 566593 390618 566829
rect 390382 566273 390618 566509
rect 396646 566593 396882 566829
rect 396646 566273 396882 566509
rect 412118 566593 412354 566829
rect 412118 566273 412354 566509
rect 418382 566593 418618 566829
rect 418382 566273 418618 566509
rect 424646 566593 424882 566829
rect 424646 566273 424882 566509
rect 440118 566593 440354 566829
rect 440118 566273 440354 566509
rect 365514 563218 365750 563454
rect 365514 562898 365750 563134
rect 387250 563218 387486 563454
rect 387250 562898 387486 563134
rect 393514 563218 393750 563454
rect 393514 562898 393750 563134
rect 415250 563218 415486 563454
rect 415250 562898 415486 563134
rect 421514 563218 421750 563454
rect 421514 562898 421750 563134
rect 443250 563218 443486 563454
rect 443250 562898 443486 563134
rect 446382 566593 446618 566829
rect 446382 566273 446618 566509
rect 452646 566593 452882 566829
rect 452646 566273 452882 566509
rect 468118 566593 468354 566829
rect 468118 566273 468354 566509
rect 474382 566593 474618 566829
rect 474382 566273 474618 566509
rect 480646 566593 480882 566829
rect 480646 566273 480882 566509
rect 496118 566593 496354 566829
rect 496118 566273 496354 566509
rect 502382 566593 502618 566829
rect 502382 566273 502618 566509
rect 508646 566593 508882 566829
rect 508646 566273 508882 566509
rect 524118 566593 524354 566829
rect 524118 566273 524354 566509
rect 530382 566593 530618 566829
rect 530382 566273 530618 566509
rect 536646 566593 536882 566829
rect 536646 566273 536882 566509
rect 552118 566593 552354 566829
rect 552118 566273 552354 566509
rect 449514 563218 449750 563454
rect 449514 562898 449750 563134
rect 471250 563218 471486 563454
rect 471250 562898 471486 563134
rect 477514 563218 477750 563454
rect 477514 562898 477750 563134
rect 499250 563218 499486 563454
rect 499250 562898 499486 563134
rect 505514 563218 505750 563454
rect 505514 562898 505750 563134
rect 527250 563218 527486 563454
rect 527250 562898 527486 563134
rect 533514 563218 533750 563454
rect 533514 562898 533750 563134
rect 555250 563218 555486 563454
rect 555250 562898 555486 563134
rect 558382 566593 558618 566829
rect 558382 566273 558618 566509
rect 564646 566593 564882 566829
rect 564646 566273 564882 566509
rect 573526 566593 573762 566829
rect 573846 566593 574082 566829
rect 573526 566273 573762 566509
rect 573846 566273 574082 566509
rect 561514 563218 561750 563454
rect 561514 562898 561750 563134
rect -1974 539593 -1738 539829
rect -1654 539593 -1418 539829
rect -1974 539273 -1738 539509
rect -1654 539273 -1418 539509
rect 20118 539593 20354 539829
rect 20118 539273 20354 539509
rect 26382 539593 26618 539829
rect 26382 539273 26618 539509
rect 32646 539593 32882 539829
rect 32646 539273 32882 539509
rect 48118 539593 48354 539829
rect 48118 539273 48354 539509
rect 54382 539593 54618 539829
rect 54382 539273 54618 539509
rect 60646 539593 60882 539829
rect 60646 539273 60882 539509
rect 76118 539593 76354 539829
rect 76118 539273 76354 539509
rect 82382 539593 82618 539829
rect 82382 539273 82618 539509
rect 88646 539593 88882 539829
rect 88646 539273 88882 539509
rect 104118 539593 104354 539829
rect 104118 539273 104354 539509
rect 110382 539593 110618 539829
rect 110382 539273 110618 539509
rect 116646 539593 116882 539829
rect 116646 539273 116882 539509
rect 23250 536218 23486 536454
rect 23250 535898 23486 536134
rect 29514 536218 29750 536454
rect 29514 535898 29750 536134
rect 51250 536218 51486 536454
rect 51250 535898 51486 536134
rect 57514 536218 57750 536454
rect 57514 535898 57750 536134
rect 79250 536218 79486 536454
rect 79250 535898 79486 536134
rect 85514 536218 85750 536454
rect 85514 535898 85750 536134
rect 107250 536218 107486 536454
rect 107250 535898 107486 536134
rect 113514 536218 113750 536454
rect 113514 535898 113750 536134
rect 132118 539593 132354 539829
rect 132118 539273 132354 539509
rect 138382 539593 138618 539829
rect 138382 539273 138618 539509
rect 144646 539593 144882 539829
rect 144646 539273 144882 539509
rect 160118 539593 160354 539829
rect 160118 539273 160354 539509
rect 166382 539593 166618 539829
rect 166382 539273 166618 539509
rect 172646 539593 172882 539829
rect 172646 539273 172882 539509
rect 188118 539593 188354 539829
rect 188118 539273 188354 539509
rect 194382 539593 194618 539829
rect 194382 539273 194618 539509
rect 135250 536218 135486 536454
rect 135250 535898 135486 536134
rect 141514 536218 141750 536454
rect 141514 535898 141750 536134
rect 163250 536218 163486 536454
rect 163250 535898 163486 536134
rect 169514 536218 169750 536454
rect 169514 535898 169750 536134
rect 191250 536218 191486 536454
rect 191250 535898 191486 536134
rect 200646 539593 200882 539829
rect 200646 539273 200882 539509
rect 216118 539593 216354 539829
rect 216118 539273 216354 539509
rect 222382 539593 222618 539829
rect 222382 539273 222618 539509
rect 228646 539593 228882 539829
rect 228646 539273 228882 539509
rect 244118 539593 244354 539829
rect 244118 539273 244354 539509
rect 250382 539593 250618 539829
rect 250382 539273 250618 539509
rect 256646 539593 256882 539829
rect 256646 539273 256882 539509
rect 272118 539593 272354 539829
rect 272118 539273 272354 539509
rect 278382 539593 278618 539829
rect 278382 539273 278618 539509
rect 284646 539593 284882 539829
rect 284646 539273 284882 539509
rect 300118 539593 300354 539829
rect 300118 539273 300354 539509
rect 306382 539593 306618 539829
rect 306382 539273 306618 539509
rect 312646 539593 312882 539829
rect 312646 539273 312882 539509
rect 328118 539593 328354 539829
rect 328118 539273 328354 539509
rect 334382 539593 334618 539829
rect 334382 539273 334618 539509
rect 340646 539593 340882 539829
rect 340646 539273 340882 539509
rect 356118 539593 356354 539829
rect 356118 539273 356354 539509
rect 362382 539593 362618 539829
rect 362382 539273 362618 539509
rect 368646 539593 368882 539829
rect 368646 539273 368882 539509
rect 384118 539593 384354 539829
rect 384118 539273 384354 539509
rect 390382 539593 390618 539829
rect 390382 539273 390618 539509
rect 197514 536218 197750 536454
rect 197514 535898 197750 536134
rect 219250 536218 219486 536454
rect 219250 535898 219486 536134
rect 225514 536218 225750 536454
rect 225514 535898 225750 536134
rect 247250 536218 247486 536454
rect 247250 535898 247486 536134
rect 253514 536218 253750 536454
rect 253514 535898 253750 536134
rect 275250 536218 275486 536454
rect 275250 535898 275486 536134
rect 281514 536218 281750 536454
rect 281514 535898 281750 536134
rect 303250 536218 303486 536454
rect 303250 535898 303486 536134
rect 309514 536218 309750 536454
rect 309514 535898 309750 536134
rect 331250 536218 331486 536454
rect 331250 535898 331486 536134
rect 337514 536218 337750 536454
rect 337514 535898 337750 536134
rect 359250 536218 359486 536454
rect 359250 535898 359486 536134
rect 365514 536218 365750 536454
rect 365514 535898 365750 536134
rect 387250 536218 387486 536454
rect 387250 535898 387486 536134
rect 396646 539593 396882 539829
rect 396646 539273 396882 539509
rect 412118 539593 412354 539829
rect 412118 539273 412354 539509
rect 418382 539593 418618 539829
rect 418382 539273 418618 539509
rect 424646 539593 424882 539829
rect 424646 539273 424882 539509
rect 440118 539593 440354 539829
rect 440118 539273 440354 539509
rect 446382 539593 446618 539829
rect 446382 539273 446618 539509
rect 452646 539593 452882 539829
rect 452646 539273 452882 539509
rect 468118 539593 468354 539829
rect 468118 539273 468354 539509
rect 474382 539593 474618 539829
rect 474382 539273 474618 539509
rect 480646 539593 480882 539829
rect 480646 539273 480882 539509
rect 496118 539593 496354 539829
rect 496118 539273 496354 539509
rect 502382 539593 502618 539829
rect 502382 539273 502618 539509
rect 508646 539593 508882 539829
rect 508646 539273 508882 539509
rect 524118 539593 524354 539829
rect 524118 539273 524354 539509
rect 530382 539593 530618 539829
rect 530382 539273 530618 539509
rect 536646 539593 536882 539829
rect 536646 539273 536882 539509
rect 552118 539593 552354 539829
rect 552118 539273 552354 539509
rect 558382 539593 558618 539829
rect 558382 539273 558618 539509
rect 564646 539593 564882 539829
rect 564646 539273 564882 539509
rect 573526 539593 573762 539829
rect 573846 539593 574082 539829
rect 573526 539273 573762 539509
rect 573846 539273 574082 539509
rect 393514 536218 393750 536454
rect 393514 535898 393750 536134
rect 415250 536218 415486 536454
rect 415250 535898 415486 536134
rect 421514 536218 421750 536454
rect 421514 535898 421750 536134
rect 443250 536218 443486 536454
rect 443250 535898 443486 536134
rect 449514 536218 449750 536454
rect 449514 535898 449750 536134
rect 471250 536218 471486 536454
rect 471250 535898 471486 536134
rect 477514 536218 477750 536454
rect 477514 535898 477750 536134
rect 499250 536218 499486 536454
rect 499250 535898 499486 536134
rect 505514 536218 505750 536454
rect 505514 535898 505750 536134
rect 527250 536218 527486 536454
rect 527250 535898 527486 536134
rect 533514 536218 533750 536454
rect 533514 535898 533750 536134
rect 555250 536218 555486 536454
rect 555250 535898 555486 536134
rect 561514 536218 561750 536454
rect 561514 535898 561750 536134
rect -1974 512593 -1738 512829
rect -1654 512593 -1418 512829
rect -1974 512273 -1738 512509
rect -1654 512273 -1418 512509
rect 20118 512593 20354 512829
rect 20118 512273 20354 512509
rect 26382 512593 26618 512829
rect 26382 512273 26618 512509
rect 32646 512593 32882 512829
rect 32646 512273 32882 512509
rect 48118 512593 48354 512829
rect 48118 512273 48354 512509
rect 54382 512593 54618 512829
rect 54382 512273 54618 512509
rect 60646 512593 60882 512829
rect 60646 512273 60882 512509
rect 76118 512593 76354 512829
rect 76118 512273 76354 512509
rect 82382 512593 82618 512829
rect 82382 512273 82618 512509
rect 88646 512593 88882 512829
rect 88646 512273 88882 512509
rect 104118 512593 104354 512829
rect 104118 512273 104354 512509
rect 110382 512593 110618 512829
rect 110382 512273 110618 512509
rect 116646 512593 116882 512829
rect 116646 512273 116882 512509
rect 132118 512593 132354 512829
rect 132118 512273 132354 512509
rect 138382 512593 138618 512829
rect 138382 512273 138618 512509
rect 144646 512593 144882 512829
rect 144646 512273 144882 512509
rect 160118 512593 160354 512829
rect 160118 512273 160354 512509
rect 23250 509218 23486 509454
rect 23250 508898 23486 509134
rect 29514 509218 29750 509454
rect 29514 508898 29750 509134
rect 51250 509218 51486 509454
rect 51250 508898 51486 509134
rect 57514 509218 57750 509454
rect 57514 508898 57750 509134
rect 79250 509218 79486 509454
rect 79250 508898 79486 509134
rect 85514 509218 85750 509454
rect 85514 508898 85750 509134
rect 107250 509218 107486 509454
rect 107250 508898 107486 509134
rect 113514 509218 113750 509454
rect 113514 508898 113750 509134
rect 135250 509218 135486 509454
rect 135250 508898 135486 509134
rect 141514 509218 141750 509454
rect 141514 508898 141750 509134
rect 163250 509218 163486 509454
rect 163250 508898 163486 509134
rect 166382 512593 166618 512829
rect 166382 512273 166618 512509
rect 172646 512593 172882 512829
rect 172646 512273 172882 512509
rect 188118 512593 188354 512829
rect 188118 512273 188354 512509
rect 194382 512593 194618 512829
rect 194382 512273 194618 512509
rect 200646 512593 200882 512829
rect 200646 512273 200882 512509
rect 216118 512593 216354 512829
rect 216118 512273 216354 512509
rect 222382 512593 222618 512829
rect 222382 512273 222618 512509
rect 228646 512593 228882 512829
rect 228646 512273 228882 512509
rect 244118 512593 244354 512829
rect 244118 512273 244354 512509
rect 250382 512593 250618 512829
rect 250382 512273 250618 512509
rect 256646 512593 256882 512829
rect 256646 512273 256882 512509
rect 169514 509218 169750 509454
rect 169514 508898 169750 509134
rect 191250 509218 191486 509454
rect 191250 508898 191486 509134
rect 197514 509218 197750 509454
rect 197514 508898 197750 509134
rect 219250 509218 219486 509454
rect 219250 508898 219486 509134
rect 225514 509218 225750 509454
rect 225514 508898 225750 509134
rect 247250 509218 247486 509454
rect 247250 508898 247486 509134
rect 253514 509218 253750 509454
rect 253514 508898 253750 509134
rect 272118 512593 272354 512829
rect 272118 512273 272354 512509
rect 278382 512593 278618 512829
rect 278382 512273 278618 512509
rect 284646 512593 284882 512829
rect 284646 512273 284882 512509
rect 300118 512593 300354 512829
rect 300118 512273 300354 512509
rect 306382 512593 306618 512829
rect 306382 512273 306618 512509
rect 312646 512593 312882 512829
rect 312646 512273 312882 512509
rect 328118 512593 328354 512829
rect 328118 512273 328354 512509
rect 334382 512593 334618 512829
rect 334382 512273 334618 512509
rect 340646 512593 340882 512829
rect 340646 512273 340882 512509
rect 356118 512593 356354 512829
rect 356118 512273 356354 512509
rect 275250 509218 275486 509454
rect 275250 508898 275486 509134
rect 281514 509218 281750 509454
rect 281514 508898 281750 509134
rect 303250 509218 303486 509454
rect 303250 508898 303486 509134
rect 309514 509218 309750 509454
rect 309514 508898 309750 509134
rect 331250 509218 331486 509454
rect 331250 508898 331486 509134
rect 337514 509218 337750 509454
rect 337514 508898 337750 509134
rect 359250 509218 359486 509454
rect 359250 508898 359486 509134
rect 362382 512593 362618 512829
rect 362382 512273 362618 512509
rect 368646 512593 368882 512829
rect 368646 512273 368882 512509
rect 384118 512593 384354 512829
rect 384118 512273 384354 512509
rect 390382 512593 390618 512829
rect 390382 512273 390618 512509
rect 396646 512593 396882 512829
rect 396646 512273 396882 512509
rect 412118 512593 412354 512829
rect 412118 512273 412354 512509
rect 418382 512593 418618 512829
rect 418382 512273 418618 512509
rect 424646 512593 424882 512829
rect 424646 512273 424882 512509
rect 440118 512593 440354 512829
rect 440118 512273 440354 512509
rect 365514 509218 365750 509454
rect 365514 508898 365750 509134
rect 387250 509218 387486 509454
rect 387250 508898 387486 509134
rect 393514 509218 393750 509454
rect 393514 508898 393750 509134
rect 415250 509218 415486 509454
rect 415250 508898 415486 509134
rect 421514 509218 421750 509454
rect 421514 508898 421750 509134
rect 443250 509218 443486 509454
rect 443250 508898 443486 509134
rect 446382 512593 446618 512829
rect 446382 512273 446618 512509
rect 452646 512593 452882 512829
rect 452646 512273 452882 512509
rect 468118 512593 468354 512829
rect 468118 512273 468354 512509
rect 474382 512593 474618 512829
rect 474382 512273 474618 512509
rect 480646 512593 480882 512829
rect 480646 512273 480882 512509
rect 496118 512593 496354 512829
rect 496118 512273 496354 512509
rect 502382 512593 502618 512829
rect 502382 512273 502618 512509
rect 508646 512593 508882 512829
rect 508646 512273 508882 512509
rect 524118 512593 524354 512829
rect 524118 512273 524354 512509
rect 530382 512593 530618 512829
rect 530382 512273 530618 512509
rect 536646 512593 536882 512829
rect 536646 512273 536882 512509
rect 552118 512593 552354 512829
rect 552118 512273 552354 512509
rect 449514 509218 449750 509454
rect 449514 508898 449750 509134
rect 471250 509218 471486 509454
rect 471250 508898 471486 509134
rect 477514 509218 477750 509454
rect 477514 508898 477750 509134
rect 499250 509218 499486 509454
rect 499250 508898 499486 509134
rect 505514 509218 505750 509454
rect 505514 508898 505750 509134
rect 527250 509218 527486 509454
rect 527250 508898 527486 509134
rect 533514 509218 533750 509454
rect 533514 508898 533750 509134
rect 555250 509218 555486 509454
rect 555250 508898 555486 509134
rect 558382 512593 558618 512829
rect 558382 512273 558618 512509
rect 564646 512593 564882 512829
rect 564646 512273 564882 512509
rect 573526 512593 573762 512829
rect 573846 512593 574082 512829
rect 573526 512273 573762 512509
rect 573846 512273 574082 512509
rect 561514 509218 561750 509454
rect 561514 508898 561750 509134
rect -1974 485593 -1738 485829
rect -1654 485593 -1418 485829
rect -1974 485273 -1738 485509
rect -1654 485273 -1418 485509
rect 20118 485593 20354 485829
rect 20118 485273 20354 485509
rect 26382 485593 26618 485829
rect 26382 485273 26618 485509
rect 32646 485593 32882 485829
rect 32646 485273 32882 485509
rect 48118 485593 48354 485829
rect 48118 485273 48354 485509
rect 54382 485593 54618 485829
rect 54382 485273 54618 485509
rect 60646 485593 60882 485829
rect 60646 485273 60882 485509
rect 76118 485593 76354 485829
rect 76118 485273 76354 485509
rect 82382 485593 82618 485829
rect 82382 485273 82618 485509
rect 88646 485593 88882 485829
rect 88646 485273 88882 485509
rect 104118 485593 104354 485829
rect 104118 485273 104354 485509
rect 110382 485593 110618 485829
rect 110382 485273 110618 485509
rect 116646 485593 116882 485829
rect 116646 485273 116882 485509
rect 23250 482218 23486 482454
rect 23250 481898 23486 482134
rect 29514 482218 29750 482454
rect 29514 481898 29750 482134
rect 51250 482218 51486 482454
rect 51250 481898 51486 482134
rect 57514 482218 57750 482454
rect 57514 481898 57750 482134
rect 79250 482218 79486 482454
rect 79250 481898 79486 482134
rect 85514 482218 85750 482454
rect 85514 481898 85750 482134
rect 107250 482218 107486 482454
rect 107250 481898 107486 482134
rect 113514 482218 113750 482454
rect 113514 481898 113750 482134
rect 132118 485593 132354 485829
rect 132118 485273 132354 485509
rect 138382 485593 138618 485829
rect 138382 485273 138618 485509
rect 144646 485593 144882 485829
rect 144646 485273 144882 485509
rect 160118 485593 160354 485829
rect 160118 485273 160354 485509
rect 166382 485593 166618 485829
rect 166382 485273 166618 485509
rect 172646 485593 172882 485829
rect 172646 485273 172882 485509
rect 188118 485593 188354 485829
rect 188118 485273 188354 485509
rect 194382 485593 194618 485829
rect 194382 485273 194618 485509
rect 135250 482218 135486 482454
rect 135250 481898 135486 482134
rect 141514 482218 141750 482454
rect 141514 481898 141750 482134
rect 163250 482218 163486 482454
rect 163250 481898 163486 482134
rect 169514 482218 169750 482454
rect 169514 481898 169750 482134
rect 191250 482218 191486 482454
rect 191250 481898 191486 482134
rect 200646 485593 200882 485829
rect 200646 485273 200882 485509
rect 216118 485593 216354 485829
rect 216118 485273 216354 485509
rect 222382 485593 222618 485829
rect 222382 485273 222618 485509
rect 228646 485593 228882 485829
rect 228646 485273 228882 485509
rect 244118 485593 244354 485829
rect 244118 485273 244354 485509
rect 250382 485593 250618 485829
rect 250382 485273 250618 485509
rect 256646 485593 256882 485829
rect 256646 485273 256882 485509
rect 272118 485593 272354 485829
rect 272118 485273 272354 485509
rect 278382 485593 278618 485829
rect 278382 485273 278618 485509
rect 284646 485593 284882 485829
rect 284646 485273 284882 485509
rect 300118 485593 300354 485829
rect 300118 485273 300354 485509
rect 306382 485593 306618 485829
rect 306382 485273 306618 485509
rect 312646 485593 312882 485829
rect 312646 485273 312882 485509
rect 328118 485593 328354 485829
rect 328118 485273 328354 485509
rect 334382 485593 334618 485829
rect 334382 485273 334618 485509
rect 340646 485593 340882 485829
rect 340646 485273 340882 485509
rect 356118 485593 356354 485829
rect 356118 485273 356354 485509
rect 362382 485593 362618 485829
rect 362382 485273 362618 485509
rect 368646 485593 368882 485829
rect 368646 485273 368882 485509
rect 384118 485593 384354 485829
rect 384118 485273 384354 485509
rect 390382 485593 390618 485829
rect 390382 485273 390618 485509
rect 197514 482218 197750 482454
rect 197514 481898 197750 482134
rect 219250 482218 219486 482454
rect 219250 481898 219486 482134
rect 225514 482218 225750 482454
rect 225514 481898 225750 482134
rect 247250 482218 247486 482454
rect 247250 481898 247486 482134
rect 253514 482218 253750 482454
rect 253514 481898 253750 482134
rect 275250 482218 275486 482454
rect 275250 481898 275486 482134
rect 281514 482218 281750 482454
rect 281514 481898 281750 482134
rect 303250 482218 303486 482454
rect 303250 481898 303486 482134
rect 309514 482218 309750 482454
rect 309514 481898 309750 482134
rect 331250 482218 331486 482454
rect 331250 481898 331486 482134
rect 337514 482218 337750 482454
rect 337514 481898 337750 482134
rect 359250 482218 359486 482454
rect 359250 481898 359486 482134
rect 365514 482218 365750 482454
rect 365514 481898 365750 482134
rect 387250 482218 387486 482454
rect 387250 481898 387486 482134
rect 396646 485593 396882 485829
rect 396646 485273 396882 485509
rect 412118 485593 412354 485829
rect 412118 485273 412354 485509
rect 418382 485593 418618 485829
rect 418382 485273 418618 485509
rect 424646 485593 424882 485829
rect 424646 485273 424882 485509
rect 440118 485593 440354 485829
rect 440118 485273 440354 485509
rect 446382 485593 446618 485829
rect 446382 485273 446618 485509
rect 452646 485593 452882 485829
rect 452646 485273 452882 485509
rect 468118 485593 468354 485829
rect 468118 485273 468354 485509
rect 474382 485593 474618 485829
rect 474382 485273 474618 485509
rect 480646 485593 480882 485829
rect 480646 485273 480882 485509
rect 496118 485593 496354 485829
rect 496118 485273 496354 485509
rect 502382 485593 502618 485829
rect 502382 485273 502618 485509
rect 508646 485593 508882 485829
rect 508646 485273 508882 485509
rect 524118 485593 524354 485829
rect 524118 485273 524354 485509
rect 530382 485593 530618 485829
rect 530382 485273 530618 485509
rect 536646 485593 536882 485829
rect 536646 485273 536882 485509
rect 552118 485593 552354 485829
rect 552118 485273 552354 485509
rect 558382 485593 558618 485829
rect 558382 485273 558618 485509
rect 564646 485593 564882 485829
rect 564646 485273 564882 485509
rect 573526 485593 573762 485829
rect 573846 485593 574082 485829
rect 573526 485273 573762 485509
rect 573846 485273 574082 485509
rect 393514 482218 393750 482454
rect 393514 481898 393750 482134
rect 415250 482218 415486 482454
rect 415250 481898 415486 482134
rect 421514 482218 421750 482454
rect 421514 481898 421750 482134
rect 443250 482218 443486 482454
rect 443250 481898 443486 482134
rect 449514 482218 449750 482454
rect 449514 481898 449750 482134
rect 471250 482218 471486 482454
rect 471250 481898 471486 482134
rect 477514 482218 477750 482454
rect 477514 481898 477750 482134
rect 499250 482218 499486 482454
rect 499250 481898 499486 482134
rect 505514 482218 505750 482454
rect 505514 481898 505750 482134
rect 527250 482218 527486 482454
rect 527250 481898 527486 482134
rect 533514 482218 533750 482454
rect 533514 481898 533750 482134
rect 555250 482218 555486 482454
rect 555250 481898 555486 482134
rect 561514 482218 561750 482454
rect 561514 481898 561750 482134
rect -1974 458593 -1738 458829
rect -1654 458593 -1418 458829
rect -1974 458273 -1738 458509
rect -1654 458273 -1418 458509
rect 20118 458593 20354 458829
rect 20118 458273 20354 458509
rect 26382 458593 26618 458829
rect 26382 458273 26618 458509
rect 32646 458593 32882 458829
rect 32646 458273 32882 458509
rect 48118 458593 48354 458829
rect 48118 458273 48354 458509
rect 54382 458593 54618 458829
rect 54382 458273 54618 458509
rect 60646 458593 60882 458829
rect 60646 458273 60882 458509
rect 76118 458593 76354 458829
rect 76118 458273 76354 458509
rect 23250 455218 23486 455454
rect 23250 454898 23486 455134
rect 29514 455218 29750 455454
rect 29514 454898 29750 455134
rect 51250 455218 51486 455454
rect 51250 454898 51486 455134
rect 57514 455218 57750 455454
rect 57514 454898 57750 455134
rect 79250 455218 79486 455454
rect 79250 454898 79486 455134
rect 82382 458593 82618 458829
rect 82382 458273 82618 458509
rect 88646 458593 88882 458829
rect 88646 458273 88882 458509
rect 104118 458593 104354 458829
rect 104118 458273 104354 458509
rect 110382 458593 110618 458829
rect 110382 458273 110618 458509
rect 116646 458593 116882 458829
rect 116646 458273 116882 458509
rect 132118 458593 132354 458829
rect 132118 458273 132354 458509
rect 138382 458593 138618 458829
rect 138382 458273 138618 458509
rect 144646 458593 144882 458829
rect 144646 458273 144882 458509
rect 160118 458593 160354 458829
rect 160118 458273 160354 458509
rect 85514 455218 85750 455454
rect 85514 454898 85750 455134
rect 107250 455218 107486 455454
rect 107250 454898 107486 455134
rect 113514 455218 113750 455454
rect 113514 454898 113750 455134
rect 135250 455218 135486 455454
rect 135250 454898 135486 455134
rect 141514 455218 141750 455454
rect 141514 454898 141750 455134
rect 163250 455218 163486 455454
rect 163250 454898 163486 455134
rect 166382 458593 166618 458829
rect 166382 458273 166618 458509
rect 172646 458593 172882 458829
rect 172646 458273 172882 458509
rect 188118 458593 188354 458829
rect 188118 458273 188354 458509
rect 194382 458593 194618 458829
rect 194382 458273 194618 458509
rect 200646 458593 200882 458829
rect 200646 458273 200882 458509
rect 216118 458593 216354 458829
rect 216118 458273 216354 458509
rect 222382 458593 222618 458829
rect 222382 458273 222618 458509
rect 228646 458593 228882 458829
rect 228646 458273 228882 458509
rect 244118 458593 244354 458829
rect 244118 458273 244354 458509
rect 250382 458593 250618 458829
rect 250382 458273 250618 458509
rect 256646 458593 256882 458829
rect 256646 458273 256882 458509
rect 169514 455218 169750 455454
rect 169514 454898 169750 455134
rect 191250 455218 191486 455454
rect 191250 454898 191486 455134
rect 197514 455218 197750 455454
rect 197514 454898 197750 455134
rect 219250 455218 219486 455454
rect 219250 454898 219486 455134
rect 225514 455218 225750 455454
rect 225514 454898 225750 455134
rect 247250 455218 247486 455454
rect 247250 454898 247486 455134
rect 253514 455218 253750 455454
rect 253514 454898 253750 455134
rect 272118 458593 272354 458829
rect 272118 458273 272354 458509
rect 278382 458593 278618 458829
rect 278382 458273 278618 458509
rect 284646 458593 284882 458829
rect 284646 458273 284882 458509
rect 300118 458593 300354 458829
rect 300118 458273 300354 458509
rect 306382 458593 306618 458829
rect 306382 458273 306618 458509
rect 312646 458593 312882 458829
rect 312646 458273 312882 458509
rect 328118 458593 328354 458829
rect 328118 458273 328354 458509
rect 334382 458593 334618 458829
rect 334382 458273 334618 458509
rect 340646 458593 340882 458829
rect 340646 458273 340882 458509
rect 356118 458593 356354 458829
rect 356118 458273 356354 458509
rect 275250 455218 275486 455454
rect 275250 454898 275486 455134
rect 281514 455218 281750 455454
rect 281514 454898 281750 455134
rect 303250 455218 303486 455454
rect 303250 454898 303486 455134
rect 309514 455218 309750 455454
rect 309514 454898 309750 455134
rect 331250 455218 331486 455454
rect 331250 454898 331486 455134
rect 337514 455218 337750 455454
rect 337514 454898 337750 455134
rect 359250 455218 359486 455454
rect 359250 454898 359486 455134
rect 362382 458593 362618 458829
rect 362382 458273 362618 458509
rect 368646 458593 368882 458829
rect 368646 458273 368882 458509
rect 384118 458593 384354 458829
rect 384118 458273 384354 458509
rect 390382 458593 390618 458829
rect 390382 458273 390618 458509
rect 396646 458593 396882 458829
rect 396646 458273 396882 458509
rect 412118 458593 412354 458829
rect 412118 458273 412354 458509
rect 418382 458593 418618 458829
rect 418382 458273 418618 458509
rect 424646 458593 424882 458829
rect 424646 458273 424882 458509
rect 440118 458593 440354 458829
rect 440118 458273 440354 458509
rect 365514 455218 365750 455454
rect 365514 454898 365750 455134
rect 387250 455218 387486 455454
rect 387250 454898 387486 455134
rect 393514 455218 393750 455454
rect 393514 454898 393750 455134
rect 415250 455218 415486 455454
rect 415250 454898 415486 455134
rect 421514 455218 421750 455454
rect 421514 454898 421750 455134
rect 443250 455218 443486 455454
rect 443250 454898 443486 455134
rect 446382 458593 446618 458829
rect 446382 458273 446618 458509
rect 452646 458593 452882 458829
rect 452646 458273 452882 458509
rect 449514 455218 449750 455454
rect 449514 454898 449750 455134
rect 468118 458593 468354 458829
rect 468118 458273 468354 458509
rect 474382 458593 474618 458829
rect 474382 458273 474618 458509
rect 480646 458593 480882 458829
rect 480646 458273 480882 458509
rect 496118 458593 496354 458829
rect 496118 458273 496354 458509
rect 502382 458593 502618 458829
rect 502382 458273 502618 458509
rect 508646 458593 508882 458829
rect 508646 458273 508882 458509
rect 524118 458593 524354 458829
rect 524118 458273 524354 458509
rect 530382 458593 530618 458829
rect 530382 458273 530618 458509
rect 536646 458593 536882 458829
rect 536646 458273 536882 458509
rect 552118 458593 552354 458829
rect 552118 458273 552354 458509
rect 471250 455218 471486 455454
rect 471250 454898 471486 455134
rect 477514 455218 477750 455454
rect 477514 454898 477750 455134
rect 499250 455218 499486 455454
rect 499250 454898 499486 455134
rect 505514 455218 505750 455454
rect 505514 454898 505750 455134
rect 527250 455218 527486 455454
rect 527250 454898 527486 455134
rect 533514 455218 533750 455454
rect 533514 454898 533750 455134
rect 555250 455218 555486 455454
rect 555250 454898 555486 455134
rect 558382 458593 558618 458829
rect 558382 458273 558618 458509
rect 564646 458593 564882 458829
rect 564646 458273 564882 458509
rect 573526 458593 573762 458829
rect 573846 458593 574082 458829
rect 573526 458273 573762 458509
rect 573846 458273 574082 458509
rect 561514 455218 561750 455454
rect 561514 454898 561750 455134
rect -1974 431593 -1738 431829
rect -1654 431593 -1418 431829
rect -1974 431273 -1738 431509
rect -1654 431273 -1418 431509
rect 20118 431593 20354 431829
rect 20118 431273 20354 431509
rect 26382 431593 26618 431829
rect 26382 431273 26618 431509
rect 32646 431593 32882 431829
rect 32646 431273 32882 431509
rect 48118 431593 48354 431829
rect 48118 431273 48354 431509
rect 54382 431593 54618 431829
rect 54382 431273 54618 431509
rect 60646 431593 60882 431829
rect 60646 431273 60882 431509
rect 76118 431593 76354 431829
rect 76118 431273 76354 431509
rect 82382 431593 82618 431829
rect 82382 431273 82618 431509
rect 88646 431593 88882 431829
rect 88646 431273 88882 431509
rect 104118 431593 104354 431829
rect 104118 431273 104354 431509
rect 110382 431593 110618 431829
rect 110382 431273 110618 431509
rect 116646 431593 116882 431829
rect 116646 431273 116882 431509
rect 23250 428218 23486 428454
rect 23250 427898 23486 428134
rect 29514 428218 29750 428454
rect 29514 427898 29750 428134
rect 51250 428218 51486 428454
rect 51250 427898 51486 428134
rect 57514 428218 57750 428454
rect 57514 427898 57750 428134
rect 79250 428218 79486 428454
rect 79250 427898 79486 428134
rect 85514 428218 85750 428454
rect 85514 427898 85750 428134
rect 107250 428218 107486 428454
rect 107250 427898 107486 428134
rect 113514 428218 113750 428454
rect 113514 427898 113750 428134
rect 132118 431593 132354 431829
rect 132118 431273 132354 431509
rect 138382 431593 138618 431829
rect 138382 431273 138618 431509
rect 144646 431593 144882 431829
rect 144646 431273 144882 431509
rect 160118 431593 160354 431829
rect 160118 431273 160354 431509
rect 166382 431593 166618 431829
rect 166382 431273 166618 431509
rect 172646 431593 172882 431829
rect 172646 431273 172882 431509
rect 188118 431593 188354 431829
rect 188118 431273 188354 431509
rect 194382 431593 194618 431829
rect 194382 431273 194618 431509
rect 135250 428218 135486 428454
rect 135250 427898 135486 428134
rect 141514 428218 141750 428454
rect 141514 427898 141750 428134
rect 163250 428218 163486 428454
rect 163250 427898 163486 428134
rect 169514 428218 169750 428454
rect 169514 427898 169750 428134
rect 191250 428218 191486 428454
rect 191250 427898 191486 428134
rect 200646 431593 200882 431829
rect 200646 431273 200882 431509
rect 216118 431593 216354 431829
rect 216118 431273 216354 431509
rect 222382 431593 222618 431829
rect 222382 431273 222618 431509
rect 228646 431593 228882 431829
rect 228646 431273 228882 431509
rect 244118 431593 244354 431829
rect 244118 431273 244354 431509
rect 250382 431593 250618 431829
rect 250382 431273 250618 431509
rect 256646 431593 256882 431829
rect 256646 431273 256882 431509
rect 272118 431593 272354 431829
rect 272118 431273 272354 431509
rect 278382 431593 278618 431829
rect 278382 431273 278618 431509
rect 284646 431593 284882 431829
rect 284646 431273 284882 431509
rect 300118 431593 300354 431829
rect 300118 431273 300354 431509
rect 306382 431593 306618 431829
rect 306382 431273 306618 431509
rect 312646 431593 312882 431829
rect 312646 431273 312882 431509
rect 328118 431593 328354 431829
rect 328118 431273 328354 431509
rect 334382 431593 334618 431829
rect 334382 431273 334618 431509
rect 340646 431593 340882 431829
rect 340646 431273 340882 431509
rect 356118 431593 356354 431829
rect 356118 431273 356354 431509
rect 362382 431593 362618 431829
rect 362382 431273 362618 431509
rect 368646 431593 368882 431829
rect 368646 431273 368882 431509
rect 384118 431593 384354 431829
rect 384118 431273 384354 431509
rect 390382 431593 390618 431829
rect 390382 431273 390618 431509
rect 197514 428218 197750 428454
rect 197514 427898 197750 428134
rect 219250 428218 219486 428454
rect 219250 427898 219486 428134
rect 225514 428218 225750 428454
rect 225514 427898 225750 428134
rect 247250 428218 247486 428454
rect 247250 427898 247486 428134
rect 253514 428218 253750 428454
rect 253514 427898 253750 428134
rect 275250 428218 275486 428454
rect 275250 427898 275486 428134
rect 281514 428218 281750 428454
rect 281514 427898 281750 428134
rect 303250 428218 303486 428454
rect 303250 427898 303486 428134
rect 309514 428218 309750 428454
rect 309514 427898 309750 428134
rect 331250 428218 331486 428454
rect 331250 427898 331486 428134
rect 337514 428218 337750 428454
rect 337514 427898 337750 428134
rect 359250 428218 359486 428454
rect 359250 427898 359486 428134
rect 365514 428218 365750 428454
rect 365514 427898 365750 428134
rect 387250 428218 387486 428454
rect 387250 427898 387486 428134
rect 396646 431593 396882 431829
rect 396646 431273 396882 431509
rect 412118 431593 412354 431829
rect 412118 431273 412354 431509
rect 418382 431593 418618 431829
rect 418382 431273 418618 431509
rect 424646 431593 424882 431829
rect 424646 431273 424882 431509
rect 440118 431593 440354 431829
rect 440118 431273 440354 431509
rect 446382 431593 446618 431829
rect 446382 431273 446618 431509
rect 452646 431593 452882 431829
rect 452646 431273 452882 431509
rect 468118 431593 468354 431829
rect 468118 431273 468354 431509
rect 474382 431593 474618 431829
rect 474382 431273 474618 431509
rect 480646 431593 480882 431829
rect 480646 431273 480882 431509
rect 496118 431593 496354 431829
rect 496118 431273 496354 431509
rect 502382 431593 502618 431829
rect 502382 431273 502618 431509
rect 508646 431593 508882 431829
rect 508646 431273 508882 431509
rect 524118 431593 524354 431829
rect 524118 431273 524354 431509
rect 530382 431593 530618 431829
rect 530382 431273 530618 431509
rect 536646 431593 536882 431829
rect 536646 431273 536882 431509
rect 552118 431593 552354 431829
rect 552118 431273 552354 431509
rect 558382 431593 558618 431829
rect 558382 431273 558618 431509
rect 564646 431593 564882 431829
rect 564646 431273 564882 431509
rect 573526 431593 573762 431829
rect 573846 431593 574082 431829
rect 573526 431273 573762 431509
rect 573846 431273 574082 431509
rect 393514 428218 393750 428454
rect 393514 427898 393750 428134
rect 415250 428218 415486 428454
rect 415250 427898 415486 428134
rect 421514 428218 421750 428454
rect 421514 427898 421750 428134
rect 443250 428218 443486 428454
rect 443250 427898 443486 428134
rect 449514 428218 449750 428454
rect 449514 427898 449750 428134
rect 471250 428218 471486 428454
rect 471250 427898 471486 428134
rect 477514 428218 477750 428454
rect 477514 427898 477750 428134
rect 499250 428218 499486 428454
rect 499250 427898 499486 428134
rect 505514 428218 505750 428454
rect 505514 427898 505750 428134
rect 527250 428218 527486 428454
rect 527250 427898 527486 428134
rect 533514 428218 533750 428454
rect 533514 427898 533750 428134
rect 555250 428218 555486 428454
rect 555250 427898 555486 428134
rect 561514 428218 561750 428454
rect 561514 427898 561750 428134
rect -1974 404593 -1738 404829
rect -1654 404593 -1418 404829
rect -1974 404273 -1738 404509
rect -1654 404273 -1418 404509
rect 20118 404593 20354 404829
rect 20118 404273 20354 404509
rect 26382 404593 26618 404829
rect 26382 404273 26618 404509
rect 32646 404593 32882 404829
rect 32646 404273 32882 404509
rect 48118 404593 48354 404829
rect 48118 404273 48354 404509
rect 54382 404593 54618 404829
rect 54382 404273 54618 404509
rect 60646 404593 60882 404829
rect 60646 404273 60882 404509
rect 76118 404593 76354 404829
rect 76118 404273 76354 404509
rect 23250 401218 23486 401454
rect 23250 400898 23486 401134
rect 29514 401218 29750 401454
rect 29514 400898 29750 401134
rect 51250 401218 51486 401454
rect 51250 400898 51486 401134
rect 57514 401218 57750 401454
rect 57514 400898 57750 401134
rect 79250 401218 79486 401454
rect 79250 400898 79486 401134
rect 82382 404593 82618 404829
rect 82382 404273 82618 404509
rect 88646 404593 88882 404829
rect 88646 404273 88882 404509
rect 104118 404593 104354 404829
rect 104118 404273 104354 404509
rect 110382 404593 110618 404829
rect 110382 404273 110618 404509
rect 116646 404593 116882 404829
rect 116646 404273 116882 404509
rect 132118 404593 132354 404829
rect 132118 404273 132354 404509
rect 138382 404593 138618 404829
rect 138382 404273 138618 404509
rect 144646 404593 144882 404829
rect 144646 404273 144882 404509
rect 160118 404593 160354 404829
rect 160118 404273 160354 404509
rect 85514 401218 85750 401454
rect 85514 400898 85750 401134
rect 107250 401218 107486 401454
rect 107250 400898 107486 401134
rect 113514 401218 113750 401454
rect 113514 400898 113750 401134
rect 135250 401218 135486 401454
rect 135250 400898 135486 401134
rect 141514 401218 141750 401454
rect 141514 400898 141750 401134
rect 163250 401218 163486 401454
rect 163250 400898 163486 401134
rect 166382 404593 166618 404829
rect 166382 404273 166618 404509
rect 172646 404593 172882 404829
rect 172646 404273 172882 404509
rect 188118 404593 188354 404829
rect 188118 404273 188354 404509
rect 194382 404593 194618 404829
rect 194382 404273 194618 404509
rect 200646 404593 200882 404829
rect 200646 404273 200882 404509
rect 216118 404593 216354 404829
rect 216118 404273 216354 404509
rect 222382 404593 222618 404829
rect 222382 404273 222618 404509
rect 228646 404593 228882 404829
rect 228646 404273 228882 404509
rect 244118 404593 244354 404829
rect 244118 404273 244354 404509
rect 250382 404593 250618 404829
rect 250382 404273 250618 404509
rect 256646 404593 256882 404829
rect 256646 404273 256882 404509
rect 169514 401218 169750 401454
rect 169514 400898 169750 401134
rect 191250 401218 191486 401454
rect 191250 400898 191486 401134
rect 197514 401218 197750 401454
rect 197514 400898 197750 401134
rect 219250 401218 219486 401454
rect 219250 400898 219486 401134
rect 225514 401218 225750 401454
rect 225514 400898 225750 401134
rect 247250 401218 247486 401454
rect 247250 400898 247486 401134
rect 253514 401218 253750 401454
rect 253514 400898 253750 401134
rect 272118 404593 272354 404829
rect 272118 404273 272354 404509
rect 278382 404593 278618 404829
rect 278382 404273 278618 404509
rect 284646 404593 284882 404829
rect 284646 404273 284882 404509
rect 300118 404593 300354 404829
rect 300118 404273 300354 404509
rect 306382 404593 306618 404829
rect 306382 404273 306618 404509
rect 312646 404593 312882 404829
rect 312646 404273 312882 404509
rect 328118 404593 328354 404829
rect 328118 404273 328354 404509
rect 334382 404593 334618 404829
rect 334382 404273 334618 404509
rect 340646 404593 340882 404829
rect 340646 404273 340882 404509
rect 356118 404593 356354 404829
rect 356118 404273 356354 404509
rect 275250 401218 275486 401454
rect 275250 400898 275486 401134
rect 281514 401218 281750 401454
rect 281514 400898 281750 401134
rect 303250 401218 303486 401454
rect 303250 400898 303486 401134
rect 309514 401218 309750 401454
rect 309514 400898 309750 401134
rect 331250 401218 331486 401454
rect 331250 400898 331486 401134
rect 337514 401218 337750 401454
rect 337514 400898 337750 401134
rect 359250 401218 359486 401454
rect 359250 400898 359486 401134
rect 362382 404593 362618 404829
rect 362382 404273 362618 404509
rect 368646 404593 368882 404829
rect 368646 404273 368882 404509
rect 384118 404593 384354 404829
rect 384118 404273 384354 404509
rect 390382 404593 390618 404829
rect 390382 404273 390618 404509
rect 396646 404593 396882 404829
rect 396646 404273 396882 404509
rect 412118 404593 412354 404829
rect 412118 404273 412354 404509
rect 418382 404593 418618 404829
rect 418382 404273 418618 404509
rect 424646 404593 424882 404829
rect 424646 404273 424882 404509
rect 440118 404593 440354 404829
rect 440118 404273 440354 404509
rect 365514 401218 365750 401454
rect 365514 400898 365750 401134
rect 387250 401218 387486 401454
rect 387250 400898 387486 401134
rect 393514 401218 393750 401454
rect 393514 400898 393750 401134
rect 415250 401218 415486 401454
rect 415250 400898 415486 401134
rect 421514 401218 421750 401454
rect 421514 400898 421750 401134
rect 443250 401218 443486 401454
rect 443250 400898 443486 401134
rect 446382 404593 446618 404829
rect 446382 404273 446618 404509
rect 452646 404593 452882 404829
rect 452646 404273 452882 404509
rect 449514 401218 449750 401454
rect 449514 400898 449750 401134
rect 468118 404593 468354 404829
rect 468118 404273 468354 404509
rect 474382 404593 474618 404829
rect 474382 404273 474618 404509
rect 480646 404593 480882 404829
rect 480646 404273 480882 404509
rect 496118 404593 496354 404829
rect 496118 404273 496354 404509
rect 502382 404593 502618 404829
rect 502382 404273 502618 404509
rect 508646 404593 508882 404829
rect 508646 404273 508882 404509
rect 524118 404593 524354 404829
rect 524118 404273 524354 404509
rect 530382 404593 530618 404829
rect 530382 404273 530618 404509
rect 536646 404593 536882 404829
rect 536646 404273 536882 404509
rect 552118 404593 552354 404829
rect 552118 404273 552354 404509
rect 471250 401218 471486 401454
rect 471250 400898 471486 401134
rect 477514 401218 477750 401454
rect 477514 400898 477750 401134
rect 499250 401218 499486 401454
rect 499250 400898 499486 401134
rect 505514 401218 505750 401454
rect 505514 400898 505750 401134
rect 527250 401218 527486 401454
rect 527250 400898 527486 401134
rect 533514 401218 533750 401454
rect 533514 400898 533750 401134
rect 555250 401218 555486 401454
rect 555250 400898 555486 401134
rect 558382 404593 558618 404829
rect 558382 404273 558618 404509
rect 564646 404593 564882 404829
rect 564646 404273 564882 404509
rect 573526 404593 573762 404829
rect 573846 404593 574082 404829
rect 573526 404273 573762 404509
rect 573846 404273 574082 404509
rect 561514 401218 561750 401454
rect 561514 400898 561750 401134
rect -1974 377593 -1738 377829
rect -1654 377593 -1418 377829
rect -1974 377273 -1738 377509
rect -1654 377273 -1418 377509
rect 20118 377593 20354 377829
rect 20118 377273 20354 377509
rect 26382 377593 26618 377829
rect 26382 377273 26618 377509
rect 32646 377593 32882 377829
rect 32646 377273 32882 377509
rect 48118 377593 48354 377829
rect 48118 377273 48354 377509
rect 54382 377593 54618 377829
rect 54382 377273 54618 377509
rect 60646 377593 60882 377829
rect 60646 377273 60882 377509
rect 76118 377593 76354 377829
rect 76118 377273 76354 377509
rect 82382 377593 82618 377829
rect 82382 377273 82618 377509
rect 88646 377593 88882 377829
rect 88646 377273 88882 377509
rect 104118 377593 104354 377829
rect 104118 377273 104354 377509
rect 110382 377593 110618 377829
rect 110382 377273 110618 377509
rect 116646 377593 116882 377829
rect 116646 377273 116882 377509
rect 23250 374218 23486 374454
rect 23250 373898 23486 374134
rect 29514 374218 29750 374454
rect 29514 373898 29750 374134
rect 51250 374218 51486 374454
rect 51250 373898 51486 374134
rect 57514 374218 57750 374454
rect 57514 373898 57750 374134
rect 79250 374218 79486 374454
rect 79250 373898 79486 374134
rect 85514 374218 85750 374454
rect 85514 373898 85750 374134
rect 107250 374218 107486 374454
rect 107250 373898 107486 374134
rect 113514 374218 113750 374454
rect 113514 373898 113750 374134
rect 132118 377593 132354 377829
rect 132118 377273 132354 377509
rect 138382 377593 138618 377829
rect 138382 377273 138618 377509
rect 144646 377593 144882 377829
rect 144646 377273 144882 377509
rect 160118 377593 160354 377829
rect 160118 377273 160354 377509
rect 166382 377593 166618 377829
rect 166382 377273 166618 377509
rect 172646 377593 172882 377829
rect 172646 377273 172882 377509
rect 188118 377593 188354 377829
rect 188118 377273 188354 377509
rect 194382 377593 194618 377829
rect 194382 377273 194618 377509
rect 135250 374218 135486 374454
rect 135250 373898 135486 374134
rect 141514 374218 141750 374454
rect 141514 373898 141750 374134
rect 163250 374218 163486 374454
rect 163250 373898 163486 374134
rect 169514 374218 169750 374454
rect 169514 373898 169750 374134
rect 191250 374218 191486 374454
rect 191250 373898 191486 374134
rect 200646 377593 200882 377829
rect 200646 377273 200882 377509
rect 216118 377593 216354 377829
rect 216118 377273 216354 377509
rect 222382 377593 222618 377829
rect 222382 377273 222618 377509
rect 228646 377593 228882 377829
rect 228646 377273 228882 377509
rect 244118 377593 244354 377829
rect 244118 377273 244354 377509
rect 250382 377593 250618 377829
rect 250382 377273 250618 377509
rect 256646 377593 256882 377829
rect 256646 377273 256882 377509
rect 272118 377593 272354 377829
rect 272118 377273 272354 377509
rect 278382 377593 278618 377829
rect 278382 377273 278618 377509
rect 284646 377593 284882 377829
rect 284646 377273 284882 377509
rect 300118 377593 300354 377829
rect 300118 377273 300354 377509
rect 306382 377593 306618 377829
rect 306382 377273 306618 377509
rect 312646 377593 312882 377829
rect 312646 377273 312882 377509
rect 328118 377593 328354 377829
rect 328118 377273 328354 377509
rect 334382 377593 334618 377829
rect 334382 377273 334618 377509
rect 340646 377593 340882 377829
rect 340646 377273 340882 377509
rect 356118 377593 356354 377829
rect 356118 377273 356354 377509
rect 362382 377593 362618 377829
rect 362382 377273 362618 377509
rect 368646 377593 368882 377829
rect 368646 377273 368882 377509
rect 384118 377593 384354 377829
rect 384118 377273 384354 377509
rect 390382 377593 390618 377829
rect 390382 377273 390618 377509
rect 197514 374218 197750 374454
rect 197514 373898 197750 374134
rect 219250 374218 219486 374454
rect 219250 373898 219486 374134
rect 225514 374218 225750 374454
rect 225514 373898 225750 374134
rect 247250 374218 247486 374454
rect 247250 373898 247486 374134
rect 253514 374218 253750 374454
rect 253514 373898 253750 374134
rect 275250 374218 275486 374454
rect 275250 373898 275486 374134
rect 281514 374218 281750 374454
rect 281514 373898 281750 374134
rect 303250 374218 303486 374454
rect 303250 373898 303486 374134
rect 309514 374218 309750 374454
rect 309514 373898 309750 374134
rect 331250 374218 331486 374454
rect 331250 373898 331486 374134
rect 337514 374218 337750 374454
rect 337514 373898 337750 374134
rect 359250 374218 359486 374454
rect 359250 373898 359486 374134
rect 365514 374218 365750 374454
rect 365514 373898 365750 374134
rect 387250 374218 387486 374454
rect 387250 373898 387486 374134
rect 396646 377593 396882 377829
rect 396646 377273 396882 377509
rect 412118 377593 412354 377829
rect 412118 377273 412354 377509
rect 418382 377593 418618 377829
rect 418382 377273 418618 377509
rect 424646 377593 424882 377829
rect 424646 377273 424882 377509
rect 440118 377593 440354 377829
rect 440118 377273 440354 377509
rect 446382 377593 446618 377829
rect 446382 377273 446618 377509
rect 452646 377593 452882 377829
rect 452646 377273 452882 377509
rect 468118 377593 468354 377829
rect 468118 377273 468354 377509
rect 474382 377593 474618 377829
rect 474382 377273 474618 377509
rect 480646 377593 480882 377829
rect 480646 377273 480882 377509
rect 496118 377593 496354 377829
rect 496118 377273 496354 377509
rect 502382 377593 502618 377829
rect 502382 377273 502618 377509
rect 508646 377593 508882 377829
rect 508646 377273 508882 377509
rect 524118 377593 524354 377829
rect 524118 377273 524354 377509
rect 530382 377593 530618 377829
rect 530382 377273 530618 377509
rect 536646 377593 536882 377829
rect 536646 377273 536882 377509
rect 552118 377593 552354 377829
rect 552118 377273 552354 377509
rect 558382 377593 558618 377829
rect 558382 377273 558618 377509
rect 564646 377593 564882 377829
rect 564646 377273 564882 377509
rect 573526 377593 573762 377829
rect 573846 377593 574082 377829
rect 573526 377273 573762 377509
rect 573846 377273 574082 377509
rect 393514 374218 393750 374454
rect 393514 373898 393750 374134
rect 415250 374218 415486 374454
rect 415250 373898 415486 374134
rect 421514 374218 421750 374454
rect 421514 373898 421750 374134
rect 443250 374218 443486 374454
rect 443250 373898 443486 374134
rect 449514 374218 449750 374454
rect 449514 373898 449750 374134
rect 471250 374218 471486 374454
rect 471250 373898 471486 374134
rect 477514 374218 477750 374454
rect 477514 373898 477750 374134
rect 499250 374218 499486 374454
rect 499250 373898 499486 374134
rect 505514 374218 505750 374454
rect 505514 373898 505750 374134
rect 527250 374218 527486 374454
rect 527250 373898 527486 374134
rect 533514 374218 533750 374454
rect 533514 373898 533750 374134
rect 555250 374218 555486 374454
rect 555250 373898 555486 374134
rect 561514 374218 561750 374454
rect 561514 373898 561750 374134
rect -1974 350593 -1738 350829
rect -1654 350593 -1418 350829
rect -1974 350273 -1738 350509
rect -1654 350273 -1418 350509
rect 20118 350593 20354 350829
rect 20118 350273 20354 350509
rect 26382 350593 26618 350829
rect 26382 350273 26618 350509
rect 32646 350593 32882 350829
rect 32646 350273 32882 350509
rect 48118 350593 48354 350829
rect 48118 350273 48354 350509
rect 54382 350593 54618 350829
rect 54382 350273 54618 350509
rect 60646 350593 60882 350829
rect 60646 350273 60882 350509
rect 76118 350593 76354 350829
rect 76118 350273 76354 350509
rect 82382 350593 82618 350829
rect 82382 350273 82618 350509
rect 88646 350593 88882 350829
rect 88646 350273 88882 350509
rect 104118 350593 104354 350829
rect 104118 350273 104354 350509
rect 110382 350593 110618 350829
rect 110382 350273 110618 350509
rect 116646 350593 116882 350829
rect 116646 350273 116882 350509
rect 132118 350593 132354 350829
rect 132118 350273 132354 350509
rect 138382 350593 138618 350829
rect 138382 350273 138618 350509
rect 144646 350593 144882 350829
rect 144646 350273 144882 350509
rect 160118 350593 160354 350829
rect 160118 350273 160354 350509
rect 23250 347218 23486 347454
rect 23250 346898 23486 347134
rect 29514 347218 29750 347454
rect 29514 346898 29750 347134
rect 51250 347218 51486 347454
rect 51250 346898 51486 347134
rect 57514 347218 57750 347454
rect 57514 346898 57750 347134
rect 79250 347218 79486 347454
rect 79250 346898 79486 347134
rect 85514 347218 85750 347454
rect 85514 346898 85750 347134
rect 107250 347218 107486 347454
rect 107250 346898 107486 347134
rect 113514 347218 113750 347454
rect 113514 346898 113750 347134
rect 135250 347218 135486 347454
rect 135250 346898 135486 347134
rect 141514 347218 141750 347454
rect 141514 346898 141750 347134
rect 163250 347218 163486 347454
rect 163250 346898 163486 347134
rect 166382 350593 166618 350829
rect 166382 350273 166618 350509
rect 172646 350593 172882 350829
rect 172646 350273 172882 350509
rect 188118 350593 188354 350829
rect 188118 350273 188354 350509
rect 194382 350593 194618 350829
rect 194382 350273 194618 350509
rect 200646 350593 200882 350829
rect 200646 350273 200882 350509
rect 216118 350593 216354 350829
rect 216118 350273 216354 350509
rect 222382 350593 222618 350829
rect 222382 350273 222618 350509
rect 228646 350593 228882 350829
rect 228646 350273 228882 350509
rect 244118 350593 244354 350829
rect 244118 350273 244354 350509
rect 250382 350593 250618 350829
rect 250382 350273 250618 350509
rect 256646 350593 256882 350829
rect 256646 350273 256882 350509
rect 169514 347218 169750 347454
rect 169514 346898 169750 347134
rect 191250 347218 191486 347454
rect 191250 346898 191486 347134
rect 197514 347218 197750 347454
rect 197514 346898 197750 347134
rect 219250 347218 219486 347454
rect 219250 346898 219486 347134
rect 225514 347218 225750 347454
rect 225514 346898 225750 347134
rect 247250 347218 247486 347454
rect 247250 346898 247486 347134
rect 253514 347218 253750 347454
rect 253514 346898 253750 347134
rect 272118 350593 272354 350829
rect 272118 350273 272354 350509
rect 278382 350593 278618 350829
rect 278382 350273 278618 350509
rect 284646 350593 284882 350829
rect 284646 350273 284882 350509
rect 300118 350593 300354 350829
rect 300118 350273 300354 350509
rect 306382 350593 306618 350829
rect 306382 350273 306618 350509
rect 312646 350593 312882 350829
rect 312646 350273 312882 350509
rect 328118 350593 328354 350829
rect 328118 350273 328354 350509
rect 334382 350593 334618 350829
rect 334382 350273 334618 350509
rect 340646 350593 340882 350829
rect 340646 350273 340882 350509
rect 356118 350593 356354 350829
rect 356118 350273 356354 350509
rect 275250 347218 275486 347454
rect 275250 346898 275486 347134
rect 281514 347218 281750 347454
rect 281514 346898 281750 347134
rect 303250 347218 303486 347454
rect 303250 346898 303486 347134
rect 309514 347218 309750 347454
rect 309514 346898 309750 347134
rect 331250 347218 331486 347454
rect 331250 346898 331486 347134
rect 337514 347218 337750 347454
rect 337514 346898 337750 347134
rect 359250 347218 359486 347454
rect 359250 346898 359486 347134
rect 362382 350593 362618 350829
rect 362382 350273 362618 350509
rect 368646 350593 368882 350829
rect 368646 350273 368882 350509
rect 384118 350593 384354 350829
rect 384118 350273 384354 350509
rect 390382 350593 390618 350829
rect 390382 350273 390618 350509
rect 396646 350593 396882 350829
rect 396646 350273 396882 350509
rect 412118 350593 412354 350829
rect 412118 350273 412354 350509
rect 418382 350593 418618 350829
rect 418382 350273 418618 350509
rect 424646 350593 424882 350829
rect 424646 350273 424882 350509
rect 440118 350593 440354 350829
rect 440118 350273 440354 350509
rect 365514 347218 365750 347454
rect 365514 346898 365750 347134
rect 387250 347218 387486 347454
rect 387250 346898 387486 347134
rect 393514 347218 393750 347454
rect 393514 346898 393750 347134
rect 415250 347218 415486 347454
rect 415250 346898 415486 347134
rect 421514 347218 421750 347454
rect 421514 346898 421750 347134
rect 443250 347218 443486 347454
rect 443250 346898 443486 347134
rect 446382 350593 446618 350829
rect 446382 350273 446618 350509
rect 452646 350593 452882 350829
rect 452646 350273 452882 350509
rect 468118 350593 468354 350829
rect 468118 350273 468354 350509
rect 474382 350593 474618 350829
rect 474382 350273 474618 350509
rect 480646 350593 480882 350829
rect 480646 350273 480882 350509
rect 496118 350593 496354 350829
rect 496118 350273 496354 350509
rect 502382 350593 502618 350829
rect 502382 350273 502618 350509
rect 508646 350593 508882 350829
rect 508646 350273 508882 350509
rect 524118 350593 524354 350829
rect 524118 350273 524354 350509
rect 530382 350593 530618 350829
rect 530382 350273 530618 350509
rect 536646 350593 536882 350829
rect 536646 350273 536882 350509
rect 552118 350593 552354 350829
rect 552118 350273 552354 350509
rect 449514 347218 449750 347454
rect 449514 346898 449750 347134
rect 471250 347218 471486 347454
rect 471250 346898 471486 347134
rect 477514 347218 477750 347454
rect 477514 346898 477750 347134
rect 499250 347218 499486 347454
rect 499250 346898 499486 347134
rect 505514 347218 505750 347454
rect 505514 346898 505750 347134
rect 527250 347218 527486 347454
rect 527250 346898 527486 347134
rect 533514 347218 533750 347454
rect 533514 346898 533750 347134
rect 555250 347218 555486 347454
rect 555250 346898 555486 347134
rect 558382 350593 558618 350829
rect 558382 350273 558618 350509
rect 564646 350593 564882 350829
rect 564646 350273 564882 350509
rect 573526 350593 573762 350829
rect 573846 350593 574082 350829
rect 573526 350273 573762 350509
rect 573846 350273 574082 350509
rect 561514 347218 561750 347454
rect 561514 346898 561750 347134
rect -1974 323593 -1738 323829
rect -1654 323593 -1418 323829
rect -1974 323273 -1738 323509
rect -1654 323273 -1418 323509
rect 20118 323593 20354 323829
rect 20118 323273 20354 323509
rect 26382 323593 26618 323829
rect 26382 323273 26618 323509
rect 32646 323593 32882 323829
rect 32646 323273 32882 323509
rect 48118 323593 48354 323829
rect 48118 323273 48354 323509
rect 54382 323593 54618 323829
rect 54382 323273 54618 323509
rect 60646 323593 60882 323829
rect 60646 323273 60882 323509
rect 76118 323593 76354 323829
rect 76118 323273 76354 323509
rect 82382 323593 82618 323829
rect 82382 323273 82618 323509
rect 88646 323593 88882 323829
rect 88646 323273 88882 323509
rect 104118 323593 104354 323829
rect 104118 323273 104354 323509
rect 110382 323593 110618 323829
rect 110382 323273 110618 323509
rect 116646 323593 116882 323829
rect 116646 323273 116882 323509
rect 23250 320218 23486 320454
rect 23250 319898 23486 320134
rect 29514 320218 29750 320454
rect 29514 319898 29750 320134
rect 51250 320218 51486 320454
rect 51250 319898 51486 320134
rect 57514 320218 57750 320454
rect 57514 319898 57750 320134
rect 79250 320218 79486 320454
rect 79250 319898 79486 320134
rect 85514 320218 85750 320454
rect 85514 319898 85750 320134
rect 107250 320218 107486 320454
rect 107250 319898 107486 320134
rect 113514 320218 113750 320454
rect 113514 319898 113750 320134
rect 132118 323593 132354 323829
rect 132118 323273 132354 323509
rect 138382 323593 138618 323829
rect 138382 323273 138618 323509
rect 144646 323593 144882 323829
rect 144646 323273 144882 323509
rect 160118 323593 160354 323829
rect 160118 323273 160354 323509
rect 166382 323593 166618 323829
rect 166382 323273 166618 323509
rect 172646 323593 172882 323829
rect 172646 323273 172882 323509
rect 188118 323593 188354 323829
rect 188118 323273 188354 323509
rect 194382 323593 194618 323829
rect 194382 323273 194618 323509
rect 135250 320218 135486 320454
rect 135250 319898 135486 320134
rect 141514 320218 141750 320454
rect 141514 319898 141750 320134
rect 163250 320218 163486 320454
rect 163250 319898 163486 320134
rect 169514 320218 169750 320454
rect 169514 319898 169750 320134
rect 191250 320218 191486 320454
rect 191250 319898 191486 320134
rect 200646 323593 200882 323829
rect 200646 323273 200882 323509
rect 216118 323593 216354 323829
rect 216118 323273 216354 323509
rect 222382 323593 222618 323829
rect 222382 323273 222618 323509
rect 228646 323593 228882 323829
rect 228646 323273 228882 323509
rect 244118 323593 244354 323829
rect 244118 323273 244354 323509
rect 250382 323593 250618 323829
rect 250382 323273 250618 323509
rect 256646 323593 256882 323829
rect 256646 323273 256882 323509
rect 272118 323593 272354 323829
rect 272118 323273 272354 323509
rect 278382 323593 278618 323829
rect 278382 323273 278618 323509
rect 284646 323593 284882 323829
rect 284646 323273 284882 323509
rect 300118 323593 300354 323829
rect 300118 323273 300354 323509
rect 306382 323593 306618 323829
rect 306382 323273 306618 323509
rect 312646 323593 312882 323829
rect 312646 323273 312882 323509
rect 328118 323593 328354 323829
rect 328118 323273 328354 323509
rect 334382 323593 334618 323829
rect 334382 323273 334618 323509
rect 340646 323593 340882 323829
rect 340646 323273 340882 323509
rect 356118 323593 356354 323829
rect 356118 323273 356354 323509
rect 362382 323593 362618 323829
rect 362382 323273 362618 323509
rect 368646 323593 368882 323829
rect 368646 323273 368882 323509
rect 384118 323593 384354 323829
rect 384118 323273 384354 323509
rect 390382 323593 390618 323829
rect 390382 323273 390618 323509
rect 197514 320218 197750 320454
rect 197514 319898 197750 320134
rect 219250 320218 219486 320454
rect 219250 319898 219486 320134
rect 225514 320218 225750 320454
rect 225514 319898 225750 320134
rect 247250 320218 247486 320454
rect 247250 319898 247486 320134
rect 253514 320218 253750 320454
rect 253514 319898 253750 320134
rect 275250 320218 275486 320454
rect 275250 319898 275486 320134
rect 281514 320218 281750 320454
rect 281514 319898 281750 320134
rect 303250 320218 303486 320454
rect 303250 319898 303486 320134
rect 309514 320218 309750 320454
rect 309514 319898 309750 320134
rect 331250 320218 331486 320454
rect 331250 319898 331486 320134
rect 337514 320218 337750 320454
rect 337514 319898 337750 320134
rect 359250 320218 359486 320454
rect 359250 319898 359486 320134
rect 365514 320218 365750 320454
rect 365514 319898 365750 320134
rect 387250 320218 387486 320454
rect 387250 319898 387486 320134
rect 396646 323593 396882 323829
rect 396646 323273 396882 323509
rect 412118 323593 412354 323829
rect 412118 323273 412354 323509
rect 418382 323593 418618 323829
rect 418382 323273 418618 323509
rect 424646 323593 424882 323829
rect 424646 323273 424882 323509
rect 440118 323593 440354 323829
rect 440118 323273 440354 323509
rect 446382 323593 446618 323829
rect 446382 323273 446618 323509
rect 452646 323593 452882 323829
rect 452646 323273 452882 323509
rect 468118 323593 468354 323829
rect 468118 323273 468354 323509
rect 474382 323593 474618 323829
rect 474382 323273 474618 323509
rect 480646 323593 480882 323829
rect 480646 323273 480882 323509
rect 496118 323593 496354 323829
rect 496118 323273 496354 323509
rect 502382 323593 502618 323829
rect 502382 323273 502618 323509
rect 508646 323593 508882 323829
rect 508646 323273 508882 323509
rect 524118 323593 524354 323829
rect 524118 323273 524354 323509
rect 530382 323593 530618 323829
rect 530382 323273 530618 323509
rect 536646 323593 536882 323829
rect 536646 323273 536882 323509
rect 552118 323593 552354 323829
rect 552118 323273 552354 323509
rect 558382 323593 558618 323829
rect 558382 323273 558618 323509
rect 564646 323593 564882 323829
rect 564646 323273 564882 323509
rect 573526 323593 573762 323829
rect 573846 323593 574082 323829
rect 393514 320218 393750 320454
rect 393514 319898 393750 320134
rect 415250 320218 415486 320454
rect 415250 319898 415486 320134
rect 421514 320218 421750 320454
rect 421514 319898 421750 320134
rect 443250 320218 443486 320454
rect 443250 319898 443486 320134
rect 449514 320218 449750 320454
rect 449514 319898 449750 320134
rect 471250 320218 471486 320454
rect 471250 319898 471486 320134
rect 477514 320218 477750 320454
rect 477514 319898 477750 320134
rect 499250 320218 499486 320454
rect 499250 319898 499486 320134
rect 505514 320218 505750 320454
rect 505514 319898 505750 320134
rect 527250 320218 527486 320454
rect 527250 319898 527486 320134
rect 533514 320218 533750 320454
rect 533514 319898 533750 320134
rect 555250 320218 555486 320454
rect 555250 319898 555486 320134
rect 561514 320218 561750 320454
rect 561514 319898 561750 320134
rect 573526 323273 573762 323509
rect 573846 323273 574082 323509
rect -1974 296593 -1738 296829
rect -1654 296593 -1418 296829
rect -1974 296273 -1738 296509
rect -1654 296273 -1418 296509
rect 20118 296593 20354 296829
rect 20118 296273 20354 296509
rect 26382 296593 26618 296829
rect 26382 296273 26618 296509
rect 32646 296593 32882 296829
rect 32646 296273 32882 296509
rect 48118 296593 48354 296829
rect 48118 296273 48354 296509
rect 54382 296593 54618 296829
rect 54382 296273 54618 296509
rect 60646 296593 60882 296829
rect 60646 296273 60882 296509
rect 76118 296593 76354 296829
rect 76118 296273 76354 296509
rect 82382 296593 82618 296829
rect 82382 296273 82618 296509
rect 88646 296593 88882 296829
rect 88646 296273 88882 296509
rect 104118 296593 104354 296829
rect 104118 296273 104354 296509
rect 110382 296593 110618 296829
rect 110382 296273 110618 296509
rect 116646 296593 116882 296829
rect 116646 296273 116882 296509
rect 132118 296593 132354 296829
rect 132118 296273 132354 296509
rect 138382 296593 138618 296829
rect 138382 296273 138618 296509
rect 144646 296593 144882 296829
rect 144646 296273 144882 296509
rect 160118 296593 160354 296829
rect 160118 296273 160354 296509
rect 23250 293218 23486 293454
rect 23250 292898 23486 293134
rect 29514 293218 29750 293454
rect 29514 292898 29750 293134
rect 51250 293218 51486 293454
rect 51250 292898 51486 293134
rect 57514 293218 57750 293454
rect 57514 292898 57750 293134
rect 79250 293218 79486 293454
rect 79250 292898 79486 293134
rect 85514 293218 85750 293454
rect 85514 292898 85750 293134
rect 107250 293218 107486 293454
rect 107250 292898 107486 293134
rect 113514 293218 113750 293454
rect 113514 292898 113750 293134
rect 135250 293218 135486 293454
rect 135250 292898 135486 293134
rect 141514 293218 141750 293454
rect 141514 292898 141750 293134
rect 163250 293218 163486 293454
rect 163250 292898 163486 293134
rect 166382 296593 166618 296829
rect 166382 296273 166618 296509
rect 172646 296593 172882 296829
rect 172646 296273 172882 296509
rect 188118 296593 188354 296829
rect 188118 296273 188354 296509
rect 194382 296593 194618 296829
rect 194382 296273 194618 296509
rect 200646 296593 200882 296829
rect 200646 296273 200882 296509
rect 216118 296593 216354 296829
rect 216118 296273 216354 296509
rect 222382 296593 222618 296829
rect 222382 296273 222618 296509
rect 228646 296593 228882 296829
rect 228646 296273 228882 296509
rect 244118 296593 244354 296829
rect 244118 296273 244354 296509
rect 250382 296593 250618 296829
rect 250382 296273 250618 296509
rect 256646 296593 256882 296829
rect 256646 296273 256882 296509
rect 169514 293218 169750 293454
rect 169514 292898 169750 293134
rect 191250 293218 191486 293454
rect 191250 292898 191486 293134
rect 197514 293218 197750 293454
rect 197514 292898 197750 293134
rect 219250 293218 219486 293454
rect 219250 292898 219486 293134
rect 225514 293218 225750 293454
rect 225514 292898 225750 293134
rect 247250 293218 247486 293454
rect 247250 292898 247486 293134
rect 253514 293218 253750 293454
rect 253514 292898 253750 293134
rect 272118 296593 272354 296829
rect 272118 296273 272354 296509
rect 278382 296593 278618 296829
rect 278382 296273 278618 296509
rect 284646 296593 284882 296829
rect 284646 296273 284882 296509
rect 300118 296593 300354 296829
rect 300118 296273 300354 296509
rect 306382 296593 306618 296829
rect 306382 296273 306618 296509
rect 312646 296593 312882 296829
rect 312646 296273 312882 296509
rect 328118 296593 328354 296829
rect 328118 296273 328354 296509
rect 334382 296593 334618 296829
rect 334382 296273 334618 296509
rect 340646 296593 340882 296829
rect 340646 296273 340882 296509
rect 356118 296593 356354 296829
rect 356118 296273 356354 296509
rect 275250 293218 275486 293454
rect 275250 292898 275486 293134
rect 281514 293218 281750 293454
rect 281514 292898 281750 293134
rect 303250 293218 303486 293454
rect 303250 292898 303486 293134
rect 309514 293218 309750 293454
rect 309514 292898 309750 293134
rect 331250 293218 331486 293454
rect 331250 292898 331486 293134
rect 337514 293218 337750 293454
rect 337514 292898 337750 293134
rect 359250 293218 359486 293454
rect 359250 292898 359486 293134
rect 362382 296593 362618 296829
rect 362382 296273 362618 296509
rect 368646 296593 368882 296829
rect 368646 296273 368882 296509
rect 384118 296593 384354 296829
rect 384118 296273 384354 296509
rect 390382 296593 390618 296829
rect 390382 296273 390618 296509
rect 396646 296593 396882 296829
rect 396646 296273 396882 296509
rect 412118 296593 412354 296829
rect 412118 296273 412354 296509
rect 418382 296593 418618 296829
rect 418382 296273 418618 296509
rect 424646 296593 424882 296829
rect 424646 296273 424882 296509
rect 440118 296593 440354 296829
rect 440118 296273 440354 296509
rect 365514 293218 365750 293454
rect 365514 292898 365750 293134
rect 387250 293218 387486 293454
rect 387250 292898 387486 293134
rect 393514 293218 393750 293454
rect 393514 292898 393750 293134
rect 415250 293218 415486 293454
rect 415250 292898 415486 293134
rect 421514 293218 421750 293454
rect 421514 292898 421750 293134
rect 443250 293218 443486 293454
rect 443250 292898 443486 293134
rect 446382 296593 446618 296829
rect 446382 296273 446618 296509
rect 452646 296593 452882 296829
rect 452646 296273 452882 296509
rect 468118 296593 468354 296829
rect 468118 296273 468354 296509
rect 474382 296593 474618 296829
rect 474382 296273 474618 296509
rect 480646 296593 480882 296829
rect 480646 296273 480882 296509
rect 496118 296593 496354 296829
rect 496118 296273 496354 296509
rect 502382 296593 502618 296829
rect 502382 296273 502618 296509
rect 508646 296593 508882 296829
rect 508646 296273 508882 296509
rect 524118 296593 524354 296829
rect 524118 296273 524354 296509
rect 530382 296593 530618 296829
rect 530382 296273 530618 296509
rect 536646 296593 536882 296829
rect 536646 296273 536882 296509
rect 552118 296593 552354 296829
rect 552118 296273 552354 296509
rect 449514 293218 449750 293454
rect 449514 292898 449750 293134
rect 471250 293218 471486 293454
rect 471250 292898 471486 293134
rect 477514 293218 477750 293454
rect 477514 292898 477750 293134
rect 499250 293218 499486 293454
rect 499250 292898 499486 293134
rect 505514 293218 505750 293454
rect 505514 292898 505750 293134
rect 527250 293218 527486 293454
rect 527250 292898 527486 293134
rect 533514 293218 533750 293454
rect 533514 292898 533750 293134
rect 555250 293218 555486 293454
rect 555250 292898 555486 293134
rect 558382 296593 558618 296829
rect 558382 296273 558618 296509
rect 564646 296593 564882 296829
rect 564646 296273 564882 296509
rect 573526 296593 573762 296829
rect 573846 296593 574082 296829
rect 573526 296273 573762 296509
rect 573846 296273 574082 296509
rect 561514 293218 561750 293454
rect 561514 292898 561750 293134
rect -1974 269593 -1738 269829
rect -1654 269593 -1418 269829
rect -1974 269273 -1738 269509
rect -1654 269273 -1418 269509
rect 20118 269593 20354 269829
rect 20118 269273 20354 269509
rect 26382 269593 26618 269829
rect 26382 269273 26618 269509
rect 32646 269593 32882 269829
rect 32646 269273 32882 269509
rect 48118 269593 48354 269829
rect 48118 269273 48354 269509
rect 54382 269593 54618 269829
rect 54382 269273 54618 269509
rect 60646 269593 60882 269829
rect 60646 269273 60882 269509
rect 76118 269593 76354 269829
rect 76118 269273 76354 269509
rect 23250 266218 23486 266454
rect 23250 265898 23486 266134
rect 29514 266218 29750 266454
rect 29514 265898 29750 266134
rect 51250 266218 51486 266454
rect 51250 265898 51486 266134
rect 57514 266218 57750 266454
rect 57514 265898 57750 266134
rect 79250 266218 79486 266454
rect 79250 265898 79486 266134
rect 82382 269593 82618 269829
rect 82382 269273 82618 269509
rect 88646 269593 88882 269829
rect 88646 269273 88882 269509
rect 104118 269593 104354 269829
rect 104118 269273 104354 269509
rect 110382 269593 110618 269829
rect 110382 269273 110618 269509
rect 116646 269593 116882 269829
rect 116646 269273 116882 269509
rect 85514 266218 85750 266454
rect 85514 265898 85750 266134
rect 107250 266218 107486 266454
rect 107250 265898 107486 266134
rect 113514 266218 113750 266454
rect 113514 265898 113750 266134
rect 132118 269593 132354 269829
rect 132118 269273 132354 269509
rect 138382 269593 138618 269829
rect 138382 269273 138618 269509
rect 144646 269593 144882 269829
rect 144646 269273 144882 269509
rect 160118 269593 160354 269829
rect 160118 269273 160354 269509
rect 166382 269593 166618 269829
rect 166382 269273 166618 269509
rect 172646 269593 172882 269829
rect 172646 269273 172882 269509
rect 188118 269593 188354 269829
rect 188118 269273 188354 269509
rect 194382 269593 194618 269829
rect 194382 269273 194618 269509
rect 135250 266218 135486 266454
rect 135250 265898 135486 266134
rect 141514 266218 141750 266454
rect 141514 265898 141750 266134
rect 163250 266218 163486 266454
rect 163250 265898 163486 266134
rect 169514 266218 169750 266454
rect 169514 265898 169750 266134
rect 191250 266218 191486 266454
rect 191250 265898 191486 266134
rect 200646 269593 200882 269829
rect 200646 269273 200882 269509
rect 216118 269593 216354 269829
rect 216118 269273 216354 269509
rect 222382 269593 222618 269829
rect 222382 269273 222618 269509
rect 228646 269593 228882 269829
rect 228646 269273 228882 269509
rect 244118 269593 244354 269829
rect 244118 269273 244354 269509
rect 250382 269593 250618 269829
rect 250382 269273 250618 269509
rect 256646 269593 256882 269829
rect 256646 269273 256882 269509
rect 272118 269593 272354 269829
rect 272118 269273 272354 269509
rect 197514 266218 197750 266454
rect 197514 265898 197750 266134
rect 219250 266218 219486 266454
rect 219250 265898 219486 266134
rect 225514 266218 225750 266454
rect 225514 265898 225750 266134
rect 247250 266218 247486 266454
rect 247250 265898 247486 266134
rect 253514 266218 253750 266454
rect 253514 265898 253750 266134
rect 275250 266218 275486 266454
rect 275250 265898 275486 266134
rect 278382 269593 278618 269829
rect 278382 269273 278618 269509
rect 284646 269593 284882 269829
rect 284646 269273 284882 269509
rect 300118 269593 300354 269829
rect 300118 269273 300354 269509
rect 306382 269593 306618 269829
rect 306382 269273 306618 269509
rect 312646 269593 312882 269829
rect 312646 269273 312882 269509
rect 328118 269593 328354 269829
rect 328118 269273 328354 269509
rect 334382 269593 334618 269829
rect 334382 269273 334618 269509
rect 340646 269593 340882 269829
rect 340646 269273 340882 269509
rect 356118 269593 356354 269829
rect 356118 269273 356354 269509
rect 362382 269593 362618 269829
rect 362382 269273 362618 269509
rect 368646 269593 368882 269829
rect 368646 269273 368882 269509
rect 384118 269593 384354 269829
rect 384118 269273 384354 269509
rect 390382 269593 390618 269829
rect 390382 269273 390618 269509
rect 281514 266218 281750 266454
rect 281514 265898 281750 266134
rect 303250 266218 303486 266454
rect 303250 265898 303486 266134
rect 309514 266218 309750 266454
rect 309514 265898 309750 266134
rect 331250 266218 331486 266454
rect 331250 265898 331486 266134
rect 337514 266218 337750 266454
rect 337514 265898 337750 266134
rect 359250 266218 359486 266454
rect 359250 265898 359486 266134
rect 365514 266218 365750 266454
rect 365514 265898 365750 266134
rect 387250 266218 387486 266454
rect 387250 265898 387486 266134
rect 396646 269593 396882 269829
rect 396646 269273 396882 269509
rect 412118 269593 412354 269829
rect 412118 269273 412354 269509
rect 418382 269593 418618 269829
rect 418382 269273 418618 269509
rect 424646 269593 424882 269829
rect 424646 269273 424882 269509
rect 440118 269593 440354 269829
rect 440118 269273 440354 269509
rect 446382 269593 446618 269829
rect 446382 269273 446618 269509
rect 452646 269593 452882 269829
rect 452646 269273 452882 269509
rect 468118 269593 468354 269829
rect 468118 269273 468354 269509
rect 393514 266218 393750 266454
rect 393514 265898 393750 266134
rect 415250 266218 415486 266454
rect 415250 265898 415486 266134
rect 421514 266218 421750 266454
rect 421514 265898 421750 266134
rect 443250 266218 443486 266454
rect 443250 265898 443486 266134
rect 449514 266218 449750 266454
rect 449514 265898 449750 266134
rect 471250 266218 471486 266454
rect 471250 265898 471486 266134
rect 474382 269593 474618 269829
rect 474382 269273 474618 269509
rect 480646 269593 480882 269829
rect 480646 269273 480882 269509
rect 496118 269593 496354 269829
rect 496118 269273 496354 269509
rect 502382 269593 502618 269829
rect 502382 269273 502618 269509
rect 508646 269593 508882 269829
rect 508646 269273 508882 269509
rect 477514 266218 477750 266454
rect 477514 265898 477750 266134
rect 499250 266218 499486 266454
rect 499250 265898 499486 266134
rect 505514 266218 505750 266454
rect 505514 265898 505750 266134
rect 524118 269593 524354 269829
rect 524118 269273 524354 269509
rect 530382 269593 530618 269829
rect 530382 269273 530618 269509
rect 536646 269593 536882 269829
rect 536646 269273 536882 269509
rect 552118 269593 552354 269829
rect 552118 269273 552354 269509
rect 558382 269593 558618 269829
rect 558382 269273 558618 269509
rect 564646 269593 564882 269829
rect 564646 269273 564882 269509
rect 573526 269593 573762 269829
rect 573846 269593 574082 269829
rect 573526 269273 573762 269509
rect 573846 269273 574082 269509
rect 527250 266218 527486 266454
rect 527250 265898 527486 266134
rect 533514 266218 533750 266454
rect 533514 265898 533750 266134
rect 555250 266218 555486 266454
rect 555250 265898 555486 266134
rect 561514 266218 561750 266454
rect 561514 265898 561750 266134
rect -1974 242593 -1738 242829
rect -1654 242593 -1418 242829
rect -1974 242273 -1738 242509
rect -1654 242273 -1418 242509
rect 20118 242593 20354 242829
rect 20118 242273 20354 242509
rect 26382 242593 26618 242829
rect 26382 242273 26618 242509
rect 32646 242593 32882 242829
rect 32646 242273 32882 242509
rect 48118 242593 48354 242829
rect 48118 242273 48354 242509
rect 54382 242593 54618 242829
rect 54382 242273 54618 242509
rect 60646 242593 60882 242829
rect 60646 242273 60882 242509
rect 76118 242593 76354 242829
rect 76118 242273 76354 242509
rect 82382 242593 82618 242829
rect 82382 242273 82618 242509
rect 88646 242593 88882 242829
rect 88646 242273 88882 242509
rect 104118 242593 104354 242829
rect 104118 242273 104354 242509
rect 110382 242593 110618 242829
rect 110382 242273 110618 242509
rect 116646 242593 116882 242829
rect 116646 242273 116882 242509
rect 132118 242593 132354 242829
rect 132118 242273 132354 242509
rect 138382 242593 138618 242829
rect 138382 242273 138618 242509
rect 144646 242593 144882 242829
rect 144646 242273 144882 242509
rect 160118 242593 160354 242829
rect 160118 242273 160354 242509
rect 23250 239218 23486 239454
rect 23250 238898 23486 239134
rect 29514 239218 29750 239454
rect 29514 238898 29750 239134
rect 51250 239218 51486 239454
rect 51250 238898 51486 239134
rect 57514 239218 57750 239454
rect 57514 238898 57750 239134
rect 79250 239218 79486 239454
rect 79250 238898 79486 239134
rect 85514 239218 85750 239454
rect 85514 238898 85750 239134
rect 107250 239218 107486 239454
rect 107250 238898 107486 239134
rect 113514 239218 113750 239454
rect 113514 238898 113750 239134
rect 135250 239218 135486 239454
rect 135250 238898 135486 239134
rect 141514 239218 141750 239454
rect 141514 238898 141750 239134
rect 163250 239218 163486 239454
rect 163250 238898 163486 239134
rect 166382 242593 166618 242829
rect 166382 242273 166618 242509
rect 172646 242593 172882 242829
rect 172646 242273 172882 242509
rect 188118 242593 188354 242829
rect 188118 242273 188354 242509
rect 194382 242593 194618 242829
rect 194382 242273 194618 242509
rect 200646 242593 200882 242829
rect 200646 242273 200882 242509
rect 216118 242593 216354 242829
rect 216118 242273 216354 242509
rect 222382 242593 222618 242829
rect 222382 242273 222618 242509
rect 228646 242593 228882 242829
rect 228646 242273 228882 242509
rect 244118 242593 244354 242829
rect 244118 242273 244354 242509
rect 250382 242593 250618 242829
rect 250382 242273 250618 242509
rect 256646 242593 256882 242829
rect 256646 242273 256882 242509
rect 169514 239218 169750 239454
rect 169514 238898 169750 239134
rect 191250 239218 191486 239454
rect 191250 238898 191486 239134
rect 197514 239218 197750 239454
rect 197514 238898 197750 239134
rect 219250 239218 219486 239454
rect 219250 238898 219486 239134
rect 225514 239218 225750 239454
rect 225514 238898 225750 239134
rect 247250 239218 247486 239454
rect 247250 238898 247486 239134
rect 253514 239218 253750 239454
rect 253514 238898 253750 239134
rect 272118 242593 272354 242829
rect 272118 242273 272354 242509
rect 278382 242593 278618 242829
rect 278382 242273 278618 242509
rect 284646 242593 284882 242829
rect 284646 242273 284882 242509
rect 300118 242593 300354 242829
rect 300118 242273 300354 242509
rect 306382 242593 306618 242829
rect 306382 242273 306618 242509
rect 312646 242593 312882 242829
rect 312646 242273 312882 242509
rect 328118 242593 328354 242829
rect 328118 242273 328354 242509
rect 334382 242593 334618 242829
rect 334382 242273 334618 242509
rect 340646 242593 340882 242829
rect 340646 242273 340882 242509
rect 356118 242593 356354 242829
rect 356118 242273 356354 242509
rect 275250 239218 275486 239454
rect 275250 238898 275486 239134
rect 281514 239218 281750 239454
rect 281514 238898 281750 239134
rect 303250 239218 303486 239454
rect 303250 238898 303486 239134
rect 309514 239218 309750 239454
rect 309514 238898 309750 239134
rect 331250 239218 331486 239454
rect 331250 238898 331486 239134
rect 337514 239218 337750 239454
rect 337514 238898 337750 239134
rect 359250 239218 359486 239454
rect 359250 238898 359486 239134
rect 362382 242593 362618 242829
rect 362382 242273 362618 242509
rect 368646 242593 368882 242829
rect 368646 242273 368882 242509
rect 384118 242593 384354 242829
rect 384118 242273 384354 242509
rect 390382 242593 390618 242829
rect 390382 242273 390618 242509
rect 396646 242593 396882 242829
rect 396646 242273 396882 242509
rect 412118 242593 412354 242829
rect 412118 242273 412354 242509
rect 418382 242593 418618 242829
rect 418382 242273 418618 242509
rect 424646 242593 424882 242829
rect 424646 242273 424882 242509
rect 440118 242593 440354 242829
rect 440118 242273 440354 242509
rect 365514 239218 365750 239454
rect 365514 238898 365750 239134
rect 387250 239218 387486 239454
rect 387250 238898 387486 239134
rect 393514 239218 393750 239454
rect 393514 238898 393750 239134
rect 415250 239218 415486 239454
rect 415250 238898 415486 239134
rect 421514 239218 421750 239454
rect 421514 238898 421750 239134
rect 443250 239218 443486 239454
rect 443250 238898 443486 239134
rect 446382 242593 446618 242829
rect 446382 242273 446618 242509
rect 452646 242593 452882 242829
rect 452646 242273 452882 242509
rect 468118 242593 468354 242829
rect 468118 242273 468354 242509
rect 474382 242593 474618 242829
rect 474382 242273 474618 242509
rect 480646 242593 480882 242829
rect 480646 242273 480882 242509
rect 496118 242593 496354 242829
rect 496118 242273 496354 242509
rect 502382 242593 502618 242829
rect 502382 242273 502618 242509
rect 508646 242593 508882 242829
rect 508646 242273 508882 242509
rect 524118 242593 524354 242829
rect 524118 242273 524354 242509
rect 530382 242593 530618 242829
rect 530382 242273 530618 242509
rect 536646 242593 536882 242829
rect 536646 242273 536882 242509
rect 552118 242593 552354 242829
rect 552118 242273 552354 242509
rect 449514 239218 449750 239454
rect 449514 238898 449750 239134
rect 471250 239218 471486 239454
rect 471250 238898 471486 239134
rect 477514 239218 477750 239454
rect 477514 238898 477750 239134
rect 499250 239218 499486 239454
rect 499250 238898 499486 239134
rect 505514 239218 505750 239454
rect 505514 238898 505750 239134
rect 527250 239218 527486 239454
rect 527250 238898 527486 239134
rect 533514 239218 533750 239454
rect 533514 238898 533750 239134
rect 555250 239218 555486 239454
rect 555250 238898 555486 239134
rect 558382 242593 558618 242829
rect 558382 242273 558618 242509
rect 564646 242593 564882 242829
rect 564646 242273 564882 242509
rect 573526 242593 573762 242829
rect 573846 242593 574082 242829
rect 573526 242273 573762 242509
rect 573846 242273 574082 242509
rect 561514 239218 561750 239454
rect 561514 238898 561750 239134
rect -1974 215593 -1738 215829
rect -1654 215593 -1418 215829
rect -1974 215273 -1738 215509
rect -1654 215273 -1418 215509
rect 20118 215593 20354 215829
rect 20118 215273 20354 215509
rect 26382 215593 26618 215829
rect 26382 215273 26618 215509
rect 32646 215593 32882 215829
rect 32646 215273 32882 215509
rect 48118 215593 48354 215829
rect 48118 215273 48354 215509
rect 54382 215593 54618 215829
rect 54382 215273 54618 215509
rect 60646 215593 60882 215829
rect 60646 215273 60882 215509
rect 76118 215593 76354 215829
rect 76118 215273 76354 215509
rect 82382 215593 82618 215829
rect 82382 215273 82618 215509
rect 88646 215593 88882 215829
rect 88646 215273 88882 215509
rect 104118 215593 104354 215829
rect 104118 215273 104354 215509
rect 110382 215593 110618 215829
rect 110382 215273 110618 215509
rect 116646 215593 116882 215829
rect 116646 215273 116882 215509
rect 23250 212218 23486 212454
rect 23250 211898 23486 212134
rect 29514 212218 29750 212454
rect 29514 211898 29750 212134
rect 51250 212218 51486 212454
rect 51250 211898 51486 212134
rect 57514 212218 57750 212454
rect 57514 211898 57750 212134
rect 79250 212218 79486 212454
rect 79250 211898 79486 212134
rect 85514 212218 85750 212454
rect 85514 211898 85750 212134
rect 107250 212218 107486 212454
rect 107250 211898 107486 212134
rect 113514 212218 113750 212454
rect 113514 211898 113750 212134
rect 132118 215593 132354 215829
rect 132118 215273 132354 215509
rect 138382 215593 138618 215829
rect 138382 215273 138618 215509
rect 144646 215593 144882 215829
rect 144646 215273 144882 215509
rect 160118 215593 160354 215829
rect 160118 215273 160354 215509
rect 166382 215593 166618 215829
rect 166382 215273 166618 215509
rect 172646 215593 172882 215829
rect 172646 215273 172882 215509
rect 187335 215593 187571 215829
rect 187335 215273 187571 215509
rect 192033 215593 192269 215829
rect 192033 215273 192269 215509
rect 135250 212218 135486 212454
rect 135250 211898 135486 212134
rect 141514 212218 141750 212454
rect 141514 211898 141750 212134
rect 163250 212218 163486 212454
rect 163250 211898 163486 212134
rect 169514 212218 169750 212454
rect 169514 211898 169750 212134
rect 189684 212218 189920 212454
rect 189684 211898 189920 212134
rect 194382 212218 194618 212454
rect 194382 211898 194618 212134
rect 196731 215593 196967 215829
rect 196731 215273 196967 215509
rect 201429 215593 201665 215829
rect 201429 215273 201665 215509
rect 215335 215593 215571 215829
rect 215335 215273 215571 215509
rect 220033 215593 220269 215829
rect 220033 215273 220269 215509
rect 224731 215593 224967 215829
rect 224731 215273 224967 215509
rect 229429 215593 229665 215829
rect 229429 215273 229665 215509
rect 243335 215593 243571 215829
rect 243335 215273 243571 215509
rect 248033 215593 248269 215829
rect 248033 215273 248269 215509
rect 252731 215593 252967 215829
rect 252731 215273 252967 215509
rect 257429 215593 257665 215829
rect 257429 215273 257665 215509
rect 271335 215593 271571 215829
rect 271335 215273 271571 215509
rect 276033 215593 276269 215829
rect 276033 215273 276269 215509
rect 280731 215593 280967 215829
rect 280731 215273 280967 215509
rect 285429 215593 285665 215829
rect 285429 215273 285665 215509
rect 299335 215593 299571 215829
rect 299335 215273 299571 215509
rect 304033 215593 304269 215829
rect 304033 215273 304269 215509
rect 308731 215593 308967 215829
rect 308731 215273 308967 215509
rect 313429 215593 313665 215829
rect 313429 215273 313665 215509
rect 328118 215593 328354 215829
rect 328118 215273 328354 215509
rect 334382 215593 334618 215829
rect 334382 215273 334618 215509
rect 340646 215593 340882 215829
rect 340646 215273 340882 215509
rect 355335 215593 355571 215829
rect 355335 215273 355571 215509
rect 360033 215593 360269 215829
rect 360033 215273 360269 215509
rect 364731 215593 364967 215829
rect 364731 215273 364967 215509
rect 369429 215593 369665 215829
rect 369429 215273 369665 215509
rect 383335 215593 383571 215829
rect 383335 215273 383571 215509
rect 388033 215593 388269 215829
rect 388033 215273 388269 215509
rect 392731 215593 392967 215829
rect 392731 215273 392967 215509
rect 397429 215593 397665 215829
rect 397429 215273 397665 215509
rect 411335 215593 411571 215829
rect 411335 215273 411571 215509
rect 416033 215593 416269 215829
rect 416033 215273 416269 215509
rect 420731 215593 420967 215829
rect 420731 215273 420967 215509
rect 425429 215593 425665 215829
rect 425429 215273 425665 215509
rect 439335 215593 439571 215829
rect 439335 215273 439571 215509
rect 444033 215593 444269 215829
rect 444033 215273 444269 215509
rect 448731 215593 448967 215829
rect 448731 215273 448967 215509
rect 453429 215593 453665 215829
rect 453429 215273 453665 215509
rect 467335 215593 467571 215829
rect 467335 215273 467571 215509
rect 472033 215593 472269 215829
rect 472033 215273 472269 215509
rect 476731 215593 476967 215829
rect 476731 215273 476967 215509
rect 481429 215593 481665 215829
rect 481429 215273 481665 215509
rect 495335 215593 495571 215829
rect 495335 215273 495571 215509
rect 500033 215593 500269 215829
rect 500033 215273 500269 215509
rect 504731 215593 504967 215829
rect 504731 215273 504967 215509
rect 509429 215593 509665 215829
rect 509429 215273 509665 215509
rect 523335 215593 523571 215829
rect 523335 215273 523571 215509
rect 528033 215593 528269 215829
rect 528033 215273 528269 215509
rect 532731 215593 532967 215829
rect 532731 215273 532967 215509
rect 537429 215593 537665 215829
rect 537429 215273 537665 215509
rect 551335 215593 551571 215829
rect 551335 215273 551571 215509
rect 556033 215593 556269 215829
rect 556033 215273 556269 215509
rect 560731 215593 560967 215829
rect 560731 215273 560967 215509
rect 565429 215593 565665 215829
rect 565429 215273 565665 215509
rect 573526 215593 573762 215829
rect 573846 215593 574082 215829
rect 573526 215273 573762 215509
rect 573846 215273 574082 215509
rect 199080 212218 199316 212454
rect 199080 211898 199316 212134
rect 217684 212218 217920 212454
rect 217684 211898 217920 212134
rect 222382 212218 222618 212454
rect 222382 211898 222618 212134
rect 227080 212218 227316 212454
rect 227080 211898 227316 212134
rect 245684 212218 245920 212454
rect 245684 211898 245920 212134
rect 250382 212218 250618 212454
rect 250382 211898 250618 212134
rect 255080 212218 255316 212454
rect 255080 211898 255316 212134
rect 273684 212218 273920 212454
rect 273684 211898 273920 212134
rect 278382 212218 278618 212454
rect 278382 211898 278618 212134
rect 283080 212218 283316 212454
rect 283080 211898 283316 212134
rect 301684 212218 301920 212454
rect 301684 211898 301920 212134
rect 306382 212218 306618 212454
rect 306382 211898 306618 212134
rect 311080 212218 311316 212454
rect 311080 211898 311316 212134
rect 331250 212218 331486 212454
rect 331250 211898 331486 212134
rect 337514 212218 337750 212454
rect 337514 211898 337750 212134
rect 357684 212218 357920 212454
rect 357684 211898 357920 212134
rect 362382 212218 362618 212454
rect 362382 211898 362618 212134
rect 367080 212218 367316 212454
rect 367080 211898 367316 212134
rect 385684 212218 385920 212454
rect 385684 211898 385920 212134
rect 390382 212218 390618 212454
rect 390382 211898 390618 212134
rect 395080 212218 395316 212454
rect 395080 211898 395316 212134
rect 413684 212218 413920 212454
rect 413684 211898 413920 212134
rect 418382 212218 418618 212454
rect 418382 211898 418618 212134
rect 423080 212218 423316 212454
rect 423080 211898 423316 212134
rect 441684 212218 441920 212454
rect 441684 211898 441920 212134
rect 446382 212218 446618 212454
rect 446382 211898 446618 212134
rect 451080 212218 451316 212454
rect 451080 211898 451316 212134
rect 469684 212218 469920 212454
rect 469684 211898 469920 212134
rect 474382 212218 474618 212454
rect 474382 211898 474618 212134
rect 479080 212218 479316 212454
rect 479080 211898 479316 212134
rect 497684 212218 497920 212454
rect 497684 211898 497920 212134
rect 502382 212218 502618 212454
rect 502382 211898 502618 212134
rect 507080 212218 507316 212454
rect 507080 211898 507316 212134
rect 525684 212218 525920 212454
rect 525684 211898 525920 212134
rect 530382 212218 530618 212454
rect 530382 211898 530618 212134
rect 535080 212218 535316 212454
rect 535080 211898 535316 212134
rect 553684 212218 553920 212454
rect 553684 211898 553920 212134
rect 558382 212218 558618 212454
rect 558382 211898 558618 212134
rect 563080 212218 563316 212454
rect 563080 211898 563316 212134
rect -1974 188593 -1738 188829
rect -1654 188593 -1418 188829
rect -1974 188273 -1738 188509
rect -1654 188273 -1418 188509
rect 19335 188593 19571 188829
rect 19335 188273 19571 188509
rect 24033 188593 24269 188829
rect 24033 188273 24269 188509
rect 28731 188593 28967 188829
rect 28731 188273 28967 188509
rect 33429 188593 33665 188829
rect 33429 188273 33665 188509
rect 47335 188593 47571 188829
rect 47335 188273 47571 188509
rect 52033 188593 52269 188829
rect 52033 188273 52269 188509
rect 56731 188593 56967 188829
rect 56731 188273 56967 188509
rect 61429 188593 61665 188829
rect 61429 188273 61665 188509
rect 21684 185218 21920 185454
rect 21684 184898 21920 185134
rect 26382 185218 26618 185454
rect 26382 184898 26618 185134
rect 31080 185218 31316 185454
rect 31080 184898 31316 185134
rect 49684 185218 49920 185454
rect 49684 184898 49920 185134
rect 54382 185218 54618 185454
rect 54382 184898 54618 185134
rect 59080 185218 59316 185454
rect 59080 184898 59316 185134
rect -1974 161593 -1738 161829
rect -1654 161593 -1418 161829
rect -1974 161273 -1738 161509
rect -1654 161273 -1418 161509
rect 19335 161593 19571 161829
rect 19335 161273 19571 161509
rect 24033 161593 24269 161829
rect 24033 161273 24269 161509
rect 28731 161593 28967 161829
rect 28731 161273 28967 161509
rect 33429 161593 33665 161829
rect 33429 161273 33665 161509
rect 47335 161593 47571 161829
rect 47335 161273 47571 161509
rect 52033 161593 52269 161829
rect 52033 161273 52269 161509
rect 56731 161593 56967 161829
rect 56731 161273 56967 161509
rect 61429 161593 61665 161829
rect 61429 161273 61665 161509
rect 21684 158218 21920 158454
rect 21684 157898 21920 158134
rect 26382 158218 26618 158454
rect 26382 157898 26618 158134
rect 31080 158218 31316 158454
rect 31080 157898 31316 158134
rect 49684 158218 49920 158454
rect 49684 157898 49920 158134
rect 54382 158218 54618 158454
rect 54382 157898 54618 158134
rect 59080 158218 59316 158454
rect 59080 157898 59316 158134
rect -1974 134593 -1738 134829
rect -1654 134593 -1418 134829
rect -1974 134273 -1738 134509
rect -1654 134273 -1418 134509
rect 19335 134593 19571 134829
rect 19335 134273 19571 134509
rect 24033 134593 24269 134829
rect 24033 134273 24269 134509
rect 28731 134593 28967 134829
rect 28731 134273 28967 134509
rect 33429 134593 33665 134829
rect 33429 134273 33665 134509
rect 47335 134593 47571 134829
rect 47335 134273 47571 134509
rect 52033 134593 52269 134829
rect 52033 134273 52269 134509
rect 56731 134593 56967 134829
rect 56731 134273 56967 134509
rect 61429 134593 61665 134829
rect 61429 134273 61665 134509
rect 21684 131218 21920 131454
rect 21684 130898 21920 131134
rect 26382 131218 26618 131454
rect 26382 130898 26618 131134
rect 31080 131218 31316 131454
rect 31080 130898 31316 131134
rect 49684 131218 49920 131454
rect 49684 130898 49920 131134
rect 54382 131218 54618 131454
rect 54382 130898 54618 131134
rect 59080 131218 59316 131454
rect 59080 130898 59316 131134
rect -1974 107593 -1738 107829
rect -1654 107593 -1418 107829
rect -1974 107273 -1738 107509
rect -1654 107273 -1418 107509
rect 19335 107593 19571 107829
rect 19335 107273 19571 107509
rect 24033 107593 24269 107829
rect 24033 107273 24269 107509
rect 28731 107593 28967 107829
rect 28731 107273 28967 107509
rect 33429 107593 33665 107829
rect 33429 107273 33665 107509
rect 47335 107593 47571 107829
rect 47335 107273 47571 107509
rect 52033 107593 52269 107829
rect 52033 107273 52269 107509
rect 56731 107593 56967 107829
rect 56731 107273 56967 107509
rect 61429 107593 61665 107829
rect 61429 107273 61665 107509
rect 21684 104218 21920 104454
rect 21684 103898 21920 104134
rect 26382 104218 26618 104454
rect 26382 103898 26618 104134
rect 31080 104218 31316 104454
rect 31080 103898 31316 104134
rect 49684 104218 49920 104454
rect 49684 103898 49920 104134
rect 54382 104218 54618 104454
rect 54382 103898 54618 104134
rect 59080 104218 59316 104454
rect 59080 103898 59316 104134
rect -1974 80593 -1738 80829
rect -1654 80593 -1418 80829
rect -1974 80273 -1738 80509
rect -1654 80273 -1418 80509
rect 20118 80593 20354 80829
rect 20118 80273 20354 80509
rect 26382 80593 26618 80829
rect 26382 80273 26618 80509
rect 32646 80593 32882 80829
rect 32646 80273 32882 80509
rect 48118 80593 48354 80829
rect 48118 80273 48354 80509
rect 54382 80593 54618 80829
rect 54382 80273 54618 80509
rect 60646 80593 60882 80829
rect 60646 80273 60882 80509
rect 23250 77218 23486 77454
rect 23250 76898 23486 77134
rect 29514 77218 29750 77454
rect 29514 76898 29750 77134
rect 51250 77218 51486 77454
rect 51250 76898 51486 77134
rect 57514 77218 57750 77454
rect 57514 76898 57750 77134
rect -1974 53593 -1738 53829
rect -1654 53593 -1418 53829
rect -1974 53273 -1738 53509
rect -1654 53273 -1418 53509
rect 20118 53593 20354 53829
rect 20118 53273 20354 53509
rect 26382 53593 26618 53829
rect 26382 53273 26618 53509
rect 32646 53593 32882 53829
rect 32646 53273 32882 53509
rect 48118 53593 48354 53829
rect 48118 53273 48354 53509
rect 54382 53593 54618 53829
rect 54382 53273 54618 53509
rect 60646 53593 60882 53829
rect 60646 53273 60882 53509
rect 23250 50218 23486 50454
rect 23250 49898 23486 50134
rect 29514 50218 29750 50454
rect 29514 49898 29750 50134
rect 51250 50218 51486 50454
rect 51250 49898 51486 50134
rect 57514 50218 57750 50454
rect 57514 49898 57750 50134
rect -1974 26593 -1738 26829
rect -1654 26593 -1418 26829
rect -1974 26273 -1738 26509
rect -1654 26273 -1418 26509
rect 22460 26593 22696 26829
rect 22460 26273 22696 26509
rect 33408 26593 33644 26829
rect 33408 26273 33644 26509
rect 44356 26593 44592 26829
rect 44356 26273 44592 26509
rect 55304 26593 55540 26829
rect 55304 26273 55540 26509
rect 27934 23218 28170 23454
rect 27934 22898 28170 23134
rect 38882 23218 39118 23454
rect 38882 22898 39118 23134
rect 49830 23218 50066 23454
rect 49830 22898 50066 23134
rect 60778 23218 61014 23454
rect 60778 22898 61014 23134
rect 75335 188593 75571 188829
rect 75335 188273 75571 188509
rect 80033 188593 80269 188829
rect 80033 188273 80269 188509
rect 84731 188593 84967 188829
rect 84731 188273 84967 188509
rect 89429 188593 89665 188829
rect 89429 188273 89665 188509
rect 103335 188593 103571 188829
rect 103335 188273 103571 188509
rect 108033 188593 108269 188829
rect 108033 188273 108269 188509
rect 112731 188593 112967 188829
rect 112731 188273 112967 188509
rect 117429 188593 117665 188829
rect 117429 188273 117665 188509
rect 131335 188593 131571 188829
rect 131335 188273 131571 188509
rect 136033 188593 136269 188829
rect 136033 188273 136269 188509
rect 140731 188593 140967 188829
rect 140731 188273 140967 188509
rect 145429 188593 145665 188829
rect 145429 188273 145665 188509
rect 159335 188593 159571 188829
rect 159335 188273 159571 188509
rect 164033 188593 164269 188829
rect 164033 188273 164269 188509
rect 168731 188593 168967 188829
rect 168731 188273 168967 188509
rect 173429 188593 173665 188829
rect 173429 188273 173665 188509
rect 187335 188593 187571 188829
rect 187335 188273 187571 188509
rect 192033 188593 192269 188829
rect 192033 188273 192269 188509
rect 196731 188593 196967 188829
rect 196731 188273 196967 188509
rect 201429 188593 201665 188829
rect 201429 188273 201665 188509
rect 215335 188593 215571 188829
rect 215335 188273 215571 188509
rect 220033 188593 220269 188829
rect 220033 188273 220269 188509
rect 224731 188593 224967 188829
rect 224731 188273 224967 188509
rect 229429 188593 229665 188829
rect 229429 188273 229665 188509
rect 243335 188593 243571 188829
rect 243335 188273 243571 188509
rect 248033 188593 248269 188829
rect 248033 188273 248269 188509
rect 252731 188593 252967 188829
rect 252731 188273 252967 188509
rect 257429 188593 257665 188829
rect 257429 188273 257665 188509
rect 77684 185218 77920 185454
rect 77684 184898 77920 185134
rect 82382 185218 82618 185454
rect 82382 184898 82618 185134
rect 87080 185218 87316 185454
rect 87080 184898 87316 185134
rect 105684 185218 105920 185454
rect 105684 184898 105920 185134
rect 110382 185218 110618 185454
rect 110382 184898 110618 185134
rect 115080 185218 115316 185454
rect 115080 184898 115316 185134
rect 133684 185218 133920 185454
rect 133684 184898 133920 185134
rect 138382 185218 138618 185454
rect 138382 184898 138618 185134
rect 143080 185218 143316 185454
rect 143080 184898 143316 185134
rect 161684 185218 161920 185454
rect 161684 184898 161920 185134
rect 166382 185218 166618 185454
rect 166382 184898 166618 185134
rect 171080 185218 171316 185454
rect 171080 184898 171316 185134
rect 189684 185218 189920 185454
rect 189684 184898 189920 185134
rect 194382 185218 194618 185454
rect 194382 184898 194618 185134
rect 199080 185218 199316 185454
rect 199080 184898 199316 185134
rect 217684 185218 217920 185454
rect 217684 184898 217920 185134
rect 222382 185218 222618 185454
rect 222382 184898 222618 185134
rect 227080 185218 227316 185454
rect 227080 184898 227316 185134
rect 245684 185218 245920 185454
rect 245684 184898 245920 185134
rect 250382 185218 250618 185454
rect 250382 184898 250618 185134
rect 255080 185218 255316 185454
rect 255080 184898 255316 185134
rect 271335 188593 271571 188829
rect 271335 188273 271571 188509
rect 276033 188593 276269 188829
rect 276033 188273 276269 188509
rect 280731 188593 280967 188829
rect 280731 188273 280967 188509
rect 285429 188593 285665 188829
rect 285429 188273 285665 188509
rect 299335 188593 299571 188829
rect 299335 188273 299571 188509
rect 304033 188593 304269 188829
rect 304033 188273 304269 188509
rect 308731 188593 308967 188829
rect 308731 188273 308967 188509
rect 313429 188593 313665 188829
rect 313429 188273 313665 188509
rect 327335 188593 327571 188829
rect 327335 188273 327571 188509
rect 332033 188593 332269 188829
rect 332033 188273 332269 188509
rect 336731 188593 336967 188829
rect 336731 188273 336967 188509
rect 341429 188593 341665 188829
rect 341429 188273 341665 188509
rect 355335 188593 355571 188829
rect 355335 188273 355571 188509
rect 360033 188593 360269 188829
rect 360033 188273 360269 188509
rect 273684 185218 273920 185454
rect 273684 184898 273920 185134
rect 278382 185218 278618 185454
rect 278382 184898 278618 185134
rect 283080 185218 283316 185454
rect 283080 184898 283316 185134
rect 301684 185218 301920 185454
rect 301684 184898 301920 185134
rect 306382 185218 306618 185454
rect 306382 184898 306618 185134
rect 311080 185218 311316 185454
rect 311080 184898 311316 185134
rect 329684 185218 329920 185454
rect 329684 184898 329920 185134
rect 334382 185218 334618 185454
rect 334382 184898 334618 185134
rect 339080 185218 339316 185454
rect 339080 184898 339316 185134
rect 357684 185218 357920 185454
rect 357684 184898 357920 185134
rect 364731 188593 364967 188829
rect 364731 188273 364967 188509
rect 369429 188593 369665 188829
rect 369429 188273 369665 188509
rect 383335 188593 383571 188829
rect 383335 188273 383571 188509
rect 388033 188593 388269 188829
rect 388033 188273 388269 188509
rect 392731 188593 392967 188829
rect 392731 188273 392967 188509
rect 397429 188593 397665 188829
rect 397429 188273 397665 188509
rect 411335 188593 411571 188829
rect 411335 188273 411571 188509
rect 416033 188593 416269 188829
rect 416033 188273 416269 188509
rect 420731 188593 420967 188829
rect 420731 188273 420967 188509
rect 425429 188593 425665 188829
rect 425429 188273 425665 188509
rect 439335 188593 439571 188829
rect 439335 188273 439571 188509
rect 444033 188593 444269 188829
rect 444033 188273 444269 188509
rect 362382 185218 362618 185454
rect 362382 184898 362618 185134
rect 367080 185218 367316 185454
rect 367080 184898 367316 185134
rect 385684 185218 385920 185454
rect 385684 184898 385920 185134
rect 390382 185218 390618 185454
rect 390382 184898 390618 185134
rect 395080 185218 395316 185454
rect 395080 184898 395316 185134
rect 413684 185218 413920 185454
rect 413684 184898 413920 185134
rect 418382 185218 418618 185454
rect 418382 184898 418618 185134
rect 423080 185218 423316 185454
rect 423080 184898 423316 185134
rect 441684 185218 441920 185454
rect 441684 184898 441920 185134
rect 448731 188593 448967 188829
rect 448731 188273 448967 188509
rect 453429 188593 453665 188829
rect 453429 188273 453665 188509
rect 467335 188593 467571 188829
rect 467335 188273 467571 188509
rect 472033 188593 472269 188829
rect 472033 188273 472269 188509
rect 476731 188593 476967 188829
rect 476731 188273 476967 188509
rect 481429 188593 481665 188829
rect 481429 188273 481665 188509
rect 495335 188593 495571 188829
rect 495335 188273 495571 188509
rect 500033 188593 500269 188829
rect 500033 188273 500269 188509
rect 504731 188593 504967 188829
rect 504731 188273 504967 188509
rect 509429 188593 509665 188829
rect 509429 188273 509665 188509
rect 523335 188593 523571 188829
rect 523335 188273 523571 188509
rect 528033 188593 528269 188829
rect 528033 188273 528269 188509
rect 532731 188593 532967 188829
rect 532731 188273 532967 188509
rect 537429 188593 537665 188829
rect 537429 188273 537665 188509
rect 551335 188593 551571 188829
rect 551335 188273 551571 188509
rect 556033 188593 556269 188829
rect 556033 188273 556269 188509
rect 560731 188593 560967 188829
rect 560731 188273 560967 188509
rect 565429 188593 565665 188829
rect 565429 188273 565665 188509
rect 573526 188593 573762 188829
rect 573846 188593 574082 188829
rect 573526 188273 573762 188509
rect 573846 188273 574082 188509
rect 446382 185218 446618 185454
rect 446382 184898 446618 185134
rect 451080 185218 451316 185454
rect 451080 184898 451316 185134
rect 469684 185218 469920 185454
rect 469684 184898 469920 185134
rect 474382 185218 474618 185454
rect 474382 184898 474618 185134
rect 479080 185218 479316 185454
rect 479080 184898 479316 185134
rect 497684 185218 497920 185454
rect 497684 184898 497920 185134
rect 502382 185218 502618 185454
rect 502382 184898 502618 185134
rect 507080 185218 507316 185454
rect 507080 184898 507316 185134
rect 525684 185218 525920 185454
rect 525684 184898 525920 185134
rect 530382 185218 530618 185454
rect 530382 184898 530618 185134
rect 535080 185218 535316 185454
rect 535080 184898 535316 185134
rect 553684 185218 553920 185454
rect 553684 184898 553920 185134
rect 558382 185218 558618 185454
rect 558382 184898 558618 185134
rect 563080 185218 563316 185454
rect 563080 184898 563316 185134
rect 75335 161593 75571 161829
rect 75335 161273 75571 161509
rect 80033 161593 80269 161829
rect 80033 161273 80269 161509
rect 84731 161593 84967 161829
rect 84731 161273 84967 161509
rect 89429 161593 89665 161829
rect 89429 161273 89665 161509
rect 103335 161593 103571 161829
rect 103335 161273 103571 161509
rect 108033 161593 108269 161829
rect 108033 161273 108269 161509
rect 112731 161593 112967 161829
rect 112731 161273 112967 161509
rect 117429 161593 117665 161829
rect 117429 161273 117665 161509
rect 131335 161593 131571 161829
rect 131335 161273 131571 161509
rect 136033 161593 136269 161829
rect 136033 161273 136269 161509
rect 140731 161593 140967 161829
rect 140731 161273 140967 161509
rect 145429 161593 145665 161829
rect 145429 161273 145665 161509
rect 159335 161593 159571 161829
rect 159335 161273 159571 161509
rect 164033 161593 164269 161829
rect 164033 161273 164269 161509
rect 168731 161593 168967 161829
rect 168731 161273 168967 161509
rect 173429 161593 173665 161829
rect 173429 161273 173665 161509
rect 187335 161593 187571 161829
rect 187335 161273 187571 161509
rect 192033 161593 192269 161829
rect 192033 161273 192269 161509
rect 196731 161593 196967 161829
rect 196731 161273 196967 161509
rect 201429 161593 201665 161829
rect 201429 161273 201665 161509
rect 215335 161593 215571 161829
rect 215335 161273 215571 161509
rect 220033 161593 220269 161829
rect 220033 161273 220269 161509
rect 224731 161593 224967 161829
rect 224731 161273 224967 161509
rect 229429 161593 229665 161829
rect 229429 161273 229665 161509
rect 243335 161593 243571 161829
rect 243335 161273 243571 161509
rect 248033 161593 248269 161829
rect 248033 161273 248269 161509
rect 252731 161593 252967 161829
rect 252731 161273 252967 161509
rect 257429 161593 257665 161829
rect 257429 161273 257665 161509
rect 271335 161593 271571 161829
rect 271335 161273 271571 161509
rect 276033 161593 276269 161829
rect 276033 161273 276269 161509
rect 280731 161593 280967 161829
rect 280731 161273 280967 161509
rect 285429 161593 285665 161829
rect 285429 161273 285665 161509
rect 299335 161593 299571 161829
rect 299335 161273 299571 161509
rect 304033 161593 304269 161829
rect 304033 161273 304269 161509
rect 308731 161593 308967 161829
rect 308731 161273 308967 161509
rect 313429 161593 313665 161829
rect 313429 161273 313665 161509
rect 327335 161593 327571 161829
rect 327335 161273 327571 161509
rect 332033 161593 332269 161829
rect 332033 161273 332269 161509
rect 336731 161593 336967 161829
rect 336731 161273 336967 161509
rect 341429 161593 341665 161829
rect 341429 161273 341665 161509
rect 355335 161593 355571 161829
rect 355335 161273 355571 161509
rect 360033 161593 360269 161829
rect 360033 161273 360269 161509
rect 364731 161593 364967 161829
rect 364731 161273 364967 161509
rect 369429 161593 369665 161829
rect 369429 161273 369665 161509
rect 383335 161593 383571 161829
rect 383335 161273 383571 161509
rect 388033 161593 388269 161829
rect 388033 161273 388269 161509
rect 392731 161593 392967 161829
rect 392731 161273 392967 161509
rect 397429 161593 397665 161829
rect 397429 161273 397665 161509
rect 411335 161593 411571 161829
rect 411335 161273 411571 161509
rect 416033 161593 416269 161829
rect 416033 161273 416269 161509
rect 420731 161593 420967 161829
rect 420731 161273 420967 161509
rect 425429 161593 425665 161829
rect 425429 161273 425665 161509
rect 439335 161593 439571 161829
rect 439335 161273 439571 161509
rect 444033 161593 444269 161829
rect 444033 161273 444269 161509
rect 448731 161593 448967 161829
rect 448731 161273 448967 161509
rect 453429 161593 453665 161829
rect 453429 161273 453665 161509
rect 467335 161593 467571 161829
rect 467335 161273 467571 161509
rect 472033 161593 472269 161829
rect 472033 161273 472269 161509
rect 476731 161593 476967 161829
rect 476731 161273 476967 161509
rect 481429 161593 481665 161829
rect 481429 161273 481665 161509
rect 495335 161593 495571 161829
rect 495335 161273 495571 161509
rect 500033 161593 500269 161829
rect 500033 161273 500269 161509
rect 504731 161593 504967 161829
rect 504731 161273 504967 161509
rect 509429 161593 509665 161829
rect 509429 161273 509665 161509
rect 523335 161593 523571 161829
rect 523335 161273 523571 161509
rect 528033 161593 528269 161829
rect 528033 161273 528269 161509
rect 532731 161593 532967 161829
rect 532731 161273 532967 161509
rect 537429 161593 537665 161829
rect 537429 161273 537665 161509
rect 551335 161593 551571 161829
rect 551335 161273 551571 161509
rect 556033 161593 556269 161829
rect 556033 161273 556269 161509
rect 560731 161593 560967 161829
rect 560731 161273 560967 161509
rect 565429 161593 565665 161829
rect 565429 161273 565665 161509
rect 573526 161593 573762 161829
rect 573846 161593 574082 161829
rect 573526 161273 573762 161509
rect 573846 161273 574082 161509
rect 77684 158218 77920 158454
rect 77684 157898 77920 158134
rect 82382 158218 82618 158454
rect 82382 157898 82618 158134
rect 87080 158218 87316 158454
rect 87080 157898 87316 158134
rect 105684 158218 105920 158454
rect 105684 157898 105920 158134
rect 110382 158218 110618 158454
rect 110382 157898 110618 158134
rect 115080 158218 115316 158454
rect 115080 157898 115316 158134
rect 133684 158218 133920 158454
rect 133684 157898 133920 158134
rect 138382 158218 138618 158454
rect 138382 157898 138618 158134
rect 143080 158218 143316 158454
rect 143080 157898 143316 158134
rect 161684 158218 161920 158454
rect 161684 157898 161920 158134
rect 166382 158218 166618 158454
rect 166382 157898 166618 158134
rect 171080 158218 171316 158454
rect 171080 157898 171316 158134
rect 189684 158218 189920 158454
rect 189684 157898 189920 158134
rect 194382 158218 194618 158454
rect 194382 157898 194618 158134
rect 199080 158218 199316 158454
rect 199080 157898 199316 158134
rect 217684 158218 217920 158454
rect 217684 157898 217920 158134
rect 222382 158218 222618 158454
rect 222382 157898 222618 158134
rect 227080 158218 227316 158454
rect 227080 157898 227316 158134
rect 245684 158218 245920 158454
rect 245684 157898 245920 158134
rect 250382 158218 250618 158454
rect 250382 157898 250618 158134
rect 255080 158218 255316 158454
rect 255080 157898 255316 158134
rect 273684 158218 273920 158454
rect 273684 157898 273920 158134
rect 278382 158218 278618 158454
rect 278382 157898 278618 158134
rect 283080 158218 283316 158454
rect 283080 157898 283316 158134
rect 301684 158218 301920 158454
rect 301684 157898 301920 158134
rect 306382 158218 306618 158454
rect 306382 157898 306618 158134
rect 311080 158218 311316 158454
rect 311080 157898 311316 158134
rect 329684 158218 329920 158454
rect 329684 157898 329920 158134
rect 334382 158218 334618 158454
rect 334382 157898 334618 158134
rect 339080 158218 339316 158454
rect 339080 157898 339316 158134
rect 357684 158218 357920 158454
rect 357684 157898 357920 158134
rect 362382 158218 362618 158454
rect 362382 157898 362618 158134
rect 367080 158218 367316 158454
rect 367080 157898 367316 158134
rect 385684 158218 385920 158454
rect 385684 157898 385920 158134
rect 390382 158218 390618 158454
rect 390382 157898 390618 158134
rect 395080 158218 395316 158454
rect 395080 157898 395316 158134
rect 413684 158218 413920 158454
rect 413684 157898 413920 158134
rect 418382 158218 418618 158454
rect 418382 157898 418618 158134
rect 423080 158218 423316 158454
rect 423080 157898 423316 158134
rect 441684 158218 441920 158454
rect 441684 157898 441920 158134
rect 446382 158218 446618 158454
rect 446382 157898 446618 158134
rect 451080 158218 451316 158454
rect 451080 157898 451316 158134
rect 469684 158218 469920 158454
rect 469684 157898 469920 158134
rect 474382 158218 474618 158454
rect 474382 157898 474618 158134
rect 479080 158218 479316 158454
rect 479080 157898 479316 158134
rect 497684 158218 497920 158454
rect 497684 157898 497920 158134
rect 502382 158218 502618 158454
rect 502382 157898 502618 158134
rect 507080 158218 507316 158454
rect 507080 157898 507316 158134
rect 525684 158218 525920 158454
rect 525684 157898 525920 158134
rect 530382 158218 530618 158454
rect 530382 157898 530618 158134
rect 535080 158218 535316 158454
rect 535080 157898 535316 158134
rect 553684 158218 553920 158454
rect 553684 157898 553920 158134
rect 558382 158218 558618 158454
rect 558382 157898 558618 158134
rect 563080 158218 563316 158454
rect 563080 157898 563316 158134
rect 75335 134593 75571 134829
rect 75335 134273 75571 134509
rect 80033 134593 80269 134829
rect 80033 134273 80269 134509
rect 84731 134593 84967 134829
rect 84731 134273 84967 134509
rect 89429 134593 89665 134829
rect 89429 134273 89665 134509
rect 103335 134593 103571 134829
rect 103335 134273 103571 134509
rect 108033 134593 108269 134829
rect 108033 134273 108269 134509
rect 112731 134593 112967 134829
rect 112731 134273 112967 134509
rect 117429 134593 117665 134829
rect 117429 134273 117665 134509
rect 131335 134593 131571 134829
rect 131335 134273 131571 134509
rect 136033 134593 136269 134829
rect 136033 134273 136269 134509
rect 140731 134593 140967 134829
rect 140731 134273 140967 134509
rect 145429 134593 145665 134829
rect 145429 134273 145665 134509
rect 159335 134593 159571 134829
rect 159335 134273 159571 134509
rect 164033 134593 164269 134829
rect 164033 134273 164269 134509
rect 168731 134593 168967 134829
rect 168731 134273 168967 134509
rect 173429 134593 173665 134829
rect 173429 134273 173665 134509
rect 187335 134593 187571 134829
rect 187335 134273 187571 134509
rect 192033 134593 192269 134829
rect 192033 134273 192269 134509
rect 196731 134593 196967 134829
rect 196731 134273 196967 134509
rect 201429 134593 201665 134829
rect 201429 134273 201665 134509
rect 215335 134593 215571 134829
rect 215335 134273 215571 134509
rect 220033 134593 220269 134829
rect 220033 134273 220269 134509
rect 224731 134593 224967 134829
rect 224731 134273 224967 134509
rect 229429 134593 229665 134829
rect 229429 134273 229665 134509
rect 243335 134593 243571 134829
rect 243335 134273 243571 134509
rect 248033 134593 248269 134829
rect 248033 134273 248269 134509
rect 252731 134593 252967 134829
rect 252731 134273 252967 134509
rect 257429 134593 257665 134829
rect 257429 134273 257665 134509
rect 271335 134593 271571 134829
rect 271335 134273 271571 134509
rect 276033 134593 276269 134829
rect 276033 134273 276269 134509
rect 280731 134593 280967 134829
rect 280731 134273 280967 134509
rect 285429 134593 285665 134829
rect 285429 134273 285665 134509
rect 299335 134593 299571 134829
rect 299335 134273 299571 134509
rect 304033 134593 304269 134829
rect 304033 134273 304269 134509
rect 308731 134593 308967 134829
rect 308731 134273 308967 134509
rect 313429 134593 313665 134829
rect 313429 134273 313665 134509
rect 327335 134593 327571 134829
rect 327335 134273 327571 134509
rect 332033 134593 332269 134829
rect 332033 134273 332269 134509
rect 336731 134593 336967 134829
rect 336731 134273 336967 134509
rect 341429 134593 341665 134829
rect 341429 134273 341665 134509
rect 355335 134593 355571 134829
rect 355335 134273 355571 134509
rect 360033 134593 360269 134829
rect 360033 134273 360269 134509
rect 77684 131218 77920 131454
rect 77684 130898 77920 131134
rect 82382 131218 82618 131454
rect 82382 130898 82618 131134
rect 87080 131218 87316 131454
rect 87080 130898 87316 131134
rect 105684 131218 105920 131454
rect 105684 130898 105920 131134
rect 110382 131218 110618 131454
rect 110382 130898 110618 131134
rect 115080 131218 115316 131454
rect 115080 130898 115316 131134
rect 133684 131218 133920 131454
rect 133684 130898 133920 131134
rect 138382 131218 138618 131454
rect 138382 130898 138618 131134
rect 143080 131218 143316 131454
rect 143080 130898 143316 131134
rect 161684 131218 161920 131454
rect 161684 130898 161920 131134
rect 166382 131218 166618 131454
rect 166382 130898 166618 131134
rect 171080 131218 171316 131454
rect 171080 130898 171316 131134
rect 189684 131218 189920 131454
rect 189684 130898 189920 131134
rect 194382 131218 194618 131454
rect 194382 130898 194618 131134
rect 199080 131218 199316 131454
rect 199080 130898 199316 131134
rect 217684 131218 217920 131454
rect 217684 130898 217920 131134
rect 222382 131218 222618 131454
rect 222382 130898 222618 131134
rect 227080 131218 227316 131454
rect 227080 130898 227316 131134
rect 245684 131218 245920 131454
rect 245684 130898 245920 131134
rect 250382 131218 250618 131454
rect 250382 130898 250618 131134
rect 255080 131218 255316 131454
rect 255080 130898 255316 131134
rect 273684 131218 273920 131454
rect 273684 130898 273920 131134
rect 278382 131218 278618 131454
rect 278382 130898 278618 131134
rect 283080 131218 283316 131454
rect 283080 130898 283316 131134
rect 301684 131218 301920 131454
rect 301684 130898 301920 131134
rect 306382 131218 306618 131454
rect 306382 130898 306618 131134
rect 311080 131218 311316 131454
rect 311080 130898 311316 131134
rect 329684 131218 329920 131454
rect 329684 130898 329920 131134
rect 334382 131218 334618 131454
rect 334382 130898 334618 131134
rect 339080 131218 339316 131454
rect 339080 130898 339316 131134
rect 357684 131218 357920 131454
rect 357684 130898 357920 131134
rect 364731 134593 364967 134829
rect 364731 134273 364967 134509
rect 369429 134593 369665 134829
rect 369429 134273 369665 134509
rect 383335 134593 383571 134829
rect 383335 134273 383571 134509
rect 388033 134593 388269 134829
rect 388033 134273 388269 134509
rect 392731 134593 392967 134829
rect 392731 134273 392967 134509
rect 397429 134593 397665 134829
rect 397429 134273 397665 134509
rect 411335 134593 411571 134829
rect 411335 134273 411571 134509
rect 416033 134593 416269 134829
rect 416033 134273 416269 134509
rect 420731 134593 420967 134829
rect 420731 134273 420967 134509
rect 425429 134593 425665 134829
rect 425429 134273 425665 134509
rect 439335 134593 439571 134829
rect 439335 134273 439571 134509
rect 444033 134593 444269 134829
rect 444033 134273 444269 134509
rect 362382 131218 362618 131454
rect 362382 130898 362618 131134
rect 367080 131218 367316 131454
rect 367080 130898 367316 131134
rect 385684 131218 385920 131454
rect 385684 130898 385920 131134
rect 390382 131218 390618 131454
rect 390382 130898 390618 131134
rect 395080 131218 395316 131454
rect 395080 130898 395316 131134
rect 413684 131218 413920 131454
rect 413684 130898 413920 131134
rect 418382 131218 418618 131454
rect 418382 130898 418618 131134
rect 423080 131218 423316 131454
rect 423080 130898 423316 131134
rect 441684 131218 441920 131454
rect 441684 130898 441920 131134
rect 448731 134593 448967 134829
rect 448731 134273 448967 134509
rect 453429 134593 453665 134829
rect 453429 134273 453665 134509
rect 467335 134593 467571 134829
rect 467335 134273 467571 134509
rect 472033 134593 472269 134829
rect 472033 134273 472269 134509
rect 476731 134593 476967 134829
rect 476731 134273 476967 134509
rect 481429 134593 481665 134829
rect 481429 134273 481665 134509
rect 495335 134593 495571 134829
rect 495335 134273 495571 134509
rect 500033 134593 500269 134829
rect 500033 134273 500269 134509
rect 504731 134593 504967 134829
rect 504731 134273 504967 134509
rect 509429 134593 509665 134829
rect 509429 134273 509665 134509
rect 523335 134593 523571 134829
rect 523335 134273 523571 134509
rect 528033 134593 528269 134829
rect 528033 134273 528269 134509
rect 532731 134593 532967 134829
rect 532731 134273 532967 134509
rect 537429 134593 537665 134829
rect 537429 134273 537665 134509
rect 551335 134593 551571 134829
rect 551335 134273 551571 134509
rect 556033 134593 556269 134829
rect 556033 134273 556269 134509
rect 560731 134593 560967 134829
rect 560731 134273 560967 134509
rect 565429 134593 565665 134829
rect 565429 134273 565665 134509
rect 573526 134593 573762 134829
rect 573846 134593 574082 134829
rect 573526 134273 573762 134509
rect 573846 134273 574082 134509
rect 446382 131218 446618 131454
rect 446382 130898 446618 131134
rect 451080 131218 451316 131454
rect 451080 130898 451316 131134
rect 469684 131218 469920 131454
rect 469684 130898 469920 131134
rect 474382 131218 474618 131454
rect 474382 130898 474618 131134
rect 479080 131218 479316 131454
rect 479080 130898 479316 131134
rect 497684 131218 497920 131454
rect 497684 130898 497920 131134
rect 502382 131218 502618 131454
rect 502382 130898 502618 131134
rect 507080 131218 507316 131454
rect 507080 130898 507316 131134
rect 525684 131218 525920 131454
rect 525684 130898 525920 131134
rect 530382 131218 530618 131454
rect 530382 130898 530618 131134
rect 535080 131218 535316 131454
rect 535080 130898 535316 131134
rect 553684 131218 553920 131454
rect 553684 130898 553920 131134
rect 558382 131218 558618 131454
rect 558382 130898 558618 131134
rect 563080 131218 563316 131454
rect 563080 130898 563316 131134
rect 75335 107593 75571 107829
rect 75335 107273 75571 107509
rect 80033 107593 80269 107829
rect 80033 107273 80269 107509
rect 84731 107593 84967 107829
rect 84731 107273 84967 107509
rect 89429 107593 89665 107829
rect 89429 107273 89665 107509
rect 103335 107593 103571 107829
rect 103335 107273 103571 107509
rect 108033 107593 108269 107829
rect 108033 107273 108269 107509
rect 112731 107593 112967 107829
rect 112731 107273 112967 107509
rect 117429 107593 117665 107829
rect 117429 107273 117665 107509
rect 131335 107593 131571 107829
rect 131335 107273 131571 107509
rect 136033 107593 136269 107829
rect 136033 107273 136269 107509
rect 140731 107593 140967 107829
rect 140731 107273 140967 107509
rect 145429 107593 145665 107829
rect 145429 107273 145665 107509
rect 159335 107593 159571 107829
rect 159335 107273 159571 107509
rect 164033 107593 164269 107829
rect 164033 107273 164269 107509
rect 168731 107593 168967 107829
rect 168731 107273 168967 107509
rect 173429 107593 173665 107829
rect 173429 107273 173665 107509
rect 187335 107593 187571 107829
rect 187335 107273 187571 107509
rect 192033 107593 192269 107829
rect 192033 107273 192269 107509
rect 77684 104218 77920 104454
rect 77684 103898 77920 104134
rect 82382 104218 82618 104454
rect 82382 103898 82618 104134
rect 87080 104218 87316 104454
rect 87080 103898 87316 104134
rect 105684 104218 105920 104454
rect 105684 103898 105920 104134
rect 110382 104218 110618 104454
rect 110382 103898 110618 104134
rect 115080 104218 115316 104454
rect 115080 103898 115316 104134
rect 133684 104218 133920 104454
rect 133684 103898 133920 104134
rect 138382 104218 138618 104454
rect 138382 103898 138618 104134
rect 143080 104218 143316 104454
rect 143080 103898 143316 104134
rect 161684 104218 161920 104454
rect 161684 103898 161920 104134
rect 166382 104218 166618 104454
rect 166382 103898 166618 104134
rect 171080 104218 171316 104454
rect 171080 103898 171316 104134
rect 189684 104218 189920 104454
rect 189684 103898 189920 104134
rect 194382 104218 194618 104454
rect 194382 103898 194618 104134
rect 196731 107593 196967 107829
rect 196731 107273 196967 107509
rect 201429 107593 201665 107829
rect 201429 107273 201665 107509
rect 215335 107593 215571 107829
rect 215335 107273 215571 107509
rect 220033 107593 220269 107829
rect 220033 107273 220269 107509
rect 224731 107593 224967 107829
rect 224731 107273 224967 107509
rect 229429 107593 229665 107829
rect 229429 107273 229665 107509
rect 244118 107593 244354 107829
rect 244118 107273 244354 107509
rect 250382 107593 250618 107829
rect 250382 107273 250618 107509
rect 256646 107593 256882 107829
rect 256646 107273 256882 107509
rect 271335 107593 271571 107829
rect 271335 107273 271571 107509
rect 276033 107593 276269 107829
rect 276033 107273 276269 107509
rect 280731 107593 280967 107829
rect 280731 107273 280967 107509
rect 285429 107593 285665 107829
rect 285429 107273 285665 107509
rect 299335 107593 299571 107829
rect 299335 107273 299571 107509
rect 304033 107593 304269 107829
rect 304033 107273 304269 107509
rect 308731 107593 308967 107829
rect 308731 107273 308967 107509
rect 313429 107593 313665 107829
rect 313429 107273 313665 107509
rect 199080 104218 199316 104454
rect 199080 103898 199316 104134
rect 217684 104218 217920 104454
rect 217684 103898 217920 104134
rect 222382 104218 222618 104454
rect 222382 103898 222618 104134
rect 227080 104218 227316 104454
rect 227080 103898 227316 104134
rect 247250 104218 247486 104454
rect 247250 103898 247486 104134
rect 253514 104218 253750 104454
rect 253514 103898 253750 104134
rect 273684 104218 273920 104454
rect 273684 103898 273920 104134
rect 278382 104218 278618 104454
rect 278382 103898 278618 104134
rect 283080 104218 283316 104454
rect 283080 103898 283316 104134
rect 301684 104218 301920 104454
rect 301684 103898 301920 104134
rect 306382 104218 306618 104454
rect 306382 103898 306618 104134
rect 311080 104218 311316 104454
rect 311080 103898 311316 104134
rect 328118 107593 328354 107829
rect 328118 107273 328354 107509
rect 334382 107593 334618 107829
rect 334382 107273 334618 107509
rect 340646 107593 340882 107829
rect 340646 107273 340882 107509
rect 355335 107593 355571 107829
rect 355335 107273 355571 107509
rect 360033 107593 360269 107829
rect 360033 107273 360269 107509
rect 364731 107593 364967 107829
rect 364731 107273 364967 107509
rect 369429 107593 369665 107829
rect 369429 107273 369665 107509
rect 383335 107593 383571 107829
rect 383335 107273 383571 107509
rect 388033 107593 388269 107829
rect 388033 107273 388269 107509
rect 392731 107593 392967 107829
rect 392731 107273 392967 107509
rect 397429 107593 397665 107829
rect 397429 107273 397665 107509
rect 411335 107593 411571 107829
rect 411335 107273 411571 107509
rect 416033 107593 416269 107829
rect 416033 107273 416269 107509
rect 420731 107593 420967 107829
rect 420731 107273 420967 107509
rect 425429 107593 425665 107829
rect 425429 107273 425665 107509
rect 439335 107593 439571 107829
rect 439335 107273 439571 107509
rect 444033 107593 444269 107829
rect 444033 107273 444269 107509
rect 448731 107593 448967 107829
rect 448731 107273 448967 107509
rect 453429 107593 453665 107829
rect 453429 107273 453665 107509
rect 467335 107593 467571 107829
rect 467335 107273 467571 107509
rect 472033 107593 472269 107829
rect 472033 107273 472269 107509
rect 476731 107593 476967 107829
rect 476731 107273 476967 107509
rect 481429 107593 481665 107829
rect 481429 107273 481665 107509
rect 495335 107593 495571 107829
rect 495335 107273 495571 107509
rect 500033 107593 500269 107829
rect 500033 107273 500269 107509
rect 504731 107593 504967 107829
rect 504731 107273 504967 107509
rect 509429 107593 509665 107829
rect 509429 107273 509665 107509
rect 523335 107593 523571 107829
rect 523335 107273 523571 107509
rect 528033 107593 528269 107829
rect 528033 107273 528269 107509
rect 532731 107593 532967 107829
rect 532731 107273 532967 107509
rect 537429 107593 537665 107829
rect 537429 107273 537665 107509
rect 551335 107593 551571 107829
rect 551335 107273 551571 107509
rect 556033 107593 556269 107829
rect 556033 107273 556269 107509
rect 560731 107593 560967 107829
rect 560731 107273 560967 107509
rect 565429 107593 565665 107829
rect 565429 107273 565665 107509
rect 573526 107593 573762 107829
rect 573846 107593 574082 107829
rect 573526 107273 573762 107509
rect 573846 107273 574082 107509
rect 331250 104218 331486 104454
rect 331250 103898 331486 104134
rect 337514 104218 337750 104454
rect 337514 103898 337750 104134
rect 357684 104218 357920 104454
rect 357684 103898 357920 104134
rect 362382 104218 362618 104454
rect 362382 103898 362618 104134
rect 367080 104218 367316 104454
rect 367080 103898 367316 104134
rect 385684 104218 385920 104454
rect 385684 103898 385920 104134
rect 390382 104218 390618 104454
rect 390382 103898 390618 104134
rect 395080 104218 395316 104454
rect 395080 103898 395316 104134
rect 413684 104218 413920 104454
rect 413684 103898 413920 104134
rect 418382 104218 418618 104454
rect 418382 103898 418618 104134
rect 423080 104218 423316 104454
rect 423080 103898 423316 104134
rect 441684 104218 441920 104454
rect 441684 103898 441920 104134
rect 446382 104218 446618 104454
rect 446382 103898 446618 104134
rect 451080 104218 451316 104454
rect 451080 103898 451316 104134
rect 469684 104218 469920 104454
rect 469684 103898 469920 104134
rect 474382 104218 474618 104454
rect 474382 103898 474618 104134
rect 479080 104218 479316 104454
rect 479080 103898 479316 104134
rect 497684 104218 497920 104454
rect 497684 103898 497920 104134
rect 502382 104218 502618 104454
rect 502382 103898 502618 104134
rect 507080 104218 507316 104454
rect 507080 103898 507316 104134
rect 525684 104218 525920 104454
rect 525684 103898 525920 104134
rect 530382 104218 530618 104454
rect 530382 103898 530618 104134
rect 535080 104218 535316 104454
rect 535080 103898 535316 104134
rect 553684 104218 553920 104454
rect 553684 103898 553920 104134
rect 558382 104218 558618 104454
rect 558382 103898 558618 104134
rect 563080 104218 563316 104454
rect 563080 103898 563316 104134
rect 76118 80593 76354 80829
rect 76118 80273 76354 80509
rect 82382 80593 82618 80829
rect 82382 80273 82618 80509
rect 88646 80593 88882 80829
rect 88646 80273 88882 80509
rect 103335 80593 103571 80829
rect 103335 80273 103571 80509
rect 108033 80593 108269 80829
rect 108033 80273 108269 80509
rect 112731 80593 112967 80829
rect 112731 80273 112967 80509
rect 117429 80593 117665 80829
rect 117429 80273 117665 80509
rect 131335 80593 131571 80829
rect 131335 80273 131571 80509
rect 136033 80593 136269 80829
rect 136033 80273 136269 80509
rect 140731 80593 140967 80829
rect 140731 80273 140967 80509
rect 145429 80593 145665 80829
rect 145429 80273 145665 80509
rect 159335 80593 159571 80829
rect 159335 80273 159571 80509
rect 164033 80593 164269 80829
rect 164033 80273 164269 80509
rect 168731 80593 168967 80829
rect 168731 80273 168967 80509
rect 173429 80593 173665 80829
rect 173429 80273 173665 80509
rect 188118 80593 188354 80829
rect 188118 80273 188354 80509
rect 194382 80593 194618 80829
rect 194382 80273 194618 80509
rect 200646 80593 200882 80829
rect 200646 80273 200882 80509
rect 216118 80593 216354 80829
rect 216118 80273 216354 80509
rect 222382 80593 222618 80829
rect 222382 80273 222618 80509
rect 228646 80593 228882 80829
rect 228646 80273 228882 80509
rect 244118 80593 244354 80829
rect 244118 80273 244354 80509
rect 250382 80593 250618 80829
rect 250382 80273 250618 80509
rect 256646 80593 256882 80829
rect 256646 80273 256882 80509
rect 272118 80593 272354 80829
rect 272118 80273 272354 80509
rect 278382 80593 278618 80829
rect 278382 80273 278618 80509
rect 284646 80593 284882 80829
rect 284646 80273 284882 80509
rect 300118 80593 300354 80829
rect 300118 80273 300354 80509
rect 306382 80593 306618 80829
rect 306382 80273 306618 80509
rect 312646 80593 312882 80829
rect 312646 80273 312882 80509
rect 328118 80593 328354 80829
rect 328118 80273 328354 80509
rect 334382 80593 334618 80829
rect 334382 80273 334618 80509
rect 340646 80593 340882 80829
rect 340646 80273 340882 80509
rect 355335 80593 355571 80829
rect 355335 80273 355571 80509
rect 360033 80593 360269 80829
rect 360033 80273 360269 80509
rect 364731 80593 364967 80829
rect 364731 80273 364967 80509
rect 369429 80593 369665 80829
rect 369429 80273 369665 80509
rect 383335 80593 383571 80829
rect 383335 80273 383571 80509
rect 388033 80593 388269 80829
rect 388033 80273 388269 80509
rect 392731 80593 392967 80829
rect 392731 80273 392967 80509
rect 397429 80593 397665 80829
rect 397429 80273 397665 80509
rect 411335 80593 411571 80829
rect 411335 80273 411571 80509
rect 416033 80593 416269 80829
rect 416033 80273 416269 80509
rect 420731 80593 420967 80829
rect 420731 80273 420967 80509
rect 425429 80593 425665 80829
rect 425429 80273 425665 80509
rect 439335 80593 439571 80829
rect 439335 80273 439571 80509
rect 444033 80593 444269 80829
rect 444033 80273 444269 80509
rect 448731 80593 448967 80829
rect 448731 80273 448967 80509
rect 453429 80593 453665 80829
rect 453429 80273 453665 80509
rect 467335 80593 467571 80829
rect 467335 80273 467571 80509
rect 472033 80593 472269 80829
rect 472033 80273 472269 80509
rect 476731 80593 476967 80829
rect 476731 80273 476967 80509
rect 481429 80593 481665 80829
rect 481429 80273 481665 80509
rect 495335 80593 495571 80829
rect 495335 80273 495571 80509
rect 500033 80593 500269 80829
rect 500033 80273 500269 80509
rect 504731 80593 504967 80829
rect 504731 80273 504967 80509
rect 509429 80593 509665 80829
rect 509429 80273 509665 80509
rect 523335 80593 523571 80829
rect 523335 80273 523571 80509
rect 528033 80593 528269 80829
rect 528033 80273 528269 80509
rect 532731 80593 532967 80829
rect 532731 80273 532967 80509
rect 537429 80593 537665 80829
rect 537429 80273 537665 80509
rect 551335 80593 551571 80829
rect 551335 80273 551571 80509
rect 556033 80593 556269 80829
rect 556033 80273 556269 80509
rect 560731 80593 560967 80829
rect 560731 80273 560967 80509
rect 565429 80593 565665 80829
rect 565429 80273 565665 80509
rect 573526 80593 573762 80829
rect 573846 80593 574082 80829
rect 573526 80273 573762 80509
rect 573846 80273 574082 80509
rect 79250 77218 79486 77454
rect 79250 76898 79486 77134
rect 85514 77218 85750 77454
rect 85514 76898 85750 77134
rect 105684 77218 105920 77454
rect 105684 76898 105920 77134
rect 110382 77218 110618 77454
rect 110382 76898 110618 77134
rect 115080 77218 115316 77454
rect 115080 76898 115316 77134
rect 133684 77218 133920 77454
rect 133684 76898 133920 77134
rect 138382 77218 138618 77454
rect 138382 76898 138618 77134
rect 143080 77218 143316 77454
rect 143080 76898 143316 77134
rect 161684 77218 161920 77454
rect 161684 76898 161920 77134
rect 166382 77218 166618 77454
rect 166382 76898 166618 77134
rect 171080 77218 171316 77454
rect 171080 76898 171316 77134
rect 191250 77218 191486 77454
rect 191250 76898 191486 77134
rect 197514 77218 197750 77454
rect 197514 76898 197750 77134
rect 219250 77218 219486 77454
rect 219250 76898 219486 77134
rect 225514 77218 225750 77454
rect 225514 76898 225750 77134
rect 247250 77218 247486 77454
rect 247250 76898 247486 77134
rect 253514 77218 253750 77454
rect 253514 76898 253750 77134
rect 275250 77218 275486 77454
rect 275250 76898 275486 77134
rect 281514 77218 281750 77454
rect 281514 76898 281750 77134
rect 303250 77218 303486 77454
rect 303250 76898 303486 77134
rect 309514 77218 309750 77454
rect 309514 76898 309750 77134
rect 331250 77218 331486 77454
rect 331250 76898 331486 77134
rect 337514 77218 337750 77454
rect 337514 76898 337750 77134
rect 357684 77218 357920 77454
rect 357684 76898 357920 77134
rect 362382 77218 362618 77454
rect 362382 76898 362618 77134
rect 367080 77218 367316 77454
rect 367080 76898 367316 77134
rect 385684 77218 385920 77454
rect 385684 76898 385920 77134
rect 390382 77218 390618 77454
rect 390382 76898 390618 77134
rect 395080 77218 395316 77454
rect 395080 76898 395316 77134
rect 413684 77218 413920 77454
rect 413684 76898 413920 77134
rect 418382 77218 418618 77454
rect 418382 76898 418618 77134
rect 423080 77218 423316 77454
rect 423080 76898 423316 77134
rect 441684 77218 441920 77454
rect 441684 76898 441920 77134
rect 446382 77218 446618 77454
rect 446382 76898 446618 77134
rect 451080 77218 451316 77454
rect 451080 76898 451316 77134
rect 469684 77218 469920 77454
rect 469684 76898 469920 77134
rect 474382 77218 474618 77454
rect 474382 76898 474618 77134
rect 479080 77218 479316 77454
rect 479080 76898 479316 77134
rect 497684 77218 497920 77454
rect 497684 76898 497920 77134
rect 502382 77218 502618 77454
rect 502382 76898 502618 77134
rect 507080 77218 507316 77454
rect 507080 76898 507316 77134
rect 525684 77218 525920 77454
rect 525684 76898 525920 77134
rect 530382 77218 530618 77454
rect 530382 76898 530618 77134
rect 535080 77218 535316 77454
rect 535080 76898 535316 77134
rect 553684 77218 553920 77454
rect 553684 76898 553920 77134
rect 558382 77218 558618 77454
rect 558382 76898 558618 77134
rect 563080 77218 563316 77454
rect 563080 76898 563316 77134
rect 76118 53593 76354 53829
rect 76118 53273 76354 53509
rect 82382 53593 82618 53829
rect 82382 53273 82618 53509
rect 88646 53593 88882 53829
rect 88646 53273 88882 53509
rect 104118 53593 104354 53829
rect 104118 53273 104354 53509
rect 110382 53593 110618 53829
rect 110382 53273 110618 53509
rect 116646 53593 116882 53829
rect 116646 53273 116882 53509
rect 132118 53593 132354 53829
rect 132118 53273 132354 53509
rect 138382 53593 138618 53829
rect 138382 53273 138618 53509
rect 144646 53593 144882 53829
rect 144646 53273 144882 53509
rect 160118 53593 160354 53829
rect 160118 53273 160354 53509
rect 166382 53593 166618 53829
rect 166382 53273 166618 53509
rect 172646 53593 172882 53829
rect 172646 53273 172882 53509
rect 188118 53593 188354 53829
rect 188118 53273 188354 53509
rect 194382 53593 194618 53829
rect 194382 53273 194618 53509
rect 200646 53593 200882 53829
rect 200646 53273 200882 53509
rect 215335 53593 215571 53829
rect 215335 53273 215571 53509
rect 220033 53593 220269 53829
rect 220033 53273 220269 53509
rect 224731 53593 224967 53829
rect 224731 53273 224967 53509
rect 229429 53593 229665 53829
rect 229429 53273 229665 53509
rect 244118 53593 244354 53829
rect 244118 53273 244354 53509
rect 250382 53593 250618 53829
rect 250382 53273 250618 53509
rect 256646 53593 256882 53829
rect 256646 53273 256882 53509
rect 272118 53593 272354 53829
rect 272118 53273 272354 53509
rect 278382 53593 278618 53829
rect 278382 53273 278618 53509
rect 284646 53593 284882 53829
rect 284646 53273 284882 53509
rect 300118 53593 300354 53829
rect 300118 53273 300354 53509
rect 306382 53593 306618 53829
rect 306382 53273 306618 53509
rect 312646 53593 312882 53829
rect 312646 53273 312882 53509
rect 327335 53593 327571 53829
rect 327335 53273 327571 53509
rect 332033 53593 332269 53829
rect 332033 53273 332269 53509
rect 336731 53593 336967 53829
rect 336731 53273 336967 53509
rect 341429 53593 341665 53829
rect 341429 53273 341665 53509
rect 356118 53593 356354 53829
rect 356118 53273 356354 53509
rect 362382 53593 362618 53829
rect 362382 53273 362618 53509
rect 368646 53593 368882 53829
rect 368646 53273 368882 53509
rect 384118 53593 384354 53829
rect 384118 53273 384354 53509
rect 390382 53593 390618 53829
rect 390382 53273 390618 53509
rect 396646 53593 396882 53829
rect 396646 53273 396882 53509
rect 412118 53593 412354 53829
rect 412118 53273 412354 53509
rect 418382 53593 418618 53829
rect 418382 53273 418618 53509
rect 424646 53593 424882 53829
rect 424646 53273 424882 53509
rect 440118 53593 440354 53829
rect 440118 53273 440354 53509
rect 446382 53593 446618 53829
rect 446382 53273 446618 53509
rect 452646 53593 452882 53829
rect 452646 53273 452882 53509
rect 468118 53593 468354 53829
rect 468118 53273 468354 53509
rect 474382 53593 474618 53829
rect 474382 53273 474618 53509
rect 480646 53593 480882 53829
rect 480646 53273 480882 53509
rect 495335 53593 495571 53829
rect 495335 53273 495571 53509
rect 500033 53593 500269 53829
rect 500033 53273 500269 53509
rect 504731 53593 504967 53829
rect 504731 53273 504967 53509
rect 509429 53593 509665 53829
rect 509429 53273 509665 53509
rect 524118 53593 524354 53829
rect 524118 53273 524354 53509
rect 530382 53593 530618 53829
rect 530382 53273 530618 53509
rect 536646 53593 536882 53829
rect 536646 53273 536882 53509
rect 552118 53593 552354 53829
rect 552118 53273 552354 53509
rect 558382 53593 558618 53829
rect 558382 53273 558618 53509
rect 564646 53593 564882 53829
rect 564646 53273 564882 53509
rect 573526 53593 573762 53829
rect 573846 53593 574082 53829
rect 573526 53273 573762 53509
rect 573846 53273 574082 53509
rect 79250 50218 79486 50454
rect 79250 49898 79486 50134
rect 85514 50218 85750 50454
rect 85514 49898 85750 50134
rect 107250 50218 107486 50454
rect 107250 49898 107486 50134
rect 113514 50218 113750 50454
rect 113514 49898 113750 50134
rect 135250 50218 135486 50454
rect 135250 49898 135486 50134
rect 141514 50218 141750 50454
rect 141514 49898 141750 50134
rect 163250 50218 163486 50454
rect 163250 49898 163486 50134
rect 169514 50218 169750 50454
rect 169514 49898 169750 50134
rect 191250 50218 191486 50454
rect 191250 49898 191486 50134
rect 197514 50218 197750 50454
rect 197514 49898 197750 50134
rect 217684 50218 217920 50454
rect 217684 49898 217920 50134
rect 222382 50218 222618 50454
rect 222382 49898 222618 50134
rect 227080 50218 227316 50454
rect 227080 49898 227316 50134
rect 247250 50218 247486 50454
rect 247250 49898 247486 50134
rect 253514 50218 253750 50454
rect 253514 49898 253750 50134
rect 275250 50218 275486 50454
rect 275250 49898 275486 50134
rect 281514 50218 281750 50454
rect 281514 49898 281750 50134
rect 303250 50218 303486 50454
rect 303250 49898 303486 50134
rect 309514 50218 309750 50454
rect 309514 49898 309750 50134
rect 329684 50218 329920 50454
rect 329684 49898 329920 50134
rect 334382 50218 334618 50454
rect 334382 49898 334618 50134
rect 339080 50218 339316 50454
rect 339080 49898 339316 50134
rect 359250 50218 359486 50454
rect 359250 49898 359486 50134
rect 365514 50218 365750 50454
rect 365514 49898 365750 50134
rect 387250 50218 387486 50454
rect 387250 49898 387486 50134
rect 393514 50218 393750 50454
rect 393514 49898 393750 50134
rect 415250 50218 415486 50454
rect 415250 49898 415486 50134
rect 421514 50218 421750 50454
rect 421514 49898 421750 50134
rect 443250 50218 443486 50454
rect 443250 49898 443486 50134
rect 449514 50218 449750 50454
rect 449514 49898 449750 50134
rect 471250 50218 471486 50454
rect 471250 49898 471486 50134
rect 477514 50218 477750 50454
rect 477514 49898 477750 50134
rect 497684 50218 497920 50454
rect 497684 49898 497920 50134
rect 502382 50218 502618 50454
rect 502382 49898 502618 50134
rect 507080 50218 507316 50454
rect 507080 49898 507316 50134
rect 527250 50218 527486 50454
rect 527250 49898 527486 50134
rect 533514 50218 533750 50454
rect 533514 49898 533750 50134
rect 555250 50218 555486 50454
rect 555250 49898 555486 50134
rect 561514 50218 561750 50454
rect 561514 49898 561750 50134
rect 76118 26593 76354 26829
rect 76118 26273 76354 26509
rect 82382 26593 82618 26829
rect 82382 26273 82618 26509
rect 88646 26593 88882 26829
rect 88646 26273 88882 26509
rect 104118 26593 104354 26829
rect 104118 26273 104354 26509
rect 110382 26593 110618 26829
rect 110382 26273 110618 26509
rect 116646 26593 116882 26829
rect 116646 26273 116882 26509
rect 132118 26593 132354 26829
rect 132118 26273 132354 26509
rect 138382 26593 138618 26829
rect 138382 26273 138618 26509
rect 144646 26593 144882 26829
rect 144646 26273 144882 26509
rect 160118 26593 160354 26829
rect 160118 26273 160354 26509
rect 166382 26593 166618 26829
rect 166382 26273 166618 26509
rect 172646 26593 172882 26829
rect 172646 26273 172882 26509
rect 188118 26593 188354 26829
rect 188118 26273 188354 26509
rect 194382 26593 194618 26829
rect 194382 26273 194618 26509
rect 200646 26593 200882 26829
rect 200646 26273 200882 26509
rect 216118 26593 216354 26829
rect 216118 26273 216354 26509
rect 222382 26593 222618 26829
rect 222382 26273 222618 26509
rect 228646 26593 228882 26829
rect 228646 26273 228882 26509
rect 244118 26593 244354 26829
rect 244118 26273 244354 26509
rect 66026 23218 66262 23454
rect 66346 23218 66582 23454
rect 66026 22898 66262 23134
rect 66346 22898 66582 23134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 79250 23218 79486 23454
rect 79250 22898 79486 23134
rect 85514 23218 85750 23454
rect 85514 22898 85750 23134
rect 107250 23218 107486 23454
rect 107250 22898 107486 23134
rect 113514 23218 113750 23454
rect 113514 22898 113750 23134
rect 135250 23218 135486 23454
rect 135250 22898 135486 23134
rect 141514 23218 141750 23454
rect 141514 22898 141750 23134
rect 163250 23218 163486 23454
rect 163250 22898 163486 23134
rect 169514 23218 169750 23454
rect 169514 22898 169750 23134
rect 191250 23218 191486 23454
rect 191250 22898 191486 23134
rect 197514 23218 197750 23454
rect 197514 22898 197750 23134
rect 219250 23218 219486 23454
rect 219250 22898 219486 23134
rect 225514 23218 225750 23454
rect 225514 22898 225750 23134
rect 247250 23218 247486 23454
rect 247250 22898 247486 23134
rect 250382 26593 250618 26829
rect 250382 26273 250618 26509
rect 256646 26593 256882 26829
rect 256646 26273 256882 26509
rect 272118 26593 272354 26829
rect 272118 26273 272354 26509
rect 278382 26593 278618 26829
rect 278382 26273 278618 26509
rect 284646 26593 284882 26829
rect 284646 26273 284882 26509
rect 300118 26593 300354 26829
rect 300118 26273 300354 26509
rect 306382 26593 306618 26829
rect 306382 26273 306618 26509
rect 312646 26593 312882 26829
rect 312646 26273 312882 26509
rect 328118 26593 328354 26829
rect 328118 26273 328354 26509
rect 334382 26593 334618 26829
rect 334382 26273 334618 26509
rect 340646 26593 340882 26829
rect 340646 26273 340882 26509
rect 355335 26593 355571 26829
rect 355335 26273 355571 26509
rect 360033 26593 360269 26829
rect 360033 26273 360269 26509
rect 364731 26593 364967 26829
rect 364731 26273 364967 26509
rect 369429 26593 369665 26829
rect 369429 26273 369665 26509
rect 384118 26593 384354 26829
rect 384118 26273 384354 26509
rect 390382 26593 390618 26829
rect 390382 26273 390618 26509
rect 396646 26593 396882 26829
rect 396646 26273 396882 26509
rect 412118 26593 412354 26829
rect 412118 26273 412354 26509
rect 418382 26593 418618 26829
rect 418382 26273 418618 26509
rect 424646 26593 424882 26829
rect 424646 26273 424882 26509
rect 440118 26593 440354 26829
rect 440118 26273 440354 26509
rect 446382 26593 446618 26829
rect 446382 26273 446618 26509
rect 452646 26593 452882 26829
rect 452646 26273 452882 26509
rect 253514 23218 253750 23454
rect 253514 22898 253750 23134
rect 275250 23218 275486 23454
rect 275250 22898 275486 23134
rect 281514 23218 281750 23454
rect 281514 22898 281750 23134
rect 303250 23218 303486 23454
rect 303250 22898 303486 23134
rect 309514 23218 309750 23454
rect 309514 22898 309750 23134
rect 331250 23218 331486 23454
rect 331250 22898 331486 23134
rect 337514 23218 337750 23454
rect 337514 22898 337750 23134
rect 357684 23218 357920 23454
rect 357684 22898 357920 23134
rect 362382 23218 362618 23454
rect 362382 22898 362618 23134
rect 367080 23218 367316 23454
rect 367080 22898 367316 23134
rect 387250 23218 387486 23454
rect 387250 22898 387486 23134
rect 393514 23218 393750 23454
rect 393514 22898 393750 23134
rect 415250 23218 415486 23454
rect 415250 22898 415486 23134
rect 421514 23218 421750 23454
rect 421514 22898 421750 23134
rect 443250 23218 443486 23454
rect 443250 22898 443486 23134
rect 449514 23218 449750 23454
rect 449514 22898 449750 23134
rect 468118 26593 468354 26829
rect 468118 26273 468354 26509
rect 474382 26593 474618 26829
rect 474382 26273 474618 26509
rect 480646 26593 480882 26829
rect 480646 26273 480882 26509
rect 496118 26593 496354 26829
rect 496118 26273 496354 26509
rect 502382 26593 502618 26829
rect 502382 26273 502618 26509
rect 508646 26593 508882 26829
rect 508646 26273 508882 26509
rect 524118 26593 524354 26829
rect 524118 26273 524354 26509
rect 530382 26593 530618 26829
rect 530382 26273 530618 26509
rect 536646 26593 536882 26829
rect 536646 26273 536882 26509
rect 552118 26593 552354 26829
rect 552118 26273 552354 26509
rect 471250 23218 471486 23454
rect 471250 22898 471486 23134
rect 477514 23218 477750 23454
rect 477514 22898 477750 23134
rect 499250 23218 499486 23454
rect 499250 22898 499486 23134
rect 505514 23218 505750 23454
rect 505514 22898 505750 23134
rect 527250 23218 527486 23454
rect 527250 22898 527486 23134
rect 533514 23218 533750 23454
rect 533514 22898 533750 23134
rect 555250 23218 555486 23454
rect 555250 22898 555486 23134
rect 558382 26593 558618 26829
rect 558382 26273 558618 26509
rect 564646 26593 564882 26829
rect 564646 26273 564882 26509
rect 585342 674593 585578 674829
rect 585662 674593 585898 674829
rect 585342 674273 585578 674509
rect 585662 674273 585898 674509
rect 573526 26593 573762 26829
rect 573846 26593 574082 26829
rect 573526 26273 573762 26509
rect 573846 26273 574082 26509
rect 561514 23218 561750 23454
rect 561514 22898 561750 23134
rect 66026 -1542 66262 -1306
rect 66346 -1542 66582 -1306
rect 66026 -1862 66262 -1626
rect 66346 -1862 66582 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 585342 647593 585578 647829
rect 585662 647593 585898 647829
rect 585342 647273 585578 647509
rect 585662 647273 585898 647509
rect 585342 620593 585578 620829
rect 585662 620593 585898 620829
rect 585342 620273 585578 620509
rect 585662 620273 585898 620509
rect 585342 593593 585578 593829
rect 585662 593593 585898 593829
rect 585342 593273 585578 593509
rect 585662 593273 585898 593509
rect 585342 566593 585578 566829
rect 585662 566593 585898 566829
rect 585342 566273 585578 566509
rect 585662 566273 585898 566509
rect 585342 539593 585578 539829
rect 585662 539593 585898 539829
rect 585342 539273 585578 539509
rect 585662 539273 585898 539509
rect 585342 512593 585578 512829
rect 585662 512593 585898 512829
rect 585342 512273 585578 512509
rect 585662 512273 585898 512509
rect 585342 485593 585578 485829
rect 585662 485593 585898 485829
rect 585342 485273 585578 485509
rect 585662 485273 585898 485509
rect 585342 458593 585578 458829
rect 585662 458593 585898 458829
rect 585342 458273 585578 458509
rect 585662 458273 585898 458509
rect 585342 431593 585578 431829
rect 585662 431593 585898 431829
rect 585342 431273 585578 431509
rect 585662 431273 585898 431509
rect 585342 404593 585578 404829
rect 585662 404593 585898 404829
rect 585342 404273 585578 404509
rect 585662 404273 585898 404509
rect 585342 377593 585578 377829
rect 585662 377593 585898 377829
rect 585342 377273 585578 377509
rect 585662 377273 585898 377509
rect 585342 350593 585578 350829
rect 585662 350593 585898 350829
rect 585342 350273 585578 350509
rect 585662 350273 585898 350509
rect 585342 323593 585578 323829
rect 585662 323593 585898 323829
rect 585342 323273 585578 323509
rect 585662 323273 585898 323509
rect 585342 296593 585578 296829
rect 585662 296593 585898 296829
rect 585342 296273 585578 296509
rect 585662 296273 585898 296509
rect 585342 269593 585578 269829
rect 585662 269593 585898 269829
rect 585342 269273 585578 269509
rect 585662 269273 585898 269509
rect 585342 242593 585578 242829
rect 585662 242593 585898 242829
rect 585342 242273 585578 242509
rect 585662 242273 585898 242509
rect 585342 215593 585578 215829
rect 585662 215593 585898 215829
rect 585342 215273 585578 215509
rect 585662 215273 585898 215509
rect 585342 188593 585578 188829
rect 585662 188593 585898 188829
rect 585342 188273 585578 188509
rect 585662 188273 585898 188509
rect 585342 161593 585578 161829
rect 585662 161593 585898 161829
rect 585342 161273 585578 161509
rect 585662 161273 585898 161509
rect 585342 134593 585578 134829
rect 585662 134593 585898 134829
rect 585342 134273 585578 134509
rect 585662 134273 585898 134509
rect 585342 107593 585578 107829
rect 585662 107593 585898 107829
rect 585342 107273 585578 107509
rect 585662 107273 585898 107509
rect 585342 80593 585578 80829
rect 585662 80593 585898 80829
rect 585342 80273 585578 80509
rect 585662 80273 585898 80509
rect 585342 53593 585578 53829
rect 585662 53593 585898 53829
rect 585342 53273 585578 53509
rect 585662 53273 585898 53509
rect 585342 26593 585578 26829
rect 585662 26593 585898 26829
rect 585342 26273 585578 26509
rect 585662 26273 585898 26509
rect 573526 -582 573762 -346
rect 573846 -582 574082 -346
rect 573526 -902 573762 -666
rect 573846 -902 574082 -666
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 698218 586538 698454
rect 586622 698218 586858 698454
rect 586302 697898 586538 698134
rect 586622 697898 586858 698134
rect 586302 671218 586538 671454
rect 586622 671218 586858 671454
rect 586302 670898 586538 671134
rect 586622 670898 586858 671134
rect 586302 644218 586538 644454
rect 586622 644218 586858 644454
rect 586302 643898 586538 644134
rect 586622 643898 586858 644134
rect 586302 617218 586538 617454
rect 586622 617218 586858 617454
rect 586302 616898 586538 617134
rect 586622 616898 586858 617134
rect 586302 590218 586538 590454
rect 586622 590218 586858 590454
rect 586302 589898 586538 590134
rect 586622 589898 586858 590134
rect 586302 563218 586538 563454
rect 586622 563218 586858 563454
rect 586302 562898 586538 563134
rect 586622 562898 586858 563134
rect 586302 536218 586538 536454
rect 586622 536218 586858 536454
rect 586302 535898 586538 536134
rect 586622 535898 586858 536134
rect 586302 509218 586538 509454
rect 586622 509218 586858 509454
rect 586302 508898 586538 509134
rect 586622 508898 586858 509134
rect 586302 482218 586538 482454
rect 586622 482218 586858 482454
rect 586302 481898 586538 482134
rect 586622 481898 586858 482134
rect 586302 455218 586538 455454
rect 586622 455218 586858 455454
rect 586302 454898 586538 455134
rect 586622 454898 586858 455134
rect 586302 428218 586538 428454
rect 586622 428218 586858 428454
rect 586302 427898 586538 428134
rect 586622 427898 586858 428134
rect 586302 401218 586538 401454
rect 586622 401218 586858 401454
rect 586302 400898 586538 401134
rect 586622 400898 586858 401134
rect 586302 374218 586538 374454
rect 586622 374218 586858 374454
rect 586302 373898 586538 374134
rect 586622 373898 586858 374134
rect 586302 347218 586538 347454
rect 586622 347218 586858 347454
rect 586302 346898 586538 347134
rect 586622 346898 586858 347134
rect 586302 320218 586538 320454
rect 586622 320218 586858 320454
rect 586302 319898 586538 320134
rect 586622 319898 586858 320134
rect 586302 293218 586538 293454
rect 586622 293218 586858 293454
rect 586302 292898 586538 293134
rect 586622 292898 586858 293134
rect 586302 266218 586538 266454
rect 586622 266218 586858 266454
rect 586302 265898 586538 266134
rect 586622 265898 586858 266134
rect 586302 239218 586538 239454
rect 586622 239218 586858 239454
rect 586302 238898 586538 239134
rect 586622 238898 586858 239134
rect 586302 212218 586538 212454
rect 586622 212218 586858 212454
rect 586302 211898 586538 212134
rect 586622 211898 586858 212134
rect 586302 185218 586538 185454
rect 586622 185218 586858 185454
rect 586302 184898 586538 185134
rect 586622 184898 586858 185134
rect 586302 158218 586538 158454
rect 586622 158218 586858 158454
rect 586302 157898 586538 158134
rect 586622 157898 586858 158134
rect 586302 131218 586538 131454
rect 586622 131218 586858 131454
rect 586302 130898 586538 131134
rect 586622 130898 586858 131134
rect 586302 104218 586538 104454
rect 586622 104218 586858 104454
rect 586302 103898 586538 104134
rect 586622 103898 586858 104134
rect 586302 77218 586538 77454
rect 586622 77218 586858 77454
rect 586302 76898 586538 77134
rect 586622 76898 586858 77134
rect 586302 50218 586538 50454
rect 586622 50218 586858 50454
rect 586302 49898 586538 50134
rect 586622 49898 586858 50134
rect 586302 23218 586538 23454
rect 586622 23218 586858 23454
rect 586302 22898 586538 23134
rect 586622 22898 586858 23134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 38026 705798
rect 38262 705562 38346 705798
rect 38582 705562 66026 705798
rect 66262 705562 66346 705798
rect 66582 705562 94026 705798
rect 94262 705562 94346 705798
rect 94582 705562 122026 705798
rect 122262 705562 122346 705798
rect 122582 705562 150026 705798
rect 150262 705562 150346 705798
rect 150582 705562 178026 705798
rect 178262 705562 178346 705798
rect 178582 705562 206026 705798
rect 206262 705562 206346 705798
rect 206582 705562 234026 705798
rect 234262 705562 234346 705798
rect 234582 705562 262026 705798
rect 262262 705562 262346 705798
rect 262582 705562 290026 705798
rect 290262 705562 290346 705798
rect 290582 705562 318026 705798
rect 318262 705562 318346 705798
rect 318582 705562 346026 705798
rect 346262 705562 346346 705798
rect 346582 705562 374026 705798
rect 374262 705562 374346 705798
rect 374582 705562 402026 705798
rect 402262 705562 402346 705798
rect 402582 705562 430026 705798
rect 430262 705562 430346 705798
rect 430582 705562 458026 705798
rect 458262 705562 458346 705798
rect 458582 705562 486026 705798
rect 486262 705562 486346 705798
rect 486582 705562 514026 705798
rect 514262 705562 514346 705798
rect 514582 705562 542026 705798
rect 542262 705562 542346 705798
rect 542582 705562 570026 705798
rect 570262 705562 570346 705798
rect 570582 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 38026 705478
rect 38262 705242 38346 705478
rect 38582 705242 66026 705478
rect 66262 705242 66346 705478
rect 66582 705242 94026 705478
rect 94262 705242 94346 705478
rect 94582 705242 122026 705478
rect 122262 705242 122346 705478
rect 122582 705242 150026 705478
rect 150262 705242 150346 705478
rect 150582 705242 178026 705478
rect 178262 705242 178346 705478
rect 178582 705242 206026 705478
rect 206262 705242 206346 705478
rect 206582 705242 234026 705478
rect 234262 705242 234346 705478
rect 234582 705242 262026 705478
rect 262262 705242 262346 705478
rect 262582 705242 290026 705478
rect 290262 705242 290346 705478
rect 290582 705242 318026 705478
rect 318262 705242 318346 705478
rect 318582 705242 346026 705478
rect 346262 705242 346346 705478
rect 346582 705242 374026 705478
rect 374262 705242 374346 705478
rect 374582 705242 402026 705478
rect 402262 705242 402346 705478
rect 402582 705242 430026 705478
rect 430262 705242 430346 705478
rect 430582 705242 458026 705478
rect 458262 705242 458346 705478
rect 458582 705242 486026 705478
rect 486262 705242 486346 705478
rect 486582 705242 514026 705478
rect 514262 705242 514346 705478
rect 514582 705242 542026 705478
rect 542262 705242 542346 705478
rect 542582 705242 570026 705478
rect 570262 705242 570346 705478
rect 570582 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 41526 704838
rect 41762 704602 41846 704838
rect 42082 704602 69526 704838
rect 69762 704602 69846 704838
rect 70082 704602 97526 704838
rect 97762 704602 97846 704838
rect 98082 704602 125526 704838
rect 125762 704602 125846 704838
rect 126082 704602 153526 704838
rect 153762 704602 153846 704838
rect 154082 704602 181526 704838
rect 181762 704602 181846 704838
rect 182082 704602 209526 704838
rect 209762 704602 209846 704838
rect 210082 704602 237526 704838
rect 237762 704602 237846 704838
rect 238082 704602 265526 704838
rect 265762 704602 265846 704838
rect 266082 704602 293526 704838
rect 293762 704602 293846 704838
rect 294082 704602 321526 704838
rect 321762 704602 321846 704838
rect 322082 704602 349526 704838
rect 349762 704602 349846 704838
rect 350082 704602 377526 704838
rect 377762 704602 377846 704838
rect 378082 704602 405526 704838
rect 405762 704602 405846 704838
rect 406082 704602 433526 704838
rect 433762 704602 433846 704838
rect 434082 704602 461526 704838
rect 461762 704602 461846 704838
rect 462082 704602 489526 704838
rect 489762 704602 489846 704838
rect 490082 704602 517526 704838
rect 517762 704602 517846 704838
rect 518082 704602 545526 704838
rect 545762 704602 545846 704838
rect 546082 704602 573526 704838
rect 573762 704602 573846 704838
rect 574082 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 41526 704518
rect 41762 704282 41846 704518
rect 42082 704282 69526 704518
rect 69762 704282 69846 704518
rect 70082 704282 97526 704518
rect 97762 704282 97846 704518
rect 98082 704282 125526 704518
rect 125762 704282 125846 704518
rect 126082 704282 153526 704518
rect 153762 704282 153846 704518
rect 154082 704282 181526 704518
rect 181762 704282 181846 704518
rect 182082 704282 209526 704518
rect 209762 704282 209846 704518
rect 210082 704282 237526 704518
rect 237762 704282 237846 704518
rect 238082 704282 265526 704518
rect 265762 704282 265846 704518
rect 266082 704282 293526 704518
rect 293762 704282 293846 704518
rect 294082 704282 321526 704518
rect 321762 704282 321846 704518
rect 322082 704282 349526 704518
rect 349762 704282 349846 704518
rect 350082 704282 377526 704518
rect 377762 704282 377846 704518
rect 378082 704282 405526 704518
rect 405762 704282 405846 704518
rect 406082 704282 433526 704518
rect 433762 704282 433846 704518
rect 434082 704282 461526 704518
rect 461762 704282 461846 704518
rect 462082 704282 489526 704518
rect 489762 704282 489846 704518
rect 490082 704282 517526 704518
rect 517762 704282 517846 704518
rect 518082 704282 545526 704518
rect 545762 704282 545846 704518
rect 546082 704282 573526 704518
rect 573762 704282 573846 704518
rect 574082 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 701829 592650 701861
rect -8726 701593 -1974 701829
rect -1738 701593 -1654 701829
rect -1418 701593 41526 701829
rect 41762 701593 41846 701829
rect 42082 701593 69526 701829
rect 69762 701593 69846 701829
rect 70082 701593 97526 701829
rect 97762 701593 97846 701829
rect 98082 701593 125526 701829
rect 125762 701593 125846 701829
rect 126082 701593 153526 701829
rect 153762 701593 153846 701829
rect 154082 701593 181526 701829
rect 181762 701593 181846 701829
rect 182082 701593 209526 701829
rect 209762 701593 209846 701829
rect 210082 701593 237526 701829
rect 237762 701593 237846 701829
rect 238082 701593 265526 701829
rect 265762 701593 265846 701829
rect 266082 701593 293526 701829
rect 293762 701593 293846 701829
rect 294082 701593 321526 701829
rect 321762 701593 321846 701829
rect 322082 701593 349526 701829
rect 349762 701593 349846 701829
rect 350082 701593 377526 701829
rect 377762 701593 377846 701829
rect 378082 701593 405526 701829
rect 405762 701593 405846 701829
rect 406082 701593 433526 701829
rect 433762 701593 433846 701829
rect 434082 701593 461526 701829
rect 461762 701593 461846 701829
rect 462082 701593 489526 701829
rect 489762 701593 489846 701829
rect 490082 701593 517526 701829
rect 517762 701593 517846 701829
rect 518082 701593 545526 701829
rect 545762 701593 545846 701829
rect 546082 701593 573526 701829
rect 573762 701593 573846 701829
rect 574082 701593 585342 701829
rect 585578 701593 585662 701829
rect 585898 701593 592650 701829
rect -8726 701509 592650 701593
rect -8726 701273 -1974 701509
rect -1738 701273 -1654 701509
rect -1418 701273 41526 701509
rect 41762 701273 41846 701509
rect 42082 701273 69526 701509
rect 69762 701273 69846 701509
rect 70082 701273 97526 701509
rect 97762 701273 97846 701509
rect 98082 701273 125526 701509
rect 125762 701273 125846 701509
rect 126082 701273 153526 701509
rect 153762 701273 153846 701509
rect 154082 701273 181526 701509
rect 181762 701273 181846 701509
rect 182082 701273 209526 701509
rect 209762 701273 209846 701509
rect 210082 701273 237526 701509
rect 237762 701273 237846 701509
rect 238082 701273 265526 701509
rect 265762 701273 265846 701509
rect 266082 701273 293526 701509
rect 293762 701273 293846 701509
rect 294082 701273 321526 701509
rect 321762 701273 321846 701509
rect 322082 701273 349526 701509
rect 349762 701273 349846 701509
rect 350082 701273 377526 701509
rect 377762 701273 377846 701509
rect 378082 701273 405526 701509
rect 405762 701273 405846 701509
rect 406082 701273 433526 701509
rect 433762 701273 433846 701509
rect 434082 701273 461526 701509
rect 461762 701273 461846 701509
rect 462082 701273 489526 701509
rect 489762 701273 489846 701509
rect 490082 701273 517526 701509
rect 517762 701273 517846 701509
rect 518082 701273 545526 701509
rect 545762 701273 545846 701509
rect 546082 701273 573526 701509
rect 573762 701273 573846 701509
rect 574082 701273 585342 701509
rect 585578 701273 585662 701509
rect 585898 701273 592650 701509
rect -8726 701241 592650 701273
rect -8726 698454 592650 698486
rect -8726 698218 -2934 698454
rect -2698 698218 -2614 698454
rect -2378 698218 38026 698454
rect 38262 698218 38346 698454
rect 38582 698218 66026 698454
rect 66262 698218 66346 698454
rect 66582 698218 94026 698454
rect 94262 698218 94346 698454
rect 94582 698218 122026 698454
rect 122262 698218 122346 698454
rect 122582 698218 150026 698454
rect 150262 698218 150346 698454
rect 150582 698218 178026 698454
rect 178262 698218 178346 698454
rect 178582 698218 206026 698454
rect 206262 698218 206346 698454
rect 206582 698218 234026 698454
rect 234262 698218 234346 698454
rect 234582 698218 262026 698454
rect 262262 698218 262346 698454
rect 262582 698218 290026 698454
rect 290262 698218 290346 698454
rect 290582 698218 318026 698454
rect 318262 698218 318346 698454
rect 318582 698218 346026 698454
rect 346262 698218 346346 698454
rect 346582 698218 374026 698454
rect 374262 698218 374346 698454
rect 374582 698218 402026 698454
rect 402262 698218 402346 698454
rect 402582 698218 430026 698454
rect 430262 698218 430346 698454
rect 430582 698218 458026 698454
rect 458262 698218 458346 698454
rect 458582 698218 486026 698454
rect 486262 698218 486346 698454
rect 486582 698218 514026 698454
rect 514262 698218 514346 698454
rect 514582 698218 542026 698454
rect 542262 698218 542346 698454
rect 542582 698218 570026 698454
rect 570262 698218 570346 698454
rect 570582 698218 586302 698454
rect 586538 698218 586622 698454
rect 586858 698218 592650 698454
rect -8726 698134 592650 698218
rect -8726 697898 -2934 698134
rect -2698 697898 -2614 698134
rect -2378 697898 38026 698134
rect 38262 697898 38346 698134
rect 38582 697898 66026 698134
rect 66262 697898 66346 698134
rect 66582 697898 94026 698134
rect 94262 697898 94346 698134
rect 94582 697898 122026 698134
rect 122262 697898 122346 698134
rect 122582 697898 150026 698134
rect 150262 697898 150346 698134
rect 150582 697898 178026 698134
rect 178262 697898 178346 698134
rect 178582 697898 206026 698134
rect 206262 697898 206346 698134
rect 206582 697898 234026 698134
rect 234262 697898 234346 698134
rect 234582 697898 262026 698134
rect 262262 697898 262346 698134
rect 262582 697898 290026 698134
rect 290262 697898 290346 698134
rect 290582 697898 318026 698134
rect 318262 697898 318346 698134
rect 318582 697898 346026 698134
rect 346262 697898 346346 698134
rect 346582 697898 374026 698134
rect 374262 697898 374346 698134
rect 374582 697898 402026 698134
rect 402262 697898 402346 698134
rect 402582 697898 430026 698134
rect 430262 697898 430346 698134
rect 430582 697898 458026 698134
rect 458262 697898 458346 698134
rect 458582 697898 486026 698134
rect 486262 697898 486346 698134
rect 486582 697898 514026 698134
rect 514262 697898 514346 698134
rect 514582 697898 542026 698134
rect 542262 697898 542346 698134
rect 542582 697898 570026 698134
rect 570262 697898 570346 698134
rect 570582 697898 586302 698134
rect 586538 697898 586622 698134
rect 586858 697898 592650 698134
rect -8726 697866 592650 697898
rect -8726 674829 592650 674861
rect -8726 674593 -1974 674829
rect -1738 674593 -1654 674829
rect -1418 674593 20118 674829
rect 20354 674593 26382 674829
rect 26618 674593 32646 674829
rect 32882 674593 48118 674829
rect 48354 674593 54382 674829
rect 54618 674593 60646 674829
rect 60882 674593 76118 674829
rect 76354 674593 82382 674829
rect 82618 674593 88646 674829
rect 88882 674593 104118 674829
rect 104354 674593 110382 674829
rect 110618 674593 116646 674829
rect 116882 674593 132118 674829
rect 132354 674593 138382 674829
rect 138618 674593 144646 674829
rect 144882 674593 160118 674829
rect 160354 674593 166382 674829
rect 166618 674593 172646 674829
rect 172882 674593 188118 674829
rect 188354 674593 194382 674829
rect 194618 674593 200646 674829
rect 200882 674593 216118 674829
rect 216354 674593 222382 674829
rect 222618 674593 228646 674829
rect 228882 674593 244118 674829
rect 244354 674593 250382 674829
rect 250618 674593 256646 674829
rect 256882 674593 272118 674829
rect 272354 674593 278382 674829
rect 278618 674593 284646 674829
rect 284882 674593 300118 674829
rect 300354 674593 306382 674829
rect 306618 674593 312646 674829
rect 312882 674593 328118 674829
rect 328354 674593 334382 674829
rect 334618 674593 340646 674829
rect 340882 674593 356118 674829
rect 356354 674593 362382 674829
rect 362618 674593 368646 674829
rect 368882 674593 384118 674829
rect 384354 674593 390382 674829
rect 390618 674593 396646 674829
rect 396882 674593 412118 674829
rect 412354 674593 418382 674829
rect 418618 674593 424646 674829
rect 424882 674593 440118 674829
rect 440354 674593 446382 674829
rect 446618 674593 452646 674829
rect 452882 674593 468118 674829
rect 468354 674593 474382 674829
rect 474618 674593 480646 674829
rect 480882 674593 496118 674829
rect 496354 674593 502382 674829
rect 502618 674593 508646 674829
rect 508882 674593 524118 674829
rect 524354 674593 530382 674829
rect 530618 674593 536646 674829
rect 536882 674593 552118 674829
rect 552354 674593 558382 674829
rect 558618 674593 564646 674829
rect 564882 674593 573526 674829
rect 573762 674593 573846 674829
rect 574082 674593 585342 674829
rect 585578 674593 585662 674829
rect 585898 674593 592650 674829
rect -8726 674509 592650 674593
rect -8726 674273 -1974 674509
rect -1738 674273 -1654 674509
rect -1418 674273 20118 674509
rect 20354 674273 26382 674509
rect 26618 674273 32646 674509
rect 32882 674273 48118 674509
rect 48354 674273 54382 674509
rect 54618 674273 60646 674509
rect 60882 674273 76118 674509
rect 76354 674273 82382 674509
rect 82618 674273 88646 674509
rect 88882 674273 104118 674509
rect 104354 674273 110382 674509
rect 110618 674273 116646 674509
rect 116882 674273 132118 674509
rect 132354 674273 138382 674509
rect 138618 674273 144646 674509
rect 144882 674273 160118 674509
rect 160354 674273 166382 674509
rect 166618 674273 172646 674509
rect 172882 674273 188118 674509
rect 188354 674273 194382 674509
rect 194618 674273 200646 674509
rect 200882 674273 216118 674509
rect 216354 674273 222382 674509
rect 222618 674273 228646 674509
rect 228882 674273 244118 674509
rect 244354 674273 250382 674509
rect 250618 674273 256646 674509
rect 256882 674273 272118 674509
rect 272354 674273 278382 674509
rect 278618 674273 284646 674509
rect 284882 674273 300118 674509
rect 300354 674273 306382 674509
rect 306618 674273 312646 674509
rect 312882 674273 328118 674509
rect 328354 674273 334382 674509
rect 334618 674273 340646 674509
rect 340882 674273 356118 674509
rect 356354 674273 362382 674509
rect 362618 674273 368646 674509
rect 368882 674273 384118 674509
rect 384354 674273 390382 674509
rect 390618 674273 396646 674509
rect 396882 674273 412118 674509
rect 412354 674273 418382 674509
rect 418618 674273 424646 674509
rect 424882 674273 440118 674509
rect 440354 674273 446382 674509
rect 446618 674273 452646 674509
rect 452882 674273 468118 674509
rect 468354 674273 474382 674509
rect 474618 674273 480646 674509
rect 480882 674273 496118 674509
rect 496354 674273 502382 674509
rect 502618 674273 508646 674509
rect 508882 674273 524118 674509
rect 524354 674273 530382 674509
rect 530618 674273 536646 674509
rect 536882 674273 552118 674509
rect 552354 674273 558382 674509
rect 558618 674273 564646 674509
rect 564882 674273 573526 674509
rect 573762 674273 573846 674509
rect 574082 674273 585342 674509
rect 585578 674273 585662 674509
rect 585898 674273 592650 674509
rect -8726 674241 592650 674273
rect -8726 671454 592650 671486
rect -8726 671218 -2934 671454
rect -2698 671218 -2614 671454
rect -2378 671218 23250 671454
rect 23486 671218 29514 671454
rect 29750 671218 51250 671454
rect 51486 671218 57514 671454
rect 57750 671218 79250 671454
rect 79486 671218 85514 671454
rect 85750 671218 107250 671454
rect 107486 671218 113514 671454
rect 113750 671218 135250 671454
rect 135486 671218 141514 671454
rect 141750 671218 163250 671454
rect 163486 671218 169514 671454
rect 169750 671218 191250 671454
rect 191486 671218 197514 671454
rect 197750 671218 219250 671454
rect 219486 671218 225514 671454
rect 225750 671218 247250 671454
rect 247486 671218 253514 671454
rect 253750 671218 275250 671454
rect 275486 671218 281514 671454
rect 281750 671218 303250 671454
rect 303486 671218 309514 671454
rect 309750 671218 331250 671454
rect 331486 671218 337514 671454
rect 337750 671218 359250 671454
rect 359486 671218 365514 671454
rect 365750 671218 387250 671454
rect 387486 671218 393514 671454
rect 393750 671218 415250 671454
rect 415486 671218 421514 671454
rect 421750 671218 443250 671454
rect 443486 671218 449514 671454
rect 449750 671218 471250 671454
rect 471486 671218 477514 671454
rect 477750 671218 499250 671454
rect 499486 671218 505514 671454
rect 505750 671218 527250 671454
rect 527486 671218 533514 671454
rect 533750 671218 555250 671454
rect 555486 671218 561514 671454
rect 561750 671218 586302 671454
rect 586538 671218 586622 671454
rect 586858 671218 592650 671454
rect -8726 671134 592650 671218
rect -8726 670898 -2934 671134
rect -2698 670898 -2614 671134
rect -2378 670898 23250 671134
rect 23486 670898 29514 671134
rect 29750 670898 51250 671134
rect 51486 670898 57514 671134
rect 57750 670898 79250 671134
rect 79486 670898 85514 671134
rect 85750 670898 107250 671134
rect 107486 670898 113514 671134
rect 113750 670898 135250 671134
rect 135486 670898 141514 671134
rect 141750 670898 163250 671134
rect 163486 670898 169514 671134
rect 169750 670898 191250 671134
rect 191486 670898 197514 671134
rect 197750 670898 219250 671134
rect 219486 670898 225514 671134
rect 225750 670898 247250 671134
rect 247486 670898 253514 671134
rect 253750 670898 275250 671134
rect 275486 670898 281514 671134
rect 281750 670898 303250 671134
rect 303486 670898 309514 671134
rect 309750 670898 331250 671134
rect 331486 670898 337514 671134
rect 337750 670898 359250 671134
rect 359486 670898 365514 671134
rect 365750 670898 387250 671134
rect 387486 670898 393514 671134
rect 393750 670898 415250 671134
rect 415486 670898 421514 671134
rect 421750 670898 443250 671134
rect 443486 670898 449514 671134
rect 449750 670898 471250 671134
rect 471486 670898 477514 671134
rect 477750 670898 499250 671134
rect 499486 670898 505514 671134
rect 505750 670898 527250 671134
rect 527486 670898 533514 671134
rect 533750 670898 555250 671134
rect 555486 670898 561514 671134
rect 561750 670898 586302 671134
rect 586538 670898 586622 671134
rect 586858 670898 592650 671134
rect -8726 670866 592650 670898
rect -8726 647829 592650 647861
rect -8726 647593 -1974 647829
rect -1738 647593 -1654 647829
rect -1418 647593 20118 647829
rect 20354 647593 26382 647829
rect 26618 647593 32646 647829
rect 32882 647593 48118 647829
rect 48354 647593 54382 647829
rect 54618 647593 60646 647829
rect 60882 647593 76118 647829
rect 76354 647593 82382 647829
rect 82618 647593 88646 647829
rect 88882 647593 104118 647829
rect 104354 647593 110382 647829
rect 110618 647593 116646 647829
rect 116882 647593 132118 647829
rect 132354 647593 138382 647829
rect 138618 647593 144646 647829
rect 144882 647593 160118 647829
rect 160354 647593 166382 647829
rect 166618 647593 172646 647829
rect 172882 647593 188118 647829
rect 188354 647593 194382 647829
rect 194618 647593 200646 647829
rect 200882 647593 216118 647829
rect 216354 647593 222382 647829
rect 222618 647593 228646 647829
rect 228882 647593 244118 647829
rect 244354 647593 250382 647829
rect 250618 647593 256646 647829
rect 256882 647593 272118 647829
rect 272354 647593 278382 647829
rect 278618 647593 284646 647829
rect 284882 647593 300118 647829
rect 300354 647593 306382 647829
rect 306618 647593 312646 647829
rect 312882 647593 328118 647829
rect 328354 647593 334382 647829
rect 334618 647593 340646 647829
rect 340882 647593 356118 647829
rect 356354 647593 362382 647829
rect 362618 647593 368646 647829
rect 368882 647593 384118 647829
rect 384354 647593 390382 647829
rect 390618 647593 396646 647829
rect 396882 647593 412118 647829
rect 412354 647593 418382 647829
rect 418618 647593 424646 647829
rect 424882 647593 440118 647829
rect 440354 647593 446382 647829
rect 446618 647593 452646 647829
rect 452882 647593 468118 647829
rect 468354 647593 474382 647829
rect 474618 647593 480646 647829
rect 480882 647593 496118 647829
rect 496354 647593 502382 647829
rect 502618 647593 508646 647829
rect 508882 647593 524118 647829
rect 524354 647593 530382 647829
rect 530618 647593 536646 647829
rect 536882 647593 552118 647829
rect 552354 647593 558382 647829
rect 558618 647593 564646 647829
rect 564882 647593 573526 647829
rect 573762 647593 573846 647829
rect 574082 647593 585342 647829
rect 585578 647593 585662 647829
rect 585898 647593 592650 647829
rect -8726 647509 592650 647593
rect -8726 647273 -1974 647509
rect -1738 647273 -1654 647509
rect -1418 647273 20118 647509
rect 20354 647273 26382 647509
rect 26618 647273 32646 647509
rect 32882 647273 48118 647509
rect 48354 647273 54382 647509
rect 54618 647273 60646 647509
rect 60882 647273 76118 647509
rect 76354 647273 82382 647509
rect 82618 647273 88646 647509
rect 88882 647273 104118 647509
rect 104354 647273 110382 647509
rect 110618 647273 116646 647509
rect 116882 647273 132118 647509
rect 132354 647273 138382 647509
rect 138618 647273 144646 647509
rect 144882 647273 160118 647509
rect 160354 647273 166382 647509
rect 166618 647273 172646 647509
rect 172882 647273 188118 647509
rect 188354 647273 194382 647509
rect 194618 647273 200646 647509
rect 200882 647273 216118 647509
rect 216354 647273 222382 647509
rect 222618 647273 228646 647509
rect 228882 647273 244118 647509
rect 244354 647273 250382 647509
rect 250618 647273 256646 647509
rect 256882 647273 272118 647509
rect 272354 647273 278382 647509
rect 278618 647273 284646 647509
rect 284882 647273 300118 647509
rect 300354 647273 306382 647509
rect 306618 647273 312646 647509
rect 312882 647273 328118 647509
rect 328354 647273 334382 647509
rect 334618 647273 340646 647509
rect 340882 647273 356118 647509
rect 356354 647273 362382 647509
rect 362618 647273 368646 647509
rect 368882 647273 384118 647509
rect 384354 647273 390382 647509
rect 390618 647273 396646 647509
rect 396882 647273 412118 647509
rect 412354 647273 418382 647509
rect 418618 647273 424646 647509
rect 424882 647273 440118 647509
rect 440354 647273 446382 647509
rect 446618 647273 452646 647509
rect 452882 647273 468118 647509
rect 468354 647273 474382 647509
rect 474618 647273 480646 647509
rect 480882 647273 496118 647509
rect 496354 647273 502382 647509
rect 502618 647273 508646 647509
rect 508882 647273 524118 647509
rect 524354 647273 530382 647509
rect 530618 647273 536646 647509
rect 536882 647273 552118 647509
rect 552354 647273 558382 647509
rect 558618 647273 564646 647509
rect 564882 647273 573526 647509
rect 573762 647273 573846 647509
rect 574082 647273 585342 647509
rect 585578 647273 585662 647509
rect 585898 647273 592650 647509
rect -8726 647241 592650 647273
rect -8726 644454 592650 644486
rect -8726 644218 -2934 644454
rect -2698 644218 -2614 644454
rect -2378 644218 23250 644454
rect 23486 644218 29514 644454
rect 29750 644218 51250 644454
rect 51486 644218 57514 644454
rect 57750 644218 79250 644454
rect 79486 644218 85514 644454
rect 85750 644218 107250 644454
rect 107486 644218 113514 644454
rect 113750 644218 135250 644454
rect 135486 644218 141514 644454
rect 141750 644218 163250 644454
rect 163486 644218 169514 644454
rect 169750 644218 191250 644454
rect 191486 644218 197514 644454
rect 197750 644218 219250 644454
rect 219486 644218 225514 644454
rect 225750 644218 247250 644454
rect 247486 644218 253514 644454
rect 253750 644218 275250 644454
rect 275486 644218 281514 644454
rect 281750 644218 303250 644454
rect 303486 644218 309514 644454
rect 309750 644218 331250 644454
rect 331486 644218 337514 644454
rect 337750 644218 359250 644454
rect 359486 644218 365514 644454
rect 365750 644218 387250 644454
rect 387486 644218 393514 644454
rect 393750 644218 415250 644454
rect 415486 644218 421514 644454
rect 421750 644218 443250 644454
rect 443486 644218 449514 644454
rect 449750 644218 471250 644454
rect 471486 644218 477514 644454
rect 477750 644218 499250 644454
rect 499486 644218 505514 644454
rect 505750 644218 527250 644454
rect 527486 644218 533514 644454
rect 533750 644218 555250 644454
rect 555486 644218 561514 644454
rect 561750 644218 586302 644454
rect 586538 644218 586622 644454
rect 586858 644218 592650 644454
rect -8726 644134 592650 644218
rect -8726 643898 -2934 644134
rect -2698 643898 -2614 644134
rect -2378 643898 23250 644134
rect 23486 643898 29514 644134
rect 29750 643898 51250 644134
rect 51486 643898 57514 644134
rect 57750 643898 79250 644134
rect 79486 643898 85514 644134
rect 85750 643898 107250 644134
rect 107486 643898 113514 644134
rect 113750 643898 135250 644134
rect 135486 643898 141514 644134
rect 141750 643898 163250 644134
rect 163486 643898 169514 644134
rect 169750 643898 191250 644134
rect 191486 643898 197514 644134
rect 197750 643898 219250 644134
rect 219486 643898 225514 644134
rect 225750 643898 247250 644134
rect 247486 643898 253514 644134
rect 253750 643898 275250 644134
rect 275486 643898 281514 644134
rect 281750 643898 303250 644134
rect 303486 643898 309514 644134
rect 309750 643898 331250 644134
rect 331486 643898 337514 644134
rect 337750 643898 359250 644134
rect 359486 643898 365514 644134
rect 365750 643898 387250 644134
rect 387486 643898 393514 644134
rect 393750 643898 415250 644134
rect 415486 643898 421514 644134
rect 421750 643898 443250 644134
rect 443486 643898 449514 644134
rect 449750 643898 471250 644134
rect 471486 643898 477514 644134
rect 477750 643898 499250 644134
rect 499486 643898 505514 644134
rect 505750 643898 527250 644134
rect 527486 643898 533514 644134
rect 533750 643898 555250 644134
rect 555486 643898 561514 644134
rect 561750 643898 586302 644134
rect 586538 643898 586622 644134
rect 586858 643898 592650 644134
rect -8726 643866 592650 643898
rect -8726 620829 592650 620861
rect -8726 620593 -1974 620829
rect -1738 620593 -1654 620829
rect -1418 620593 20118 620829
rect 20354 620593 26382 620829
rect 26618 620593 32646 620829
rect 32882 620593 48118 620829
rect 48354 620593 54382 620829
rect 54618 620593 60646 620829
rect 60882 620593 76118 620829
rect 76354 620593 82382 620829
rect 82618 620593 88646 620829
rect 88882 620593 104118 620829
rect 104354 620593 110382 620829
rect 110618 620593 116646 620829
rect 116882 620593 132118 620829
rect 132354 620593 138382 620829
rect 138618 620593 144646 620829
rect 144882 620593 160118 620829
rect 160354 620593 166382 620829
rect 166618 620593 172646 620829
rect 172882 620593 188118 620829
rect 188354 620593 194382 620829
rect 194618 620593 200646 620829
rect 200882 620593 216118 620829
rect 216354 620593 222382 620829
rect 222618 620593 228646 620829
rect 228882 620593 244118 620829
rect 244354 620593 250382 620829
rect 250618 620593 256646 620829
rect 256882 620593 272118 620829
rect 272354 620593 278382 620829
rect 278618 620593 284646 620829
rect 284882 620593 300118 620829
rect 300354 620593 306382 620829
rect 306618 620593 312646 620829
rect 312882 620593 328118 620829
rect 328354 620593 334382 620829
rect 334618 620593 340646 620829
rect 340882 620593 356118 620829
rect 356354 620593 362382 620829
rect 362618 620593 368646 620829
rect 368882 620593 384118 620829
rect 384354 620593 390382 620829
rect 390618 620593 396646 620829
rect 396882 620593 412118 620829
rect 412354 620593 418382 620829
rect 418618 620593 424646 620829
rect 424882 620593 440118 620829
rect 440354 620593 446382 620829
rect 446618 620593 452646 620829
rect 452882 620593 468118 620829
rect 468354 620593 474382 620829
rect 474618 620593 480646 620829
rect 480882 620593 496118 620829
rect 496354 620593 502382 620829
rect 502618 620593 508646 620829
rect 508882 620593 524118 620829
rect 524354 620593 530382 620829
rect 530618 620593 536646 620829
rect 536882 620593 552118 620829
rect 552354 620593 558382 620829
rect 558618 620593 564646 620829
rect 564882 620593 573526 620829
rect 573762 620593 573846 620829
rect 574082 620593 585342 620829
rect 585578 620593 585662 620829
rect 585898 620593 592650 620829
rect -8726 620509 592650 620593
rect -8726 620273 -1974 620509
rect -1738 620273 -1654 620509
rect -1418 620273 20118 620509
rect 20354 620273 26382 620509
rect 26618 620273 32646 620509
rect 32882 620273 48118 620509
rect 48354 620273 54382 620509
rect 54618 620273 60646 620509
rect 60882 620273 76118 620509
rect 76354 620273 82382 620509
rect 82618 620273 88646 620509
rect 88882 620273 104118 620509
rect 104354 620273 110382 620509
rect 110618 620273 116646 620509
rect 116882 620273 132118 620509
rect 132354 620273 138382 620509
rect 138618 620273 144646 620509
rect 144882 620273 160118 620509
rect 160354 620273 166382 620509
rect 166618 620273 172646 620509
rect 172882 620273 188118 620509
rect 188354 620273 194382 620509
rect 194618 620273 200646 620509
rect 200882 620273 216118 620509
rect 216354 620273 222382 620509
rect 222618 620273 228646 620509
rect 228882 620273 244118 620509
rect 244354 620273 250382 620509
rect 250618 620273 256646 620509
rect 256882 620273 272118 620509
rect 272354 620273 278382 620509
rect 278618 620273 284646 620509
rect 284882 620273 300118 620509
rect 300354 620273 306382 620509
rect 306618 620273 312646 620509
rect 312882 620273 328118 620509
rect 328354 620273 334382 620509
rect 334618 620273 340646 620509
rect 340882 620273 356118 620509
rect 356354 620273 362382 620509
rect 362618 620273 368646 620509
rect 368882 620273 384118 620509
rect 384354 620273 390382 620509
rect 390618 620273 396646 620509
rect 396882 620273 412118 620509
rect 412354 620273 418382 620509
rect 418618 620273 424646 620509
rect 424882 620273 440118 620509
rect 440354 620273 446382 620509
rect 446618 620273 452646 620509
rect 452882 620273 468118 620509
rect 468354 620273 474382 620509
rect 474618 620273 480646 620509
rect 480882 620273 496118 620509
rect 496354 620273 502382 620509
rect 502618 620273 508646 620509
rect 508882 620273 524118 620509
rect 524354 620273 530382 620509
rect 530618 620273 536646 620509
rect 536882 620273 552118 620509
rect 552354 620273 558382 620509
rect 558618 620273 564646 620509
rect 564882 620273 573526 620509
rect 573762 620273 573846 620509
rect 574082 620273 585342 620509
rect 585578 620273 585662 620509
rect 585898 620273 592650 620509
rect -8726 620241 592650 620273
rect -8726 617454 592650 617486
rect -8726 617218 -2934 617454
rect -2698 617218 -2614 617454
rect -2378 617218 23250 617454
rect 23486 617218 29514 617454
rect 29750 617218 51250 617454
rect 51486 617218 57514 617454
rect 57750 617218 79250 617454
rect 79486 617218 85514 617454
rect 85750 617218 107250 617454
rect 107486 617218 113514 617454
rect 113750 617218 135250 617454
rect 135486 617218 141514 617454
rect 141750 617218 163250 617454
rect 163486 617218 169514 617454
rect 169750 617218 191250 617454
rect 191486 617218 197514 617454
rect 197750 617218 219250 617454
rect 219486 617218 225514 617454
rect 225750 617218 247250 617454
rect 247486 617218 253514 617454
rect 253750 617218 275250 617454
rect 275486 617218 281514 617454
rect 281750 617218 303250 617454
rect 303486 617218 309514 617454
rect 309750 617218 331250 617454
rect 331486 617218 337514 617454
rect 337750 617218 359250 617454
rect 359486 617218 365514 617454
rect 365750 617218 387250 617454
rect 387486 617218 393514 617454
rect 393750 617218 415250 617454
rect 415486 617218 421514 617454
rect 421750 617218 443250 617454
rect 443486 617218 449514 617454
rect 449750 617218 471250 617454
rect 471486 617218 477514 617454
rect 477750 617218 499250 617454
rect 499486 617218 505514 617454
rect 505750 617218 527250 617454
rect 527486 617218 533514 617454
rect 533750 617218 555250 617454
rect 555486 617218 561514 617454
rect 561750 617218 586302 617454
rect 586538 617218 586622 617454
rect 586858 617218 592650 617454
rect -8726 617134 592650 617218
rect -8726 616898 -2934 617134
rect -2698 616898 -2614 617134
rect -2378 616898 23250 617134
rect 23486 616898 29514 617134
rect 29750 616898 51250 617134
rect 51486 616898 57514 617134
rect 57750 616898 79250 617134
rect 79486 616898 85514 617134
rect 85750 616898 107250 617134
rect 107486 616898 113514 617134
rect 113750 616898 135250 617134
rect 135486 616898 141514 617134
rect 141750 616898 163250 617134
rect 163486 616898 169514 617134
rect 169750 616898 191250 617134
rect 191486 616898 197514 617134
rect 197750 616898 219250 617134
rect 219486 616898 225514 617134
rect 225750 616898 247250 617134
rect 247486 616898 253514 617134
rect 253750 616898 275250 617134
rect 275486 616898 281514 617134
rect 281750 616898 303250 617134
rect 303486 616898 309514 617134
rect 309750 616898 331250 617134
rect 331486 616898 337514 617134
rect 337750 616898 359250 617134
rect 359486 616898 365514 617134
rect 365750 616898 387250 617134
rect 387486 616898 393514 617134
rect 393750 616898 415250 617134
rect 415486 616898 421514 617134
rect 421750 616898 443250 617134
rect 443486 616898 449514 617134
rect 449750 616898 471250 617134
rect 471486 616898 477514 617134
rect 477750 616898 499250 617134
rect 499486 616898 505514 617134
rect 505750 616898 527250 617134
rect 527486 616898 533514 617134
rect 533750 616898 555250 617134
rect 555486 616898 561514 617134
rect 561750 616898 586302 617134
rect 586538 616898 586622 617134
rect 586858 616898 592650 617134
rect -8726 616866 592650 616898
rect -8726 593829 592650 593861
rect -8726 593593 -1974 593829
rect -1738 593593 -1654 593829
rect -1418 593593 20118 593829
rect 20354 593593 26382 593829
rect 26618 593593 32646 593829
rect 32882 593593 48118 593829
rect 48354 593593 54382 593829
rect 54618 593593 60646 593829
rect 60882 593593 76118 593829
rect 76354 593593 82382 593829
rect 82618 593593 88646 593829
rect 88882 593593 104118 593829
rect 104354 593593 110382 593829
rect 110618 593593 116646 593829
rect 116882 593593 132118 593829
rect 132354 593593 138382 593829
rect 138618 593593 144646 593829
rect 144882 593593 160118 593829
rect 160354 593593 166382 593829
rect 166618 593593 172646 593829
rect 172882 593593 188118 593829
rect 188354 593593 194382 593829
rect 194618 593593 200646 593829
rect 200882 593593 216118 593829
rect 216354 593593 222382 593829
rect 222618 593593 228646 593829
rect 228882 593593 244118 593829
rect 244354 593593 250382 593829
rect 250618 593593 256646 593829
rect 256882 593593 272118 593829
rect 272354 593593 278382 593829
rect 278618 593593 284646 593829
rect 284882 593593 300118 593829
rect 300354 593593 306382 593829
rect 306618 593593 312646 593829
rect 312882 593593 328118 593829
rect 328354 593593 334382 593829
rect 334618 593593 340646 593829
rect 340882 593593 356118 593829
rect 356354 593593 362382 593829
rect 362618 593593 368646 593829
rect 368882 593593 384118 593829
rect 384354 593593 390382 593829
rect 390618 593593 396646 593829
rect 396882 593593 412118 593829
rect 412354 593593 418382 593829
rect 418618 593593 424646 593829
rect 424882 593593 440118 593829
rect 440354 593593 446382 593829
rect 446618 593593 452646 593829
rect 452882 593593 468118 593829
rect 468354 593593 474382 593829
rect 474618 593593 480646 593829
rect 480882 593593 496118 593829
rect 496354 593593 502382 593829
rect 502618 593593 508646 593829
rect 508882 593593 524118 593829
rect 524354 593593 530382 593829
rect 530618 593593 536646 593829
rect 536882 593593 552118 593829
rect 552354 593593 558382 593829
rect 558618 593593 564646 593829
rect 564882 593593 573526 593829
rect 573762 593593 573846 593829
rect 574082 593593 585342 593829
rect 585578 593593 585662 593829
rect 585898 593593 592650 593829
rect -8726 593509 592650 593593
rect -8726 593273 -1974 593509
rect -1738 593273 -1654 593509
rect -1418 593273 20118 593509
rect 20354 593273 26382 593509
rect 26618 593273 32646 593509
rect 32882 593273 48118 593509
rect 48354 593273 54382 593509
rect 54618 593273 60646 593509
rect 60882 593273 76118 593509
rect 76354 593273 82382 593509
rect 82618 593273 88646 593509
rect 88882 593273 104118 593509
rect 104354 593273 110382 593509
rect 110618 593273 116646 593509
rect 116882 593273 132118 593509
rect 132354 593273 138382 593509
rect 138618 593273 144646 593509
rect 144882 593273 160118 593509
rect 160354 593273 166382 593509
rect 166618 593273 172646 593509
rect 172882 593273 188118 593509
rect 188354 593273 194382 593509
rect 194618 593273 200646 593509
rect 200882 593273 216118 593509
rect 216354 593273 222382 593509
rect 222618 593273 228646 593509
rect 228882 593273 244118 593509
rect 244354 593273 250382 593509
rect 250618 593273 256646 593509
rect 256882 593273 272118 593509
rect 272354 593273 278382 593509
rect 278618 593273 284646 593509
rect 284882 593273 300118 593509
rect 300354 593273 306382 593509
rect 306618 593273 312646 593509
rect 312882 593273 328118 593509
rect 328354 593273 334382 593509
rect 334618 593273 340646 593509
rect 340882 593273 356118 593509
rect 356354 593273 362382 593509
rect 362618 593273 368646 593509
rect 368882 593273 384118 593509
rect 384354 593273 390382 593509
rect 390618 593273 396646 593509
rect 396882 593273 412118 593509
rect 412354 593273 418382 593509
rect 418618 593273 424646 593509
rect 424882 593273 440118 593509
rect 440354 593273 446382 593509
rect 446618 593273 452646 593509
rect 452882 593273 468118 593509
rect 468354 593273 474382 593509
rect 474618 593273 480646 593509
rect 480882 593273 496118 593509
rect 496354 593273 502382 593509
rect 502618 593273 508646 593509
rect 508882 593273 524118 593509
rect 524354 593273 530382 593509
rect 530618 593273 536646 593509
rect 536882 593273 552118 593509
rect 552354 593273 558382 593509
rect 558618 593273 564646 593509
rect 564882 593273 573526 593509
rect 573762 593273 573846 593509
rect 574082 593273 585342 593509
rect 585578 593273 585662 593509
rect 585898 593273 592650 593509
rect -8726 593241 592650 593273
rect -8726 590454 592650 590486
rect -8726 590218 -2934 590454
rect -2698 590218 -2614 590454
rect -2378 590218 23250 590454
rect 23486 590218 29514 590454
rect 29750 590218 51250 590454
rect 51486 590218 57514 590454
rect 57750 590218 79250 590454
rect 79486 590218 85514 590454
rect 85750 590218 107250 590454
rect 107486 590218 113514 590454
rect 113750 590218 135250 590454
rect 135486 590218 141514 590454
rect 141750 590218 163250 590454
rect 163486 590218 169514 590454
rect 169750 590218 191250 590454
rect 191486 590218 197514 590454
rect 197750 590218 219250 590454
rect 219486 590218 225514 590454
rect 225750 590218 247250 590454
rect 247486 590218 253514 590454
rect 253750 590218 275250 590454
rect 275486 590218 281514 590454
rect 281750 590218 303250 590454
rect 303486 590218 309514 590454
rect 309750 590218 331250 590454
rect 331486 590218 337514 590454
rect 337750 590218 359250 590454
rect 359486 590218 365514 590454
rect 365750 590218 387250 590454
rect 387486 590218 393514 590454
rect 393750 590218 415250 590454
rect 415486 590218 421514 590454
rect 421750 590218 443250 590454
rect 443486 590218 449514 590454
rect 449750 590218 471250 590454
rect 471486 590218 477514 590454
rect 477750 590218 499250 590454
rect 499486 590218 505514 590454
rect 505750 590218 527250 590454
rect 527486 590218 533514 590454
rect 533750 590218 555250 590454
rect 555486 590218 561514 590454
rect 561750 590218 586302 590454
rect 586538 590218 586622 590454
rect 586858 590218 592650 590454
rect -8726 590134 592650 590218
rect -8726 589898 -2934 590134
rect -2698 589898 -2614 590134
rect -2378 589898 23250 590134
rect 23486 589898 29514 590134
rect 29750 589898 51250 590134
rect 51486 589898 57514 590134
rect 57750 589898 79250 590134
rect 79486 589898 85514 590134
rect 85750 589898 107250 590134
rect 107486 589898 113514 590134
rect 113750 589898 135250 590134
rect 135486 589898 141514 590134
rect 141750 589898 163250 590134
rect 163486 589898 169514 590134
rect 169750 589898 191250 590134
rect 191486 589898 197514 590134
rect 197750 589898 219250 590134
rect 219486 589898 225514 590134
rect 225750 589898 247250 590134
rect 247486 589898 253514 590134
rect 253750 589898 275250 590134
rect 275486 589898 281514 590134
rect 281750 589898 303250 590134
rect 303486 589898 309514 590134
rect 309750 589898 331250 590134
rect 331486 589898 337514 590134
rect 337750 589898 359250 590134
rect 359486 589898 365514 590134
rect 365750 589898 387250 590134
rect 387486 589898 393514 590134
rect 393750 589898 415250 590134
rect 415486 589898 421514 590134
rect 421750 589898 443250 590134
rect 443486 589898 449514 590134
rect 449750 589898 471250 590134
rect 471486 589898 477514 590134
rect 477750 589898 499250 590134
rect 499486 589898 505514 590134
rect 505750 589898 527250 590134
rect 527486 589898 533514 590134
rect 533750 589898 555250 590134
rect 555486 589898 561514 590134
rect 561750 589898 586302 590134
rect 586538 589898 586622 590134
rect 586858 589898 592650 590134
rect -8726 589866 592650 589898
rect -8726 566829 592650 566861
rect -8726 566593 -1974 566829
rect -1738 566593 -1654 566829
rect -1418 566593 20118 566829
rect 20354 566593 26382 566829
rect 26618 566593 32646 566829
rect 32882 566593 48118 566829
rect 48354 566593 54382 566829
rect 54618 566593 60646 566829
rect 60882 566593 76118 566829
rect 76354 566593 82382 566829
rect 82618 566593 88646 566829
rect 88882 566593 104118 566829
rect 104354 566593 110382 566829
rect 110618 566593 116646 566829
rect 116882 566593 132118 566829
rect 132354 566593 138382 566829
rect 138618 566593 144646 566829
rect 144882 566593 160118 566829
rect 160354 566593 166382 566829
rect 166618 566593 172646 566829
rect 172882 566593 188118 566829
rect 188354 566593 194382 566829
rect 194618 566593 200646 566829
rect 200882 566593 216118 566829
rect 216354 566593 222382 566829
rect 222618 566593 228646 566829
rect 228882 566593 244118 566829
rect 244354 566593 250382 566829
rect 250618 566593 256646 566829
rect 256882 566593 272118 566829
rect 272354 566593 278382 566829
rect 278618 566593 284646 566829
rect 284882 566593 300118 566829
rect 300354 566593 306382 566829
rect 306618 566593 312646 566829
rect 312882 566593 328118 566829
rect 328354 566593 334382 566829
rect 334618 566593 340646 566829
rect 340882 566593 356118 566829
rect 356354 566593 362382 566829
rect 362618 566593 368646 566829
rect 368882 566593 384118 566829
rect 384354 566593 390382 566829
rect 390618 566593 396646 566829
rect 396882 566593 412118 566829
rect 412354 566593 418382 566829
rect 418618 566593 424646 566829
rect 424882 566593 440118 566829
rect 440354 566593 446382 566829
rect 446618 566593 452646 566829
rect 452882 566593 468118 566829
rect 468354 566593 474382 566829
rect 474618 566593 480646 566829
rect 480882 566593 496118 566829
rect 496354 566593 502382 566829
rect 502618 566593 508646 566829
rect 508882 566593 524118 566829
rect 524354 566593 530382 566829
rect 530618 566593 536646 566829
rect 536882 566593 552118 566829
rect 552354 566593 558382 566829
rect 558618 566593 564646 566829
rect 564882 566593 573526 566829
rect 573762 566593 573846 566829
rect 574082 566593 585342 566829
rect 585578 566593 585662 566829
rect 585898 566593 592650 566829
rect -8726 566509 592650 566593
rect -8726 566273 -1974 566509
rect -1738 566273 -1654 566509
rect -1418 566273 20118 566509
rect 20354 566273 26382 566509
rect 26618 566273 32646 566509
rect 32882 566273 48118 566509
rect 48354 566273 54382 566509
rect 54618 566273 60646 566509
rect 60882 566273 76118 566509
rect 76354 566273 82382 566509
rect 82618 566273 88646 566509
rect 88882 566273 104118 566509
rect 104354 566273 110382 566509
rect 110618 566273 116646 566509
rect 116882 566273 132118 566509
rect 132354 566273 138382 566509
rect 138618 566273 144646 566509
rect 144882 566273 160118 566509
rect 160354 566273 166382 566509
rect 166618 566273 172646 566509
rect 172882 566273 188118 566509
rect 188354 566273 194382 566509
rect 194618 566273 200646 566509
rect 200882 566273 216118 566509
rect 216354 566273 222382 566509
rect 222618 566273 228646 566509
rect 228882 566273 244118 566509
rect 244354 566273 250382 566509
rect 250618 566273 256646 566509
rect 256882 566273 272118 566509
rect 272354 566273 278382 566509
rect 278618 566273 284646 566509
rect 284882 566273 300118 566509
rect 300354 566273 306382 566509
rect 306618 566273 312646 566509
rect 312882 566273 328118 566509
rect 328354 566273 334382 566509
rect 334618 566273 340646 566509
rect 340882 566273 356118 566509
rect 356354 566273 362382 566509
rect 362618 566273 368646 566509
rect 368882 566273 384118 566509
rect 384354 566273 390382 566509
rect 390618 566273 396646 566509
rect 396882 566273 412118 566509
rect 412354 566273 418382 566509
rect 418618 566273 424646 566509
rect 424882 566273 440118 566509
rect 440354 566273 446382 566509
rect 446618 566273 452646 566509
rect 452882 566273 468118 566509
rect 468354 566273 474382 566509
rect 474618 566273 480646 566509
rect 480882 566273 496118 566509
rect 496354 566273 502382 566509
rect 502618 566273 508646 566509
rect 508882 566273 524118 566509
rect 524354 566273 530382 566509
rect 530618 566273 536646 566509
rect 536882 566273 552118 566509
rect 552354 566273 558382 566509
rect 558618 566273 564646 566509
rect 564882 566273 573526 566509
rect 573762 566273 573846 566509
rect 574082 566273 585342 566509
rect 585578 566273 585662 566509
rect 585898 566273 592650 566509
rect -8726 566241 592650 566273
rect -8726 563454 592650 563486
rect -8726 563218 -2934 563454
rect -2698 563218 -2614 563454
rect -2378 563218 23250 563454
rect 23486 563218 29514 563454
rect 29750 563218 51250 563454
rect 51486 563218 57514 563454
rect 57750 563218 79250 563454
rect 79486 563218 85514 563454
rect 85750 563218 107250 563454
rect 107486 563218 113514 563454
rect 113750 563218 135250 563454
rect 135486 563218 141514 563454
rect 141750 563218 163250 563454
rect 163486 563218 169514 563454
rect 169750 563218 191250 563454
rect 191486 563218 197514 563454
rect 197750 563218 219250 563454
rect 219486 563218 225514 563454
rect 225750 563218 247250 563454
rect 247486 563218 253514 563454
rect 253750 563218 275250 563454
rect 275486 563218 281514 563454
rect 281750 563218 303250 563454
rect 303486 563218 309514 563454
rect 309750 563218 331250 563454
rect 331486 563218 337514 563454
rect 337750 563218 359250 563454
rect 359486 563218 365514 563454
rect 365750 563218 387250 563454
rect 387486 563218 393514 563454
rect 393750 563218 415250 563454
rect 415486 563218 421514 563454
rect 421750 563218 443250 563454
rect 443486 563218 449514 563454
rect 449750 563218 471250 563454
rect 471486 563218 477514 563454
rect 477750 563218 499250 563454
rect 499486 563218 505514 563454
rect 505750 563218 527250 563454
rect 527486 563218 533514 563454
rect 533750 563218 555250 563454
rect 555486 563218 561514 563454
rect 561750 563218 586302 563454
rect 586538 563218 586622 563454
rect 586858 563218 592650 563454
rect -8726 563134 592650 563218
rect -8726 562898 -2934 563134
rect -2698 562898 -2614 563134
rect -2378 562898 23250 563134
rect 23486 562898 29514 563134
rect 29750 562898 51250 563134
rect 51486 562898 57514 563134
rect 57750 562898 79250 563134
rect 79486 562898 85514 563134
rect 85750 562898 107250 563134
rect 107486 562898 113514 563134
rect 113750 562898 135250 563134
rect 135486 562898 141514 563134
rect 141750 562898 163250 563134
rect 163486 562898 169514 563134
rect 169750 562898 191250 563134
rect 191486 562898 197514 563134
rect 197750 562898 219250 563134
rect 219486 562898 225514 563134
rect 225750 562898 247250 563134
rect 247486 562898 253514 563134
rect 253750 562898 275250 563134
rect 275486 562898 281514 563134
rect 281750 562898 303250 563134
rect 303486 562898 309514 563134
rect 309750 562898 331250 563134
rect 331486 562898 337514 563134
rect 337750 562898 359250 563134
rect 359486 562898 365514 563134
rect 365750 562898 387250 563134
rect 387486 562898 393514 563134
rect 393750 562898 415250 563134
rect 415486 562898 421514 563134
rect 421750 562898 443250 563134
rect 443486 562898 449514 563134
rect 449750 562898 471250 563134
rect 471486 562898 477514 563134
rect 477750 562898 499250 563134
rect 499486 562898 505514 563134
rect 505750 562898 527250 563134
rect 527486 562898 533514 563134
rect 533750 562898 555250 563134
rect 555486 562898 561514 563134
rect 561750 562898 586302 563134
rect 586538 562898 586622 563134
rect 586858 562898 592650 563134
rect -8726 562866 592650 562898
rect -8726 539829 592650 539861
rect -8726 539593 -1974 539829
rect -1738 539593 -1654 539829
rect -1418 539593 20118 539829
rect 20354 539593 26382 539829
rect 26618 539593 32646 539829
rect 32882 539593 48118 539829
rect 48354 539593 54382 539829
rect 54618 539593 60646 539829
rect 60882 539593 76118 539829
rect 76354 539593 82382 539829
rect 82618 539593 88646 539829
rect 88882 539593 104118 539829
rect 104354 539593 110382 539829
rect 110618 539593 116646 539829
rect 116882 539593 132118 539829
rect 132354 539593 138382 539829
rect 138618 539593 144646 539829
rect 144882 539593 160118 539829
rect 160354 539593 166382 539829
rect 166618 539593 172646 539829
rect 172882 539593 188118 539829
rect 188354 539593 194382 539829
rect 194618 539593 200646 539829
rect 200882 539593 216118 539829
rect 216354 539593 222382 539829
rect 222618 539593 228646 539829
rect 228882 539593 244118 539829
rect 244354 539593 250382 539829
rect 250618 539593 256646 539829
rect 256882 539593 272118 539829
rect 272354 539593 278382 539829
rect 278618 539593 284646 539829
rect 284882 539593 300118 539829
rect 300354 539593 306382 539829
rect 306618 539593 312646 539829
rect 312882 539593 328118 539829
rect 328354 539593 334382 539829
rect 334618 539593 340646 539829
rect 340882 539593 356118 539829
rect 356354 539593 362382 539829
rect 362618 539593 368646 539829
rect 368882 539593 384118 539829
rect 384354 539593 390382 539829
rect 390618 539593 396646 539829
rect 396882 539593 412118 539829
rect 412354 539593 418382 539829
rect 418618 539593 424646 539829
rect 424882 539593 440118 539829
rect 440354 539593 446382 539829
rect 446618 539593 452646 539829
rect 452882 539593 468118 539829
rect 468354 539593 474382 539829
rect 474618 539593 480646 539829
rect 480882 539593 496118 539829
rect 496354 539593 502382 539829
rect 502618 539593 508646 539829
rect 508882 539593 524118 539829
rect 524354 539593 530382 539829
rect 530618 539593 536646 539829
rect 536882 539593 552118 539829
rect 552354 539593 558382 539829
rect 558618 539593 564646 539829
rect 564882 539593 573526 539829
rect 573762 539593 573846 539829
rect 574082 539593 585342 539829
rect 585578 539593 585662 539829
rect 585898 539593 592650 539829
rect -8726 539509 592650 539593
rect -8726 539273 -1974 539509
rect -1738 539273 -1654 539509
rect -1418 539273 20118 539509
rect 20354 539273 26382 539509
rect 26618 539273 32646 539509
rect 32882 539273 48118 539509
rect 48354 539273 54382 539509
rect 54618 539273 60646 539509
rect 60882 539273 76118 539509
rect 76354 539273 82382 539509
rect 82618 539273 88646 539509
rect 88882 539273 104118 539509
rect 104354 539273 110382 539509
rect 110618 539273 116646 539509
rect 116882 539273 132118 539509
rect 132354 539273 138382 539509
rect 138618 539273 144646 539509
rect 144882 539273 160118 539509
rect 160354 539273 166382 539509
rect 166618 539273 172646 539509
rect 172882 539273 188118 539509
rect 188354 539273 194382 539509
rect 194618 539273 200646 539509
rect 200882 539273 216118 539509
rect 216354 539273 222382 539509
rect 222618 539273 228646 539509
rect 228882 539273 244118 539509
rect 244354 539273 250382 539509
rect 250618 539273 256646 539509
rect 256882 539273 272118 539509
rect 272354 539273 278382 539509
rect 278618 539273 284646 539509
rect 284882 539273 300118 539509
rect 300354 539273 306382 539509
rect 306618 539273 312646 539509
rect 312882 539273 328118 539509
rect 328354 539273 334382 539509
rect 334618 539273 340646 539509
rect 340882 539273 356118 539509
rect 356354 539273 362382 539509
rect 362618 539273 368646 539509
rect 368882 539273 384118 539509
rect 384354 539273 390382 539509
rect 390618 539273 396646 539509
rect 396882 539273 412118 539509
rect 412354 539273 418382 539509
rect 418618 539273 424646 539509
rect 424882 539273 440118 539509
rect 440354 539273 446382 539509
rect 446618 539273 452646 539509
rect 452882 539273 468118 539509
rect 468354 539273 474382 539509
rect 474618 539273 480646 539509
rect 480882 539273 496118 539509
rect 496354 539273 502382 539509
rect 502618 539273 508646 539509
rect 508882 539273 524118 539509
rect 524354 539273 530382 539509
rect 530618 539273 536646 539509
rect 536882 539273 552118 539509
rect 552354 539273 558382 539509
rect 558618 539273 564646 539509
rect 564882 539273 573526 539509
rect 573762 539273 573846 539509
rect 574082 539273 585342 539509
rect 585578 539273 585662 539509
rect 585898 539273 592650 539509
rect -8726 539241 592650 539273
rect -8726 536454 592650 536486
rect -8726 536218 -2934 536454
rect -2698 536218 -2614 536454
rect -2378 536218 23250 536454
rect 23486 536218 29514 536454
rect 29750 536218 51250 536454
rect 51486 536218 57514 536454
rect 57750 536218 79250 536454
rect 79486 536218 85514 536454
rect 85750 536218 107250 536454
rect 107486 536218 113514 536454
rect 113750 536218 135250 536454
rect 135486 536218 141514 536454
rect 141750 536218 163250 536454
rect 163486 536218 169514 536454
rect 169750 536218 191250 536454
rect 191486 536218 197514 536454
rect 197750 536218 219250 536454
rect 219486 536218 225514 536454
rect 225750 536218 247250 536454
rect 247486 536218 253514 536454
rect 253750 536218 275250 536454
rect 275486 536218 281514 536454
rect 281750 536218 303250 536454
rect 303486 536218 309514 536454
rect 309750 536218 331250 536454
rect 331486 536218 337514 536454
rect 337750 536218 359250 536454
rect 359486 536218 365514 536454
rect 365750 536218 387250 536454
rect 387486 536218 393514 536454
rect 393750 536218 415250 536454
rect 415486 536218 421514 536454
rect 421750 536218 443250 536454
rect 443486 536218 449514 536454
rect 449750 536218 471250 536454
rect 471486 536218 477514 536454
rect 477750 536218 499250 536454
rect 499486 536218 505514 536454
rect 505750 536218 527250 536454
rect 527486 536218 533514 536454
rect 533750 536218 555250 536454
rect 555486 536218 561514 536454
rect 561750 536218 586302 536454
rect 586538 536218 586622 536454
rect 586858 536218 592650 536454
rect -8726 536134 592650 536218
rect -8726 535898 -2934 536134
rect -2698 535898 -2614 536134
rect -2378 535898 23250 536134
rect 23486 535898 29514 536134
rect 29750 535898 51250 536134
rect 51486 535898 57514 536134
rect 57750 535898 79250 536134
rect 79486 535898 85514 536134
rect 85750 535898 107250 536134
rect 107486 535898 113514 536134
rect 113750 535898 135250 536134
rect 135486 535898 141514 536134
rect 141750 535898 163250 536134
rect 163486 535898 169514 536134
rect 169750 535898 191250 536134
rect 191486 535898 197514 536134
rect 197750 535898 219250 536134
rect 219486 535898 225514 536134
rect 225750 535898 247250 536134
rect 247486 535898 253514 536134
rect 253750 535898 275250 536134
rect 275486 535898 281514 536134
rect 281750 535898 303250 536134
rect 303486 535898 309514 536134
rect 309750 535898 331250 536134
rect 331486 535898 337514 536134
rect 337750 535898 359250 536134
rect 359486 535898 365514 536134
rect 365750 535898 387250 536134
rect 387486 535898 393514 536134
rect 393750 535898 415250 536134
rect 415486 535898 421514 536134
rect 421750 535898 443250 536134
rect 443486 535898 449514 536134
rect 449750 535898 471250 536134
rect 471486 535898 477514 536134
rect 477750 535898 499250 536134
rect 499486 535898 505514 536134
rect 505750 535898 527250 536134
rect 527486 535898 533514 536134
rect 533750 535898 555250 536134
rect 555486 535898 561514 536134
rect 561750 535898 586302 536134
rect 586538 535898 586622 536134
rect 586858 535898 592650 536134
rect -8726 535866 592650 535898
rect -8726 512829 592650 512861
rect -8726 512593 -1974 512829
rect -1738 512593 -1654 512829
rect -1418 512593 20118 512829
rect 20354 512593 26382 512829
rect 26618 512593 32646 512829
rect 32882 512593 48118 512829
rect 48354 512593 54382 512829
rect 54618 512593 60646 512829
rect 60882 512593 76118 512829
rect 76354 512593 82382 512829
rect 82618 512593 88646 512829
rect 88882 512593 104118 512829
rect 104354 512593 110382 512829
rect 110618 512593 116646 512829
rect 116882 512593 132118 512829
rect 132354 512593 138382 512829
rect 138618 512593 144646 512829
rect 144882 512593 160118 512829
rect 160354 512593 166382 512829
rect 166618 512593 172646 512829
rect 172882 512593 188118 512829
rect 188354 512593 194382 512829
rect 194618 512593 200646 512829
rect 200882 512593 216118 512829
rect 216354 512593 222382 512829
rect 222618 512593 228646 512829
rect 228882 512593 244118 512829
rect 244354 512593 250382 512829
rect 250618 512593 256646 512829
rect 256882 512593 272118 512829
rect 272354 512593 278382 512829
rect 278618 512593 284646 512829
rect 284882 512593 300118 512829
rect 300354 512593 306382 512829
rect 306618 512593 312646 512829
rect 312882 512593 328118 512829
rect 328354 512593 334382 512829
rect 334618 512593 340646 512829
rect 340882 512593 356118 512829
rect 356354 512593 362382 512829
rect 362618 512593 368646 512829
rect 368882 512593 384118 512829
rect 384354 512593 390382 512829
rect 390618 512593 396646 512829
rect 396882 512593 412118 512829
rect 412354 512593 418382 512829
rect 418618 512593 424646 512829
rect 424882 512593 440118 512829
rect 440354 512593 446382 512829
rect 446618 512593 452646 512829
rect 452882 512593 468118 512829
rect 468354 512593 474382 512829
rect 474618 512593 480646 512829
rect 480882 512593 496118 512829
rect 496354 512593 502382 512829
rect 502618 512593 508646 512829
rect 508882 512593 524118 512829
rect 524354 512593 530382 512829
rect 530618 512593 536646 512829
rect 536882 512593 552118 512829
rect 552354 512593 558382 512829
rect 558618 512593 564646 512829
rect 564882 512593 573526 512829
rect 573762 512593 573846 512829
rect 574082 512593 585342 512829
rect 585578 512593 585662 512829
rect 585898 512593 592650 512829
rect -8726 512509 592650 512593
rect -8726 512273 -1974 512509
rect -1738 512273 -1654 512509
rect -1418 512273 20118 512509
rect 20354 512273 26382 512509
rect 26618 512273 32646 512509
rect 32882 512273 48118 512509
rect 48354 512273 54382 512509
rect 54618 512273 60646 512509
rect 60882 512273 76118 512509
rect 76354 512273 82382 512509
rect 82618 512273 88646 512509
rect 88882 512273 104118 512509
rect 104354 512273 110382 512509
rect 110618 512273 116646 512509
rect 116882 512273 132118 512509
rect 132354 512273 138382 512509
rect 138618 512273 144646 512509
rect 144882 512273 160118 512509
rect 160354 512273 166382 512509
rect 166618 512273 172646 512509
rect 172882 512273 188118 512509
rect 188354 512273 194382 512509
rect 194618 512273 200646 512509
rect 200882 512273 216118 512509
rect 216354 512273 222382 512509
rect 222618 512273 228646 512509
rect 228882 512273 244118 512509
rect 244354 512273 250382 512509
rect 250618 512273 256646 512509
rect 256882 512273 272118 512509
rect 272354 512273 278382 512509
rect 278618 512273 284646 512509
rect 284882 512273 300118 512509
rect 300354 512273 306382 512509
rect 306618 512273 312646 512509
rect 312882 512273 328118 512509
rect 328354 512273 334382 512509
rect 334618 512273 340646 512509
rect 340882 512273 356118 512509
rect 356354 512273 362382 512509
rect 362618 512273 368646 512509
rect 368882 512273 384118 512509
rect 384354 512273 390382 512509
rect 390618 512273 396646 512509
rect 396882 512273 412118 512509
rect 412354 512273 418382 512509
rect 418618 512273 424646 512509
rect 424882 512273 440118 512509
rect 440354 512273 446382 512509
rect 446618 512273 452646 512509
rect 452882 512273 468118 512509
rect 468354 512273 474382 512509
rect 474618 512273 480646 512509
rect 480882 512273 496118 512509
rect 496354 512273 502382 512509
rect 502618 512273 508646 512509
rect 508882 512273 524118 512509
rect 524354 512273 530382 512509
rect 530618 512273 536646 512509
rect 536882 512273 552118 512509
rect 552354 512273 558382 512509
rect 558618 512273 564646 512509
rect 564882 512273 573526 512509
rect 573762 512273 573846 512509
rect 574082 512273 585342 512509
rect 585578 512273 585662 512509
rect 585898 512273 592650 512509
rect -8726 512241 592650 512273
rect -8726 509454 592650 509486
rect -8726 509218 -2934 509454
rect -2698 509218 -2614 509454
rect -2378 509218 23250 509454
rect 23486 509218 29514 509454
rect 29750 509218 51250 509454
rect 51486 509218 57514 509454
rect 57750 509218 79250 509454
rect 79486 509218 85514 509454
rect 85750 509218 107250 509454
rect 107486 509218 113514 509454
rect 113750 509218 135250 509454
rect 135486 509218 141514 509454
rect 141750 509218 163250 509454
rect 163486 509218 169514 509454
rect 169750 509218 191250 509454
rect 191486 509218 197514 509454
rect 197750 509218 219250 509454
rect 219486 509218 225514 509454
rect 225750 509218 247250 509454
rect 247486 509218 253514 509454
rect 253750 509218 275250 509454
rect 275486 509218 281514 509454
rect 281750 509218 303250 509454
rect 303486 509218 309514 509454
rect 309750 509218 331250 509454
rect 331486 509218 337514 509454
rect 337750 509218 359250 509454
rect 359486 509218 365514 509454
rect 365750 509218 387250 509454
rect 387486 509218 393514 509454
rect 393750 509218 415250 509454
rect 415486 509218 421514 509454
rect 421750 509218 443250 509454
rect 443486 509218 449514 509454
rect 449750 509218 471250 509454
rect 471486 509218 477514 509454
rect 477750 509218 499250 509454
rect 499486 509218 505514 509454
rect 505750 509218 527250 509454
rect 527486 509218 533514 509454
rect 533750 509218 555250 509454
rect 555486 509218 561514 509454
rect 561750 509218 586302 509454
rect 586538 509218 586622 509454
rect 586858 509218 592650 509454
rect -8726 509134 592650 509218
rect -8726 508898 -2934 509134
rect -2698 508898 -2614 509134
rect -2378 508898 23250 509134
rect 23486 508898 29514 509134
rect 29750 508898 51250 509134
rect 51486 508898 57514 509134
rect 57750 508898 79250 509134
rect 79486 508898 85514 509134
rect 85750 508898 107250 509134
rect 107486 508898 113514 509134
rect 113750 508898 135250 509134
rect 135486 508898 141514 509134
rect 141750 508898 163250 509134
rect 163486 508898 169514 509134
rect 169750 508898 191250 509134
rect 191486 508898 197514 509134
rect 197750 508898 219250 509134
rect 219486 508898 225514 509134
rect 225750 508898 247250 509134
rect 247486 508898 253514 509134
rect 253750 508898 275250 509134
rect 275486 508898 281514 509134
rect 281750 508898 303250 509134
rect 303486 508898 309514 509134
rect 309750 508898 331250 509134
rect 331486 508898 337514 509134
rect 337750 508898 359250 509134
rect 359486 508898 365514 509134
rect 365750 508898 387250 509134
rect 387486 508898 393514 509134
rect 393750 508898 415250 509134
rect 415486 508898 421514 509134
rect 421750 508898 443250 509134
rect 443486 508898 449514 509134
rect 449750 508898 471250 509134
rect 471486 508898 477514 509134
rect 477750 508898 499250 509134
rect 499486 508898 505514 509134
rect 505750 508898 527250 509134
rect 527486 508898 533514 509134
rect 533750 508898 555250 509134
rect 555486 508898 561514 509134
rect 561750 508898 586302 509134
rect 586538 508898 586622 509134
rect 586858 508898 592650 509134
rect -8726 508866 592650 508898
rect -8726 485829 592650 485861
rect -8726 485593 -1974 485829
rect -1738 485593 -1654 485829
rect -1418 485593 20118 485829
rect 20354 485593 26382 485829
rect 26618 485593 32646 485829
rect 32882 485593 48118 485829
rect 48354 485593 54382 485829
rect 54618 485593 60646 485829
rect 60882 485593 76118 485829
rect 76354 485593 82382 485829
rect 82618 485593 88646 485829
rect 88882 485593 104118 485829
rect 104354 485593 110382 485829
rect 110618 485593 116646 485829
rect 116882 485593 132118 485829
rect 132354 485593 138382 485829
rect 138618 485593 144646 485829
rect 144882 485593 160118 485829
rect 160354 485593 166382 485829
rect 166618 485593 172646 485829
rect 172882 485593 188118 485829
rect 188354 485593 194382 485829
rect 194618 485593 200646 485829
rect 200882 485593 216118 485829
rect 216354 485593 222382 485829
rect 222618 485593 228646 485829
rect 228882 485593 244118 485829
rect 244354 485593 250382 485829
rect 250618 485593 256646 485829
rect 256882 485593 272118 485829
rect 272354 485593 278382 485829
rect 278618 485593 284646 485829
rect 284882 485593 300118 485829
rect 300354 485593 306382 485829
rect 306618 485593 312646 485829
rect 312882 485593 328118 485829
rect 328354 485593 334382 485829
rect 334618 485593 340646 485829
rect 340882 485593 356118 485829
rect 356354 485593 362382 485829
rect 362618 485593 368646 485829
rect 368882 485593 384118 485829
rect 384354 485593 390382 485829
rect 390618 485593 396646 485829
rect 396882 485593 412118 485829
rect 412354 485593 418382 485829
rect 418618 485593 424646 485829
rect 424882 485593 440118 485829
rect 440354 485593 446382 485829
rect 446618 485593 452646 485829
rect 452882 485593 468118 485829
rect 468354 485593 474382 485829
rect 474618 485593 480646 485829
rect 480882 485593 496118 485829
rect 496354 485593 502382 485829
rect 502618 485593 508646 485829
rect 508882 485593 524118 485829
rect 524354 485593 530382 485829
rect 530618 485593 536646 485829
rect 536882 485593 552118 485829
rect 552354 485593 558382 485829
rect 558618 485593 564646 485829
rect 564882 485593 573526 485829
rect 573762 485593 573846 485829
rect 574082 485593 585342 485829
rect 585578 485593 585662 485829
rect 585898 485593 592650 485829
rect -8726 485509 592650 485593
rect -8726 485273 -1974 485509
rect -1738 485273 -1654 485509
rect -1418 485273 20118 485509
rect 20354 485273 26382 485509
rect 26618 485273 32646 485509
rect 32882 485273 48118 485509
rect 48354 485273 54382 485509
rect 54618 485273 60646 485509
rect 60882 485273 76118 485509
rect 76354 485273 82382 485509
rect 82618 485273 88646 485509
rect 88882 485273 104118 485509
rect 104354 485273 110382 485509
rect 110618 485273 116646 485509
rect 116882 485273 132118 485509
rect 132354 485273 138382 485509
rect 138618 485273 144646 485509
rect 144882 485273 160118 485509
rect 160354 485273 166382 485509
rect 166618 485273 172646 485509
rect 172882 485273 188118 485509
rect 188354 485273 194382 485509
rect 194618 485273 200646 485509
rect 200882 485273 216118 485509
rect 216354 485273 222382 485509
rect 222618 485273 228646 485509
rect 228882 485273 244118 485509
rect 244354 485273 250382 485509
rect 250618 485273 256646 485509
rect 256882 485273 272118 485509
rect 272354 485273 278382 485509
rect 278618 485273 284646 485509
rect 284882 485273 300118 485509
rect 300354 485273 306382 485509
rect 306618 485273 312646 485509
rect 312882 485273 328118 485509
rect 328354 485273 334382 485509
rect 334618 485273 340646 485509
rect 340882 485273 356118 485509
rect 356354 485273 362382 485509
rect 362618 485273 368646 485509
rect 368882 485273 384118 485509
rect 384354 485273 390382 485509
rect 390618 485273 396646 485509
rect 396882 485273 412118 485509
rect 412354 485273 418382 485509
rect 418618 485273 424646 485509
rect 424882 485273 440118 485509
rect 440354 485273 446382 485509
rect 446618 485273 452646 485509
rect 452882 485273 468118 485509
rect 468354 485273 474382 485509
rect 474618 485273 480646 485509
rect 480882 485273 496118 485509
rect 496354 485273 502382 485509
rect 502618 485273 508646 485509
rect 508882 485273 524118 485509
rect 524354 485273 530382 485509
rect 530618 485273 536646 485509
rect 536882 485273 552118 485509
rect 552354 485273 558382 485509
rect 558618 485273 564646 485509
rect 564882 485273 573526 485509
rect 573762 485273 573846 485509
rect 574082 485273 585342 485509
rect 585578 485273 585662 485509
rect 585898 485273 592650 485509
rect -8726 485241 592650 485273
rect -8726 482454 592650 482486
rect -8726 482218 -2934 482454
rect -2698 482218 -2614 482454
rect -2378 482218 23250 482454
rect 23486 482218 29514 482454
rect 29750 482218 51250 482454
rect 51486 482218 57514 482454
rect 57750 482218 79250 482454
rect 79486 482218 85514 482454
rect 85750 482218 107250 482454
rect 107486 482218 113514 482454
rect 113750 482218 135250 482454
rect 135486 482218 141514 482454
rect 141750 482218 163250 482454
rect 163486 482218 169514 482454
rect 169750 482218 191250 482454
rect 191486 482218 197514 482454
rect 197750 482218 219250 482454
rect 219486 482218 225514 482454
rect 225750 482218 247250 482454
rect 247486 482218 253514 482454
rect 253750 482218 275250 482454
rect 275486 482218 281514 482454
rect 281750 482218 303250 482454
rect 303486 482218 309514 482454
rect 309750 482218 331250 482454
rect 331486 482218 337514 482454
rect 337750 482218 359250 482454
rect 359486 482218 365514 482454
rect 365750 482218 387250 482454
rect 387486 482218 393514 482454
rect 393750 482218 415250 482454
rect 415486 482218 421514 482454
rect 421750 482218 443250 482454
rect 443486 482218 449514 482454
rect 449750 482218 471250 482454
rect 471486 482218 477514 482454
rect 477750 482218 499250 482454
rect 499486 482218 505514 482454
rect 505750 482218 527250 482454
rect 527486 482218 533514 482454
rect 533750 482218 555250 482454
rect 555486 482218 561514 482454
rect 561750 482218 586302 482454
rect 586538 482218 586622 482454
rect 586858 482218 592650 482454
rect -8726 482134 592650 482218
rect -8726 481898 -2934 482134
rect -2698 481898 -2614 482134
rect -2378 481898 23250 482134
rect 23486 481898 29514 482134
rect 29750 481898 51250 482134
rect 51486 481898 57514 482134
rect 57750 481898 79250 482134
rect 79486 481898 85514 482134
rect 85750 481898 107250 482134
rect 107486 481898 113514 482134
rect 113750 481898 135250 482134
rect 135486 481898 141514 482134
rect 141750 481898 163250 482134
rect 163486 481898 169514 482134
rect 169750 481898 191250 482134
rect 191486 481898 197514 482134
rect 197750 481898 219250 482134
rect 219486 481898 225514 482134
rect 225750 481898 247250 482134
rect 247486 481898 253514 482134
rect 253750 481898 275250 482134
rect 275486 481898 281514 482134
rect 281750 481898 303250 482134
rect 303486 481898 309514 482134
rect 309750 481898 331250 482134
rect 331486 481898 337514 482134
rect 337750 481898 359250 482134
rect 359486 481898 365514 482134
rect 365750 481898 387250 482134
rect 387486 481898 393514 482134
rect 393750 481898 415250 482134
rect 415486 481898 421514 482134
rect 421750 481898 443250 482134
rect 443486 481898 449514 482134
rect 449750 481898 471250 482134
rect 471486 481898 477514 482134
rect 477750 481898 499250 482134
rect 499486 481898 505514 482134
rect 505750 481898 527250 482134
rect 527486 481898 533514 482134
rect 533750 481898 555250 482134
rect 555486 481898 561514 482134
rect 561750 481898 586302 482134
rect 586538 481898 586622 482134
rect 586858 481898 592650 482134
rect -8726 481866 592650 481898
rect -8726 458829 592650 458861
rect -8726 458593 -1974 458829
rect -1738 458593 -1654 458829
rect -1418 458593 20118 458829
rect 20354 458593 26382 458829
rect 26618 458593 32646 458829
rect 32882 458593 48118 458829
rect 48354 458593 54382 458829
rect 54618 458593 60646 458829
rect 60882 458593 76118 458829
rect 76354 458593 82382 458829
rect 82618 458593 88646 458829
rect 88882 458593 104118 458829
rect 104354 458593 110382 458829
rect 110618 458593 116646 458829
rect 116882 458593 132118 458829
rect 132354 458593 138382 458829
rect 138618 458593 144646 458829
rect 144882 458593 160118 458829
rect 160354 458593 166382 458829
rect 166618 458593 172646 458829
rect 172882 458593 188118 458829
rect 188354 458593 194382 458829
rect 194618 458593 200646 458829
rect 200882 458593 216118 458829
rect 216354 458593 222382 458829
rect 222618 458593 228646 458829
rect 228882 458593 244118 458829
rect 244354 458593 250382 458829
rect 250618 458593 256646 458829
rect 256882 458593 272118 458829
rect 272354 458593 278382 458829
rect 278618 458593 284646 458829
rect 284882 458593 300118 458829
rect 300354 458593 306382 458829
rect 306618 458593 312646 458829
rect 312882 458593 328118 458829
rect 328354 458593 334382 458829
rect 334618 458593 340646 458829
rect 340882 458593 356118 458829
rect 356354 458593 362382 458829
rect 362618 458593 368646 458829
rect 368882 458593 384118 458829
rect 384354 458593 390382 458829
rect 390618 458593 396646 458829
rect 396882 458593 412118 458829
rect 412354 458593 418382 458829
rect 418618 458593 424646 458829
rect 424882 458593 440118 458829
rect 440354 458593 446382 458829
rect 446618 458593 452646 458829
rect 452882 458593 468118 458829
rect 468354 458593 474382 458829
rect 474618 458593 480646 458829
rect 480882 458593 496118 458829
rect 496354 458593 502382 458829
rect 502618 458593 508646 458829
rect 508882 458593 524118 458829
rect 524354 458593 530382 458829
rect 530618 458593 536646 458829
rect 536882 458593 552118 458829
rect 552354 458593 558382 458829
rect 558618 458593 564646 458829
rect 564882 458593 573526 458829
rect 573762 458593 573846 458829
rect 574082 458593 585342 458829
rect 585578 458593 585662 458829
rect 585898 458593 592650 458829
rect -8726 458509 592650 458593
rect -8726 458273 -1974 458509
rect -1738 458273 -1654 458509
rect -1418 458273 20118 458509
rect 20354 458273 26382 458509
rect 26618 458273 32646 458509
rect 32882 458273 48118 458509
rect 48354 458273 54382 458509
rect 54618 458273 60646 458509
rect 60882 458273 76118 458509
rect 76354 458273 82382 458509
rect 82618 458273 88646 458509
rect 88882 458273 104118 458509
rect 104354 458273 110382 458509
rect 110618 458273 116646 458509
rect 116882 458273 132118 458509
rect 132354 458273 138382 458509
rect 138618 458273 144646 458509
rect 144882 458273 160118 458509
rect 160354 458273 166382 458509
rect 166618 458273 172646 458509
rect 172882 458273 188118 458509
rect 188354 458273 194382 458509
rect 194618 458273 200646 458509
rect 200882 458273 216118 458509
rect 216354 458273 222382 458509
rect 222618 458273 228646 458509
rect 228882 458273 244118 458509
rect 244354 458273 250382 458509
rect 250618 458273 256646 458509
rect 256882 458273 272118 458509
rect 272354 458273 278382 458509
rect 278618 458273 284646 458509
rect 284882 458273 300118 458509
rect 300354 458273 306382 458509
rect 306618 458273 312646 458509
rect 312882 458273 328118 458509
rect 328354 458273 334382 458509
rect 334618 458273 340646 458509
rect 340882 458273 356118 458509
rect 356354 458273 362382 458509
rect 362618 458273 368646 458509
rect 368882 458273 384118 458509
rect 384354 458273 390382 458509
rect 390618 458273 396646 458509
rect 396882 458273 412118 458509
rect 412354 458273 418382 458509
rect 418618 458273 424646 458509
rect 424882 458273 440118 458509
rect 440354 458273 446382 458509
rect 446618 458273 452646 458509
rect 452882 458273 468118 458509
rect 468354 458273 474382 458509
rect 474618 458273 480646 458509
rect 480882 458273 496118 458509
rect 496354 458273 502382 458509
rect 502618 458273 508646 458509
rect 508882 458273 524118 458509
rect 524354 458273 530382 458509
rect 530618 458273 536646 458509
rect 536882 458273 552118 458509
rect 552354 458273 558382 458509
rect 558618 458273 564646 458509
rect 564882 458273 573526 458509
rect 573762 458273 573846 458509
rect 574082 458273 585342 458509
rect 585578 458273 585662 458509
rect 585898 458273 592650 458509
rect -8726 458241 592650 458273
rect -8726 455454 592650 455486
rect -8726 455218 -2934 455454
rect -2698 455218 -2614 455454
rect -2378 455218 23250 455454
rect 23486 455218 29514 455454
rect 29750 455218 51250 455454
rect 51486 455218 57514 455454
rect 57750 455218 79250 455454
rect 79486 455218 85514 455454
rect 85750 455218 107250 455454
rect 107486 455218 113514 455454
rect 113750 455218 135250 455454
rect 135486 455218 141514 455454
rect 141750 455218 163250 455454
rect 163486 455218 169514 455454
rect 169750 455218 191250 455454
rect 191486 455218 197514 455454
rect 197750 455218 219250 455454
rect 219486 455218 225514 455454
rect 225750 455218 247250 455454
rect 247486 455218 253514 455454
rect 253750 455218 275250 455454
rect 275486 455218 281514 455454
rect 281750 455218 303250 455454
rect 303486 455218 309514 455454
rect 309750 455218 331250 455454
rect 331486 455218 337514 455454
rect 337750 455218 359250 455454
rect 359486 455218 365514 455454
rect 365750 455218 387250 455454
rect 387486 455218 393514 455454
rect 393750 455218 415250 455454
rect 415486 455218 421514 455454
rect 421750 455218 443250 455454
rect 443486 455218 449514 455454
rect 449750 455218 471250 455454
rect 471486 455218 477514 455454
rect 477750 455218 499250 455454
rect 499486 455218 505514 455454
rect 505750 455218 527250 455454
rect 527486 455218 533514 455454
rect 533750 455218 555250 455454
rect 555486 455218 561514 455454
rect 561750 455218 586302 455454
rect 586538 455218 586622 455454
rect 586858 455218 592650 455454
rect -8726 455134 592650 455218
rect -8726 454898 -2934 455134
rect -2698 454898 -2614 455134
rect -2378 454898 23250 455134
rect 23486 454898 29514 455134
rect 29750 454898 51250 455134
rect 51486 454898 57514 455134
rect 57750 454898 79250 455134
rect 79486 454898 85514 455134
rect 85750 454898 107250 455134
rect 107486 454898 113514 455134
rect 113750 454898 135250 455134
rect 135486 454898 141514 455134
rect 141750 454898 163250 455134
rect 163486 454898 169514 455134
rect 169750 454898 191250 455134
rect 191486 454898 197514 455134
rect 197750 454898 219250 455134
rect 219486 454898 225514 455134
rect 225750 454898 247250 455134
rect 247486 454898 253514 455134
rect 253750 454898 275250 455134
rect 275486 454898 281514 455134
rect 281750 454898 303250 455134
rect 303486 454898 309514 455134
rect 309750 454898 331250 455134
rect 331486 454898 337514 455134
rect 337750 454898 359250 455134
rect 359486 454898 365514 455134
rect 365750 454898 387250 455134
rect 387486 454898 393514 455134
rect 393750 454898 415250 455134
rect 415486 454898 421514 455134
rect 421750 454898 443250 455134
rect 443486 454898 449514 455134
rect 449750 454898 471250 455134
rect 471486 454898 477514 455134
rect 477750 454898 499250 455134
rect 499486 454898 505514 455134
rect 505750 454898 527250 455134
rect 527486 454898 533514 455134
rect 533750 454898 555250 455134
rect 555486 454898 561514 455134
rect 561750 454898 586302 455134
rect 586538 454898 586622 455134
rect 586858 454898 592650 455134
rect -8726 454866 592650 454898
rect -8726 431829 592650 431861
rect -8726 431593 -1974 431829
rect -1738 431593 -1654 431829
rect -1418 431593 20118 431829
rect 20354 431593 26382 431829
rect 26618 431593 32646 431829
rect 32882 431593 48118 431829
rect 48354 431593 54382 431829
rect 54618 431593 60646 431829
rect 60882 431593 76118 431829
rect 76354 431593 82382 431829
rect 82618 431593 88646 431829
rect 88882 431593 104118 431829
rect 104354 431593 110382 431829
rect 110618 431593 116646 431829
rect 116882 431593 132118 431829
rect 132354 431593 138382 431829
rect 138618 431593 144646 431829
rect 144882 431593 160118 431829
rect 160354 431593 166382 431829
rect 166618 431593 172646 431829
rect 172882 431593 188118 431829
rect 188354 431593 194382 431829
rect 194618 431593 200646 431829
rect 200882 431593 216118 431829
rect 216354 431593 222382 431829
rect 222618 431593 228646 431829
rect 228882 431593 244118 431829
rect 244354 431593 250382 431829
rect 250618 431593 256646 431829
rect 256882 431593 272118 431829
rect 272354 431593 278382 431829
rect 278618 431593 284646 431829
rect 284882 431593 300118 431829
rect 300354 431593 306382 431829
rect 306618 431593 312646 431829
rect 312882 431593 328118 431829
rect 328354 431593 334382 431829
rect 334618 431593 340646 431829
rect 340882 431593 356118 431829
rect 356354 431593 362382 431829
rect 362618 431593 368646 431829
rect 368882 431593 384118 431829
rect 384354 431593 390382 431829
rect 390618 431593 396646 431829
rect 396882 431593 412118 431829
rect 412354 431593 418382 431829
rect 418618 431593 424646 431829
rect 424882 431593 440118 431829
rect 440354 431593 446382 431829
rect 446618 431593 452646 431829
rect 452882 431593 468118 431829
rect 468354 431593 474382 431829
rect 474618 431593 480646 431829
rect 480882 431593 496118 431829
rect 496354 431593 502382 431829
rect 502618 431593 508646 431829
rect 508882 431593 524118 431829
rect 524354 431593 530382 431829
rect 530618 431593 536646 431829
rect 536882 431593 552118 431829
rect 552354 431593 558382 431829
rect 558618 431593 564646 431829
rect 564882 431593 573526 431829
rect 573762 431593 573846 431829
rect 574082 431593 585342 431829
rect 585578 431593 585662 431829
rect 585898 431593 592650 431829
rect -8726 431509 592650 431593
rect -8726 431273 -1974 431509
rect -1738 431273 -1654 431509
rect -1418 431273 20118 431509
rect 20354 431273 26382 431509
rect 26618 431273 32646 431509
rect 32882 431273 48118 431509
rect 48354 431273 54382 431509
rect 54618 431273 60646 431509
rect 60882 431273 76118 431509
rect 76354 431273 82382 431509
rect 82618 431273 88646 431509
rect 88882 431273 104118 431509
rect 104354 431273 110382 431509
rect 110618 431273 116646 431509
rect 116882 431273 132118 431509
rect 132354 431273 138382 431509
rect 138618 431273 144646 431509
rect 144882 431273 160118 431509
rect 160354 431273 166382 431509
rect 166618 431273 172646 431509
rect 172882 431273 188118 431509
rect 188354 431273 194382 431509
rect 194618 431273 200646 431509
rect 200882 431273 216118 431509
rect 216354 431273 222382 431509
rect 222618 431273 228646 431509
rect 228882 431273 244118 431509
rect 244354 431273 250382 431509
rect 250618 431273 256646 431509
rect 256882 431273 272118 431509
rect 272354 431273 278382 431509
rect 278618 431273 284646 431509
rect 284882 431273 300118 431509
rect 300354 431273 306382 431509
rect 306618 431273 312646 431509
rect 312882 431273 328118 431509
rect 328354 431273 334382 431509
rect 334618 431273 340646 431509
rect 340882 431273 356118 431509
rect 356354 431273 362382 431509
rect 362618 431273 368646 431509
rect 368882 431273 384118 431509
rect 384354 431273 390382 431509
rect 390618 431273 396646 431509
rect 396882 431273 412118 431509
rect 412354 431273 418382 431509
rect 418618 431273 424646 431509
rect 424882 431273 440118 431509
rect 440354 431273 446382 431509
rect 446618 431273 452646 431509
rect 452882 431273 468118 431509
rect 468354 431273 474382 431509
rect 474618 431273 480646 431509
rect 480882 431273 496118 431509
rect 496354 431273 502382 431509
rect 502618 431273 508646 431509
rect 508882 431273 524118 431509
rect 524354 431273 530382 431509
rect 530618 431273 536646 431509
rect 536882 431273 552118 431509
rect 552354 431273 558382 431509
rect 558618 431273 564646 431509
rect 564882 431273 573526 431509
rect 573762 431273 573846 431509
rect 574082 431273 585342 431509
rect 585578 431273 585662 431509
rect 585898 431273 592650 431509
rect -8726 431241 592650 431273
rect -8726 428454 592650 428486
rect -8726 428218 -2934 428454
rect -2698 428218 -2614 428454
rect -2378 428218 23250 428454
rect 23486 428218 29514 428454
rect 29750 428218 51250 428454
rect 51486 428218 57514 428454
rect 57750 428218 79250 428454
rect 79486 428218 85514 428454
rect 85750 428218 107250 428454
rect 107486 428218 113514 428454
rect 113750 428218 135250 428454
rect 135486 428218 141514 428454
rect 141750 428218 163250 428454
rect 163486 428218 169514 428454
rect 169750 428218 191250 428454
rect 191486 428218 197514 428454
rect 197750 428218 219250 428454
rect 219486 428218 225514 428454
rect 225750 428218 247250 428454
rect 247486 428218 253514 428454
rect 253750 428218 275250 428454
rect 275486 428218 281514 428454
rect 281750 428218 303250 428454
rect 303486 428218 309514 428454
rect 309750 428218 331250 428454
rect 331486 428218 337514 428454
rect 337750 428218 359250 428454
rect 359486 428218 365514 428454
rect 365750 428218 387250 428454
rect 387486 428218 393514 428454
rect 393750 428218 415250 428454
rect 415486 428218 421514 428454
rect 421750 428218 443250 428454
rect 443486 428218 449514 428454
rect 449750 428218 471250 428454
rect 471486 428218 477514 428454
rect 477750 428218 499250 428454
rect 499486 428218 505514 428454
rect 505750 428218 527250 428454
rect 527486 428218 533514 428454
rect 533750 428218 555250 428454
rect 555486 428218 561514 428454
rect 561750 428218 586302 428454
rect 586538 428218 586622 428454
rect 586858 428218 592650 428454
rect -8726 428134 592650 428218
rect -8726 427898 -2934 428134
rect -2698 427898 -2614 428134
rect -2378 427898 23250 428134
rect 23486 427898 29514 428134
rect 29750 427898 51250 428134
rect 51486 427898 57514 428134
rect 57750 427898 79250 428134
rect 79486 427898 85514 428134
rect 85750 427898 107250 428134
rect 107486 427898 113514 428134
rect 113750 427898 135250 428134
rect 135486 427898 141514 428134
rect 141750 427898 163250 428134
rect 163486 427898 169514 428134
rect 169750 427898 191250 428134
rect 191486 427898 197514 428134
rect 197750 427898 219250 428134
rect 219486 427898 225514 428134
rect 225750 427898 247250 428134
rect 247486 427898 253514 428134
rect 253750 427898 275250 428134
rect 275486 427898 281514 428134
rect 281750 427898 303250 428134
rect 303486 427898 309514 428134
rect 309750 427898 331250 428134
rect 331486 427898 337514 428134
rect 337750 427898 359250 428134
rect 359486 427898 365514 428134
rect 365750 427898 387250 428134
rect 387486 427898 393514 428134
rect 393750 427898 415250 428134
rect 415486 427898 421514 428134
rect 421750 427898 443250 428134
rect 443486 427898 449514 428134
rect 449750 427898 471250 428134
rect 471486 427898 477514 428134
rect 477750 427898 499250 428134
rect 499486 427898 505514 428134
rect 505750 427898 527250 428134
rect 527486 427898 533514 428134
rect 533750 427898 555250 428134
rect 555486 427898 561514 428134
rect 561750 427898 586302 428134
rect 586538 427898 586622 428134
rect 586858 427898 592650 428134
rect -8726 427866 592650 427898
rect -8726 404829 592650 404861
rect -8726 404593 -1974 404829
rect -1738 404593 -1654 404829
rect -1418 404593 20118 404829
rect 20354 404593 26382 404829
rect 26618 404593 32646 404829
rect 32882 404593 48118 404829
rect 48354 404593 54382 404829
rect 54618 404593 60646 404829
rect 60882 404593 76118 404829
rect 76354 404593 82382 404829
rect 82618 404593 88646 404829
rect 88882 404593 104118 404829
rect 104354 404593 110382 404829
rect 110618 404593 116646 404829
rect 116882 404593 132118 404829
rect 132354 404593 138382 404829
rect 138618 404593 144646 404829
rect 144882 404593 160118 404829
rect 160354 404593 166382 404829
rect 166618 404593 172646 404829
rect 172882 404593 188118 404829
rect 188354 404593 194382 404829
rect 194618 404593 200646 404829
rect 200882 404593 216118 404829
rect 216354 404593 222382 404829
rect 222618 404593 228646 404829
rect 228882 404593 244118 404829
rect 244354 404593 250382 404829
rect 250618 404593 256646 404829
rect 256882 404593 272118 404829
rect 272354 404593 278382 404829
rect 278618 404593 284646 404829
rect 284882 404593 300118 404829
rect 300354 404593 306382 404829
rect 306618 404593 312646 404829
rect 312882 404593 328118 404829
rect 328354 404593 334382 404829
rect 334618 404593 340646 404829
rect 340882 404593 356118 404829
rect 356354 404593 362382 404829
rect 362618 404593 368646 404829
rect 368882 404593 384118 404829
rect 384354 404593 390382 404829
rect 390618 404593 396646 404829
rect 396882 404593 412118 404829
rect 412354 404593 418382 404829
rect 418618 404593 424646 404829
rect 424882 404593 440118 404829
rect 440354 404593 446382 404829
rect 446618 404593 452646 404829
rect 452882 404593 468118 404829
rect 468354 404593 474382 404829
rect 474618 404593 480646 404829
rect 480882 404593 496118 404829
rect 496354 404593 502382 404829
rect 502618 404593 508646 404829
rect 508882 404593 524118 404829
rect 524354 404593 530382 404829
rect 530618 404593 536646 404829
rect 536882 404593 552118 404829
rect 552354 404593 558382 404829
rect 558618 404593 564646 404829
rect 564882 404593 573526 404829
rect 573762 404593 573846 404829
rect 574082 404593 585342 404829
rect 585578 404593 585662 404829
rect 585898 404593 592650 404829
rect -8726 404509 592650 404593
rect -8726 404273 -1974 404509
rect -1738 404273 -1654 404509
rect -1418 404273 20118 404509
rect 20354 404273 26382 404509
rect 26618 404273 32646 404509
rect 32882 404273 48118 404509
rect 48354 404273 54382 404509
rect 54618 404273 60646 404509
rect 60882 404273 76118 404509
rect 76354 404273 82382 404509
rect 82618 404273 88646 404509
rect 88882 404273 104118 404509
rect 104354 404273 110382 404509
rect 110618 404273 116646 404509
rect 116882 404273 132118 404509
rect 132354 404273 138382 404509
rect 138618 404273 144646 404509
rect 144882 404273 160118 404509
rect 160354 404273 166382 404509
rect 166618 404273 172646 404509
rect 172882 404273 188118 404509
rect 188354 404273 194382 404509
rect 194618 404273 200646 404509
rect 200882 404273 216118 404509
rect 216354 404273 222382 404509
rect 222618 404273 228646 404509
rect 228882 404273 244118 404509
rect 244354 404273 250382 404509
rect 250618 404273 256646 404509
rect 256882 404273 272118 404509
rect 272354 404273 278382 404509
rect 278618 404273 284646 404509
rect 284882 404273 300118 404509
rect 300354 404273 306382 404509
rect 306618 404273 312646 404509
rect 312882 404273 328118 404509
rect 328354 404273 334382 404509
rect 334618 404273 340646 404509
rect 340882 404273 356118 404509
rect 356354 404273 362382 404509
rect 362618 404273 368646 404509
rect 368882 404273 384118 404509
rect 384354 404273 390382 404509
rect 390618 404273 396646 404509
rect 396882 404273 412118 404509
rect 412354 404273 418382 404509
rect 418618 404273 424646 404509
rect 424882 404273 440118 404509
rect 440354 404273 446382 404509
rect 446618 404273 452646 404509
rect 452882 404273 468118 404509
rect 468354 404273 474382 404509
rect 474618 404273 480646 404509
rect 480882 404273 496118 404509
rect 496354 404273 502382 404509
rect 502618 404273 508646 404509
rect 508882 404273 524118 404509
rect 524354 404273 530382 404509
rect 530618 404273 536646 404509
rect 536882 404273 552118 404509
rect 552354 404273 558382 404509
rect 558618 404273 564646 404509
rect 564882 404273 573526 404509
rect 573762 404273 573846 404509
rect 574082 404273 585342 404509
rect 585578 404273 585662 404509
rect 585898 404273 592650 404509
rect -8726 404241 592650 404273
rect -8726 401454 592650 401486
rect -8726 401218 -2934 401454
rect -2698 401218 -2614 401454
rect -2378 401218 23250 401454
rect 23486 401218 29514 401454
rect 29750 401218 51250 401454
rect 51486 401218 57514 401454
rect 57750 401218 79250 401454
rect 79486 401218 85514 401454
rect 85750 401218 107250 401454
rect 107486 401218 113514 401454
rect 113750 401218 135250 401454
rect 135486 401218 141514 401454
rect 141750 401218 163250 401454
rect 163486 401218 169514 401454
rect 169750 401218 191250 401454
rect 191486 401218 197514 401454
rect 197750 401218 219250 401454
rect 219486 401218 225514 401454
rect 225750 401218 247250 401454
rect 247486 401218 253514 401454
rect 253750 401218 275250 401454
rect 275486 401218 281514 401454
rect 281750 401218 303250 401454
rect 303486 401218 309514 401454
rect 309750 401218 331250 401454
rect 331486 401218 337514 401454
rect 337750 401218 359250 401454
rect 359486 401218 365514 401454
rect 365750 401218 387250 401454
rect 387486 401218 393514 401454
rect 393750 401218 415250 401454
rect 415486 401218 421514 401454
rect 421750 401218 443250 401454
rect 443486 401218 449514 401454
rect 449750 401218 471250 401454
rect 471486 401218 477514 401454
rect 477750 401218 499250 401454
rect 499486 401218 505514 401454
rect 505750 401218 527250 401454
rect 527486 401218 533514 401454
rect 533750 401218 555250 401454
rect 555486 401218 561514 401454
rect 561750 401218 586302 401454
rect 586538 401218 586622 401454
rect 586858 401218 592650 401454
rect -8726 401134 592650 401218
rect -8726 400898 -2934 401134
rect -2698 400898 -2614 401134
rect -2378 400898 23250 401134
rect 23486 400898 29514 401134
rect 29750 400898 51250 401134
rect 51486 400898 57514 401134
rect 57750 400898 79250 401134
rect 79486 400898 85514 401134
rect 85750 400898 107250 401134
rect 107486 400898 113514 401134
rect 113750 400898 135250 401134
rect 135486 400898 141514 401134
rect 141750 400898 163250 401134
rect 163486 400898 169514 401134
rect 169750 400898 191250 401134
rect 191486 400898 197514 401134
rect 197750 400898 219250 401134
rect 219486 400898 225514 401134
rect 225750 400898 247250 401134
rect 247486 400898 253514 401134
rect 253750 400898 275250 401134
rect 275486 400898 281514 401134
rect 281750 400898 303250 401134
rect 303486 400898 309514 401134
rect 309750 400898 331250 401134
rect 331486 400898 337514 401134
rect 337750 400898 359250 401134
rect 359486 400898 365514 401134
rect 365750 400898 387250 401134
rect 387486 400898 393514 401134
rect 393750 400898 415250 401134
rect 415486 400898 421514 401134
rect 421750 400898 443250 401134
rect 443486 400898 449514 401134
rect 449750 400898 471250 401134
rect 471486 400898 477514 401134
rect 477750 400898 499250 401134
rect 499486 400898 505514 401134
rect 505750 400898 527250 401134
rect 527486 400898 533514 401134
rect 533750 400898 555250 401134
rect 555486 400898 561514 401134
rect 561750 400898 586302 401134
rect 586538 400898 586622 401134
rect 586858 400898 592650 401134
rect -8726 400866 592650 400898
rect -8726 377829 592650 377861
rect -8726 377593 -1974 377829
rect -1738 377593 -1654 377829
rect -1418 377593 20118 377829
rect 20354 377593 26382 377829
rect 26618 377593 32646 377829
rect 32882 377593 48118 377829
rect 48354 377593 54382 377829
rect 54618 377593 60646 377829
rect 60882 377593 76118 377829
rect 76354 377593 82382 377829
rect 82618 377593 88646 377829
rect 88882 377593 104118 377829
rect 104354 377593 110382 377829
rect 110618 377593 116646 377829
rect 116882 377593 132118 377829
rect 132354 377593 138382 377829
rect 138618 377593 144646 377829
rect 144882 377593 160118 377829
rect 160354 377593 166382 377829
rect 166618 377593 172646 377829
rect 172882 377593 188118 377829
rect 188354 377593 194382 377829
rect 194618 377593 200646 377829
rect 200882 377593 216118 377829
rect 216354 377593 222382 377829
rect 222618 377593 228646 377829
rect 228882 377593 244118 377829
rect 244354 377593 250382 377829
rect 250618 377593 256646 377829
rect 256882 377593 272118 377829
rect 272354 377593 278382 377829
rect 278618 377593 284646 377829
rect 284882 377593 300118 377829
rect 300354 377593 306382 377829
rect 306618 377593 312646 377829
rect 312882 377593 328118 377829
rect 328354 377593 334382 377829
rect 334618 377593 340646 377829
rect 340882 377593 356118 377829
rect 356354 377593 362382 377829
rect 362618 377593 368646 377829
rect 368882 377593 384118 377829
rect 384354 377593 390382 377829
rect 390618 377593 396646 377829
rect 396882 377593 412118 377829
rect 412354 377593 418382 377829
rect 418618 377593 424646 377829
rect 424882 377593 440118 377829
rect 440354 377593 446382 377829
rect 446618 377593 452646 377829
rect 452882 377593 468118 377829
rect 468354 377593 474382 377829
rect 474618 377593 480646 377829
rect 480882 377593 496118 377829
rect 496354 377593 502382 377829
rect 502618 377593 508646 377829
rect 508882 377593 524118 377829
rect 524354 377593 530382 377829
rect 530618 377593 536646 377829
rect 536882 377593 552118 377829
rect 552354 377593 558382 377829
rect 558618 377593 564646 377829
rect 564882 377593 573526 377829
rect 573762 377593 573846 377829
rect 574082 377593 585342 377829
rect 585578 377593 585662 377829
rect 585898 377593 592650 377829
rect -8726 377509 592650 377593
rect -8726 377273 -1974 377509
rect -1738 377273 -1654 377509
rect -1418 377273 20118 377509
rect 20354 377273 26382 377509
rect 26618 377273 32646 377509
rect 32882 377273 48118 377509
rect 48354 377273 54382 377509
rect 54618 377273 60646 377509
rect 60882 377273 76118 377509
rect 76354 377273 82382 377509
rect 82618 377273 88646 377509
rect 88882 377273 104118 377509
rect 104354 377273 110382 377509
rect 110618 377273 116646 377509
rect 116882 377273 132118 377509
rect 132354 377273 138382 377509
rect 138618 377273 144646 377509
rect 144882 377273 160118 377509
rect 160354 377273 166382 377509
rect 166618 377273 172646 377509
rect 172882 377273 188118 377509
rect 188354 377273 194382 377509
rect 194618 377273 200646 377509
rect 200882 377273 216118 377509
rect 216354 377273 222382 377509
rect 222618 377273 228646 377509
rect 228882 377273 244118 377509
rect 244354 377273 250382 377509
rect 250618 377273 256646 377509
rect 256882 377273 272118 377509
rect 272354 377273 278382 377509
rect 278618 377273 284646 377509
rect 284882 377273 300118 377509
rect 300354 377273 306382 377509
rect 306618 377273 312646 377509
rect 312882 377273 328118 377509
rect 328354 377273 334382 377509
rect 334618 377273 340646 377509
rect 340882 377273 356118 377509
rect 356354 377273 362382 377509
rect 362618 377273 368646 377509
rect 368882 377273 384118 377509
rect 384354 377273 390382 377509
rect 390618 377273 396646 377509
rect 396882 377273 412118 377509
rect 412354 377273 418382 377509
rect 418618 377273 424646 377509
rect 424882 377273 440118 377509
rect 440354 377273 446382 377509
rect 446618 377273 452646 377509
rect 452882 377273 468118 377509
rect 468354 377273 474382 377509
rect 474618 377273 480646 377509
rect 480882 377273 496118 377509
rect 496354 377273 502382 377509
rect 502618 377273 508646 377509
rect 508882 377273 524118 377509
rect 524354 377273 530382 377509
rect 530618 377273 536646 377509
rect 536882 377273 552118 377509
rect 552354 377273 558382 377509
rect 558618 377273 564646 377509
rect 564882 377273 573526 377509
rect 573762 377273 573846 377509
rect 574082 377273 585342 377509
rect 585578 377273 585662 377509
rect 585898 377273 592650 377509
rect -8726 377241 592650 377273
rect -8726 374454 592650 374486
rect -8726 374218 -2934 374454
rect -2698 374218 -2614 374454
rect -2378 374218 23250 374454
rect 23486 374218 29514 374454
rect 29750 374218 51250 374454
rect 51486 374218 57514 374454
rect 57750 374218 79250 374454
rect 79486 374218 85514 374454
rect 85750 374218 107250 374454
rect 107486 374218 113514 374454
rect 113750 374218 135250 374454
rect 135486 374218 141514 374454
rect 141750 374218 163250 374454
rect 163486 374218 169514 374454
rect 169750 374218 191250 374454
rect 191486 374218 197514 374454
rect 197750 374218 219250 374454
rect 219486 374218 225514 374454
rect 225750 374218 247250 374454
rect 247486 374218 253514 374454
rect 253750 374218 275250 374454
rect 275486 374218 281514 374454
rect 281750 374218 303250 374454
rect 303486 374218 309514 374454
rect 309750 374218 331250 374454
rect 331486 374218 337514 374454
rect 337750 374218 359250 374454
rect 359486 374218 365514 374454
rect 365750 374218 387250 374454
rect 387486 374218 393514 374454
rect 393750 374218 415250 374454
rect 415486 374218 421514 374454
rect 421750 374218 443250 374454
rect 443486 374218 449514 374454
rect 449750 374218 471250 374454
rect 471486 374218 477514 374454
rect 477750 374218 499250 374454
rect 499486 374218 505514 374454
rect 505750 374218 527250 374454
rect 527486 374218 533514 374454
rect 533750 374218 555250 374454
rect 555486 374218 561514 374454
rect 561750 374218 586302 374454
rect 586538 374218 586622 374454
rect 586858 374218 592650 374454
rect -8726 374134 592650 374218
rect -8726 373898 -2934 374134
rect -2698 373898 -2614 374134
rect -2378 373898 23250 374134
rect 23486 373898 29514 374134
rect 29750 373898 51250 374134
rect 51486 373898 57514 374134
rect 57750 373898 79250 374134
rect 79486 373898 85514 374134
rect 85750 373898 107250 374134
rect 107486 373898 113514 374134
rect 113750 373898 135250 374134
rect 135486 373898 141514 374134
rect 141750 373898 163250 374134
rect 163486 373898 169514 374134
rect 169750 373898 191250 374134
rect 191486 373898 197514 374134
rect 197750 373898 219250 374134
rect 219486 373898 225514 374134
rect 225750 373898 247250 374134
rect 247486 373898 253514 374134
rect 253750 373898 275250 374134
rect 275486 373898 281514 374134
rect 281750 373898 303250 374134
rect 303486 373898 309514 374134
rect 309750 373898 331250 374134
rect 331486 373898 337514 374134
rect 337750 373898 359250 374134
rect 359486 373898 365514 374134
rect 365750 373898 387250 374134
rect 387486 373898 393514 374134
rect 393750 373898 415250 374134
rect 415486 373898 421514 374134
rect 421750 373898 443250 374134
rect 443486 373898 449514 374134
rect 449750 373898 471250 374134
rect 471486 373898 477514 374134
rect 477750 373898 499250 374134
rect 499486 373898 505514 374134
rect 505750 373898 527250 374134
rect 527486 373898 533514 374134
rect 533750 373898 555250 374134
rect 555486 373898 561514 374134
rect 561750 373898 586302 374134
rect 586538 373898 586622 374134
rect 586858 373898 592650 374134
rect -8726 373866 592650 373898
rect -8726 350829 592650 350861
rect -8726 350593 -1974 350829
rect -1738 350593 -1654 350829
rect -1418 350593 20118 350829
rect 20354 350593 26382 350829
rect 26618 350593 32646 350829
rect 32882 350593 48118 350829
rect 48354 350593 54382 350829
rect 54618 350593 60646 350829
rect 60882 350593 76118 350829
rect 76354 350593 82382 350829
rect 82618 350593 88646 350829
rect 88882 350593 104118 350829
rect 104354 350593 110382 350829
rect 110618 350593 116646 350829
rect 116882 350593 132118 350829
rect 132354 350593 138382 350829
rect 138618 350593 144646 350829
rect 144882 350593 160118 350829
rect 160354 350593 166382 350829
rect 166618 350593 172646 350829
rect 172882 350593 188118 350829
rect 188354 350593 194382 350829
rect 194618 350593 200646 350829
rect 200882 350593 216118 350829
rect 216354 350593 222382 350829
rect 222618 350593 228646 350829
rect 228882 350593 244118 350829
rect 244354 350593 250382 350829
rect 250618 350593 256646 350829
rect 256882 350593 272118 350829
rect 272354 350593 278382 350829
rect 278618 350593 284646 350829
rect 284882 350593 300118 350829
rect 300354 350593 306382 350829
rect 306618 350593 312646 350829
rect 312882 350593 328118 350829
rect 328354 350593 334382 350829
rect 334618 350593 340646 350829
rect 340882 350593 356118 350829
rect 356354 350593 362382 350829
rect 362618 350593 368646 350829
rect 368882 350593 384118 350829
rect 384354 350593 390382 350829
rect 390618 350593 396646 350829
rect 396882 350593 412118 350829
rect 412354 350593 418382 350829
rect 418618 350593 424646 350829
rect 424882 350593 440118 350829
rect 440354 350593 446382 350829
rect 446618 350593 452646 350829
rect 452882 350593 468118 350829
rect 468354 350593 474382 350829
rect 474618 350593 480646 350829
rect 480882 350593 496118 350829
rect 496354 350593 502382 350829
rect 502618 350593 508646 350829
rect 508882 350593 524118 350829
rect 524354 350593 530382 350829
rect 530618 350593 536646 350829
rect 536882 350593 552118 350829
rect 552354 350593 558382 350829
rect 558618 350593 564646 350829
rect 564882 350593 573526 350829
rect 573762 350593 573846 350829
rect 574082 350593 585342 350829
rect 585578 350593 585662 350829
rect 585898 350593 592650 350829
rect -8726 350509 592650 350593
rect -8726 350273 -1974 350509
rect -1738 350273 -1654 350509
rect -1418 350273 20118 350509
rect 20354 350273 26382 350509
rect 26618 350273 32646 350509
rect 32882 350273 48118 350509
rect 48354 350273 54382 350509
rect 54618 350273 60646 350509
rect 60882 350273 76118 350509
rect 76354 350273 82382 350509
rect 82618 350273 88646 350509
rect 88882 350273 104118 350509
rect 104354 350273 110382 350509
rect 110618 350273 116646 350509
rect 116882 350273 132118 350509
rect 132354 350273 138382 350509
rect 138618 350273 144646 350509
rect 144882 350273 160118 350509
rect 160354 350273 166382 350509
rect 166618 350273 172646 350509
rect 172882 350273 188118 350509
rect 188354 350273 194382 350509
rect 194618 350273 200646 350509
rect 200882 350273 216118 350509
rect 216354 350273 222382 350509
rect 222618 350273 228646 350509
rect 228882 350273 244118 350509
rect 244354 350273 250382 350509
rect 250618 350273 256646 350509
rect 256882 350273 272118 350509
rect 272354 350273 278382 350509
rect 278618 350273 284646 350509
rect 284882 350273 300118 350509
rect 300354 350273 306382 350509
rect 306618 350273 312646 350509
rect 312882 350273 328118 350509
rect 328354 350273 334382 350509
rect 334618 350273 340646 350509
rect 340882 350273 356118 350509
rect 356354 350273 362382 350509
rect 362618 350273 368646 350509
rect 368882 350273 384118 350509
rect 384354 350273 390382 350509
rect 390618 350273 396646 350509
rect 396882 350273 412118 350509
rect 412354 350273 418382 350509
rect 418618 350273 424646 350509
rect 424882 350273 440118 350509
rect 440354 350273 446382 350509
rect 446618 350273 452646 350509
rect 452882 350273 468118 350509
rect 468354 350273 474382 350509
rect 474618 350273 480646 350509
rect 480882 350273 496118 350509
rect 496354 350273 502382 350509
rect 502618 350273 508646 350509
rect 508882 350273 524118 350509
rect 524354 350273 530382 350509
rect 530618 350273 536646 350509
rect 536882 350273 552118 350509
rect 552354 350273 558382 350509
rect 558618 350273 564646 350509
rect 564882 350273 573526 350509
rect 573762 350273 573846 350509
rect 574082 350273 585342 350509
rect 585578 350273 585662 350509
rect 585898 350273 592650 350509
rect -8726 350241 592650 350273
rect -8726 347454 592650 347486
rect -8726 347218 -2934 347454
rect -2698 347218 -2614 347454
rect -2378 347218 23250 347454
rect 23486 347218 29514 347454
rect 29750 347218 51250 347454
rect 51486 347218 57514 347454
rect 57750 347218 79250 347454
rect 79486 347218 85514 347454
rect 85750 347218 107250 347454
rect 107486 347218 113514 347454
rect 113750 347218 135250 347454
rect 135486 347218 141514 347454
rect 141750 347218 163250 347454
rect 163486 347218 169514 347454
rect 169750 347218 191250 347454
rect 191486 347218 197514 347454
rect 197750 347218 219250 347454
rect 219486 347218 225514 347454
rect 225750 347218 247250 347454
rect 247486 347218 253514 347454
rect 253750 347218 275250 347454
rect 275486 347218 281514 347454
rect 281750 347218 303250 347454
rect 303486 347218 309514 347454
rect 309750 347218 331250 347454
rect 331486 347218 337514 347454
rect 337750 347218 359250 347454
rect 359486 347218 365514 347454
rect 365750 347218 387250 347454
rect 387486 347218 393514 347454
rect 393750 347218 415250 347454
rect 415486 347218 421514 347454
rect 421750 347218 443250 347454
rect 443486 347218 449514 347454
rect 449750 347218 471250 347454
rect 471486 347218 477514 347454
rect 477750 347218 499250 347454
rect 499486 347218 505514 347454
rect 505750 347218 527250 347454
rect 527486 347218 533514 347454
rect 533750 347218 555250 347454
rect 555486 347218 561514 347454
rect 561750 347218 586302 347454
rect 586538 347218 586622 347454
rect 586858 347218 592650 347454
rect -8726 347134 592650 347218
rect -8726 346898 -2934 347134
rect -2698 346898 -2614 347134
rect -2378 346898 23250 347134
rect 23486 346898 29514 347134
rect 29750 346898 51250 347134
rect 51486 346898 57514 347134
rect 57750 346898 79250 347134
rect 79486 346898 85514 347134
rect 85750 346898 107250 347134
rect 107486 346898 113514 347134
rect 113750 346898 135250 347134
rect 135486 346898 141514 347134
rect 141750 346898 163250 347134
rect 163486 346898 169514 347134
rect 169750 346898 191250 347134
rect 191486 346898 197514 347134
rect 197750 346898 219250 347134
rect 219486 346898 225514 347134
rect 225750 346898 247250 347134
rect 247486 346898 253514 347134
rect 253750 346898 275250 347134
rect 275486 346898 281514 347134
rect 281750 346898 303250 347134
rect 303486 346898 309514 347134
rect 309750 346898 331250 347134
rect 331486 346898 337514 347134
rect 337750 346898 359250 347134
rect 359486 346898 365514 347134
rect 365750 346898 387250 347134
rect 387486 346898 393514 347134
rect 393750 346898 415250 347134
rect 415486 346898 421514 347134
rect 421750 346898 443250 347134
rect 443486 346898 449514 347134
rect 449750 346898 471250 347134
rect 471486 346898 477514 347134
rect 477750 346898 499250 347134
rect 499486 346898 505514 347134
rect 505750 346898 527250 347134
rect 527486 346898 533514 347134
rect 533750 346898 555250 347134
rect 555486 346898 561514 347134
rect 561750 346898 586302 347134
rect 586538 346898 586622 347134
rect 586858 346898 592650 347134
rect -8726 346866 592650 346898
rect -8726 323829 592650 323861
rect -8726 323593 -1974 323829
rect -1738 323593 -1654 323829
rect -1418 323593 20118 323829
rect 20354 323593 26382 323829
rect 26618 323593 32646 323829
rect 32882 323593 48118 323829
rect 48354 323593 54382 323829
rect 54618 323593 60646 323829
rect 60882 323593 76118 323829
rect 76354 323593 82382 323829
rect 82618 323593 88646 323829
rect 88882 323593 104118 323829
rect 104354 323593 110382 323829
rect 110618 323593 116646 323829
rect 116882 323593 132118 323829
rect 132354 323593 138382 323829
rect 138618 323593 144646 323829
rect 144882 323593 160118 323829
rect 160354 323593 166382 323829
rect 166618 323593 172646 323829
rect 172882 323593 188118 323829
rect 188354 323593 194382 323829
rect 194618 323593 200646 323829
rect 200882 323593 216118 323829
rect 216354 323593 222382 323829
rect 222618 323593 228646 323829
rect 228882 323593 244118 323829
rect 244354 323593 250382 323829
rect 250618 323593 256646 323829
rect 256882 323593 272118 323829
rect 272354 323593 278382 323829
rect 278618 323593 284646 323829
rect 284882 323593 300118 323829
rect 300354 323593 306382 323829
rect 306618 323593 312646 323829
rect 312882 323593 328118 323829
rect 328354 323593 334382 323829
rect 334618 323593 340646 323829
rect 340882 323593 356118 323829
rect 356354 323593 362382 323829
rect 362618 323593 368646 323829
rect 368882 323593 384118 323829
rect 384354 323593 390382 323829
rect 390618 323593 396646 323829
rect 396882 323593 412118 323829
rect 412354 323593 418382 323829
rect 418618 323593 424646 323829
rect 424882 323593 440118 323829
rect 440354 323593 446382 323829
rect 446618 323593 452646 323829
rect 452882 323593 468118 323829
rect 468354 323593 474382 323829
rect 474618 323593 480646 323829
rect 480882 323593 496118 323829
rect 496354 323593 502382 323829
rect 502618 323593 508646 323829
rect 508882 323593 524118 323829
rect 524354 323593 530382 323829
rect 530618 323593 536646 323829
rect 536882 323593 552118 323829
rect 552354 323593 558382 323829
rect 558618 323593 564646 323829
rect 564882 323593 573526 323829
rect 573762 323593 573846 323829
rect 574082 323593 585342 323829
rect 585578 323593 585662 323829
rect 585898 323593 592650 323829
rect -8726 323509 592650 323593
rect -8726 323273 -1974 323509
rect -1738 323273 -1654 323509
rect -1418 323273 20118 323509
rect 20354 323273 26382 323509
rect 26618 323273 32646 323509
rect 32882 323273 48118 323509
rect 48354 323273 54382 323509
rect 54618 323273 60646 323509
rect 60882 323273 76118 323509
rect 76354 323273 82382 323509
rect 82618 323273 88646 323509
rect 88882 323273 104118 323509
rect 104354 323273 110382 323509
rect 110618 323273 116646 323509
rect 116882 323273 132118 323509
rect 132354 323273 138382 323509
rect 138618 323273 144646 323509
rect 144882 323273 160118 323509
rect 160354 323273 166382 323509
rect 166618 323273 172646 323509
rect 172882 323273 188118 323509
rect 188354 323273 194382 323509
rect 194618 323273 200646 323509
rect 200882 323273 216118 323509
rect 216354 323273 222382 323509
rect 222618 323273 228646 323509
rect 228882 323273 244118 323509
rect 244354 323273 250382 323509
rect 250618 323273 256646 323509
rect 256882 323273 272118 323509
rect 272354 323273 278382 323509
rect 278618 323273 284646 323509
rect 284882 323273 300118 323509
rect 300354 323273 306382 323509
rect 306618 323273 312646 323509
rect 312882 323273 328118 323509
rect 328354 323273 334382 323509
rect 334618 323273 340646 323509
rect 340882 323273 356118 323509
rect 356354 323273 362382 323509
rect 362618 323273 368646 323509
rect 368882 323273 384118 323509
rect 384354 323273 390382 323509
rect 390618 323273 396646 323509
rect 396882 323273 412118 323509
rect 412354 323273 418382 323509
rect 418618 323273 424646 323509
rect 424882 323273 440118 323509
rect 440354 323273 446382 323509
rect 446618 323273 452646 323509
rect 452882 323273 468118 323509
rect 468354 323273 474382 323509
rect 474618 323273 480646 323509
rect 480882 323273 496118 323509
rect 496354 323273 502382 323509
rect 502618 323273 508646 323509
rect 508882 323273 524118 323509
rect 524354 323273 530382 323509
rect 530618 323273 536646 323509
rect 536882 323273 552118 323509
rect 552354 323273 558382 323509
rect 558618 323273 564646 323509
rect 564882 323273 573526 323509
rect 573762 323273 573846 323509
rect 574082 323273 585342 323509
rect 585578 323273 585662 323509
rect 585898 323273 592650 323509
rect -8726 323241 592650 323273
rect -8726 320454 592650 320486
rect -8726 320218 -2934 320454
rect -2698 320218 -2614 320454
rect -2378 320218 23250 320454
rect 23486 320218 29514 320454
rect 29750 320218 51250 320454
rect 51486 320218 57514 320454
rect 57750 320218 79250 320454
rect 79486 320218 85514 320454
rect 85750 320218 107250 320454
rect 107486 320218 113514 320454
rect 113750 320218 135250 320454
rect 135486 320218 141514 320454
rect 141750 320218 163250 320454
rect 163486 320218 169514 320454
rect 169750 320218 191250 320454
rect 191486 320218 197514 320454
rect 197750 320218 219250 320454
rect 219486 320218 225514 320454
rect 225750 320218 247250 320454
rect 247486 320218 253514 320454
rect 253750 320218 275250 320454
rect 275486 320218 281514 320454
rect 281750 320218 303250 320454
rect 303486 320218 309514 320454
rect 309750 320218 331250 320454
rect 331486 320218 337514 320454
rect 337750 320218 359250 320454
rect 359486 320218 365514 320454
rect 365750 320218 387250 320454
rect 387486 320218 393514 320454
rect 393750 320218 415250 320454
rect 415486 320218 421514 320454
rect 421750 320218 443250 320454
rect 443486 320218 449514 320454
rect 449750 320218 471250 320454
rect 471486 320218 477514 320454
rect 477750 320218 499250 320454
rect 499486 320218 505514 320454
rect 505750 320218 527250 320454
rect 527486 320218 533514 320454
rect 533750 320218 555250 320454
rect 555486 320218 561514 320454
rect 561750 320218 586302 320454
rect 586538 320218 586622 320454
rect 586858 320218 592650 320454
rect -8726 320134 592650 320218
rect -8726 319898 -2934 320134
rect -2698 319898 -2614 320134
rect -2378 319898 23250 320134
rect 23486 319898 29514 320134
rect 29750 319898 51250 320134
rect 51486 319898 57514 320134
rect 57750 319898 79250 320134
rect 79486 319898 85514 320134
rect 85750 319898 107250 320134
rect 107486 319898 113514 320134
rect 113750 319898 135250 320134
rect 135486 319898 141514 320134
rect 141750 319898 163250 320134
rect 163486 319898 169514 320134
rect 169750 319898 191250 320134
rect 191486 319898 197514 320134
rect 197750 319898 219250 320134
rect 219486 319898 225514 320134
rect 225750 319898 247250 320134
rect 247486 319898 253514 320134
rect 253750 319898 275250 320134
rect 275486 319898 281514 320134
rect 281750 319898 303250 320134
rect 303486 319898 309514 320134
rect 309750 319898 331250 320134
rect 331486 319898 337514 320134
rect 337750 319898 359250 320134
rect 359486 319898 365514 320134
rect 365750 319898 387250 320134
rect 387486 319898 393514 320134
rect 393750 319898 415250 320134
rect 415486 319898 421514 320134
rect 421750 319898 443250 320134
rect 443486 319898 449514 320134
rect 449750 319898 471250 320134
rect 471486 319898 477514 320134
rect 477750 319898 499250 320134
rect 499486 319898 505514 320134
rect 505750 319898 527250 320134
rect 527486 319898 533514 320134
rect 533750 319898 555250 320134
rect 555486 319898 561514 320134
rect 561750 319898 586302 320134
rect 586538 319898 586622 320134
rect 586858 319898 592650 320134
rect -8726 319866 592650 319898
rect -8726 296829 592650 296861
rect -8726 296593 -1974 296829
rect -1738 296593 -1654 296829
rect -1418 296593 20118 296829
rect 20354 296593 26382 296829
rect 26618 296593 32646 296829
rect 32882 296593 48118 296829
rect 48354 296593 54382 296829
rect 54618 296593 60646 296829
rect 60882 296593 76118 296829
rect 76354 296593 82382 296829
rect 82618 296593 88646 296829
rect 88882 296593 104118 296829
rect 104354 296593 110382 296829
rect 110618 296593 116646 296829
rect 116882 296593 132118 296829
rect 132354 296593 138382 296829
rect 138618 296593 144646 296829
rect 144882 296593 160118 296829
rect 160354 296593 166382 296829
rect 166618 296593 172646 296829
rect 172882 296593 188118 296829
rect 188354 296593 194382 296829
rect 194618 296593 200646 296829
rect 200882 296593 216118 296829
rect 216354 296593 222382 296829
rect 222618 296593 228646 296829
rect 228882 296593 244118 296829
rect 244354 296593 250382 296829
rect 250618 296593 256646 296829
rect 256882 296593 272118 296829
rect 272354 296593 278382 296829
rect 278618 296593 284646 296829
rect 284882 296593 300118 296829
rect 300354 296593 306382 296829
rect 306618 296593 312646 296829
rect 312882 296593 328118 296829
rect 328354 296593 334382 296829
rect 334618 296593 340646 296829
rect 340882 296593 356118 296829
rect 356354 296593 362382 296829
rect 362618 296593 368646 296829
rect 368882 296593 384118 296829
rect 384354 296593 390382 296829
rect 390618 296593 396646 296829
rect 396882 296593 412118 296829
rect 412354 296593 418382 296829
rect 418618 296593 424646 296829
rect 424882 296593 440118 296829
rect 440354 296593 446382 296829
rect 446618 296593 452646 296829
rect 452882 296593 468118 296829
rect 468354 296593 474382 296829
rect 474618 296593 480646 296829
rect 480882 296593 496118 296829
rect 496354 296593 502382 296829
rect 502618 296593 508646 296829
rect 508882 296593 524118 296829
rect 524354 296593 530382 296829
rect 530618 296593 536646 296829
rect 536882 296593 552118 296829
rect 552354 296593 558382 296829
rect 558618 296593 564646 296829
rect 564882 296593 573526 296829
rect 573762 296593 573846 296829
rect 574082 296593 585342 296829
rect 585578 296593 585662 296829
rect 585898 296593 592650 296829
rect -8726 296509 592650 296593
rect -8726 296273 -1974 296509
rect -1738 296273 -1654 296509
rect -1418 296273 20118 296509
rect 20354 296273 26382 296509
rect 26618 296273 32646 296509
rect 32882 296273 48118 296509
rect 48354 296273 54382 296509
rect 54618 296273 60646 296509
rect 60882 296273 76118 296509
rect 76354 296273 82382 296509
rect 82618 296273 88646 296509
rect 88882 296273 104118 296509
rect 104354 296273 110382 296509
rect 110618 296273 116646 296509
rect 116882 296273 132118 296509
rect 132354 296273 138382 296509
rect 138618 296273 144646 296509
rect 144882 296273 160118 296509
rect 160354 296273 166382 296509
rect 166618 296273 172646 296509
rect 172882 296273 188118 296509
rect 188354 296273 194382 296509
rect 194618 296273 200646 296509
rect 200882 296273 216118 296509
rect 216354 296273 222382 296509
rect 222618 296273 228646 296509
rect 228882 296273 244118 296509
rect 244354 296273 250382 296509
rect 250618 296273 256646 296509
rect 256882 296273 272118 296509
rect 272354 296273 278382 296509
rect 278618 296273 284646 296509
rect 284882 296273 300118 296509
rect 300354 296273 306382 296509
rect 306618 296273 312646 296509
rect 312882 296273 328118 296509
rect 328354 296273 334382 296509
rect 334618 296273 340646 296509
rect 340882 296273 356118 296509
rect 356354 296273 362382 296509
rect 362618 296273 368646 296509
rect 368882 296273 384118 296509
rect 384354 296273 390382 296509
rect 390618 296273 396646 296509
rect 396882 296273 412118 296509
rect 412354 296273 418382 296509
rect 418618 296273 424646 296509
rect 424882 296273 440118 296509
rect 440354 296273 446382 296509
rect 446618 296273 452646 296509
rect 452882 296273 468118 296509
rect 468354 296273 474382 296509
rect 474618 296273 480646 296509
rect 480882 296273 496118 296509
rect 496354 296273 502382 296509
rect 502618 296273 508646 296509
rect 508882 296273 524118 296509
rect 524354 296273 530382 296509
rect 530618 296273 536646 296509
rect 536882 296273 552118 296509
rect 552354 296273 558382 296509
rect 558618 296273 564646 296509
rect 564882 296273 573526 296509
rect 573762 296273 573846 296509
rect 574082 296273 585342 296509
rect 585578 296273 585662 296509
rect 585898 296273 592650 296509
rect -8726 296241 592650 296273
rect -8726 293454 592650 293486
rect -8726 293218 -2934 293454
rect -2698 293218 -2614 293454
rect -2378 293218 23250 293454
rect 23486 293218 29514 293454
rect 29750 293218 51250 293454
rect 51486 293218 57514 293454
rect 57750 293218 79250 293454
rect 79486 293218 85514 293454
rect 85750 293218 107250 293454
rect 107486 293218 113514 293454
rect 113750 293218 135250 293454
rect 135486 293218 141514 293454
rect 141750 293218 163250 293454
rect 163486 293218 169514 293454
rect 169750 293218 191250 293454
rect 191486 293218 197514 293454
rect 197750 293218 219250 293454
rect 219486 293218 225514 293454
rect 225750 293218 247250 293454
rect 247486 293218 253514 293454
rect 253750 293218 275250 293454
rect 275486 293218 281514 293454
rect 281750 293218 303250 293454
rect 303486 293218 309514 293454
rect 309750 293218 331250 293454
rect 331486 293218 337514 293454
rect 337750 293218 359250 293454
rect 359486 293218 365514 293454
rect 365750 293218 387250 293454
rect 387486 293218 393514 293454
rect 393750 293218 415250 293454
rect 415486 293218 421514 293454
rect 421750 293218 443250 293454
rect 443486 293218 449514 293454
rect 449750 293218 471250 293454
rect 471486 293218 477514 293454
rect 477750 293218 499250 293454
rect 499486 293218 505514 293454
rect 505750 293218 527250 293454
rect 527486 293218 533514 293454
rect 533750 293218 555250 293454
rect 555486 293218 561514 293454
rect 561750 293218 586302 293454
rect 586538 293218 586622 293454
rect 586858 293218 592650 293454
rect -8726 293134 592650 293218
rect -8726 292898 -2934 293134
rect -2698 292898 -2614 293134
rect -2378 292898 23250 293134
rect 23486 292898 29514 293134
rect 29750 292898 51250 293134
rect 51486 292898 57514 293134
rect 57750 292898 79250 293134
rect 79486 292898 85514 293134
rect 85750 292898 107250 293134
rect 107486 292898 113514 293134
rect 113750 292898 135250 293134
rect 135486 292898 141514 293134
rect 141750 292898 163250 293134
rect 163486 292898 169514 293134
rect 169750 292898 191250 293134
rect 191486 292898 197514 293134
rect 197750 292898 219250 293134
rect 219486 292898 225514 293134
rect 225750 292898 247250 293134
rect 247486 292898 253514 293134
rect 253750 292898 275250 293134
rect 275486 292898 281514 293134
rect 281750 292898 303250 293134
rect 303486 292898 309514 293134
rect 309750 292898 331250 293134
rect 331486 292898 337514 293134
rect 337750 292898 359250 293134
rect 359486 292898 365514 293134
rect 365750 292898 387250 293134
rect 387486 292898 393514 293134
rect 393750 292898 415250 293134
rect 415486 292898 421514 293134
rect 421750 292898 443250 293134
rect 443486 292898 449514 293134
rect 449750 292898 471250 293134
rect 471486 292898 477514 293134
rect 477750 292898 499250 293134
rect 499486 292898 505514 293134
rect 505750 292898 527250 293134
rect 527486 292898 533514 293134
rect 533750 292898 555250 293134
rect 555486 292898 561514 293134
rect 561750 292898 586302 293134
rect 586538 292898 586622 293134
rect 586858 292898 592650 293134
rect -8726 292866 592650 292898
rect -8726 269829 592650 269861
rect -8726 269593 -1974 269829
rect -1738 269593 -1654 269829
rect -1418 269593 20118 269829
rect 20354 269593 26382 269829
rect 26618 269593 32646 269829
rect 32882 269593 48118 269829
rect 48354 269593 54382 269829
rect 54618 269593 60646 269829
rect 60882 269593 76118 269829
rect 76354 269593 82382 269829
rect 82618 269593 88646 269829
rect 88882 269593 104118 269829
rect 104354 269593 110382 269829
rect 110618 269593 116646 269829
rect 116882 269593 132118 269829
rect 132354 269593 138382 269829
rect 138618 269593 144646 269829
rect 144882 269593 160118 269829
rect 160354 269593 166382 269829
rect 166618 269593 172646 269829
rect 172882 269593 188118 269829
rect 188354 269593 194382 269829
rect 194618 269593 200646 269829
rect 200882 269593 216118 269829
rect 216354 269593 222382 269829
rect 222618 269593 228646 269829
rect 228882 269593 244118 269829
rect 244354 269593 250382 269829
rect 250618 269593 256646 269829
rect 256882 269593 272118 269829
rect 272354 269593 278382 269829
rect 278618 269593 284646 269829
rect 284882 269593 300118 269829
rect 300354 269593 306382 269829
rect 306618 269593 312646 269829
rect 312882 269593 328118 269829
rect 328354 269593 334382 269829
rect 334618 269593 340646 269829
rect 340882 269593 356118 269829
rect 356354 269593 362382 269829
rect 362618 269593 368646 269829
rect 368882 269593 384118 269829
rect 384354 269593 390382 269829
rect 390618 269593 396646 269829
rect 396882 269593 412118 269829
rect 412354 269593 418382 269829
rect 418618 269593 424646 269829
rect 424882 269593 440118 269829
rect 440354 269593 446382 269829
rect 446618 269593 452646 269829
rect 452882 269593 468118 269829
rect 468354 269593 474382 269829
rect 474618 269593 480646 269829
rect 480882 269593 496118 269829
rect 496354 269593 502382 269829
rect 502618 269593 508646 269829
rect 508882 269593 524118 269829
rect 524354 269593 530382 269829
rect 530618 269593 536646 269829
rect 536882 269593 552118 269829
rect 552354 269593 558382 269829
rect 558618 269593 564646 269829
rect 564882 269593 573526 269829
rect 573762 269593 573846 269829
rect 574082 269593 585342 269829
rect 585578 269593 585662 269829
rect 585898 269593 592650 269829
rect -8726 269509 592650 269593
rect -8726 269273 -1974 269509
rect -1738 269273 -1654 269509
rect -1418 269273 20118 269509
rect 20354 269273 26382 269509
rect 26618 269273 32646 269509
rect 32882 269273 48118 269509
rect 48354 269273 54382 269509
rect 54618 269273 60646 269509
rect 60882 269273 76118 269509
rect 76354 269273 82382 269509
rect 82618 269273 88646 269509
rect 88882 269273 104118 269509
rect 104354 269273 110382 269509
rect 110618 269273 116646 269509
rect 116882 269273 132118 269509
rect 132354 269273 138382 269509
rect 138618 269273 144646 269509
rect 144882 269273 160118 269509
rect 160354 269273 166382 269509
rect 166618 269273 172646 269509
rect 172882 269273 188118 269509
rect 188354 269273 194382 269509
rect 194618 269273 200646 269509
rect 200882 269273 216118 269509
rect 216354 269273 222382 269509
rect 222618 269273 228646 269509
rect 228882 269273 244118 269509
rect 244354 269273 250382 269509
rect 250618 269273 256646 269509
rect 256882 269273 272118 269509
rect 272354 269273 278382 269509
rect 278618 269273 284646 269509
rect 284882 269273 300118 269509
rect 300354 269273 306382 269509
rect 306618 269273 312646 269509
rect 312882 269273 328118 269509
rect 328354 269273 334382 269509
rect 334618 269273 340646 269509
rect 340882 269273 356118 269509
rect 356354 269273 362382 269509
rect 362618 269273 368646 269509
rect 368882 269273 384118 269509
rect 384354 269273 390382 269509
rect 390618 269273 396646 269509
rect 396882 269273 412118 269509
rect 412354 269273 418382 269509
rect 418618 269273 424646 269509
rect 424882 269273 440118 269509
rect 440354 269273 446382 269509
rect 446618 269273 452646 269509
rect 452882 269273 468118 269509
rect 468354 269273 474382 269509
rect 474618 269273 480646 269509
rect 480882 269273 496118 269509
rect 496354 269273 502382 269509
rect 502618 269273 508646 269509
rect 508882 269273 524118 269509
rect 524354 269273 530382 269509
rect 530618 269273 536646 269509
rect 536882 269273 552118 269509
rect 552354 269273 558382 269509
rect 558618 269273 564646 269509
rect 564882 269273 573526 269509
rect 573762 269273 573846 269509
rect 574082 269273 585342 269509
rect 585578 269273 585662 269509
rect 585898 269273 592650 269509
rect -8726 269241 592650 269273
rect -8726 266454 592650 266486
rect -8726 266218 -2934 266454
rect -2698 266218 -2614 266454
rect -2378 266218 23250 266454
rect 23486 266218 29514 266454
rect 29750 266218 51250 266454
rect 51486 266218 57514 266454
rect 57750 266218 79250 266454
rect 79486 266218 85514 266454
rect 85750 266218 107250 266454
rect 107486 266218 113514 266454
rect 113750 266218 135250 266454
rect 135486 266218 141514 266454
rect 141750 266218 163250 266454
rect 163486 266218 169514 266454
rect 169750 266218 191250 266454
rect 191486 266218 197514 266454
rect 197750 266218 219250 266454
rect 219486 266218 225514 266454
rect 225750 266218 247250 266454
rect 247486 266218 253514 266454
rect 253750 266218 275250 266454
rect 275486 266218 281514 266454
rect 281750 266218 303250 266454
rect 303486 266218 309514 266454
rect 309750 266218 331250 266454
rect 331486 266218 337514 266454
rect 337750 266218 359250 266454
rect 359486 266218 365514 266454
rect 365750 266218 387250 266454
rect 387486 266218 393514 266454
rect 393750 266218 415250 266454
rect 415486 266218 421514 266454
rect 421750 266218 443250 266454
rect 443486 266218 449514 266454
rect 449750 266218 471250 266454
rect 471486 266218 477514 266454
rect 477750 266218 499250 266454
rect 499486 266218 505514 266454
rect 505750 266218 527250 266454
rect 527486 266218 533514 266454
rect 533750 266218 555250 266454
rect 555486 266218 561514 266454
rect 561750 266218 586302 266454
rect 586538 266218 586622 266454
rect 586858 266218 592650 266454
rect -8726 266134 592650 266218
rect -8726 265898 -2934 266134
rect -2698 265898 -2614 266134
rect -2378 265898 23250 266134
rect 23486 265898 29514 266134
rect 29750 265898 51250 266134
rect 51486 265898 57514 266134
rect 57750 265898 79250 266134
rect 79486 265898 85514 266134
rect 85750 265898 107250 266134
rect 107486 265898 113514 266134
rect 113750 265898 135250 266134
rect 135486 265898 141514 266134
rect 141750 265898 163250 266134
rect 163486 265898 169514 266134
rect 169750 265898 191250 266134
rect 191486 265898 197514 266134
rect 197750 265898 219250 266134
rect 219486 265898 225514 266134
rect 225750 265898 247250 266134
rect 247486 265898 253514 266134
rect 253750 265898 275250 266134
rect 275486 265898 281514 266134
rect 281750 265898 303250 266134
rect 303486 265898 309514 266134
rect 309750 265898 331250 266134
rect 331486 265898 337514 266134
rect 337750 265898 359250 266134
rect 359486 265898 365514 266134
rect 365750 265898 387250 266134
rect 387486 265898 393514 266134
rect 393750 265898 415250 266134
rect 415486 265898 421514 266134
rect 421750 265898 443250 266134
rect 443486 265898 449514 266134
rect 449750 265898 471250 266134
rect 471486 265898 477514 266134
rect 477750 265898 499250 266134
rect 499486 265898 505514 266134
rect 505750 265898 527250 266134
rect 527486 265898 533514 266134
rect 533750 265898 555250 266134
rect 555486 265898 561514 266134
rect 561750 265898 586302 266134
rect 586538 265898 586622 266134
rect 586858 265898 592650 266134
rect -8726 265866 592650 265898
rect -8726 242829 592650 242861
rect -8726 242593 -1974 242829
rect -1738 242593 -1654 242829
rect -1418 242593 20118 242829
rect 20354 242593 26382 242829
rect 26618 242593 32646 242829
rect 32882 242593 48118 242829
rect 48354 242593 54382 242829
rect 54618 242593 60646 242829
rect 60882 242593 76118 242829
rect 76354 242593 82382 242829
rect 82618 242593 88646 242829
rect 88882 242593 104118 242829
rect 104354 242593 110382 242829
rect 110618 242593 116646 242829
rect 116882 242593 132118 242829
rect 132354 242593 138382 242829
rect 138618 242593 144646 242829
rect 144882 242593 160118 242829
rect 160354 242593 166382 242829
rect 166618 242593 172646 242829
rect 172882 242593 188118 242829
rect 188354 242593 194382 242829
rect 194618 242593 200646 242829
rect 200882 242593 216118 242829
rect 216354 242593 222382 242829
rect 222618 242593 228646 242829
rect 228882 242593 244118 242829
rect 244354 242593 250382 242829
rect 250618 242593 256646 242829
rect 256882 242593 272118 242829
rect 272354 242593 278382 242829
rect 278618 242593 284646 242829
rect 284882 242593 300118 242829
rect 300354 242593 306382 242829
rect 306618 242593 312646 242829
rect 312882 242593 328118 242829
rect 328354 242593 334382 242829
rect 334618 242593 340646 242829
rect 340882 242593 356118 242829
rect 356354 242593 362382 242829
rect 362618 242593 368646 242829
rect 368882 242593 384118 242829
rect 384354 242593 390382 242829
rect 390618 242593 396646 242829
rect 396882 242593 412118 242829
rect 412354 242593 418382 242829
rect 418618 242593 424646 242829
rect 424882 242593 440118 242829
rect 440354 242593 446382 242829
rect 446618 242593 452646 242829
rect 452882 242593 468118 242829
rect 468354 242593 474382 242829
rect 474618 242593 480646 242829
rect 480882 242593 496118 242829
rect 496354 242593 502382 242829
rect 502618 242593 508646 242829
rect 508882 242593 524118 242829
rect 524354 242593 530382 242829
rect 530618 242593 536646 242829
rect 536882 242593 552118 242829
rect 552354 242593 558382 242829
rect 558618 242593 564646 242829
rect 564882 242593 573526 242829
rect 573762 242593 573846 242829
rect 574082 242593 585342 242829
rect 585578 242593 585662 242829
rect 585898 242593 592650 242829
rect -8726 242509 592650 242593
rect -8726 242273 -1974 242509
rect -1738 242273 -1654 242509
rect -1418 242273 20118 242509
rect 20354 242273 26382 242509
rect 26618 242273 32646 242509
rect 32882 242273 48118 242509
rect 48354 242273 54382 242509
rect 54618 242273 60646 242509
rect 60882 242273 76118 242509
rect 76354 242273 82382 242509
rect 82618 242273 88646 242509
rect 88882 242273 104118 242509
rect 104354 242273 110382 242509
rect 110618 242273 116646 242509
rect 116882 242273 132118 242509
rect 132354 242273 138382 242509
rect 138618 242273 144646 242509
rect 144882 242273 160118 242509
rect 160354 242273 166382 242509
rect 166618 242273 172646 242509
rect 172882 242273 188118 242509
rect 188354 242273 194382 242509
rect 194618 242273 200646 242509
rect 200882 242273 216118 242509
rect 216354 242273 222382 242509
rect 222618 242273 228646 242509
rect 228882 242273 244118 242509
rect 244354 242273 250382 242509
rect 250618 242273 256646 242509
rect 256882 242273 272118 242509
rect 272354 242273 278382 242509
rect 278618 242273 284646 242509
rect 284882 242273 300118 242509
rect 300354 242273 306382 242509
rect 306618 242273 312646 242509
rect 312882 242273 328118 242509
rect 328354 242273 334382 242509
rect 334618 242273 340646 242509
rect 340882 242273 356118 242509
rect 356354 242273 362382 242509
rect 362618 242273 368646 242509
rect 368882 242273 384118 242509
rect 384354 242273 390382 242509
rect 390618 242273 396646 242509
rect 396882 242273 412118 242509
rect 412354 242273 418382 242509
rect 418618 242273 424646 242509
rect 424882 242273 440118 242509
rect 440354 242273 446382 242509
rect 446618 242273 452646 242509
rect 452882 242273 468118 242509
rect 468354 242273 474382 242509
rect 474618 242273 480646 242509
rect 480882 242273 496118 242509
rect 496354 242273 502382 242509
rect 502618 242273 508646 242509
rect 508882 242273 524118 242509
rect 524354 242273 530382 242509
rect 530618 242273 536646 242509
rect 536882 242273 552118 242509
rect 552354 242273 558382 242509
rect 558618 242273 564646 242509
rect 564882 242273 573526 242509
rect 573762 242273 573846 242509
rect 574082 242273 585342 242509
rect 585578 242273 585662 242509
rect 585898 242273 592650 242509
rect -8726 242241 592650 242273
rect -8726 239454 592650 239486
rect -8726 239218 -2934 239454
rect -2698 239218 -2614 239454
rect -2378 239218 23250 239454
rect 23486 239218 29514 239454
rect 29750 239218 51250 239454
rect 51486 239218 57514 239454
rect 57750 239218 79250 239454
rect 79486 239218 85514 239454
rect 85750 239218 107250 239454
rect 107486 239218 113514 239454
rect 113750 239218 135250 239454
rect 135486 239218 141514 239454
rect 141750 239218 163250 239454
rect 163486 239218 169514 239454
rect 169750 239218 191250 239454
rect 191486 239218 197514 239454
rect 197750 239218 219250 239454
rect 219486 239218 225514 239454
rect 225750 239218 247250 239454
rect 247486 239218 253514 239454
rect 253750 239218 275250 239454
rect 275486 239218 281514 239454
rect 281750 239218 303250 239454
rect 303486 239218 309514 239454
rect 309750 239218 331250 239454
rect 331486 239218 337514 239454
rect 337750 239218 359250 239454
rect 359486 239218 365514 239454
rect 365750 239218 387250 239454
rect 387486 239218 393514 239454
rect 393750 239218 415250 239454
rect 415486 239218 421514 239454
rect 421750 239218 443250 239454
rect 443486 239218 449514 239454
rect 449750 239218 471250 239454
rect 471486 239218 477514 239454
rect 477750 239218 499250 239454
rect 499486 239218 505514 239454
rect 505750 239218 527250 239454
rect 527486 239218 533514 239454
rect 533750 239218 555250 239454
rect 555486 239218 561514 239454
rect 561750 239218 586302 239454
rect 586538 239218 586622 239454
rect 586858 239218 592650 239454
rect -8726 239134 592650 239218
rect -8726 238898 -2934 239134
rect -2698 238898 -2614 239134
rect -2378 238898 23250 239134
rect 23486 238898 29514 239134
rect 29750 238898 51250 239134
rect 51486 238898 57514 239134
rect 57750 238898 79250 239134
rect 79486 238898 85514 239134
rect 85750 238898 107250 239134
rect 107486 238898 113514 239134
rect 113750 238898 135250 239134
rect 135486 238898 141514 239134
rect 141750 238898 163250 239134
rect 163486 238898 169514 239134
rect 169750 238898 191250 239134
rect 191486 238898 197514 239134
rect 197750 238898 219250 239134
rect 219486 238898 225514 239134
rect 225750 238898 247250 239134
rect 247486 238898 253514 239134
rect 253750 238898 275250 239134
rect 275486 238898 281514 239134
rect 281750 238898 303250 239134
rect 303486 238898 309514 239134
rect 309750 238898 331250 239134
rect 331486 238898 337514 239134
rect 337750 238898 359250 239134
rect 359486 238898 365514 239134
rect 365750 238898 387250 239134
rect 387486 238898 393514 239134
rect 393750 238898 415250 239134
rect 415486 238898 421514 239134
rect 421750 238898 443250 239134
rect 443486 238898 449514 239134
rect 449750 238898 471250 239134
rect 471486 238898 477514 239134
rect 477750 238898 499250 239134
rect 499486 238898 505514 239134
rect 505750 238898 527250 239134
rect 527486 238898 533514 239134
rect 533750 238898 555250 239134
rect 555486 238898 561514 239134
rect 561750 238898 586302 239134
rect 586538 238898 586622 239134
rect 586858 238898 592650 239134
rect -8726 238866 592650 238898
rect -8726 215829 592650 215861
rect -8726 215593 -1974 215829
rect -1738 215593 -1654 215829
rect -1418 215593 20118 215829
rect 20354 215593 26382 215829
rect 26618 215593 32646 215829
rect 32882 215593 48118 215829
rect 48354 215593 54382 215829
rect 54618 215593 60646 215829
rect 60882 215593 76118 215829
rect 76354 215593 82382 215829
rect 82618 215593 88646 215829
rect 88882 215593 104118 215829
rect 104354 215593 110382 215829
rect 110618 215593 116646 215829
rect 116882 215593 132118 215829
rect 132354 215593 138382 215829
rect 138618 215593 144646 215829
rect 144882 215593 160118 215829
rect 160354 215593 166382 215829
rect 166618 215593 172646 215829
rect 172882 215593 187335 215829
rect 187571 215593 192033 215829
rect 192269 215593 196731 215829
rect 196967 215593 201429 215829
rect 201665 215593 215335 215829
rect 215571 215593 220033 215829
rect 220269 215593 224731 215829
rect 224967 215593 229429 215829
rect 229665 215593 243335 215829
rect 243571 215593 248033 215829
rect 248269 215593 252731 215829
rect 252967 215593 257429 215829
rect 257665 215593 271335 215829
rect 271571 215593 276033 215829
rect 276269 215593 280731 215829
rect 280967 215593 285429 215829
rect 285665 215593 299335 215829
rect 299571 215593 304033 215829
rect 304269 215593 308731 215829
rect 308967 215593 313429 215829
rect 313665 215593 328118 215829
rect 328354 215593 334382 215829
rect 334618 215593 340646 215829
rect 340882 215593 355335 215829
rect 355571 215593 360033 215829
rect 360269 215593 364731 215829
rect 364967 215593 369429 215829
rect 369665 215593 383335 215829
rect 383571 215593 388033 215829
rect 388269 215593 392731 215829
rect 392967 215593 397429 215829
rect 397665 215593 411335 215829
rect 411571 215593 416033 215829
rect 416269 215593 420731 215829
rect 420967 215593 425429 215829
rect 425665 215593 439335 215829
rect 439571 215593 444033 215829
rect 444269 215593 448731 215829
rect 448967 215593 453429 215829
rect 453665 215593 467335 215829
rect 467571 215593 472033 215829
rect 472269 215593 476731 215829
rect 476967 215593 481429 215829
rect 481665 215593 495335 215829
rect 495571 215593 500033 215829
rect 500269 215593 504731 215829
rect 504967 215593 509429 215829
rect 509665 215593 523335 215829
rect 523571 215593 528033 215829
rect 528269 215593 532731 215829
rect 532967 215593 537429 215829
rect 537665 215593 551335 215829
rect 551571 215593 556033 215829
rect 556269 215593 560731 215829
rect 560967 215593 565429 215829
rect 565665 215593 573526 215829
rect 573762 215593 573846 215829
rect 574082 215593 585342 215829
rect 585578 215593 585662 215829
rect 585898 215593 592650 215829
rect -8726 215509 592650 215593
rect -8726 215273 -1974 215509
rect -1738 215273 -1654 215509
rect -1418 215273 20118 215509
rect 20354 215273 26382 215509
rect 26618 215273 32646 215509
rect 32882 215273 48118 215509
rect 48354 215273 54382 215509
rect 54618 215273 60646 215509
rect 60882 215273 76118 215509
rect 76354 215273 82382 215509
rect 82618 215273 88646 215509
rect 88882 215273 104118 215509
rect 104354 215273 110382 215509
rect 110618 215273 116646 215509
rect 116882 215273 132118 215509
rect 132354 215273 138382 215509
rect 138618 215273 144646 215509
rect 144882 215273 160118 215509
rect 160354 215273 166382 215509
rect 166618 215273 172646 215509
rect 172882 215273 187335 215509
rect 187571 215273 192033 215509
rect 192269 215273 196731 215509
rect 196967 215273 201429 215509
rect 201665 215273 215335 215509
rect 215571 215273 220033 215509
rect 220269 215273 224731 215509
rect 224967 215273 229429 215509
rect 229665 215273 243335 215509
rect 243571 215273 248033 215509
rect 248269 215273 252731 215509
rect 252967 215273 257429 215509
rect 257665 215273 271335 215509
rect 271571 215273 276033 215509
rect 276269 215273 280731 215509
rect 280967 215273 285429 215509
rect 285665 215273 299335 215509
rect 299571 215273 304033 215509
rect 304269 215273 308731 215509
rect 308967 215273 313429 215509
rect 313665 215273 328118 215509
rect 328354 215273 334382 215509
rect 334618 215273 340646 215509
rect 340882 215273 355335 215509
rect 355571 215273 360033 215509
rect 360269 215273 364731 215509
rect 364967 215273 369429 215509
rect 369665 215273 383335 215509
rect 383571 215273 388033 215509
rect 388269 215273 392731 215509
rect 392967 215273 397429 215509
rect 397665 215273 411335 215509
rect 411571 215273 416033 215509
rect 416269 215273 420731 215509
rect 420967 215273 425429 215509
rect 425665 215273 439335 215509
rect 439571 215273 444033 215509
rect 444269 215273 448731 215509
rect 448967 215273 453429 215509
rect 453665 215273 467335 215509
rect 467571 215273 472033 215509
rect 472269 215273 476731 215509
rect 476967 215273 481429 215509
rect 481665 215273 495335 215509
rect 495571 215273 500033 215509
rect 500269 215273 504731 215509
rect 504967 215273 509429 215509
rect 509665 215273 523335 215509
rect 523571 215273 528033 215509
rect 528269 215273 532731 215509
rect 532967 215273 537429 215509
rect 537665 215273 551335 215509
rect 551571 215273 556033 215509
rect 556269 215273 560731 215509
rect 560967 215273 565429 215509
rect 565665 215273 573526 215509
rect 573762 215273 573846 215509
rect 574082 215273 585342 215509
rect 585578 215273 585662 215509
rect 585898 215273 592650 215509
rect -8726 215241 592650 215273
rect -8726 212454 592650 212486
rect -8726 212218 -2934 212454
rect -2698 212218 -2614 212454
rect -2378 212218 23250 212454
rect 23486 212218 29514 212454
rect 29750 212218 51250 212454
rect 51486 212218 57514 212454
rect 57750 212218 79250 212454
rect 79486 212218 85514 212454
rect 85750 212218 107250 212454
rect 107486 212218 113514 212454
rect 113750 212218 135250 212454
rect 135486 212218 141514 212454
rect 141750 212218 163250 212454
rect 163486 212218 169514 212454
rect 169750 212218 189684 212454
rect 189920 212218 194382 212454
rect 194618 212218 199080 212454
rect 199316 212218 217684 212454
rect 217920 212218 222382 212454
rect 222618 212218 227080 212454
rect 227316 212218 245684 212454
rect 245920 212218 250382 212454
rect 250618 212218 255080 212454
rect 255316 212218 273684 212454
rect 273920 212218 278382 212454
rect 278618 212218 283080 212454
rect 283316 212218 301684 212454
rect 301920 212218 306382 212454
rect 306618 212218 311080 212454
rect 311316 212218 331250 212454
rect 331486 212218 337514 212454
rect 337750 212218 357684 212454
rect 357920 212218 362382 212454
rect 362618 212218 367080 212454
rect 367316 212218 385684 212454
rect 385920 212218 390382 212454
rect 390618 212218 395080 212454
rect 395316 212218 413684 212454
rect 413920 212218 418382 212454
rect 418618 212218 423080 212454
rect 423316 212218 441684 212454
rect 441920 212218 446382 212454
rect 446618 212218 451080 212454
rect 451316 212218 469684 212454
rect 469920 212218 474382 212454
rect 474618 212218 479080 212454
rect 479316 212218 497684 212454
rect 497920 212218 502382 212454
rect 502618 212218 507080 212454
rect 507316 212218 525684 212454
rect 525920 212218 530382 212454
rect 530618 212218 535080 212454
rect 535316 212218 553684 212454
rect 553920 212218 558382 212454
rect 558618 212218 563080 212454
rect 563316 212218 586302 212454
rect 586538 212218 586622 212454
rect 586858 212218 592650 212454
rect -8726 212134 592650 212218
rect -8726 211898 -2934 212134
rect -2698 211898 -2614 212134
rect -2378 211898 23250 212134
rect 23486 211898 29514 212134
rect 29750 211898 51250 212134
rect 51486 211898 57514 212134
rect 57750 211898 79250 212134
rect 79486 211898 85514 212134
rect 85750 211898 107250 212134
rect 107486 211898 113514 212134
rect 113750 211898 135250 212134
rect 135486 211898 141514 212134
rect 141750 211898 163250 212134
rect 163486 211898 169514 212134
rect 169750 211898 189684 212134
rect 189920 211898 194382 212134
rect 194618 211898 199080 212134
rect 199316 211898 217684 212134
rect 217920 211898 222382 212134
rect 222618 211898 227080 212134
rect 227316 211898 245684 212134
rect 245920 211898 250382 212134
rect 250618 211898 255080 212134
rect 255316 211898 273684 212134
rect 273920 211898 278382 212134
rect 278618 211898 283080 212134
rect 283316 211898 301684 212134
rect 301920 211898 306382 212134
rect 306618 211898 311080 212134
rect 311316 211898 331250 212134
rect 331486 211898 337514 212134
rect 337750 211898 357684 212134
rect 357920 211898 362382 212134
rect 362618 211898 367080 212134
rect 367316 211898 385684 212134
rect 385920 211898 390382 212134
rect 390618 211898 395080 212134
rect 395316 211898 413684 212134
rect 413920 211898 418382 212134
rect 418618 211898 423080 212134
rect 423316 211898 441684 212134
rect 441920 211898 446382 212134
rect 446618 211898 451080 212134
rect 451316 211898 469684 212134
rect 469920 211898 474382 212134
rect 474618 211898 479080 212134
rect 479316 211898 497684 212134
rect 497920 211898 502382 212134
rect 502618 211898 507080 212134
rect 507316 211898 525684 212134
rect 525920 211898 530382 212134
rect 530618 211898 535080 212134
rect 535316 211898 553684 212134
rect 553920 211898 558382 212134
rect 558618 211898 563080 212134
rect 563316 211898 586302 212134
rect 586538 211898 586622 212134
rect 586858 211898 592650 212134
rect -8726 211866 592650 211898
rect -8726 188829 592650 188861
rect -8726 188593 -1974 188829
rect -1738 188593 -1654 188829
rect -1418 188593 19335 188829
rect 19571 188593 24033 188829
rect 24269 188593 28731 188829
rect 28967 188593 33429 188829
rect 33665 188593 47335 188829
rect 47571 188593 52033 188829
rect 52269 188593 56731 188829
rect 56967 188593 61429 188829
rect 61665 188593 75335 188829
rect 75571 188593 80033 188829
rect 80269 188593 84731 188829
rect 84967 188593 89429 188829
rect 89665 188593 103335 188829
rect 103571 188593 108033 188829
rect 108269 188593 112731 188829
rect 112967 188593 117429 188829
rect 117665 188593 131335 188829
rect 131571 188593 136033 188829
rect 136269 188593 140731 188829
rect 140967 188593 145429 188829
rect 145665 188593 159335 188829
rect 159571 188593 164033 188829
rect 164269 188593 168731 188829
rect 168967 188593 173429 188829
rect 173665 188593 187335 188829
rect 187571 188593 192033 188829
rect 192269 188593 196731 188829
rect 196967 188593 201429 188829
rect 201665 188593 215335 188829
rect 215571 188593 220033 188829
rect 220269 188593 224731 188829
rect 224967 188593 229429 188829
rect 229665 188593 243335 188829
rect 243571 188593 248033 188829
rect 248269 188593 252731 188829
rect 252967 188593 257429 188829
rect 257665 188593 271335 188829
rect 271571 188593 276033 188829
rect 276269 188593 280731 188829
rect 280967 188593 285429 188829
rect 285665 188593 299335 188829
rect 299571 188593 304033 188829
rect 304269 188593 308731 188829
rect 308967 188593 313429 188829
rect 313665 188593 327335 188829
rect 327571 188593 332033 188829
rect 332269 188593 336731 188829
rect 336967 188593 341429 188829
rect 341665 188593 355335 188829
rect 355571 188593 360033 188829
rect 360269 188593 364731 188829
rect 364967 188593 369429 188829
rect 369665 188593 383335 188829
rect 383571 188593 388033 188829
rect 388269 188593 392731 188829
rect 392967 188593 397429 188829
rect 397665 188593 411335 188829
rect 411571 188593 416033 188829
rect 416269 188593 420731 188829
rect 420967 188593 425429 188829
rect 425665 188593 439335 188829
rect 439571 188593 444033 188829
rect 444269 188593 448731 188829
rect 448967 188593 453429 188829
rect 453665 188593 467335 188829
rect 467571 188593 472033 188829
rect 472269 188593 476731 188829
rect 476967 188593 481429 188829
rect 481665 188593 495335 188829
rect 495571 188593 500033 188829
rect 500269 188593 504731 188829
rect 504967 188593 509429 188829
rect 509665 188593 523335 188829
rect 523571 188593 528033 188829
rect 528269 188593 532731 188829
rect 532967 188593 537429 188829
rect 537665 188593 551335 188829
rect 551571 188593 556033 188829
rect 556269 188593 560731 188829
rect 560967 188593 565429 188829
rect 565665 188593 573526 188829
rect 573762 188593 573846 188829
rect 574082 188593 585342 188829
rect 585578 188593 585662 188829
rect 585898 188593 592650 188829
rect -8726 188509 592650 188593
rect -8726 188273 -1974 188509
rect -1738 188273 -1654 188509
rect -1418 188273 19335 188509
rect 19571 188273 24033 188509
rect 24269 188273 28731 188509
rect 28967 188273 33429 188509
rect 33665 188273 47335 188509
rect 47571 188273 52033 188509
rect 52269 188273 56731 188509
rect 56967 188273 61429 188509
rect 61665 188273 75335 188509
rect 75571 188273 80033 188509
rect 80269 188273 84731 188509
rect 84967 188273 89429 188509
rect 89665 188273 103335 188509
rect 103571 188273 108033 188509
rect 108269 188273 112731 188509
rect 112967 188273 117429 188509
rect 117665 188273 131335 188509
rect 131571 188273 136033 188509
rect 136269 188273 140731 188509
rect 140967 188273 145429 188509
rect 145665 188273 159335 188509
rect 159571 188273 164033 188509
rect 164269 188273 168731 188509
rect 168967 188273 173429 188509
rect 173665 188273 187335 188509
rect 187571 188273 192033 188509
rect 192269 188273 196731 188509
rect 196967 188273 201429 188509
rect 201665 188273 215335 188509
rect 215571 188273 220033 188509
rect 220269 188273 224731 188509
rect 224967 188273 229429 188509
rect 229665 188273 243335 188509
rect 243571 188273 248033 188509
rect 248269 188273 252731 188509
rect 252967 188273 257429 188509
rect 257665 188273 271335 188509
rect 271571 188273 276033 188509
rect 276269 188273 280731 188509
rect 280967 188273 285429 188509
rect 285665 188273 299335 188509
rect 299571 188273 304033 188509
rect 304269 188273 308731 188509
rect 308967 188273 313429 188509
rect 313665 188273 327335 188509
rect 327571 188273 332033 188509
rect 332269 188273 336731 188509
rect 336967 188273 341429 188509
rect 341665 188273 355335 188509
rect 355571 188273 360033 188509
rect 360269 188273 364731 188509
rect 364967 188273 369429 188509
rect 369665 188273 383335 188509
rect 383571 188273 388033 188509
rect 388269 188273 392731 188509
rect 392967 188273 397429 188509
rect 397665 188273 411335 188509
rect 411571 188273 416033 188509
rect 416269 188273 420731 188509
rect 420967 188273 425429 188509
rect 425665 188273 439335 188509
rect 439571 188273 444033 188509
rect 444269 188273 448731 188509
rect 448967 188273 453429 188509
rect 453665 188273 467335 188509
rect 467571 188273 472033 188509
rect 472269 188273 476731 188509
rect 476967 188273 481429 188509
rect 481665 188273 495335 188509
rect 495571 188273 500033 188509
rect 500269 188273 504731 188509
rect 504967 188273 509429 188509
rect 509665 188273 523335 188509
rect 523571 188273 528033 188509
rect 528269 188273 532731 188509
rect 532967 188273 537429 188509
rect 537665 188273 551335 188509
rect 551571 188273 556033 188509
rect 556269 188273 560731 188509
rect 560967 188273 565429 188509
rect 565665 188273 573526 188509
rect 573762 188273 573846 188509
rect 574082 188273 585342 188509
rect 585578 188273 585662 188509
rect 585898 188273 592650 188509
rect -8726 188241 592650 188273
rect -8726 185454 592650 185486
rect -8726 185218 -2934 185454
rect -2698 185218 -2614 185454
rect -2378 185218 21684 185454
rect 21920 185218 26382 185454
rect 26618 185218 31080 185454
rect 31316 185218 49684 185454
rect 49920 185218 54382 185454
rect 54618 185218 59080 185454
rect 59316 185218 77684 185454
rect 77920 185218 82382 185454
rect 82618 185218 87080 185454
rect 87316 185218 105684 185454
rect 105920 185218 110382 185454
rect 110618 185218 115080 185454
rect 115316 185218 133684 185454
rect 133920 185218 138382 185454
rect 138618 185218 143080 185454
rect 143316 185218 161684 185454
rect 161920 185218 166382 185454
rect 166618 185218 171080 185454
rect 171316 185218 189684 185454
rect 189920 185218 194382 185454
rect 194618 185218 199080 185454
rect 199316 185218 217684 185454
rect 217920 185218 222382 185454
rect 222618 185218 227080 185454
rect 227316 185218 245684 185454
rect 245920 185218 250382 185454
rect 250618 185218 255080 185454
rect 255316 185218 273684 185454
rect 273920 185218 278382 185454
rect 278618 185218 283080 185454
rect 283316 185218 301684 185454
rect 301920 185218 306382 185454
rect 306618 185218 311080 185454
rect 311316 185218 329684 185454
rect 329920 185218 334382 185454
rect 334618 185218 339080 185454
rect 339316 185218 357684 185454
rect 357920 185218 362382 185454
rect 362618 185218 367080 185454
rect 367316 185218 385684 185454
rect 385920 185218 390382 185454
rect 390618 185218 395080 185454
rect 395316 185218 413684 185454
rect 413920 185218 418382 185454
rect 418618 185218 423080 185454
rect 423316 185218 441684 185454
rect 441920 185218 446382 185454
rect 446618 185218 451080 185454
rect 451316 185218 469684 185454
rect 469920 185218 474382 185454
rect 474618 185218 479080 185454
rect 479316 185218 497684 185454
rect 497920 185218 502382 185454
rect 502618 185218 507080 185454
rect 507316 185218 525684 185454
rect 525920 185218 530382 185454
rect 530618 185218 535080 185454
rect 535316 185218 553684 185454
rect 553920 185218 558382 185454
rect 558618 185218 563080 185454
rect 563316 185218 586302 185454
rect 586538 185218 586622 185454
rect 586858 185218 592650 185454
rect -8726 185134 592650 185218
rect -8726 184898 -2934 185134
rect -2698 184898 -2614 185134
rect -2378 184898 21684 185134
rect 21920 184898 26382 185134
rect 26618 184898 31080 185134
rect 31316 184898 49684 185134
rect 49920 184898 54382 185134
rect 54618 184898 59080 185134
rect 59316 184898 77684 185134
rect 77920 184898 82382 185134
rect 82618 184898 87080 185134
rect 87316 184898 105684 185134
rect 105920 184898 110382 185134
rect 110618 184898 115080 185134
rect 115316 184898 133684 185134
rect 133920 184898 138382 185134
rect 138618 184898 143080 185134
rect 143316 184898 161684 185134
rect 161920 184898 166382 185134
rect 166618 184898 171080 185134
rect 171316 184898 189684 185134
rect 189920 184898 194382 185134
rect 194618 184898 199080 185134
rect 199316 184898 217684 185134
rect 217920 184898 222382 185134
rect 222618 184898 227080 185134
rect 227316 184898 245684 185134
rect 245920 184898 250382 185134
rect 250618 184898 255080 185134
rect 255316 184898 273684 185134
rect 273920 184898 278382 185134
rect 278618 184898 283080 185134
rect 283316 184898 301684 185134
rect 301920 184898 306382 185134
rect 306618 184898 311080 185134
rect 311316 184898 329684 185134
rect 329920 184898 334382 185134
rect 334618 184898 339080 185134
rect 339316 184898 357684 185134
rect 357920 184898 362382 185134
rect 362618 184898 367080 185134
rect 367316 184898 385684 185134
rect 385920 184898 390382 185134
rect 390618 184898 395080 185134
rect 395316 184898 413684 185134
rect 413920 184898 418382 185134
rect 418618 184898 423080 185134
rect 423316 184898 441684 185134
rect 441920 184898 446382 185134
rect 446618 184898 451080 185134
rect 451316 184898 469684 185134
rect 469920 184898 474382 185134
rect 474618 184898 479080 185134
rect 479316 184898 497684 185134
rect 497920 184898 502382 185134
rect 502618 184898 507080 185134
rect 507316 184898 525684 185134
rect 525920 184898 530382 185134
rect 530618 184898 535080 185134
rect 535316 184898 553684 185134
rect 553920 184898 558382 185134
rect 558618 184898 563080 185134
rect 563316 184898 586302 185134
rect 586538 184898 586622 185134
rect 586858 184898 592650 185134
rect -8726 184866 592650 184898
rect -8726 161829 592650 161861
rect -8726 161593 -1974 161829
rect -1738 161593 -1654 161829
rect -1418 161593 19335 161829
rect 19571 161593 24033 161829
rect 24269 161593 28731 161829
rect 28967 161593 33429 161829
rect 33665 161593 47335 161829
rect 47571 161593 52033 161829
rect 52269 161593 56731 161829
rect 56967 161593 61429 161829
rect 61665 161593 75335 161829
rect 75571 161593 80033 161829
rect 80269 161593 84731 161829
rect 84967 161593 89429 161829
rect 89665 161593 103335 161829
rect 103571 161593 108033 161829
rect 108269 161593 112731 161829
rect 112967 161593 117429 161829
rect 117665 161593 131335 161829
rect 131571 161593 136033 161829
rect 136269 161593 140731 161829
rect 140967 161593 145429 161829
rect 145665 161593 159335 161829
rect 159571 161593 164033 161829
rect 164269 161593 168731 161829
rect 168967 161593 173429 161829
rect 173665 161593 187335 161829
rect 187571 161593 192033 161829
rect 192269 161593 196731 161829
rect 196967 161593 201429 161829
rect 201665 161593 215335 161829
rect 215571 161593 220033 161829
rect 220269 161593 224731 161829
rect 224967 161593 229429 161829
rect 229665 161593 243335 161829
rect 243571 161593 248033 161829
rect 248269 161593 252731 161829
rect 252967 161593 257429 161829
rect 257665 161593 271335 161829
rect 271571 161593 276033 161829
rect 276269 161593 280731 161829
rect 280967 161593 285429 161829
rect 285665 161593 299335 161829
rect 299571 161593 304033 161829
rect 304269 161593 308731 161829
rect 308967 161593 313429 161829
rect 313665 161593 327335 161829
rect 327571 161593 332033 161829
rect 332269 161593 336731 161829
rect 336967 161593 341429 161829
rect 341665 161593 355335 161829
rect 355571 161593 360033 161829
rect 360269 161593 364731 161829
rect 364967 161593 369429 161829
rect 369665 161593 383335 161829
rect 383571 161593 388033 161829
rect 388269 161593 392731 161829
rect 392967 161593 397429 161829
rect 397665 161593 411335 161829
rect 411571 161593 416033 161829
rect 416269 161593 420731 161829
rect 420967 161593 425429 161829
rect 425665 161593 439335 161829
rect 439571 161593 444033 161829
rect 444269 161593 448731 161829
rect 448967 161593 453429 161829
rect 453665 161593 467335 161829
rect 467571 161593 472033 161829
rect 472269 161593 476731 161829
rect 476967 161593 481429 161829
rect 481665 161593 495335 161829
rect 495571 161593 500033 161829
rect 500269 161593 504731 161829
rect 504967 161593 509429 161829
rect 509665 161593 523335 161829
rect 523571 161593 528033 161829
rect 528269 161593 532731 161829
rect 532967 161593 537429 161829
rect 537665 161593 551335 161829
rect 551571 161593 556033 161829
rect 556269 161593 560731 161829
rect 560967 161593 565429 161829
rect 565665 161593 573526 161829
rect 573762 161593 573846 161829
rect 574082 161593 585342 161829
rect 585578 161593 585662 161829
rect 585898 161593 592650 161829
rect -8726 161509 592650 161593
rect -8726 161273 -1974 161509
rect -1738 161273 -1654 161509
rect -1418 161273 19335 161509
rect 19571 161273 24033 161509
rect 24269 161273 28731 161509
rect 28967 161273 33429 161509
rect 33665 161273 47335 161509
rect 47571 161273 52033 161509
rect 52269 161273 56731 161509
rect 56967 161273 61429 161509
rect 61665 161273 75335 161509
rect 75571 161273 80033 161509
rect 80269 161273 84731 161509
rect 84967 161273 89429 161509
rect 89665 161273 103335 161509
rect 103571 161273 108033 161509
rect 108269 161273 112731 161509
rect 112967 161273 117429 161509
rect 117665 161273 131335 161509
rect 131571 161273 136033 161509
rect 136269 161273 140731 161509
rect 140967 161273 145429 161509
rect 145665 161273 159335 161509
rect 159571 161273 164033 161509
rect 164269 161273 168731 161509
rect 168967 161273 173429 161509
rect 173665 161273 187335 161509
rect 187571 161273 192033 161509
rect 192269 161273 196731 161509
rect 196967 161273 201429 161509
rect 201665 161273 215335 161509
rect 215571 161273 220033 161509
rect 220269 161273 224731 161509
rect 224967 161273 229429 161509
rect 229665 161273 243335 161509
rect 243571 161273 248033 161509
rect 248269 161273 252731 161509
rect 252967 161273 257429 161509
rect 257665 161273 271335 161509
rect 271571 161273 276033 161509
rect 276269 161273 280731 161509
rect 280967 161273 285429 161509
rect 285665 161273 299335 161509
rect 299571 161273 304033 161509
rect 304269 161273 308731 161509
rect 308967 161273 313429 161509
rect 313665 161273 327335 161509
rect 327571 161273 332033 161509
rect 332269 161273 336731 161509
rect 336967 161273 341429 161509
rect 341665 161273 355335 161509
rect 355571 161273 360033 161509
rect 360269 161273 364731 161509
rect 364967 161273 369429 161509
rect 369665 161273 383335 161509
rect 383571 161273 388033 161509
rect 388269 161273 392731 161509
rect 392967 161273 397429 161509
rect 397665 161273 411335 161509
rect 411571 161273 416033 161509
rect 416269 161273 420731 161509
rect 420967 161273 425429 161509
rect 425665 161273 439335 161509
rect 439571 161273 444033 161509
rect 444269 161273 448731 161509
rect 448967 161273 453429 161509
rect 453665 161273 467335 161509
rect 467571 161273 472033 161509
rect 472269 161273 476731 161509
rect 476967 161273 481429 161509
rect 481665 161273 495335 161509
rect 495571 161273 500033 161509
rect 500269 161273 504731 161509
rect 504967 161273 509429 161509
rect 509665 161273 523335 161509
rect 523571 161273 528033 161509
rect 528269 161273 532731 161509
rect 532967 161273 537429 161509
rect 537665 161273 551335 161509
rect 551571 161273 556033 161509
rect 556269 161273 560731 161509
rect 560967 161273 565429 161509
rect 565665 161273 573526 161509
rect 573762 161273 573846 161509
rect 574082 161273 585342 161509
rect 585578 161273 585662 161509
rect 585898 161273 592650 161509
rect -8726 161241 592650 161273
rect -8726 158454 592650 158486
rect -8726 158218 -2934 158454
rect -2698 158218 -2614 158454
rect -2378 158218 21684 158454
rect 21920 158218 26382 158454
rect 26618 158218 31080 158454
rect 31316 158218 49684 158454
rect 49920 158218 54382 158454
rect 54618 158218 59080 158454
rect 59316 158218 77684 158454
rect 77920 158218 82382 158454
rect 82618 158218 87080 158454
rect 87316 158218 105684 158454
rect 105920 158218 110382 158454
rect 110618 158218 115080 158454
rect 115316 158218 133684 158454
rect 133920 158218 138382 158454
rect 138618 158218 143080 158454
rect 143316 158218 161684 158454
rect 161920 158218 166382 158454
rect 166618 158218 171080 158454
rect 171316 158218 189684 158454
rect 189920 158218 194382 158454
rect 194618 158218 199080 158454
rect 199316 158218 217684 158454
rect 217920 158218 222382 158454
rect 222618 158218 227080 158454
rect 227316 158218 245684 158454
rect 245920 158218 250382 158454
rect 250618 158218 255080 158454
rect 255316 158218 273684 158454
rect 273920 158218 278382 158454
rect 278618 158218 283080 158454
rect 283316 158218 301684 158454
rect 301920 158218 306382 158454
rect 306618 158218 311080 158454
rect 311316 158218 329684 158454
rect 329920 158218 334382 158454
rect 334618 158218 339080 158454
rect 339316 158218 357684 158454
rect 357920 158218 362382 158454
rect 362618 158218 367080 158454
rect 367316 158218 385684 158454
rect 385920 158218 390382 158454
rect 390618 158218 395080 158454
rect 395316 158218 413684 158454
rect 413920 158218 418382 158454
rect 418618 158218 423080 158454
rect 423316 158218 441684 158454
rect 441920 158218 446382 158454
rect 446618 158218 451080 158454
rect 451316 158218 469684 158454
rect 469920 158218 474382 158454
rect 474618 158218 479080 158454
rect 479316 158218 497684 158454
rect 497920 158218 502382 158454
rect 502618 158218 507080 158454
rect 507316 158218 525684 158454
rect 525920 158218 530382 158454
rect 530618 158218 535080 158454
rect 535316 158218 553684 158454
rect 553920 158218 558382 158454
rect 558618 158218 563080 158454
rect 563316 158218 586302 158454
rect 586538 158218 586622 158454
rect 586858 158218 592650 158454
rect -8726 158134 592650 158218
rect -8726 157898 -2934 158134
rect -2698 157898 -2614 158134
rect -2378 157898 21684 158134
rect 21920 157898 26382 158134
rect 26618 157898 31080 158134
rect 31316 157898 49684 158134
rect 49920 157898 54382 158134
rect 54618 157898 59080 158134
rect 59316 157898 77684 158134
rect 77920 157898 82382 158134
rect 82618 157898 87080 158134
rect 87316 157898 105684 158134
rect 105920 157898 110382 158134
rect 110618 157898 115080 158134
rect 115316 157898 133684 158134
rect 133920 157898 138382 158134
rect 138618 157898 143080 158134
rect 143316 157898 161684 158134
rect 161920 157898 166382 158134
rect 166618 157898 171080 158134
rect 171316 157898 189684 158134
rect 189920 157898 194382 158134
rect 194618 157898 199080 158134
rect 199316 157898 217684 158134
rect 217920 157898 222382 158134
rect 222618 157898 227080 158134
rect 227316 157898 245684 158134
rect 245920 157898 250382 158134
rect 250618 157898 255080 158134
rect 255316 157898 273684 158134
rect 273920 157898 278382 158134
rect 278618 157898 283080 158134
rect 283316 157898 301684 158134
rect 301920 157898 306382 158134
rect 306618 157898 311080 158134
rect 311316 157898 329684 158134
rect 329920 157898 334382 158134
rect 334618 157898 339080 158134
rect 339316 157898 357684 158134
rect 357920 157898 362382 158134
rect 362618 157898 367080 158134
rect 367316 157898 385684 158134
rect 385920 157898 390382 158134
rect 390618 157898 395080 158134
rect 395316 157898 413684 158134
rect 413920 157898 418382 158134
rect 418618 157898 423080 158134
rect 423316 157898 441684 158134
rect 441920 157898 446382 158134
rect 446618 157898 451080 158134
rect 451316 157898 469684 158134
rect 469920 157898 474382 158134
rect 474618 157898 479080 158134
rect 479316 157898 497684 158134
rect 497920 157898 502382 158134
rect 502618 157898 507080 158134
rect 507316 157898 525684 158134
rect 525920 157898 530382 158134
rect 530618 157898 535080 158134
rect 535316 157898 553684 158134
rect 553920 157898 558382 158134
rect 558618 157898 563080 158134
rect 563316 157898 586302 158134
rect 586538 157898 586622 158134
rect 586858 157898 592650 158134
rect -8726 157866 592650 157898
rect -8726 134829 592650 134861
rect -8726 134593 -1974 134829
rect -1738 134593 -1654 134829
rect -1418 134593 19335 134829
rect 19571 134593 24033 134829
rect 24269 134593 28731 134829
rect 28967 134593 33429 134829
rect 33665 134593 47335 134829
rect 47571 134593 52033 134829
rect 52269 134593 56731 134829
rect 56967 134593 61429 134829
rect 61665 134593 75335 134829
rect 75571 134593 80033 134829
rect 80269 134593 84731 134829
rect 84967 134593 89429 134829
rect 89665 134593 103335 134829
rect 103571 134593 108033 134829
rect 108269 134593 112731 134829
rect 112967 134593 117429 134829
rect 117665 134593 131335 134829
rect 131571 134593 136033 134829
rect 136269 134593 140731 134829
rect 140967 134593 145429 134829
rect 145665 134593 159335 134829
rect 159571 134593 164033 134829
rect 164269 134593 168731 134829
rect 168967 134593 173429 134829
rect 173665 134593 187335 134829
rect 187571 134593 192033 134829
rect 192269 134593 196731 134829
rect 196967 134593 201429 134829
rect 201665 134593 215335 134829
rect 215571 134593 220033 134829
rect 220269 134593 224731 134829
rect 224967 134593 229429 134829
rect 229665 134593 243335 134829
rect 243571 134593 248033 134829
rect 248269 134593 252731 134829
rect 252967 134593 257429 134829
rect 257665 134593 271335 134829
rect 271571 134593 276033 134829
rect 276269 134593 280731 134829
rect 280967 134593 285429 134829
rect 285665 134593 299335 134829
rect 299571 134593 304033 134829
rect 304269 134593 308731 134829
rect 308967 134593 313429 134829
rect 313665 134593 327335 134829
rect 327571 134593 332033 134829
rect 332269 134593 336731 134829
rect 336967 134593 341429 134829
rect 341665 134593 355335 134829
rect 355571 134593 360033 134829
rect 360269 134593 364731 134829
rect 364967 134593 369429 134829
rect 369665 134593 383335 134829
rect 383571 134593 388033 134829
rect 388269 134593 392731 134829
rect 392967 134593 397429 134829
rect 397665 134593 411335 134829
rect 411571 134593 416033 134829
rect 416269 134593 420731 134829
rect 420967 134593 425429 134829
rect 425665 134593 439335 134829
rect 439571 134593 444033 134829
rect 444269 134593 448731 134829
rect 448967 134593 453429 134829
rect 453665 134593 467335 134829
rect 467571 134593 472033 134829
rect 472269 134593 476731 134829
rect 476967 134593 481429 134829
rect 481665 134593 495335 134829
rect 495571 134593 500033 134829
rect 500269 134593 504731 134829
rect 504967 134593 509429 134829
rect 509665 134593 523335 134829
rect 523571 134593 528033 134829
rect 528269 134593 532731 134829
rect 532967 134593 537429 134829
rect 537665 134593 551335 134829
rect 551571 134593 556033 134829
rect 556269 134593 560731 134829
rect 560967 134593 565429 134829
rect 565665 134593 573526 134829
rect 573762 134593 573846 134829
rect 574082 134593 585342 134829
rect 585578 134593 585662 134829
rect 585898 134593 592650 134829
rect -8726 134509 592650 134593
rect -8726 134273 -1974 134509
rect -1738 134273 -1654 134509
rect -1418 134273 19335 134509
rect 19571 134273 24033 134509
rect 24269 134273 28731 134509
rect 28967 134273 33429 134509
rect 33665 134273 47335 134509
rect 47571 134273 52033 134509
rect 52269 134273 56731 134509
rect 56967 134273 61429 134509
rect 61665 134273 75335 134509
rect 75571 134273 80033 134509
rect 80269 134273 84731 134509
rect 84967 134273 89429 134509
rect 89665 134273 103335 134509
rect 103571 134273 108033 134509
rect 108269 134273 112731 134509
rect 112967 134273 117429 134509
rect 117665 134273 131335 134509
rect 131571 134273 136033 134509
rect 136269 134273 140731 134509
rect 140967 134273 145429 134509
rect 145665 134273 159335 134509
rect 159571 134273 164033 134509
rect 164269 134273 168731 134509
rect 168967 134273 173429 134509
rect 173665 134273 187335 134509
rect 187571 134273 192033 134509
rect 192269 134273 196731 134509
rect 196967 134273 201429 134509
rect 201665 134273 215335 134509
rect 215571 134273 220033 134509
rect 220269 134273 224731 134509
rect 224967 134273 229429 134509
rect 229665 134273 243335 134509
rect 243571 134273 248033 134509
rect 248269 134273 252731 134509
rect 252967 134273 257429 134509
rect 257665 134273 271335 134509
rect 271571 134273 276033 134509
rect 276269 134273 280731 134509
rect 280967 134273 285429 134509
rect 285665 134273 299335 134509
rect 299571 134273 304033 134509
rect 304269 134273 308731 134509
rect 308967 134273 313429 134509
rect 313665 134273 327335 134509
rect 327571 134273 332033 134509
rect 332269 134273 336731 134509
rect 336967 134273 341429 134509
rect 341665 134273 355335 134509
rect 355571 134273 360033 134509
rect 360269 134273 364731 134509
rect 364967 134273 369429 134509
rect 369665 134273 383335 134509
rect 383571 134273 388033 134509
rect 388269 134273 392731 134509
rect 392967 134273 397429 134509
rect 397665 134273 411335 134509
rect 411571 134273 416033 134509
rect 416269 134273 420731 134509
rect 420967 134273 425429 134509
rect 425665 134273 439335 134509
rect 439571 134273 444033 134509
rect 444269 134273 448731 134509
rect 448967 134273 453429 134509
rect 453665 134273 467335 134509
rect 467571 134273 472033 134509
rect 472269 134273 476731 134509
rect 476967 134273 481429 134509
rect 481665 134273 495335 134509
rect 495571 134273 500033 134509
rect 500269 134273 504731 134509
rect 504967 134273 509429 134509
rect 509665 134273 523335 134509
rect 523571 134273 528033 134509
rect 528269 134273 532731 134509
rect 532967 134273 537429 134509
rect 537665 134273 551335 134509
rect 551571 134273 556033 134509
rect 556269 134273 560731 134509
rect 560967 134273 565429 134509
rect 565665 134273 573526 134509
rect 573762 134273 573846 134509
rect 574082 134273 585342 134509
rect 585578 134273 585662 134509
rect 585898 134273 592650 134509
rect -8726 134241 592650 134273
rect -8726 131454 592650 131486
rect -8726 131218 -2934 131454
rect -2698 131218 -2614 131454
rect -2378 131218 21684 131454
rect 21920 131218 26382 131454
rect 26618 131218 31080 131454
rect 31316 131218 49684 131454
rect 49920 131218 54382 131454
rect 54618 131218 59080 131454
rect 59316 131218 77684 131454
rect 77920 131218 82382 131454
rect 82618 131218 87080 131454
rect 87316 131218 105684 131454
rect 105920 131218 110382 131454
rect 110618 131218 115080 131454
rect 115316 131218 133684 131454
rect 133920 131218 138382 131454
rect 138618 131218 143080 131454
rect 143316 131218 161684 131454
rect 161920 131218 166382 131454
rect 166618 131218 171080 131454
rect 171316 131218 189684 131454
rect 189920 131218 194382 131454
rect 194618 131218 199080 131454
rect 199316 131218 217684 131454
rect 217920 131218 222382 131454
rect 222618 131218 227080 131454
rect 227316 131218 245684 131454
rect 245920 131218 250382 131454
rect 250618 131218 255080 131454
rect 255316 131218 273684 131454
rect 273920 131218 278382 131454
rect 278618 131218 283080 131454
rect 283316 131218 301684 131454
rect 301920 131218 306382 131454
rect 306618 131218 311080 131454
rect 311316 131218 329684 131454
rect 329920 131218 334382 131454
rect 334618 131218 339080 131454
rect 339316 131218 357684 131454
rect 357920 131218 362382 131454
rect 362618 131218 367080 131454
rect 367316 131218 385684 131454
rect 385920 131218 390382 131454
rect 390618 131218 395080 131454
rect 395316 131218 413684 131454
rect 413920 131218 418382 131454
rect 418618 131218 423080 131454
rect 423316 131218 441684 131454
rect 441920 131218 446382 131454
rect 446618 131218 451080 131454
rect 451316 131218 469684 131454
rect 469920 131218 474382 131454
rect 474618 131218 479080 131454
rect 479316 131218 497684 131454
rect 497920 131218 502382 131454
rect 502618 131218 507080 131454
rect 507316 131218 525684 131454
rect 525920 131218 530382 131454
rect 530618 131218 535080 131454
rect 535316 131218 553684 131454
rect 553920 131218 558382 131454
rect 558618 131218 563080 131454
rect 563316 131218 586302 131454
rect 586538 131218 586622 131454
rect 586858 131218 592650 131454
rect -8726 131134 592650 131218
rect -8726 130898 -2934 131134
rect -2698 130898 -2614 131134
rect -2378 130898 21684 131134
rect 21920 130898 26382 131134
rect 26618 130898 31080 131134
rect 31316 130898 49684 131134
rect 49920 130898 54382 131134
rect 54618 130898 59080 131134
rect 59316 130898 77684 131134
rect 77920 130898 82382 131134
rect 82618 130898 87080 131134
rect 87316 130898 105684 131134
rect 105920 130898 110382 131134
rect 110618 130898 115080 131134
rect 115316 130898 133684 131134
rect 133920 130898 138382 131134
rect 138618 130898 143080 131134
rect 143316 130898 161684 131134
rect 161920 130898 166382 131134
rect 166618 130898 171080 131134
rect 171316 130898 189684 131134
rect 189920 130898 194382 131134
rect 194618 130898 199080 131134
rect 199316 130898 217684 131134
rect 217920 130898 222382 131134
rect 222618 130898 227080 131134
rect 227316 130898 245684 131134
rect 245920 130898 250382 131134
rect 250618 130898 255080 131134
rect 255316 130898 273684 131134
rect 273920 130898 278382 131134
rect 278618 130898 283080 131134
rect 283316 130898 301684 131134
rect 301920 130898 306382 131134
rect 306618 130898 311080 131134
rect 311316 130898 329684 131134
rect 329920 130898 334382 131134
rect 334618 130898 339080 131134
rect 339316 130898 357684 131134
rect 357920 130898 362382 131134
rect 362618 130898 367080 131134
rect 367316 130898 385684 131134
rect 385920 130898 390382 131134
rect 390618 130898 395080 131134
rect 395316 130898 413684 131134
rect 413920 130898 418382 131134
rect 418618 130898 423080 131134
rect 423316 130898 441684 131134
rect 441920 130898 446382 131134
rect 446618 130898 451080 131134
rect 451316 130898 469684 131134
rect 469920 130898 474382 131134
rect 474618 130898 479080 131134
rect 479316 130898 497684 131134
rect 497920 130898 502382 131134
rect 502618 130898 507080 131134
rect 507316 130898 525684 131134
rect 525920 130898 530382 131134
rect 530618 130898 535080 131134
rect 535316 130898 553684 131134
rect 553920 130898 558382 131134
rect 558618 130898 563080 131134
rect 563316 130898 586302 131134
rect 586538 130898 586622 131134
rect 586858 130898 592650 131134
rect -8726 130866 592650 130898
rect -8726 107829 592650 107861
rect -8726 107593 -1974 107829
rect -1738 107593 -1654 107829
rect -1418 107593 19335 107829
rect 19571 107593 24033 107829
rect 24269 107593 28731 107829
rect 28967 107593 33429 107829
rect 33665 107593 47335 107829
rect 47571 107593 52033 107829
rect 52269 107593 56731 107829
rect 56967 107593 61429 107829
rect 61665 107593 75335 107829
rect 75571 107593 80033 107829
rect 80269 107593 84731 107829
rect 84967 107593 89429 107829
rect 89665 107593 103335 107829
rect 103571 107593 108033 107829
rect 108269 107593 112731 107829
rect 112967 107593 117429 107829
rect 117665 107593 131335 107829
rect 131571 107593 136033 107829
rect 136269 107593 140731 107829
rect 140967 107593 145429 107829
rect 145665 107593 159335 107829
rect 159571 107593 164033 107829
rect 164269 107593 168731 107829
rect 168967 107593 173429 107829
rect 173665 107593 187335 107829
rect 187571 107593 192033 107829
rect 192269 107593 196731 107829
rect 196967 107593 201429 107829
rect 201665 107593 215335 107829
rect 215571 107593 220033 107829
rect 220269 107593 224731 107829
rect 224967 107593 229429 107829
rect 229665 107593 244118 107829
rect 244354 107593 250382 107829
rect 250618 107593 256646 107829
rect 256882 107593 271335 107829
rect 271571 107593 276033 107829
rect 276269 107593 280731 107829
rect 280967 107593 285429 107829
rect 285665 107593 299335 107829
rect 299571 107593 304033 107829
rect 304269 107593 308731 107829
rect 308967 107593 313429 107829
rect 313665 107593 328118 107829
rect 328354 107593 334382 107829
rect 334618 107593 340646 107829
rect 340882 107593 355335 107829
rect 355571 107593 360033 107829
rect 360269 107593 364731 107829
rect 364967 107593 369429 107829
rect 369665 107593 383335 107829
rect 383571 107593 388033 107829
rect 388269 107593 392731 107829
rect 392967 107593 397429 107829
rect 397665 107593 411335 107829
rect 411571 107593 416033 107829
rect 416269 107593 420731 107829
rect 420967 107593 425429 107829
rect 425665 107593 439335 107829
rect 439571 107593 444033 107829
rect 444269 107593 448731 107829
rect 448967 107593 453429 107829
rect 453665 107593 467335 107829
rect 467571 107593 472033 107829
rect 472269 107593 476731 107829
rect 476967 107593 481429 107829
rect 481665 107593 495335 107829
rect 495571 107593 500033 107829
rect 500269 107593 504731 107829
rect 504967 107593 509429 107829
rect 509665 107593 523335 107829
rect 523571 107593 528033 107829
rect 528269 107593 532731 107829
rect 532967 107593 537429 107829
rect 537665 107593 551335 107829
rect 551571 107593 556033 107829
rect 556269 107593 560731 107829
rect 560967 107593 565429 107829
rect 565665 107593 573526 107829
rect 573762 107593 573846 107829
rect 574082 107593 585342 107829
rect 585578 107593 585662 107829
rect 585898 107593 592650 107829
rect -8726 107509 592650 107593
rect -8726 107273 -1974 107509
rect -1738 107273 -1654 107509
rect -1418 107273 19335 107509
rect 19571 107273 24033 107509
rect 24269 107273 28731 107509
rect 28967 107273 33429 107509
rect 33665 107273 47335 107509
rect 47571 107273 52033 107509
rect 52269 107273 56731 107509
rect 56967 107273 61429 107509
rect 61665 107273 75335 107509
rect 75571 107273 80033 107509
rect 80269 107273 84731 107509
rect 84967 107273 89429 107509
rect 89665 107273 103335 107509
rect 103571 107273 108033 107509
rect 108269 107273 112731 107509
rect 112967 107273 117429 107509
rect 117665 107273 131335 107509
rect 131571 107273 136033 107509
rect 136269 107273 140731 107509
rect 140967 107273 145429 107509
rect 145665 107273 159335 107509
rect 159571 107273 164033 107509
rect 164269 107273 168731 107509
rect 168967 107273 173429 107509
rect 173665 107273 187335 107509
rect 187571 107273 192033 107509
rect 192269 107273 196731 107509
rect 196967 107273 201429 107509
rect 201665 107273 215335 107509
rect 215571 107273 220033 107509
rect 220269 107273 224731 107509
rect 224967 107273 229429 107509
rect 229665 107273 244118 107509
rect 244354 107273 250382 107509
rect 250618 107273 256646 107509
rect 256882 107273 271335 107509
rect 271571 107273 276033 107509
rect 276269 107273 280731 107509
rect 280967 107273 285429 107509
rect 285665 107273 299335 107509
rect 299571 107273 304033 107509
rect 304269 107273 308731 107509
rect 308967 107273 313429 107509
rect 313665 107273 328118 107509
rect 328354 107273 334382 107509
rect 334618 107273 340646 107509
rect 340882 107273 355335 107509
rect 355571 107273 360033 107509
rect 360269 107273 364731 107509
rect 364967 107273 369429 107509
rect 369665 107273 383335 107509
rect 383571 107273 388033 107509
rect 388269 107273 392731 107509
rect 392967 107273 397429 107509
rect 397665 107273 411335 107509
rect 411571 107273 416033 107509
rect 416269 107273 420731 107509
rect 420967 107273 425429 107509
rect 425665 107273 439335 107509
rect 439571 107273 444033 107509
rect 444269 107273 448731 107509
rect 448967 107273 453429 107509
rect 453665 107273 467335 107509
rect 467571 107273 472033 107509
rect 472269 107273 476731 107509
rect 476967 107273 481429 107509
rect 481665 107273 495335 107509
rect 495571 107273 500033 107509
rect 500269 107273 504731 107509
rect 504967 107273 509429 107509
rect 509665 107273 523335 107509
rect 523571 107273 528033 107509
rect 528269 107273 532731 107509
rect 532967 107273 537429 107509
rect 537665 107273 551335 107509
rect 551571 107273 556033 107509
rect 556269 107273 560731 107509
rect 560967 107273 565429 107509
rect 565665 107273 573526 107509
rect 573762 107273 573846 107509
rect 574082 107273 585342 107509
rect 585578 107273 585662 107509
rect 585898 107273 592650 107509
rect -8726 107241 592650 107273
rect -8726 104454 592650 104486
rect -8726 104218 -2934 104454
rect -2698 104218 -2614 104454
rect -2378 104218 21684 104454
rect 21920 104218 26382 104454
rect 26618 104218 31080 104454
rect 31316 104218 49684 104454
rect 49920 104218 54382 104454
rect 54618 104218 59080 104454
rect 59316 104218 77684 104454
rect 77920 104218 82382 104454
rect 82618 104218 87080 104454
rect 87316 104218 105684 104454
rect 105920 104218 110382 104454
rect 110618 104218 115080 104454
rect 115316 104218 133684 104454
rect 133920 104218 138382 104454
rect 138618 104218 143080 104454
rect 143316 104218 161684 104454
rect 161920 104218 166382 104454
rect 166618 104218 171080 104454
rect 171316 104218 189684 104454
rect 189920 104218 194382 104454
rect 194618 104218 199080 104454
rect 199316 104218 217684 104454
rect 217920 104218 222382 104454
rect 222618 104218 227080 104454
rect 227316 104218 247250 104454
rect 247486 104218 253514 104454
rect 253750 104218 273684 104454
rect 273920 104218 278382 104454
rect 278618 104218 283080 104454
rect 283316 104218 301684 104454
rect 301920 104218 306382 104454
rect 306618 104218 311080 104454
rect 311316 104218 331250 104454
rect 331486 104218 337514 104454
rect 337750 104218 357684 104454
rect 357920 104218 362382 104454
rect 362618 104218 367080 104454
rect 367316 104218 385684 104454
rect 385920 104218 390382 104454
rect 390618 104218 395080 104454
rect 395316 104218 413684 104454
rect 413920 104218 418382 104454
rect 418618 104218 423080 104454
rect 423316 104218 441684 104454
rect 441920 104218 446382 104454
rect 446618 104218 451080 104454
rect 451316 104218 469684 104454
rect 469920 104218 474382 104454
rect 474618 104218 479080 104454
rect 479316 104218 497684 104454
rect 497920 104218 502382 104454
rect 502618 104218 507080 104454
rect 507316 104218 525684 104454
rect 525920 104218 530382 104454
rect 530618 104218 535080 104454
rect 535316 104218 553684 104454
rect 553920 104218 558382 104454
rect 558618 104218 563080 104454
rect 563316 104218 586302 104454
rect 586538 104218 586622 104454
rect 586858 104218 592650 104454
rect -8726 104134 592650 104218
rect -8726 103898 -2934 104134
rect -2698 103898 -2614 104134
rect -2378 103898 21684 104134
rect 21920 103898 26382 104134
rect 26618 103898 31080 104134
rect 31316 103898 49684 104134
rect 49920 103898 54382 104134
rect 54618 103898 59080 104134
rect 59316 103898 77684 104134
rect 77920 103898 82382 104134
rect 82618 103898 87080 104134
rect 87316 103898 105684 104134
rect 105920 103898 110382 104134
rect 110618 103898 115080 104134
rect 115316 103898 133684 104134
rect 133920 103898 138382 104134
rect 138618 103898 143080 104134
rect 143316 103898 161684 104134
rect 161920 103898 166382 104134
rect 166618 103898 171080 104134
rect 171316 103898 189684 104134
rect 189920 103898 194382 104134
rect 194618 103898 199080 104134
rect 199316 103898 217684 104134
rect 217920 103898 222382 104134
rect 222618 103898 227080 104134
rect 227316 103898 247250 104134
rect 247486 103898 253514 104134
rect 253750 103898 273684 104134
rect 273920 103898 278382 104134
rect 278618 103898 283080 104134
rect 283316 103898 301684 104134
rect 301920 103898 306382 104134
rect 306618 103898 311080 104134
rect 311316 103898 331250 104134
rect 331486 103898 337514 104134
rect 337750 103898 357684 104134
rect 357920 103898 362382 104134
rect 362618 103898 367080 104134
rect 367316 103898 385684 104134
rect 385920 103898 390382 104134
rect 390618 103898 395080 104134
rect 395316 103898 413684 104134
rect 413920 103898 418382 104134
rect 418618 103898 423080 104134
rect 423316 103898 441684 104134
rect 441920 103898 446382 104134
rect 446618 103898 451080 104134
rect 451316 103898 469684 104134
rect 469920 103898 474382 104134
rect 474618 103898 479080 104134
rect 479316 103898 497684 104134
rect 497920 103898 502382 104134
rect 502618 103898 507080 104134
rect 507316 103898 525684 104134
rect 525920 103898 530382 104134
rect 530618 103898 535080 104134
rect 535316 103898 553684 104134
rect 553920 103898 558382 104134
rect 558618 103898 563080 104134
rect 563316 103898 586302 104134
rect 586538 103898 586622 104134
rect 586858 103898 592650 104134
rect -8726 103866 592650 103898
rect -8726 80829 592650 80861
rect -8726 80593 -1974 80829
rect -1738 80593 -1654 80829
rect -1418 80593 20118 80829
rect 20354 80593 26382 80829
rect 26618 80593 32646 80829
rect 32882 80593 48118 80829
rect 48354 80593 54382 80829
rect 54618 80593 60646 80829
rect 60882 80593 76118 80829
rect 76354 80593 82382 80829
rect 82618 80593 88646 80829
rect 88882 80593 103335 80829
rect 103571 80593 108033 80829
rect 108269 80593 112731 80829
rect 112967 80593 117429 80829
rect 117665 80593 131335 80829
rect 131571 80593 136033 80829
rect 136269 80593 140731 80829
rect 140967 80593 145429 80829
rect 145665 80593 159335 80829
rect 159571 80593 164033 80829
rect 164269 80593 168731 80829
rect 168967 80593 173429 80829
rect 173665 80593 188118 80829
rect 188354 80593 194382 80829
rect 194618 80593 200646 80829
rect 200882 80593 216118 80829
rect 216354 80593 222382 80829
rect 222618 80593 228646 80829
rect 228882 80593 244118 80829
rect 244354 80593 250382 80829
rect 250618 80593 256646 80829
rect 256882 80593 272118 80829
rect 272354 80593 278382 80829
rect 278618 80593 284646 80829
rect 284882 80593 300118 80829
rect 300354 80593 306382 80829
rect 306618 80593 312646 80829
rect 312882 80593 328118 80829
rect 328354 80593 334382 80829
rect 334618 80593 340646 80829
rect 340882 80593 355335 80829
rect 355571 80593 360033 80829
rect 360269 80593 364731 80829
rect 364967 80593 369429 80829
rect 369665 80593 383335 80829
rect 383571 80593 388033 80829
rect 388269 80593 392731 80829
rect 392967 80593 397429 80829
rect 397665 80593 411335 80829
rect 411571 80593 416033 80829
rect 416269 80593 420731 80829
rect 420967 80593 425429 80829
rect 425665 80593 439335 80829
rect 439571 80593 444033 80829
rect 444269 80593 448731 80829
rect 448967 80593 453429 80829
rect 453665 80593 467335 80829
rect 467571 80593 472033 80829
rect 472269 80593 476731 80829
rect 476967 80593 481429 80829
rect 481665 80593 495335 80829
rect 495571 80593 500033 80829
rect 500269 80593 504731 80829
rect 504967 80593 509429 80829
rect 509665 80593 523335 80829
rect 523571 80593 528033 80829
rect 528269 80593 532731 80829
rect 532967 80593 537429 80829
rect 537665 80593 551335 80829
rect 551571 80593 556033 80829
rect 556269 80593 560731 80829
rect 560967 80593 565429 80829
rect 565665 80593 573526 80829
rect 573762 80593 573846 80829
rect 574082 80593 585342 80829
rect 585578 80593 585662 80829
rect 585898 80593 592650 80829
rect -8726 80509 592650 80593
rect -8726 80273 -1974 80509
rect -1738 80273 -1654 80509
rect -1418 80273 20118 80509
rect 20354 80273 26382 80509
rect 26618 80273 32646 80509
rect 32882 80273 48118 80509
rect 48354 80273 54382 80509
rect 54618 80273 60646 80509
rect 60882 80273 76118 80509
rect 76354 80273 82382 80509
rect 82618 80273 88646 80509
rect 88882 80273 103335 80509
rect 103571 80273 108033 80509
rect 108269 80273 112731 80509
rect 112967 80273 117429 80509
rect 117665 80273 131335 80509
rect 131571 80273 136033 80509
rect 136269 80273 140731 80509
rect 140967 80273 145429 80509
rect 145665 80273 159335 80509
rect 159571 80273 164033 80509
rect 164269 80273 168731 80509
rect 168967 80273 173429 80509
rect 173665 80273 188118 80509
rect 188354 80273 194382 80509
rect 194618 80273 200646 80509
rect 200882 80273 216118 80509
rect 216354 80273 222382 80509
rect 222618 80273 228646 80509
rect 228882 80273 244118 80509
rect 244354 80273 250382 80509
rect 250618 80273 256646 80509
rect 256882 80273 272118 80509
rect 272354 80273 278382 80509
rect 278618 80273 284646 80509
rect 284882 80273 300118 80509
rect 300354 80273 306382 80509
rect 306618 80273 312646 80509
rect 312882 80273 328118 80509
rect 328354 80273 334382 80509
rect 334618 80273 340646 80509
rect 340882 80273 355335 80509
rect 355571 80273 360033 80509
rect 360269 80273 364731 80509
rect 364967 80273 369429 80509
rect 369665 80273 383335 80509
rect 383571 80273 388033 80509
rect 388269 80273 392731 80509
rect 392967 80273 397429 80509
rect 397665 80273 411335 80509
rect 411571 80273 416033 80509
rect 416269 80273 420731 80509
rect 420967 80273 425429 80509
rect 425665 80273 439335 80509
rect 439571 80273 444033 80509
rect 444269 80273 448731 80509
rect 448967 80273 453429 80509
rect 453665 80273 467335 80509
rect 467571 80273 472033 80509
rect 472269 80273 476731 80509
rect 476967 80273 481429 80509
rect 481665 80273 495335 80509
rect 495571 80273 500033 80509
rect 500269 80273 504731 80509
rect 504967 80273 509429 80509
rect 509665 80273 523335 80509
rect 523571 80273 528033 80509
rect 528269 80273 532731 80509
rect 532967 80273 537429 80509
rect 537665 80273 551335 80509
rect 551571 80273 556033 80509
rect 556269 80273 560731 80509
rect 560967 80273 565429 80509
rect 565665 80273 573526 80509
rect 573762 80273 573846 80509
rect 574082 80273 585342 80509
rect 585578 80273 585662 80509
rect 585898 80273 592650 80509
rect -8726 80241 592650 80273
rect -8726 77454 592650 77486
rect -8726 77218 -2934 77454
rect -2698 77218 -2614 77454
rect -2378 77218 23250 77454
rect 23486 77218 29514 77454
rect 29750 77218 51250 77454
rect 51486 77218 57514 77454
rect 57750 77218 79250 77454
rect 79486 77218 85514 77454
rect 85750 77218 105684 77454
rect 105920 77218 110382 77454
rect 110618 77218 115080 77454
rect 115316 77218 133684 77454
rect 133920 77218 138382 77454
rect 138618 77218 143080 77454
rect 143316 77218 161684 77454
rect 161920 77218 166382 77454
rect 166618 77218 171080 77454
rect 171316 77218 191250 77454
rect 191486 77218 197514 77454
rect 197750 77218 219250 77454
rect 219486 77218 225514 77454
rect 225750 77218 247250 77454
rect 247486 77218 253514 77454
rect 253750 77218 275250 77454
rect 275486 77218 281514 77454
rect 281750 77218 303250 77454
rect 303486 77218 309514 77454
rect 309750 77218 331250 77454
rect 331486 77218 337514 77454
rect 337750 77218 357684 77454
rect 357920 77218 362382 77454
rect 362618 77218 367080 77454
rect 367316 77218 385684 77454
rect 385920 77218 390382 77454
rect 390618 77218 395080 77454
rect 395316 77218 413684 77454
rect 413920 77218 418382 77454
rect 418618 77218 423080 77454
rect 423316 77218 441684 77454
rect 441920 77218 446382 77454
rect 446618 77218 451080 77454
rect 451316 77218 469684 77454
rect 469920 77218 474382 77454
rect 474618 77218 479080 77454
rect 479316 77218 497684 77454
rect 497920 77218 502382 77454
rect 502618 77218 507080 77454
rect 507316 77218 525684 77454
rect 525920 77218 530382 77454
rect 530618 77218 535080 77454
rect 535316 77218 553684 77454
rect 553920 77218 558382 77454
rect 558618 77218 563080 77454
rect 563316 77218 586302 77454
rect 586538 77218 586622 77454
rect 586858 77218 592650 77454
rect -8726 77134 592650 77218
rect -8726 76898 -2934 77134
rect -2698 76898 -2614 77134
rect -2378 76898 23250 77134
rect 23486 76898 29514 77134
rect 29750 76898 51250 77134
rect 51486 76898 57514 77134
rect 57750 76898 79250 77134
rect 79486 76898 85514 77134
rect 85750 76898 105684 77134
rect 105920 76898 110382 77134
rect 110618 76898 115080 77134
rect 115316 76898 133684 77134
rect 133920 76898 138382 77134
rect 138618 76898 143080 77134
rect 143316 76898 161684 77134
rect 161920 76898 166382 77134
rect 166618 76898 171080 77134
rect 171316 76898 191250 77134
rect 191486 76898 197514 77134
rect 197750 76898 219250 77134
rect 219486 76898 225514 77134
rect 225750 76898 247250 77134
rect 247486 76898 253514 77134
rect 253750 76898 275250 77134
rect 275486 76898 281514 77134
rect 281750 76898 303250 77134
rect 303486 76898 309514 77134
rect 309750 76898 331250 77134
rect 331486 76898 337514 77134
rect 337750 76898 357684 77134
rect 357920 76898 362382 77134
rect 362618 76898 367080 77134
rect 367316 76898 385684 77134
rect 385920 76898 390382 77134
rect 390618 76898 395080 77134
rect 395316 76898 413684 77134
rect 413920 76898 418382 77134
rect 418618 76898 423080 77134
rect 423316 76898 441684 77134
rect 441920 76898 446382 77134
rect 446618 76898 451080 77134
rect 451316 76898 469684 77134
rect 469920 76898 474382 77134
rect 474618 76898 479080 77134
rect 479316 76898 497684 77134
rect 497920 76898 502382 77134
rect 502618 76898 507080 77134
rect 507316 76898 525684 77134
rect 525920 76898 530382 77134
rect 530618 76898 535080 77134
rect 535316 76898 553684 77134
rect 553920 76898 558382 77134
rect 558618 76898 563080 77134
rect 563316 76898 586302 77134
rect 586538 76898 586622 77134
rect 586858 76898 592650 77134
rect -8726 76866 592650 76898
rect -8726 53829 592650 53861
rect -8726 53593 -1974 53829
rect -1738 53593 -1654 53829
rect -1418 53593 20118 53829
rect 20354 53593 26382 53829
rect 26618 53593 32646 53829
rect 32882 53593 48118 53829
rect 48354 53593 54382 53829
rect 54618 53593 60646 53829
rect 60882 53593 76118 53829
rect 76354 53593 82382 53829
rect 82618 53593 88646 53829
rect 88882 53593 104118 53829
rect 104354 53593 110382 53829
rect 110618 53593 116646 53829
rect 116882 53593 132118 53829
rect 132354 53593 138382 53829
rect 138618 53593 144646 53829
rect 144882 53593 160118 53829
rect 160354 53593 166382 53829
rect 166618 53593 172646 53829
rect 172882 53593 188118 53829
rect 188354 53593 194382 53829
rect 194618 53593 200646 53829
rect 200882 53593 215335 53829
rect 215571 53593 220033 53829
rect 220269 53593 224731 53829
rect 224967 53593 229429 53829
rect 229665 53593 244118 53829
rect 244354 53593 250382 53829
rect 250618 53593 256646 53829
rect 256882 53593 272118 53829
rect 272354 53593 278382 53829
rect 278618 53593 284646 53829
rect 284882 53593 300118 53829
rect 300354 53593 306382 53829
rect 306618 53593 312646 53829
rect 312882 53593 327335 53829
rect 327571 53593 332033 53829
rect 332269 53593 336731 53829
rect 336967 53593 341429 53829
rect 341665 53593 356118 53829
rect 356354 53593 362382 53829
rect 362618 53593 368646 53829
rect 368882 53593 384118 53829
rect 384354 53593 390382 53829
rect 390618 53593 396646 53829
rect 396882 53593 412118 53829
rect 412354 53593 418382 53829
rect 418618 53593 424646 53829
rect 424882 53593 440118 53829
rect 440354 53593 446382 53829
rect 446618 53593 452646 53829
rect 452882 53593 468118 53829
rect 468354 53593 474382 53829
rect 474618 53593 480646 53829
rect 480882 53593 495335 53829
rect 495571 53593 500033 53829
rect 500269 53593 504731 53829
rect 504967 53593 509429 53829
rect 509665 53593 524118 53829
rect 524354 53593 530382 53829
rect 530618 53593 536646 53829
rect 536882 53593 552118 53829
rect 552354 53593 558382 53829
rect 558618 53593 564646 53829
rect 564882 53593 573526 53829
rect 573762 53593 573846 53829
rect 574082 53593 585342 53829
rect 585578 53593 585662 53829
rect 585898 53593 592650 53829
rect -8726 53509 592650 53593
rect -8726 53273 -1974 53509
rect -1738 53273 -1654 53509
rect -1418 53273 20118 53509
rect 20354 53273 26382 53509
rect 26618 53273 32646 53509
rect 32882 53273 48118 53509
rect 48354 53273 54382 53509
rect 54618 53273 60646 53509
rect 60882 53273 76118 53509
rect 76354 53273 82382 53509
rect 82618 53273 88646 53509
rect 88882 53273 104118 53509
rect 104354 53273 110382 53509
rect 110618 53273 116646 53509
rect 116882 53273 132118 53509
rect 132354 53273 138382 53509
rect 138618 53273 144646 53509
rect 144882 53273 160118 53509
rect 160354 53273 166382 53509
rect 166618 53273 172646 53509
rect 172882 53273 188118 53509
rect 188354 53273 194382 53509
rect 194618 53273 200646 53509
rect 200882 53273 215335 53509
rect 215571 53273 220033 53509
rect 220269 53273 224731 53509
rect 224967 53273 229429 53509
rect 229665 53273 244118 53509
rect 244354 53273 250382 53509
rect 250618 53273 256646 53509
rect 256882 53273 272118 53509
rect 272354 53273 278382 53509
rect 278618 53273 284646 53509
rect 284882 53273 300118 53509
rect 300354 53273 306382 53509
rect 306618 53273 312646 53509
rect 312882 53273 327335 53509
rect 327571 53273 332033 53509
rect 332269 53273 336731 53509
rect 336967 53273 341429 53509
rect 341665 53273 356118 53509
rect 356354 53273 362382 53509
rect 362618 53273 368646 53509
rect 368882 53273 384118 53509
rect 384354 53273 390382 53509
rect 390618 53273 396646 53509
rect 396882 53273 412118 53509
rect 412354 53273 418382 53509
rect 418618 53273 424646 53509
rect 424882 53273 440118 53509
rect 440354 53273 446382 53509
rect 446618 53273 452646 53509
rect 452882 53273 468118 53509
rect 468354 53273 474382 53509
rect 474618 53273 480646 53509
rect 480882 53273 495335 53509
rect 495571 53273 500033 53509
rect 500269 53273 504731 53509
rect 504967 53273 509429 53509
rect 509665 53273 524118 53509
rect 524354 53273 530382 53509
rect 530618 53273 536646 53509
rect 536882 53273 552118 53509
rect 552354 53273 558382 53509
rect 558618 53273 564646 53509
rect 564882 53273 573526 53509
rect 573762 53273 573846 53509
rect 574082 53273 585342 53509
rect 585578 53273 585662 53509
rect 585898 53273 592650 53509
rect -8726 53241 592650 53273
rect -8726 50454 592650 50486
rect -8726 50218 -2934 50454
rect -2698 50218 -2614 50454
rect -2378 50218 23250 50454
rect 23486 50218 29514 50454
rect 29750 50218 51250 50454
rect 51486 50218 57514 50454
rect 57750 50218 79250 50454
rect 79486 50218 85514 50454
rect 85750 50218 107250 50454
rect 107486 50218 113514 50454
rect 113750 50218 135250 50454
rect 135486 50218 141514 50454
rect 141750 50218 163250 50454
rect 163486 50218 169514 50454
rect 169750 50218 191250 50454
rect 191486 50218 197514 50454
rect 197750 50218 217684 50454
rect 217920 50218 222382 50454
rect 222618 50218 227080 50454
rect 227316 50218 247250 50454
rect 247486 50218 253514 50454
rect 253750 50218 275250 50454
rect 275486 50218 281514 50454
rect 281750 50218 303250 50454
rect 303486 50218 309514 50454
rect 309750 50218 329684 50454
rect 329920 50218 334382 50454
rect 334618 50218 339080 50454
rect 339316 50218 359250 50454
rect 359486 50218 365514 50454
rect 365750 50218 387250 50454
rect 387486 50218 393514 50454
rect 393750 50218 415250 50454
rect 415486 50218 421514 50454
rect 421750 50218 443250 50454
rect 443486 50218 449514 50454
rect 449750 50218 471250 50454
rect 471486 50218 477514 50454
rect 477750 50218 497684 50454
rect 497920 50218 502382 50454
rect 502618 50218 507080 50454
rect 507316 50218 527250 50454
rect 527486 50218 533514 50454
rect 533750 50218 555250 50454
rect 555486 50218 561514 50454
rect 561750 50218 586302 50454
rect 586538 50218 586622 50454
rect 586858 50218 592650 50454
rect -8726 50134 592650 50218
rect -8726 49898 -2934 50134
rect -2698 49898 -2614 50134
rect -2378 49898 23250 50134
rect 23486 49898 29514 50134
rect 29750 49898 51250 50134
rect 51486 49898 57514 50134
rect 57750 49898 79250 50134
rect 79486 49898 85514 50134
rect 85750 49898 107250 50134
rect 107486 49898 113514 50134
rect 113750 49898 135250 50134
rect 135486 49898 141514 50134
rect 141750 49898 163250 50134
rect 163486 49898 169514 50134
rect 169750 49898 191250 50134
rect 191486 49898 197514 50134
rect 197750 49898 217684 50134
rect 217920 49898 222382 50134
rect 222618 49898 227080 50134
rect 227316 49898 247250 50134
rect 247486 49898 253514 50134
rect 253750 49898 275250 50134
rect 275486 49898 281514 50134
rect 281750 49898 303250 50134
rect 303486 49898 309514 50134
rect 309750 49898 329684 50134
rect 329920 49898 334382 50134
rect 334618 49898 339080 50134
rect 339316 49898 359250 50134
rect 359486 49898 365514 50134
rect 365750 49898 387250 50134
rect 387486 49898 393514 50134
rect 393750 49898 415250 50134
rect 415486 49898 421514 50134
rect 421750 49898 443250 50134
rect 443486 49898 449514 50134
rect 449750 49898 471250 50134
rect 471486 49898 477514 50134
rect 477750 49898 497684 50134
rect 497920 49898 502382 50134
rect 502618 49898 507080 50134
rect 507316 49898 527250 50134
rect 527486 49898 533514 50134
rect 533750 49898 555250 50134
rect 555486 49898 561514 50134
rect 561750 49898 586302 50134
rect 586538 49898 586622 50134
rect 586858 49898 592650 50134
rect -8726 49866 592650 49898
rect -8726 26829 592650 26861
rect -8726 26593 -1974 26829
rect -1738 26593 -1654 26829
rect -1418 26593 22460 26829
rect 22696 26593 33408 26829
rect 33644 26593 44356 26829
rect 44592 26593 55304 26829
rect 55540 26593 76118 26829
rect 76354 26593 82382 26829
rect 82618 26593 88646 26829
rect 88882 26593 104118 26829
rect 104354 26593 110382 26829
rect 110618 26593 116646 26829
rect 116882 26593 132118 26829
rect 132354 26593 138382 26829
rect 138618 26593 144646 26829
rect 144882 26593 160118 26829
rect 160354 26593 166382 26829
rect 166618 26593 172646 26829
rect 172882 26593 188118 26829
rect 188354 26593 194382 26829
rect 194618 26593 200646 26829
rect 200882 26593 216118 26829
rect 216354 26593 222382 26829
rect 222618 26593 228646 26829
rect 228882 26593 244118 26829
rect 244354 26593 250382 26829
rect 250618 26593 256646 26829
rect 256882 26593 272118 26829
rect 272354 26593 278382 26829
rect 278618 26593 284646 26829
rect 284882 26593 300118 26829
rect 300354 26593 306382 26829
rect 306618 26593 312646 26829
rect 312882 26593 328118 26829
rect 328354 26593 334382 26829
rect 334618 26593 340646 26829
rect 340882 26593 355335 26829
rect 355571 26593 360033 26829
rect 360269 26593 364731 26829
rect 364967 26593 369429 26829
rect 369665 26593 384118 26829
rect 384354 26593 390382 26829
rect 390618 26593 396646 26829
rect 396882 26593 412118 26829
rect 412354 26593 418382 26829
rect 418618 26593 424646 26829
rect 424882 26593 440118 26829
rect 440354 26593 446382 26829
rect 446618 26593 452646 26829
rect 452882 26593 468118 26829
rect 468354 26593 474382 26829
rect 474618 26593 480646 26829
rect 480882 26593 496118 26829
rect 496354 26593 502382 26829
rect 502618 26593 508646 26829
rect 508882 26593 524118 26829
rect 524354 26593 530382 26829
rect 530618 26593 536646 26829
rect 536882 26593 552118 26829
rect 552354 26593 558382 26829
rect 558618 26593 564646 26829
rect 564882 26593 573526 26829
rect 573762 26593 573846 26829
rect 574082 26593 585342 26829
rect 585578 26593 585662 26829
rect 585898 26593 592650 26829
rect -8726 26509 592650 26593
rect -8726 26273 -1974 26509
rect -1738 26273 -1654 26509
rect -1418 26273 22460 26509
rect 22696 26273 33408 26509
rect 33644 26273 44356 26509
rect 44592 26273 55304 26509
rect 55540 26273 76118 26509
rect 76354 26273 82382 26509
rect 82618 26273 88646 26509
rect 88882 26273 104118 26509
rect 104354 26273 110382 26509
rect 110618 26273 116646 26509
rect 116882 26273 132118 26509
rect 132354 26273 138382 26509
rect 138618 26273 144646 26509
rect 144882 26273 160118 26509
rect 160354 26273 166382 26509
rect 166618 26273 172646 26509
rect 172882 26273 188118 26509
rect 188354 26273 194382 26509
rect 194618 26273 200646 26509
rect 200882 26273 216118 26509
rect 216354 26273 222382 26509
rect 222618 26273 228646 26509
rect 228882 26273 244118 26509
rect 244354 26273 250382 26509
rect 250618 26273 256646 26509
rect 256882 26273 272118 26509
rect 272354 26273 278382 26509
rect 278618 26273 284646 26509
rect 284882 26273 300118 26509
rect 300354 26273 306382 26509
rect 306618 26273 312646 26509
rect 312882 26273 328118 26509
rect 328354 26273 334382 26509
rect 334618 26273 340646 26509
rect 340882 26273 355335 26509
rect 355571 26273 360033 26509
rect 360269 26273 364731 26509
rect 364967 26273 369429 26509
rect 369665 26273 384118 26509
rect 384354 26273 390382 26509
rect 390618 26273 396646 26509
rect 396882 26273 412118 26509
rect 412354 26273 418382 26509
rect 418618 26273 424646 26509
rect 424882 26273 440118 26509
rect 440354 26273 446382 26509
rect 446618 26273 452646 26509
rect 452882 26273 468118 26509
rect 468354 26273 474382 26509
rect 474618 26273 480646 26509
rect 480882 26273 496118 26509
rect 496354 26273 502382 26509
rect 502618 26273 508646 26509
rect 508882 26273 524118 26509
rect 524354 26273 530382 26509
rect 530618 26273 536646 26509
rect 536882 26273 552118 26509
rect 552354 26273 558382 26509
rect 558618 26273 564646 26509
rect 564882 26273 573526 26509
rect 573762 26273 573846 26509
rect 574082 26273 585342 26509
rect 585578 26273 585662 26509
rect 585898 26273 592650 26509
rect -8726 26241 592650 26273
rect -8726 23454 592650 23486
rect -8726 23218 -2934 23454
rect -2698 23218 -2614 23454
rect -2378 23218 27934 23454
rect 28170 23218 38882 23454
rect 39118 23218 49830 23454
rect 50066 23218 60778 23454
rect 61014 23218 66026 23454
rect 66262 23218 66346 23454
rect 66582 23218 79250 23454
rect 79486 23218 85514 23454
rect 85750 23218 107250 23454
rect 107486 23218 113514 23454
rect 113750 23218 135250 23454
rect 135486 23218 141514 23454
rect 141750 23218 163250 23454
rect 163486 23218 169514 23454
rect 169750 23218 191250 23454
rect 191486 23218 197514 23454
rect 197750 23218 219250 23454
rect 219486 23218 225514 23454
rect 225750 23218 247250 23454
rect 247486 23218 253514 23454
rect 253750 23218 275250 23454
rect 275486 23218 281514 23454
rect 281750 23218 303250 23454
rect 303486 23218 309514 23454
rect 309750 23218 331250 23454
rect 331486 23218 337514 23454
rect 337750 23218 357684 23454
rect 357920 23218 362382 23454
rect 362618 23218 367080 23454
rect 367316 23218 387250 23454
rect 387486 23218 393514 23454
rect 393750 23218 415250 23454
rect 415486 23218 421514 23454
rect 421750 23218 443250 23454
rect 443486 23218 449514 23454
rect 449750 23218 471250 23454
rect 471486 23218 477514 23454
rect 477750 23218 499250 23454
rect 499486 23218 505514 23454
rect 505750 23218 527250 23454
rect 527486 23218 533514 23454
rect 533750 23218 555250 23454
rect 555486 23218 561514 23454
rect 561750 23218 586302 23454
rect 586538 23218 586622 23454
rect 586858 23218 592650 23454
rect -8726 23134 592650 23218
rect -8726 22898 -2934 23134
rect -2698 22898 -2614 23134
rect -2378 22898 27934 23134
rect 28170 22898 38882 23134
rect 39118 22898 49830 23134
rect 50066 22898 60778 23134
rect 61014 22898 66026 23134
rect 66262 22898 66346 23134
rect 66582 22898 79250 23134
rect 79486 22898 85514 23134
rect 85750 22898 107250 23134
rect 107486 22898 113514 23134
rect 113750 22898 135250 23134
rect 135486 22898 141514 23134
rect 141750 22898 163250 23134
rect 163486 22898 169514 23134
rect 169750 22898 191250 23134
rect 191486 22898 197514 23134
rect 197750 22898 219250 23134
rect 219486 22898 225514 23134
rect 225750 22898 247250 23134
rect 247486 22898 253514 23134
rect 253750 22898 275250 23134
rect 275486 22898 281514 23134
rect 281750 22898 303250 23134
rect 303486 22898 309514 23134
rect 309750 22898 331250 23134
rect 331486 22898 337514 23134
rect 337750 22898 357684 23134
rect 357920 22898 362382 23134
rect 362618 22898 367080 23134
rect 367316 22898 387250 23134
rect 387486 22898 393514 23134
rect 393750 22898 415250 23134
rect 415486 22898 421514 23134
rect 421750 22898 443250 23134
rect 443486 22898 449514 23134
rect 449750 22898 471250 23134
rect 471486 22898 477514 23134
rect 477750 22898 499250 23134
rect 499486 22898 505514 23134
rect 505750 22898 527250 23134
rect 527486 22898 533514 23134
rect 533750 22898 555250 23134
rect 555486 22898 561514 23134
rect 561750 22898 586302 23134
rect 586538 22898 586622 23134
rect 586858 22898 592650 23134
rect -8726 22866 592650 22898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 573526 -346
rect 573762 -582 573846 -346
rect 574082 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 573526 -666
rect 573762 -902 573846 -666
rect 574082 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 66026 -1306
rect 66262 -1542 66346 -1306
rect 66582 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 66026 -1626
rect 66262 -1862 66346 -1626
rect 66582 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use scan_controller  scan_controller
timestamp 0
transform 1 0 16000 0 1 16000
box -10 0 46000 20000
use scan_wrapper_1f985e14df1ed789231bb6e0189d6e39  scan_wrapper_1f985e14df1ed789231bb6e0189d6e39_44
timestamp 0
transform 1 0 184000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_019235602376235615  scan_wrapper_019235602376235615_77
timestamp 0
transform -1 0 37000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_0
timestamp 0
transform 1 0 72000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_152
timestamp 0
transform -1 0 177000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_153
timestamp 0
transform -1 0 149000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_154
timestamp 0
transform -1 0 121000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_155
timestamp 0
transform -1 0 93000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_156
timestamp 0
transform -1 0 65000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_157
timestamp 0
transform -1 0 37000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_158
timestamp 0
transform 1 0 16000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_159
timestamp 0
transform 1 0 44000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_160
timestamp 0
transform 1 0 72000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_161
timestamp 0
transform 1 0 100000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_162
timestamp 0
transform 1 0 128000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_163
timestamp 0
transform 1 0 156000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_164
timestamp 0
transform 1 0 184000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_165
timestamp 0
transform 1 0 212000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_166
timestamp 0
transform 1 0 240000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_167
timestamp 0
transform 1 0 268000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_168
timestamp 0
transform 1 0 296000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_169
timestamp 0
transform 1 0 324000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_170
timestamp 0
transform 1 0 352000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_171
timestamp 0
transform 1 0 380000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_172
timestamp 0
transform 1 0 408000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_173
timestamp 0
transform 1 0 436000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_174
timestamp 0
transform 1 0 464000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_175
timestamp 0
transform 1 0 492000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_176
timestamp 0
transform 1 0 520000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_177
timestamp 0
transform 1 0 548000 0 1 232000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_178
timestamp 0
transform -1 0 569000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_179
timestamp 0
transform -1 0 541000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_180
timestamp 0
transform -1 0 513000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_181
timestamp 0
transform -1 0 485000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_182
timestamp 0
transform -1 0 457000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_183
timestamp 0
transform -1 0 429000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_184
timestamp 0
transform -1 0 401000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_185
timestamp 0
transform -1 0 373000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_186
timestamp 0
transform -1 0 345000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_187
timestamp 0
transform -1 0 317000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_188
timestamp 0
transform -1 0 289000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_189
timestamp 0
transform -1 0 261000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_190
timestamp 0
transform -1 0 233000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_191
timestamp 0
transform -1 0 205000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_192
timestamp 0
transform -1 0 177000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_193
timestamp 0
transform -1 0 149000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_194
timestamp 0
transform -1 0 121000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_195
timestamp 0
transform -1 0 93000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_196
timestamp 0
transform -1 0 65000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_197
timestamp 0
transform -1 0 37000 0 -1 280000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_198
timestamp 0
transform 1 0 16000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_199
timestamp 0
transform 1 0 44000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_200
timestamp 0
transform 1 0 72000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_201
timestamp 0
transform 1 0 100000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_202
timestamp 0
transform 1 0 128000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_203
timestamp 0
transform 1 0 156000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_204
timestamp 0
transform 1 0 184000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_205
timestamp 0
transform 1 0 212000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_206
timestamp 0
transform 1 0 240000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_207
timestamp 0
transform 1 0 268000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_208
timestamp 0
transform 1 0 296000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_209
timestamp 0
transform 1 0 324000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_210
timestamp 0
transform 1 0 352000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_211
timestamp 0
transform 1 0 380000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_212
timestamp 0
transform 1 0 408000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_213
timestamp 0
transform 1 0 436000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_214
timestamp 0
transform 1 0 464000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_215
timestamp 0
transform 1 0 492000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_216
timestamp 0
transform 1 0 520000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_217
timestamp 0
transform 1 0 548000 0 1 286000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_218
timestamp 0
transform -1 0 569000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_219
timestamp 0
transform -1 0 541000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_220
timestamp 0
transform -1 0 513000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_221
timestamp 0
transform -1 0 485000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_222
timestamp 0
transform -1 0 457000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_223
timestamp 0
transform -1 0 429000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_224
timestamp 0
transform -1 0 401000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_225
timestamp 0
transform -1 0 373000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_226
timestamp 0
transform -1 0 345000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_227
timestamp 0
transform -1 0 317000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_228
timestamp 0
transform -1 0 289000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_229
timestamp 0
transform -1 0 261000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_230
timestamp 0
transform -1 0 233000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_231
timestamp 0
transform -1 0 205000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_232
timestamp 0
transform -1 0 177000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_233
timestamp 0
transform -1 0 149000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_234
timestamp 0
transform -1 0 121000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_235
timestamp 0
transform -1 0 93000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_236
timestamp 0
transform -1 0 65000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_237
timestamp 0
transform -1 0 37000 0 -1 334000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_238
timestamp 0
transform 1 0 16000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_239
timestamp 0
transform 1 0 44000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_240
timestamp 0
transform 1 0 72000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_241
timestamp 0
transform 1 0 100000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_242
timestamp 0
transform 1 0 128000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_243
timestamp 0
transform 1 0 156000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_244
timestamp 0
transform 1 0 184000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_245
timestamp 0
transform 1 0 212000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_246
timestamp 0
transform 1 0 240000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_247
timestamp 0
transform 1 0 268000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_248
timestamp 0
transform 1 0 296000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_249
timestamp 0
transform 1 0 324000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_250
timestamp 0
transform 1 0 352000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_251
timestamp 0
transform 1 0 380000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_252
timestamp 0
transform 1 0 408000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_253
timestamp 0
transform 1 0 436000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_254
timestamp 0
transform 1 0 464000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_255
timestamp 0
transform 1 0 492000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_256
timestamp 0
transform 1 0 520000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_257
timestamp 0
transform 1 0 548000 0 1 340000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_258
timestamp 0
transform -1 0 569000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_259
timestamp 0
transform -1 0 541000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_260
timestamp 0
transform -1 0 513000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_261
timestamp 0
transform -1 0 485000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_262
timestamp 0
transform -1 0 457000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_263
timestamp 0
transform -1 0 429000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_264
timestamp 0
transform -1 0 401000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_265
timestamp 0
transform -1 0 373000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_266
timestamp 0
transform -1 0 345000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_267
timestamp 0
transform -1 0 317000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_268
timestamp 0
transform -1 0 289000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_269
timestamp 0
transform -1 0 261000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_270
timestamp 0
transform -1 0 233000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_271
timestamp 0
transform -1 0 205000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_272
timestamp 0
transform -1 0 177000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_273
timestamp 0
transform -1 0 149000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_274
timestamp 0
transform -1 0 121000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_275
timestamp 0
transform -1 0 93000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_276
timestamp 0
transform -1 0 65000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_277
timestamp 0
transform -1 0 37000 0 -1 388000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_278
timestamp 0
transform 1 0 16000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_279
timestamp 0
transform 1 0 44000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_280
timestamp 0
transform 1 0 72000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_281
timestamp 0
transform 1 0 100000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_282
timestamp 0
transform 1 0 128000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_283
timestamp 0
transform 1 0 156000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_284
timestamp 0
transform 1 0 184000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_285
timestamp 0
transform 1 0 212000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_286
timestamp 0
transform 1 0 240000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_287
timestamp 0
transform 1 0 268000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_288
timestamp 0
transform 1 0 296000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_289
timestamp 0
transform 1 0 324000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_290
timestamp 0
transform 1 0 352000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_291
timestamp 0
transform 1 0 380000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_292
timestamp 0
transform 1 0 408000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_293
timestamp 0
transform 1 0 436000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_294
timestamp 0
transform 1 0 464000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_295
timestamp 0
transform 1 0 492000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_296
timestamp 0
transform 1 0 520000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_297
timestamp 0
transform 1 0 548000 0 1 394000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_298
timestamp 0
transform -1 0 569000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_299
timestamp 0
transform -1 0 541000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_300
timestamp 0
transform -1 0 513000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_301
timestamp 0
transform -1 0 485000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_302
timestamp 0
transform -1 0 457000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_303
timestamp 0
transform -1 0 429000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_304
timestamp 0
transform -1 0 401000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_305
timestamp 0
transform -1 0 373000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_306
timestamp 0
transform -1 0 345000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_307
timestamp 0
transform -1 0 317000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_308
timestamp 0
transform -1 0 289000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_309
timestamp 0
transform -1 0 261000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_310
timestamp 0
transform -1 0 233000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_311
timestamp 0
transform -1 0 205000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_312
timestamp 0
transform -1 0 177000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_313
timestamp 0
transform -1 0 149000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_314
timestamp 0
transform -1 0 121000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_315
timestamp 0
transform -1 0 93000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_316
timestamp 0
transform -1 0 65000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_317
timestamp 0
transform -1 0 37000 0 -1 442000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_318
timestamp 0
transform 1 0 16000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_319
timestamp 0
transform 1 0 44000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_320
timestamp 0
transform 1 0 72000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_321
timestamp 0
transform 1 0 100000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_322
timestamp 0
transform 1 0 128000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_323
timestamp 0
transform 1 0 156000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_324
timestamp 0
transform 1 0 184000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_325
timestamp 0
transform 1 0 212000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_326
timestamp 0
transform 1 0 240000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_327
timestamp 0
transform 1 0 268000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_328
timestamp 0
transform 1 0 296000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_329
timestamp 0
transform 1 0 324000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_330
timestamp 0
transform 1 0 352000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_331
timestamp 0
transform 1 0 380000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_332
timestamp 0
transform 1 0 408000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_333
timestamp 0
transform 1 0 436000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_334
timestamp 0
transform 1 0 464000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_335
timestamp 0
transform 1 0 492000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_336
timestamp 0
transform 1 0 520000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_337
timestamp 0
transform 1 0 548000 0 1 448000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_338
timestamp 0
transform -1 0 569000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_339
timestamp 0
transform -1 0 541000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_340
timestamp 0
transform -1 0 513000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_341
timestamp 0
transform -1 0 485000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_342
timestamp 0
transform -1 0 457000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_343
timestamp 0
transform -1 0 429000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_344
timestamp 0
transform -1 0 401000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_345
timestamp 0
transform -1 0 373000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_346
timestamp 0
transform -1 0 345000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_347
timestamp 0
transform -1 0 317000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_348
timestamp 0
transform -1 0 289000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_349
timestamp 0
transform -1 0 261000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_350
timestamp 0
transform -1 0 233000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_351
timestamp 0
transform -1 0 205000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_352
timestamp 0
transform -1 0 177000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_353
timestamp 0
transform -1 0 149000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_354
timestamp 0
transform -1 0 121000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_355
timestamp 0
transform -1 0 93000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_356
timestamp 0
transform -1 0 65000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_357
timestamp 0
transform -1 0 37000 0 -1 496000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_358
timestamp 0
transform 1 0 16000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_359
timestamp 0
transform 1 0 44000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_360
timestamp 0
transform 1 0 72000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_361
timestamp 0
transform 1 0 100000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_362
timestamp 0
transform 1 0 128000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_363
timestamp 0
transform 1 0 156000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_364
timestamp 0
transform 1 0 184000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_365
timestamp 0
transform 1 0 212000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_366
timestamp 0
transform 1 0 240000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_367
timestamp 0
transform 1 0 268000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_368
timestamp 0
transform 1 0 296000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_369
timestamp 0
transform 1 0 324000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_370
timestamp 0
transform 1 0 352000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_371
timestamp 0
transform 1 0 380000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_372
timestamp 0
transform 1 0 408000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_373
timestamp 0
transform 1 0 436000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_374
timestamp 0
transform 1 0 464000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_375
timestamp 0
transform 1 0 492000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_376
timestamp 0
transform 1 0 520000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_377
timestamp 0
transform 1 0 548000 0 1 502000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_378
timestamp 0
transform -1 0 569000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_379
timestamp 0
transform -1 0 541000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_380
timestamp 0
transform -1 0 513000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_381
timestamp 0
transform -1 0 485000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_382
timestamp 0
transform -1 0 457000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_383
timestamp 0
transform -1 0 429000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_384
timestamp 0
transform -1 0 401000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_385
timestamp 0
transform -1 0 373000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_386
timestamp 0
transform -1 0 345000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_387
timestamp 0
transform -1 0 317000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_388
timestamp 0
transform -1 0 289000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_389
timestamp 0
transform -1 0 261000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_390
timestamp 0
transform -1 0 233000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_391
timestamp 0
transform -1 0 205000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_392
timestamp 0
transform -1 0 177000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_393
timestamp 0
transform -1 0 149000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_394
timestamp 0
transform -1 0 121000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_395
timestamp 0
transform -1 0 93000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_396
timestamp 0
transform -1 0 65000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_397
timestamp 0
transform -1 0 37000 0 -1 550000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_398
timestamp 0
transform 1 0 16000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_399
timestamp 0
transform 1 0 44000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_400
timestamp 0
transform 1 0 72000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_401
timestamp 0
transform 1 0 100000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_402
timestamp 0
transform 1 0 128000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_403
timestamp 0
transform 1 0 156000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_404
timestamp 0
transform 1 0 184000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_405
timestamp 0
transform 1 0 212000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_406
timestamp 0
transform 1 0 240000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_407
timestamp 0
transform 1 0 268000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_408
timestamp 0
transform 1 0 296000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_409
timestamp 0
transform 1 0 324000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_410
timestamp 0
transform 1 0 352000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_411
timestamp 0
transform 1 0 380000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_412
timestamp 0
transform 1 0 408000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_413
timestamp 0
transform 1 0 436000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_414
timestamp 0
transform 1 0 464000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_415
timestamp 0
transform 1 0 492000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_416
timestamp 0
transform 1 0 520000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_417
timestamp 0
transform 1 0 548000 0 1 556000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_418
timestamp 0
transform -1 0 569000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_419
timestamp 0
transform -1 0 541000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_420
timestamp 0
transform -1 0 513000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_421
timestamp 0
transform -1 0 485000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_422
timestamp 0
transform -1 0 457000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_423
timestamp 0
transform -1 0 429000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_424
timestamp 0
transform -1 0 401000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_425
timestamp 0
transform -1 0 373000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_426
timestamp 0
transform -1 0 345000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_427
timestamp 0
transform -1 0 317000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_428
timestamp 0
transform -1 0 289000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_429
timestamp 0
transform -1 0 261000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_430
timestamp 0
transform -1 0 233000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_431
timestamp 0
transform -1 0 205000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_432
timestamp 0
transform -1 0 177000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_433
timestamp 0
transform -1 0 149000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_434
timestamp 0
transform -1 0 121000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_435
timestamp 0
transform -1 0 93000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_436
timestamp 0
transform -1 0 65000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_437
timestamp 0
transform -1 0 37000 0 -1 604000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_438
timestamp 0
transform 1 0 16000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_439
timestamp 0
transform 1 0 44000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_440
timestamp 0
transform 1 0 72000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_441
timestamp 0
transform 1 0 100000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_442
timestamp 0
transform 1 0 128000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_443
timestamp 0
transform 1 0 156000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_444
timestamp 0
transform 1 0 184000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_445
timestamp 0
transform 1 0 212000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_446
timestamp 0
transform 1 0 240000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_447
timestamp 0
transform 1 0 268000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_448
timestamp 0
transform 1 0 296000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_449
timestamp 0
transform 1 0 324000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_450
timestamp 0
transform 1 0 352000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_451
timestamp 0
transform 1 0 380000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_452
timestamp 0
transform 1 0 408000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_453
timestamp 0
transform 1 0 436000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_454
timestamp 0
transform 1 0 464000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_455
timestamp 0
transform 1 0 492000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_456
timestamp 0
transform 1 0 520000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_457
timestamp 0
transform 1 0 548000 0 1 610000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_458
timestamp 0
transform -1 0 569000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_459
timestamp 0
transform -1 0 541000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_460
timestamp 0
transform -1 0 513000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_461
timestamp 0
transform -1 0 485000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_462
timestamp 0
transform -1 0 457000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_463
timestamp 0
transform -1 0 429000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_464
timestamp 0
transform -1 0 401000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_465
timestamp 0
transform -1 0 373000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_466
timestamp 0
transform -1 0 345000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_467
timestamp 0
transform -1 0 317000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_468
timestamp 0
transform -1 0 289000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_469
timestamp 0
transform -1 0 261000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_470
timestamp 0
transform -1 0 233000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_471
timestamp 0
transform -1 0 205000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_472
timestamp 0
transform -1 0 177000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_473
timestamp 0
transform -1 0 149000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_474
timestamp 0
transform -1 0 121000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_475
timestamp 0
transform -1 0 93000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_476
timestamp 0
transform -1 0 65000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_477
timestamp 0
transform -1 0 37000 0 -1 658000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_478
timestamp 0
transform 1 0 16000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_479
timestamp 0
transform 1 0 44000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_480
timestamp 0
transform 1 0 72000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_481
timestamp 0
transform 1 0 100000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_482
timestamp 0
transform 1 0 128000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_483
timestamp 0
transform 1 0 156000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_484
timestamp 0
transform 1 0 184000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_485
timestamp 0
transform 1 0 212000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_486
timestamp 0
transform 1 0 240000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_487
timestamp 0
transform 1 0 268000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_488
timestamp 0
transform 1 0 296000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_489
timestamp 0
transform 1 0 324000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_490
timestamp 0
transform 1 0 352000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_491
timestamp 0
transform 1 0 380000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_492
timestamp 0
transform 1 0 408000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_493
timestamp 0
transform 1 0 436000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_494
timestamp 0
transform 1 0 464000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_495
timestamp 0
transform 1 0 492000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_496
timestamp 0
transform 1 0 520000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_497
timestamp 0
transform 1 0 548000 0 1 664000
box 0 0 21000 21000
use scan_wrapper_339688086163161683  scan_wrapper_339688086163161683_1
timestamp 0
transform 1 0 100000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_339800239192932947  scan_wrapper_339800239192932947_7
timestamp 0
transform 1 0 268000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_340067262721426004  scan_wrapper_340067262721426004_96
timestamp 0
transform 1 0 520000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_340218629792465491  scan_wrapper_340218629792465491_2
timestamp 0
transform 1 0 128000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_340285391309374034  scan_wrapper_340285391309374034_4
timestamp 0
transform 1 0 184000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_340318610245288530  scan_wrapper_340318610245288530_3
timestamp 0
transform 1 0 156000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_340579111348994642  scan_wrapper_340579111348994642_30
timestamp 0
transform -1 0 233000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_340596276030603858  scan_wrapper_340596276030603858_150
timestamp 0
transform -1 0 233000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_340661930553246290  scan_wrapper_340661930553246290_5
timestamp 0
transform 1 0 212000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_340979268609638995  scan_wrapper_340979268609638995_116
timestamp 0
transform -1 0 65000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341063825089364563  scan_wrapper_341063825089364563_68
timestamp 0
transform -1 0 289000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341136771628663380  scan_wrapper_341136771628663380_6
timestamp 0
transform 1 0 240000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_341152580068442706  scan_wrapper_341152580068442706_15
timestamp 0
transform 1 0 492000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_341154068332282450  scan_wrapper_341154068332282450_10
timestamp 0
transform 1 0 352000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_341154161238213203  scan_wrapper_341154161238213203_8
timestamp 0
transform 1 0 296000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_341155178824598098  scan_wrapper_341155178824598098_16
timestamp 0
transform 1 0 520000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_341159915403870803  scan_wrapper_341159915403870803_9
timestamp 0
transform 1 0 324000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_341160201697624660  scan_wrapper_341160201697624660_11
timestamp 0
transform 1 0 380000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_341160271679586899  scan_wrapper_341160271679586899_13
timestamp 0
transform 1 0 436000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_341161378978988626  scan_wrapper_341161378978988626_14
timestamp 0
transform 1 0 464000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_341162950004834900  scan_wrapper_341162950004834900_25
timestamp 0
transform -1 0 373000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341163800289870419  scan_wrapper_341163800289870419_12
timestamp 0
transform 1 0 408000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_341164228775772755  scan_wrapper_341164228775772755_38
timestamp 0
transform 1 0 16000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341164910646919762  scan_wrapper_341164910646919762_34
timestamp 0
transform -1 0 121000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341167691532337747  scan_wrapper_341167691532337747_17
timestamp 0
transform 1 0 548000 0 1 16000
box 0 0 21000 21000
use scan_wrapper_341174480471589458  scan_wrapper_341174480471589458_69
timestamp 0
transform -1 0 261000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341174563322724948  scan_wrapper_341174563322724948_40
timestamp 0
transform 1 0 72000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341176884318437971  scan_wrapper_341176884318437971_20
timestamp 0
transform -1 0 513000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341178154799333971  scan_wrapper_341178154799333971_18
timestamp 0
transform -1 0 569000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341178296293130834  scan_wrapper_341178296293130834_43
timestamp 0
transform 1 0 156000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341178481588044372  scan_wrapper_341178481588044372_19
timestamp 0
transform -1 0 541000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341182944314917460  scan_wrapper_341182944314917460_21
timestamp 0
transform -1 0 485000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341188777753969234  scan_wrapper_341188777753969234_22
timestamp 0
transform -1 0 457000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341191836498395731  scan_wrapper_341191836498395731_27
timestamp 0
transform -1 0 317000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341192113929585235  scan_wrapper_341192113929585235_28
timestamp 0
transform -1 0 289000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341192621088047698  scan_wrapper_341192621088047698_29
timestamp 0
transform -1 0 261000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341193419111006803  scan_wrapper_341193419111006803_56
timestamp 0
transform 1 0 520000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341194143598379604  scan_wrapper_341194143598379604_23
timestamp 0
transform -1 0 429000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341202178192441940  scan_wrapper_341202178192441940_26
timestamp 0
transform -1 0 345000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341205508016833108  scan_wrapper_341205508016833108_24
timestamp 0
transform -1 0 401000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341224613878956628  scan_wrapper_341224613878956628_31
timestamp 0
transform -1 0 205000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341233739099013714  scan_wrapper_341233739099013714_35
timestamp 0
transform -1 0 93000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341235575572922964  scan_wrapper_341235575572922964_33
timestamp 0
transform -1 0 149000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341235973870322258  scan_wrapper_341235973870322258_32
timestamp 0
transform -1 0 177000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341240110454407762  scan_wrapper_341240110454407762_36
timestamp 0
transform -1 0 65000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341243232292700755  scan_wrapper_341243232292700755_102
timestamp 0
transform -1 0 457000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341259651269001812  scan_wrapper_341259651269001812_53
timestamp 0
transform 1 0 436000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341262321634509394  scan_wrapper_341262321634509394_39
timestamp 0
transform 1 0 44000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341263346544149074  scan_wrapper_341263346544149074_46
timestamp 0
transform 1 0 240000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341264068701586004  scan_wrapper_341264068701586004_37
timestamp 0
transform -1 0 37000 0 -1 64000
box 0 0 21000 21000
use scan_wrapper_341266732010177108  scan_wrapper_341266732010177108_57
timestamp 0
transform 1 0 548000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341271902949474898  scan_wrapper_341271902949474898_41
timestamp 0
transform 1 0 100000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341277789473735250  scan_wrapper_341277789473735250_45
timestamp 0
transform 1 0 212000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341279123277087315  scan_wrapper_341279123277087315_62
timestamp 0
transform -1 0 457000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341296149788885588  scan_wrapper_341296149788885588_47
timestamp 0
transform 1 0 268000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341315210433266259  scan_wrapper_341315210433266259_60
timestamp 0
transform -1 0 513000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341332847867462227  scan_wrapper_341332847867462227_48
timestamp 0
transform 1 0 296000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341337976625693266  scan_wrapper_341337976625693266_49
timestamp 0
transform 1 0 324000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341339883600609876  scan_wrapper_341339883600609876_50
timestamp 0
transform 1 0 352000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341342096033055316  scan_wrapper_341342096033055316_52
timestamp 0
transform 1 0 408000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341344337258349139  scan_wrapper_341344337258349139_51
timestamp 0
transform 1 0 380000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341353777861755476  scan_wrapper_341353777861755476_58
timestamp 0
transform -1 0 569000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341353780122485332  scan_wrapper_341353780122485332_55
timestamp 0
transform 1 0 492000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341353928049295956  scan_wrapper_341353928049295956_54
timestamp 0
transform 1 0 464000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_341359404107432531  scan_wrapper_341359404107432531_59
timestamp 0
transform -1 0 541000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341360223723717202  scan_wrapper_341360223723717202_114
timestamp 0
transform -1 0 121000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341364381657858642  scan_wrapper_341364381657858642_61
timestamp 0
transform -1 0 485000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341382703379120723  scan_wrapper_341382703379120723_64
timestamp 0
transform -1 0 401000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341389786199622227  scan_wrapper_341389786199622227_65
timestamp 0
transform -1 0 373000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341399568412312147  scan_wrapper_341399568412312147_82
timestamp 0
transform 1 0 128000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341404507891040852  scan_wrapper_341404507891040852_66
timestamp 0
transform -1 0 345000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341410909669818963  scan_wrapper_341410909669818963_67
timestamp 0
transform -1 0 317000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341419328215712339  scan_wrapper_341419328215712339_70
timestamp 0
transform -1 0 233000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341423712597181012  scan_wrapper_341423712597181012_99
timestamp 0
transform -1 0 541000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341424636358034002  scan_wrapper_341424636358034002_110
timestamp 0
transform -1 0 233000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341426151397261906  scan_wrapper_341426151397261906_146
timestamp 0
transform -1 0 345000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_341431339142087251  scan_wrapper_341431339142087251_71
timestamp 0
transform -1 0 205000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341431502448362067  scan_wrapper_341431502448362067_107
timestamp 0
transform -1 0 317000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341432030163108435  scan_wrapper_341432030163108435_72
timestamp 0
transform -1 0 177000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341432284947153491  scan_wrapper_341432284947153491_80
timestamp 0
transform 1 0 72000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341438392303616596  scan_wrapper_341438392303616596_79
timestamp 0
transform 1 0 44000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341440114308678227  scan_wrapper_341440114308678227_73
timestamp 0
transform -1 0 149000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341440781874102868  scan_wrapper_341440781874102868_75
timestamp 0
transform -1 0 93000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341444501414347346  scan_wrapper_341444501414347346_76
timestamp 0
transform -1 0 65000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341446083683025490  scan_wrapper_341446083683025490_104
timestamp 0
transform -1 0 401000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341449297858921043  scan_wrapper_341449297858921043_94
timestamp 0
transform 1 0 464000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341450853309219412  scan_wrapper_341450853309219412_78
timestamp 0
transform 1 0 16000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341452019534398035  scan_wrapper_341452019534398035_86
timestamp 0
transform 1 0 240000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341457494561784402  scan_wrapper_341457494561784402_127
timestamp 0
transform 1 0 268000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341457971277988435  scan_wrapper_341457971277988435_81
timestamp 0
transform 1 0 100000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341462925422101075  scan_wrapper_341462925422101075_97
timestamp 0
transform 1 0 548000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341464767397888596  scan_wrapper_341464767397888596_83
timestamp 0
transform 1 0 156000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341473139924927058  scan_wrapper_341473139924927058_108
timestamp 0
transform -1 0 289000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341476989274686036  scan_wrapper_341476989274686036_84
timestamp 0
transform 1 0 184000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341482086419399252  scan_wrapper_341482086419399252_85
timestamp 0
transform 1 0 212000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341490465660469844  scan_wrapper_341490465660469844_125
timestamp 0
transform 1 0 212000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341493393195532884  scan_wrapper_341493393195532884_92
timestamp 0
transform 1 0 408000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341496918381167187  scan_wrapper_341496918381167187_74
timestamp 0
transform -1 0 121000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_341497938559631956  scan_wrapper_341497938559631956_89
timestamp 0
transform 1 0 324000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341497964482527828  scan_wrapper_341497964482527828_88
timestamp 0
transform 1 0 296000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341497971083313748  scan_wrapper_341497971083313748_87
timestamp 0
transform 1 0 268000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341499976001520211  scan_wrapper_341499976001520211_90
timestamp 0
transform 1 0 352000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341500800901579348  scan_wrapper_341500800901579348_91
timestamp 0
transform 1 0 380000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341506274933867090  scan_wrapper_341506274933867090_93
timestamp 0
transform 1 0 436000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341516949939814994  scan_wrapper_341516949939814994_100
timestamp 0
transform -1 0 513000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341519170869920338  scan_wrapper_341519170869920338_103
timestamp 0
transform -1 0 429000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341520747710120530  scan_wrapper_341520747710120530_98
timestamp 0
transform -1 0 569000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341521390605697619  scan_wrapper_341521390605697619_101
timestamp 0
transform -1 0 485000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341524192738411090  scan_wrapper_341524192738411090_105
timestamp 0
transform -1 0 373000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341528610027340372  scan_wrapper_341528610027340372_109
timestamp 0
transform -1 0 261000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341533740987581011  scan_wrapper_341533740987581011_106
timestamp 0
transform -1 0 345000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341538994733974098  scan_wrapper_341538994733974098_120
timestamp 0
transform 1 0 72000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341541108650607187  scan_wrapper_341541108650607187_113
timestamp 0
transform -1 0 149000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341542971476279892  scan_wrapper_341542971476279892_117
timestamp 0
transform -1 0 37000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341546888233747026  scan_wrapper_341546888233747026_115
timestamp 0
transform -1 0 93000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341556236196512338  scan_wrapper_341556236196512338_118
timestamp 0
transform 1 0 16000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341557831870186068  scan_wrapper_341557831870186068_121
timestamp 0
transform 1 0 100000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341558189536313940  scan_wrapper_341558189536313940_119
timestamp 0
transform 1 0 44000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341567111632519764  scan_wrapper_341567111632519764_140
timestamp 0
transform -1 0 513000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_341569483755749970  scan_wrapper_341569483755749970_122
timestamp 0
transform 1 0 128000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341571228858843732  scan_wrapper_341571228858843732_124
timestamp 0
transform 1 0 184000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341573751072096850  scan_wrapper_341573751072096850_123
timestamp 0
transform 1 0 156000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341581732833657427  scan_wrapper_341581732833657427_126
timestamp 0
transform 1 0 240000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341589685194195540  scan_wrapper_341589685194195540_129
timestamp 0
transform 1 0 324000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341590933015364178  scan_wrapper_341590933015364178_128
timestamp 0
transform 1 0 296000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341608297106768466  scan_wrapper_341608297106768466_131
timestamp 0
transform 1 0 380000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341608574336631379  scan_wrapper_341608574336631379_130
timestamp 0
transform 1 0 352000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341609034095264340  scan_wrapper_341609034095264340_133
timestamp 0
transform 1 0 436000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341613097060926036  scan_wrapper_341613097060926036_135
timestamp 0
transform 1 0 492000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341614346808328788  scan_wrapper_341614346808328788_136
timestamp 0
transform 1 0 520000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341614536664547922  scan_wrapper_341614536664547922_139
timestamp 0
transform -1 0 541000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_341617722294010450  scan_wrapper_341617722294010450_134
timestamp 0
transform 1 0 464000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341620484740219475  scan_wrapper_341620484740219475_137
timestamp 0
transform 1 0 548000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341624400621077076  scan_wrapper_341624400621077076_138
timestamp 0
transform -1 0 569000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_341628725785264722  scan_wrapper_341628725785264722_144
timestamp 0
transform -1 0 401000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_341629415144292948  scan_wrapper_341629415144292948_147
timestamp 0
transform -1 0 317000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_341631485498884690  scan_wrapper_341631485498884690_142
timestamp 0
transform -1 0 457000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_341631511790879314  scan_wrapper_341631511790879314_145
timestamp 0
transform -1 0 373000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_341631644820570706  scan_wrapper_341631644820570706_149
timestamp 0
transform -1 0 261000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_341632596577354323  scan_wrapper_341632596577354323_143
timestamp 0
transform -1 0 429000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_341637831098106450  scan_wrapper_341637831098106450_148
timestamp 0
transform -1 0 289000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_341678527574180436  scan_wrapper_341678527574180436_151
timestamp 0
transform -1 0 205000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_341710255833481812  scan_wrapper_341710255833481812_95
timestamp 0
transform 1 0 492000 0 1 124000
box 0 0 21000 21000
use scan_wrapper_341717091617866324  scan_wrapper_341717091617866324_111
timestamp 0
transform -1 0 205000 0 -1 172000
box 0 0 21000 21000
use scan_wrapper_341802448429515346  scan_wrapper_341802448429515346_132
timestamp 0
transform 1 0 408000 0 1 178000
box 0 0 21000 21000
use scan_wrapper_341802655228625490  scan_wrapper_341802655228625490_63
timestamp 0
transform -1 0 429000 0 -1 118000
box 0 0 21000 21000
use scan_wrapper_3398002391929329472  scan_wrapper_3398002391929329472_141
timestamp 0
transform -1 0 485000 0 -1 226000
box 0 0 21000 21000
use scan_wrapper_bc4d7220e4fdbf20a574d56ea112a8e1  scan_wrapper_bc4d7220e4fdbf20a574d56ea112a8e1_42
timestamp 0
transform 1 0 128000 0 1 70000
box 0 0 21000 21000
use scan_wrapper_hamming74  scan_wrapper_hamming74_112
timestamp 0
transform -1 0 177000 0 -1 172000
box 0 0 21000 21000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 41494 687000 42114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 69494 687000 70114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 97494 687000 98114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 125494 687000 126114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 153494 687000 154114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181494 687000 182114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 209494 687000 210114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 237494 687000 238114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 265494 687000 266114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 293494 687000 294114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 321494 687000 322114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 349494 687000 350114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 377494 687000 378114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 405494 687000 406114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433494 687000 434114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 461494 687000 462114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 489494 687000 490114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 517494 687000 518114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 545494 687000 546114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 573494 -7654 574114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 26241 592650 26861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 53241 592650 53861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 80241 592650 80861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 107241 592650 107861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 134241 592650 134861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 161241 592650 161861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 188241 592650 188861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 215241 592650 215861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 242241 592650 242861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 269241 592650 269861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 296241 592650 296861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 323241 592650 323861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 350241 592650 350861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 377241 592650 377861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 404241 592650 404861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 431241 592650 431861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 458241 592650 458861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 485241 592650 485861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 512241 592650 512861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 539241 592650 539861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 566241 592650 566861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 593241 592650 593861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 620241 592650 620861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 647241 592650 647861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 674241 592650 674861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 701241 592650 701861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 37994 687000 38614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 65994 -7654 66614 41000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 65994 687000 66614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 93994 687000 94614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 121994 687000 122614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149994 687000 150614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 177994 687000 178614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 205994 687000 206614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 233994 687000 234614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 261994 687000 262614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 289994 687000 290614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 317994 687000 318614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 345994 687000 346614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 373994 687000 374614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401994 687000 402614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 429994 687000 430614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 457994 687000 458614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 485994 687000 486614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 513994 687000 514614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 541994 687000 542614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 569994 687000 570614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 22866 592650 23486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 49866 592650 50486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 76866 592650 77486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 103866 592650 104486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 130866 592650 131486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 157866 592650 158486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 184866 592650 185486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 211866 592650 212486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 238866 592650 239486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 265866 592650 266486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 292866 592650 293486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 319866 592650 320486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 346866 592650 347486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 373866 592650 374486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 400866 592650 401486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 427866 592650 428486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 454866 592650 455486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 481866 592650 482486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 508866 592650 509486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 535866 592650 536486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 562866 592650 563486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 589866 592650 590486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 616866 592650 617486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 643866 592650 644486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 670866 592650 671486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 697866 592650 698486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
