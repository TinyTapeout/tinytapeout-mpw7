// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_project_wrapper
 *
 * This wrapper enumerates all of the pins available to the
 * user for the user project.
 *
 * An example user project is provided in this wrapper.  The
 * example should be removed and replaced with the actual
 * user project.
 *
 * THIS FILE HAS BEEN GENERATED USING multi_tools_project CODEGEN
 * IF YOU NEED TO MAKE EDITS TO IT, EDIT codegen/caravel_iface_header.txt
 *
 *-------------------------------------------------------------
 */

module user_project_wrapper #(
    parameter BITS = 32
)(
`ifdef USE_POWER_PINS
    inout vdda1,       // User area 1 3.3V supply
    inout vdda2,       // User area 2 3.3V supply
    inout vssa1,       // User area 1 analog ground
    inout vssa2,       // User area 2 analog ground
    inout vccd1,       // User area 1 1.8V supply
    inout vccd2,       // User area 2 1.8v supply
    inout vssd1,       // User area 1 digital ground
    inout vssd2,       // User area 2 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // Analog (direct connection to GPIO pad---use with caution)
    // Note that analog I/O is not available on the 7 lowest-numbered
    // GPIO pads, and so the analog_io indexing is offset from the
    // GPIO indexing by 7 (also upper 2 GPIOs do not have analog_io).
    inout [`MPRJ_IO_PADS-10:0] analog_io,

    // Independent clock (on independent integer divider)
    input   user_clock2,

    // User maskable interrupt signals
    output [2:0] user_irq
);

    // start of module instantiation

        localparam NUM_MACROS = 498;
        wire [NUM_MACROS:0] data, scan, latch, clk;
        
        scan_controller #(.NUM_DESIGNS(NUM_MACROS)) scan_controller(
            .clk                    (wb_clk_i),
            .reset                  (wb_rst_i),
            .active_select          (io_in[20:12]),
            .inputs                 (io_in[28:21]),
            .outputs                (io_out[36:29]),
            .ready                  (io_out[37]),
            .slow_clk               (io_out[10]),
            .set_clk_div            (io_in[11]),

            .scan_clk_out           (clk[0]),
            .scan_clk_in            (clk[NUM_MACROS]),
            .scan_data_out          (data[0]),
            .scan_data_in           (data[NUM_MACROS]),
            .scan_select            (scan[0]),
            .scan_latch_en          (latch[0]),

            .la_scan_clk_in         (la_data_in[0]),
            .la_scan_data_in        (la_data_in[1]),
            .la_scan_data_out       (la_data_out[0]),
            .la_scan_select         (la_data_in[2]),
            .la_scan_latch_en       (la_data_in[3]),

            .driver_sel             (io_in[9:8]),

            .oeb                    (io_oeb)
        );

        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_0 (
            .clk_in          (clk  [0]),
            .data_in         (data [0]),
            .scan_select_in  (scan [0]),
            .latch_enable_in (latch[0]),
            .clk_out         (clk  [1]),
            .data_out        (data [1]),
            .scan_select_out (scan [1]),
            .latch_enable_out(latch[1])
            );
        
        // https://github.com/mattvenn/tinytapeout_m_segments
        scan_wrapper_339688086163161683 #(.NUM_IOS(8)) scan_wrapper_339688086163161683_1 (
            .clk_in          (clk  [1]),
            .data_in         (data [1]),
            .scan_select_in  (scan [1]),
            .latch_enable_in (latch[1]),
            .clk_out         (clk  [2]),
            .data_out        (data [2]),
            .scan_select_out (scan [2]),
            .latch_enable_out(latch[2])
            );
        
        // https://github.com/gregdavill/tinytapeout_spin0
        scan_wrapper_340218629792465491 #(.NUM_IOS(8)) scan_wrapper_340218629792465491_2 (
            .clk_in          (clk  [2]),
            .data_in         (data [2]),
            .scan_select_in  (scan [2]),
            .latch_enable_in (latch[2]),
            .clk_out         (clk  [3]),
            .data_out        (data [3]),
            .scan_select_out (scan [3]),
            .latch_enable_out(latch[3])
            );
        
        // https://github.com/mole99/wokwi-1bit-alu
        scan_wrapper_340318610245288530 #(.NUM_IOS(8)) scan_wrapper_340318610245288530_3 (
            .clk_in          (clk  [3]),
            .data_in         (data [3]),
            .scan_select_in  (scan [3]),
            .latch_enable_in (latch[3]),
            .clk_out         (clk  [4]),
            .data_out        (data [4]),
            .scan_select_out (scan [4]),
            .latch_enable_out(latch[4])
            );
        
        // https://github.com/ericsmi/tinytapeout_popcnt.git
        scan_wrapper_340285391309374034 #(.NUM_IOS(8)) scan_wrapper_340285391309374034_4 (
            .clk_in          (clk  [4]),
            .data_in         (data [4]),
            .scan_select_in  (scan [4]),
            .latch_enable_in (latch[4]),
            .clk_out         (clk  [5]),
            .data_out        (data [5]),
            .scan_select_out (scan [5]),
            .latch_enable_out(latch[5])
            );
        
        // https://github.com/krasin/wokwi-guess-my-number
        scan_wrapper_340661930553246290 #(.NUM_IOS(8)) scan_wrapper_340661930553246290_5 (
            .clk_in          (clk  [5]),
            .data_in         (data [5]),
            .scan_select_in  (scan [5]),
            .latch_enable_in (latch[5]),
            .clk_out         (clk  [6]),
            .data_out        (data [6]),
            .scan_select_out (scan [6]),
            .latch_enable_out(latch[6])
            );
        
        // https://github.com/johshoff/barrelshifter-wokwi-gds
        scan_wrapper_341136771628663380 #(.NUM_IOS(8)) scan_wrapper_341136771628663380_6 (
            .clk_in          (clk  [6]),
            .data_in         (data [6]),
            .scan_select_in  (scan [6]),
            .latch_enable_in (latch[6]),
            .clk_out         (clk  [7]),
            .data_out        (data [7]),
            .scan_select_out (scan [7]),
            .latch_enable_out(latch[7])
            );
        
        // https://github.com/pretentious7/tinytapeout
        scan_wrapper_339800239192932947 #(.NUM_IOS(8)) scan_wrapper_339800239192932947_7 (
            .clk_in          (clk  [7]),
            .data_in         (data [7]),
            .scan_select_in  (scan [7]),
            .latch_enable_in (latch[7]),
            .clk_out         (clk  [8]),
            .data_out        (data [8]),
            .scan_select_out (scan [8]),
            .latch_enable_out(latch[8])
            );
        
        // https://github.com/GuzTech/wokwi-ripple-carry-adder
        scan_wrapper_341154161238213203 #(.NUM_IOS(8)) scan_wrapper_341154161238213203_8 (
            .clk_in          (clk  [8]),
            .data_in         (data [8]),
            .scan_select_in  (scan [8]),
            .latch_enable_in (latch[8]),
            .clk_out         (clk  [9]),
            .data_out        (data [9]),
            .scan_select_out (scan [9]),
            .latch_enable_out(latch[9])
            );
        
        // https://github.com/kbeckmann/tinytapeout_kbeckmann1
        scan_wrapper_341159915403870803 #(.NUM_IOS(8)) scan_wrapper_341159915403870803_9 (
            .clk_in          (clk  [9]),
            .data_in         (data [9]),
            .scan_select_in  (scan [9]),
            .latch_enable_in (latch[9]),
            .clk_out         (clk  [10]),
            .data_out        (data [10]),
            .scan_select_out (scan [10]),
            .latch_enable_out(latch[10])
            );
        
        // https://github.com/H-S-S-11/tinytapeout-verilog-test
        scan_wrapper_341154068332282450 #(.NUM_IOS(8)) scan_wrapper_341154068332282450_10 (
            .clk_in          (clk  [10]),
            .data_in         (data [10]),
            .scan_select_in  (scan [10]),
            .latch_enable_in (latch[10]),
            .clk_out         (clk  [11]),
            .data_out        (data [11]),
            .scan_select_out (scan [11]),
            .latch_enable_out(latch[11])
            );
        
        // https://github.com/skerr92/tinytapeout_frequency_div
        scan_wrapper_341160201697624660 #(.NUM_IOS(8)) scan_wrapper_341160201697624660_11 (
            .clk_in          (clk  [11]),
            .data_in         (data [11]),
            .scan_select_in  (scan [11]),
            .latch_enable_in (latch[11]),
            .clk_out         (clk  [12]),
            .data_out        (data [12]),
            .scan_select_out (scan [12]),
            .latch_enable_out(latch[12])
            );
        
        // https://github.com/argunda/tinytapeout_dualedgedetector
        scan_wrapper_341163800289870419 #(.NUM_IOS(8)) scan_wrapper_341163800289870419_12 (
            .clk_in          (clk  [12]),
            .data_in         (data [12]),
            .scan_select_in  (scan [12]),
            .latch_enable_in (latch[12]),
            .clk_out         (clk  [13]),
            .data_out        (data [13]),
            .scan_select_out (scan [13]),
            .latch_enable_out(latch[13])
            );
        
        // https://github.com/libokuohai/tinytapeout-2022-08
        scan_wrapper_341160271679586899 #(.NUM_IOS(8)) scan_wrapper_341160271679586899_13 (
            .clk_in          (clk  [13]),
            .data_in         (data [13]),
            .scan_select_in  (scan [13]),
            .latch_enable_in (latch[13]),
            .clk_out         (clk  [14]),
            .data_out        (data [14]),
            .scan_select_out (scan [14]),
            .latch_enable_out(latch[14])
            );
        
        // https://github.com/jglim/tinytapeout_bcd-dec
        scan_wrapper_341161378978988626 #(.NUM_IOS(8)) scan_wrapper_341161378978988626_14 (
            .clk_in          (clk  [14]),
            .data_in         (data [14]),
            .scan_select_in  (scan [14]),
            .latch_enable_in (latch[14]),
            .clk_out         (clk  [15]),
            .data_out        (data [15]),
            .scan_select_out (scan [15]),
            .latch_enable_out(latch[15])
            );
        
        // https://github.com/jglim/tinytapeout_bcd-7seg
        scan_wrapper_341152580068442706 #(.NUM_IOS(8)) scan_wrapper_341152580068442706_15 (
            .clk_in          (clk  [15]),
            .data_in         (data [15]),
            .scan_select_in  (scan [15]),
            .latch_enable_in (latch[15]),
            .clk_out         (clk  [16]),
            .data_out        (data [16]),
            .scan_select_out (scan [16]),
            .latch_enable_out(latch[16])
            );
        
        // https://github.com/tkuester/wokwi-directghost
        scan_wrapper_341155178824598098 #(.NUM_IOS(8)) scan_wrapper_341155178824598098_16 (
            .clk_in          (clk  [16]),
            .data_in         (data [16]),
            .scan_select_in  (scan [16]),
            .latch_enable_in (latch[16]),
            .clk_out         (clk  [17]),
            .data_out        (data [17]),
            .scan_select_out (scan [17]),
            .latch_enable_out(latch[17])
            );
        
        // https://github.com/shahzaibk23/tinytapeout-barrel-shifter
        scan_wrapper_341167691532337747 #(.NUM_IOS(8)) scan_wrapper_341167691532337747_17 (
            .clk_in          (clk  [17]),
            .data_in         (data [17]),
            .scan_select_in  (scan [17]),
            .latch_enable_in (latch[17]),
            .clk_out         (clk  [18]),
            .data_out        (data [18]),
            .scan_select_out (scan [18]),
            .latch_enable_out(latch[18])
            );
        
        // https://github.com/tcptomato/tinytapeout
        scan_wrapper_341178154799333971 #(.NUM_IOS(8)) scan_wrapper_341178154799333971_18 (
            .clk_in          (clk  [18]),
            .data_in         (data [18]),
            .scan_select_in  (scan [18]),
            .latch_enable_in (latch[18]),
            .clk_out         (clk  [19]),
            .data_out        (data [19]),
            .scan_select_out (scan [19]),
            .latch_enable_out(latch[19])
            );
        
        // https://github.com/DaveyPocket/chaser
        scan_wrapper_341178481588044372 #(.NUM_IOS(8)) scan_wrapper_341178481588044372_19 (
            .clk_in          (clk  [19]),
            .data_in         (data [19]),
            .scan_select_in  (scan [19]),
            .latch_enable_in (latch[19]),
            .clk_out         (clk  [20]),
            .data_out        (data [20]),
            .scan_select_out (scan [20]),
            .latch_enable_out(latch[20])
            );
        
        // https://github.com/GuzTech/tinytapeout-4x4-multiplier
        scan_wrapper_341176884318437971 #(.NUM_IOS(8)) scan_wrapper_341176884318437971_20 (
            .clk_in          (clk  [20]),
            .data_in         (data [20]),
            .scan_select_in  (scan [20]),
            .latch_enable_in (latch[20]),
            .clk_out         (clk  [21]),
            .data_out        (data [21]),
            .scan_select_out (scan [21]),
            .latch_enable_out(latch[21])
            );
        
        // https://github.com/derhexenmeister/tinytapeout_nco
        scan_wrapper_341182944314917460 #(.NUM_IOS(8)) scan_wrapper_341182944314917460_21 (
            .clk_in          (clk  [21]),
            .data_in         (data [21]),
            .scan_select_in  (scan [21]),
            .latch_enable_in (latch[21]),
            .clk_out         (clk  [22]),
            .data_out        (data [22]),
            .scan_select_out (scan [22]),
            .latch_enable_out(latch[22])
            );
        
        // https://github.com/mbalestrini/tinytapeout_rgb_lut_test
        scan_wrapper_341188777753969234 #(.NUM_IOS(8)) scan_wrapper_341188777753969234_22 (
            .clk_in          (clk  [22]),
            .data_in         (data [22]),
            .scan_select_in  (scan [22]),
            .latch_enable_in (latch[22]),
            .clk_out         (clk  [23]),
            .data_out        (data [23]),
            .scan_select_out (scan [23]),
            .latch_enable_out(latch[23])
            );
        
        // https://github.com/derhexenmeister/tinytapeout_updwnbcd
        scan_wrapper_341194143598379604 #(.NUM_IOS(8)) scan_wrapper_341194143598379604_23 (
            .clk_in          (clk  [23]),
            .data_in         (data [23]),
            .scan_select_in  (scan [23]),
            .latch_enable_in (latch[23]),
            .clk_out         (clk  [24]),
            .data_out        (data [24]),
            .scan_select_out (scan [24]),
            .latch_enable_out(latch[24])
            );
        
        // https://github.com/bradysalz/pll_tiny_tapeout_demo
        scan_wrapper_341205508016833108 #(.NUM_IOS(8)) scan_wrapper_341205508016833108_24 (
            .clk_in          (clk  [24]),
            .data_in         (data [24]),
            .scan_select_in  (scan [24]),
            .latch_enable_in (latch[24]),
            .clk_out         (clk  [25]),
            .data_out        (data [25]),
            .scan_select_out (scan [25]),
            .latch_enable_out(latch[25])
            );
        
        // https://github.com/pramitpal/tinytapeout_pramit
        scan_wrapper_341162950004834900 #(.NUM_IOS(8)) scan_wrapper_341162950004834900_25 (
            .clk_in          (clk  [25]),
            .data_in         (data [25]),
            .scan_select_in  (scan [25]),
            .latch_enable_in (latch[25]),
            .clk_out         (clk  [26]),
            .data_out        (data [26]),
            .scan_select_out (scan [26]),
            .latch_enable_out(latch[26])
            );
        
        // https://github.com/gregdavill/tinytapeout-verilog-fifo
        scan_wrapper_341202178192441940 #(.NUM_IOS(8)) scan_wrapper_341202178192441940_26 (
            .clk_in          (clk  [26]),
            .data_in         (data [26]),
            .scan_select_in  (scan [26]),
            .latch_enable_in (latch[26]),
            .clk_out         (clk  [27]),
            .data_out        (data [27]),
            .scan_select_out (scan [27]),
            .latch_enable_out(latch[27])
            );
        
        // https://github.com/gregdavill/tinytapeout-wokwi-74x1G00
        scan_wrapper_341191836498395731 #(.NUM_IOS(8)) scan_wrapper_341191836498395731_27 (
            .clk_in          (clk  [27]),
            .data_in         (data [27]),
            .scan_select_in  (scan [27]),
            .latch_enable_in (latch[27]),
            .clk_out         (clk  [28]),
            .data_out        (data [28]),
            .scan_select_out (scan [28]),
            .latch_enable_out(latch[28])
            );
        
        // https://github.com/gregdavill/tinytapeout-wokwi-74x1G02
        scan_wrapper_341192113929585235 #(.NUM_IOS(8)) scan_wrapper_341192113929585235_28 (
            .clk_in          (clk  [28]),
            .data_in         (data [28]),
            .scan_select_in  (scan [28]),
            .latch_enable_in (latch[28]),
            .clk_out         (clk  [29]),
            .data_out        (data [29]),
            .scan_select_out (scan [29]),
            .latch_enable_out(latch[29])
            );
        
        // https://github.com/gregdavill/tinytapeout-wokwi-74xG198
        scan_wrapper_341192621088047698 #(.NUM_IOS(8)) scan_wrapper_341192621088047698_29 (
            .clk_in          (clk  [29]),
            .data_in         (data [29]),
            .scan_select_in  (scan [29]),
            .latch_enable_in (latch[29]),
            .clk_out         (clk  [30]),
            .data_out        (data [30]),
            .scan_select_out (scan [30]),
            .latch_enable_out(latch[30])
            );
        
        // https://github.com/gregdavill/tinytapeout-verilog-7seg-clock
        scan_wrapper_340579111348994642 #(.NUM_IOS(8)) scan_wrapper_340579111348994642_30 (
            .clk_in          (clk  [30]),
            .data_in         (data [30]),
            .scan_select_in  (scan [30]),
            .latch_enable_in (latch[30]),
            .clk_out         (clk  [31]),
            .data_out        (data [31]),
            .scan_select_out (scan [31]),
            .latch_enable_out(latch[31])
            );
        
        // https://github.com/alanvgreen/tinytapeout4bitadder
        scan_wrapper_341224613878956628 #(.NUM_IOS(8)) scan_wrapper_341224613878956628_31 (
            .clk_in          (clk  [31]),
            .data_in         (data [31]),
            .scan_select_in  (scan [31]),
            .latch_enable_in (latch[31]),
            .clk_out         (clk  [32]),
            .data_out        (data [32]),
            .scan_select_out (scan [32]),
            .latch_enable_out(latch[32])
            );
        
        // https://github.com/benlaurie/twistedringcounter
        scan_wrapper_341235973870322258 #(.NUM_IOS(8)) scan_wrapper_341235973870322258_32 (
            .clk_in          (clk  [32]),
            .data_in         (data [32]),
            .scan_select_in  (scan [32]),
            .latch_enable_in (latch[32]),
            .clk_out         (clk  [33]),
            .data_out        (data [33]),
            .scan_select_out (scan [33]),
            .latch_enable_out(latch[33])
            );
        
        // https://github.com/sureshsugumar/tinytapeout_counter
        scan_wrapper_341235575572922964 #(.NUM_IOS(8)) scan_wrapper_341235575572922964_33 (
            .clk_in          (clk  [33]),
            .data_in         (data [33]),
            .scan_select_in  (scan [33]),
            .latch_enable_in (latch[33]),
            .clk_out         (clk  [34]),
            .data_out        (data [34]),
            .scan_select_out (scan [34]),
            .latch_enable_out(latch[34])
            );
        
        // https://github.com/daniestevez/tinytapeout-verilog
        scan_wrapper_341164910646919762 #(.NUM_IOS(8)) scan_wrapper_341164910646919762_34 (
            .clk_in          (clk  [34]),
            .data_in         (data [34]),
            .scan_select_in  (scan [34]),
            .latch_enable_in (latch[34]),
            .clk_out         (clk  [35]),
            .data_out        (data [35]),
            .scan_select_out (scan [35]),
            .latch_enable_out(latch[35])
            );
        
        // https://github.com/pkuligowski/tinytapeout_tmr
        scan_wrapper_341233739099013714 #(.NUM_IOS(8)) scan_wrapper_341233739099013714_35 (
            .clk_in          (clk  [35]),
            .data_in         (data [35]),
            .scan_select_in  (scan [35]),
            .latch_enable_in (latch[35]),
            .clk_out         (clk  [36]),
            .data_out        (data [36]),
            .scan_select_out (scan [36]),
            .latch_enable_out(latch[36])
            );
        
        // https://github.com/chiplet/tinytapeout-snake
        scan_wrapper_341240110454407762 #(.NUM_IOS(8)) scan_wrapper_341240110454407762_36 (
            .clk_in          (clk  [36]),
            .data_in         (data [36]),
            .scan_select_in  (scan [36]),
            .latch_enable_in (latch[36]),
            .clk_out         (clk  [37]),
            .data_out        (data [37]),
            .scan_select_out (scan [37]),
            .latch_enable_out(latch[37])
            );
        
        // https://github.com/derhexenmeister/tinytapeout_pwm
        scan_wrapper_341264068701586004 #(.NUM_IOS(8)) scan_wrapper_341264068701586004_37 (
            .clk_in          (clk  [37]),
            .data_in         (data [37]),
            .scan_select_in  (scan [37]),
            .latch_enable_in (latch[37]),
            .clk_out         (clk  [38]),
            .data_out        (data [38]),
            .scan_select_out (scan [38]),
            .latch_enable_out(latch[38])
            );
        
        // https://github.com/raha96/tinycharacters-locked
        scan_wrapper_341164228775772755 #(.NUM_IOS(8)) scan_wrapper_341164228775772755_38 (
            .clk_in          (clk  [38]),
            .data_in         (data [38]),
            .scan_select_in  (scan [38]),
            .latch_enable_in (latch[38]),
            .clk_out         (clk  [39]),
            .data_out        (data [39]),
            .scan_select_out (scan [39]),
            .latch_enable_out(latch[39])
            );
        
        // https://github.com/nathancheek/tinytapeout-loop
        scan_wrapper_341262321634509394 #(.NUM_IOS(8)) scan_wrapper_341262321634509394_39 (
            .clk_in          (clk  [39]),
            .data_in         (data [39]),
            .scan_select_in  (scan [39]),
            .latch_enable_in (latch[39]),
            .clk_out         (clk  [40]),
            .data_out        (data [40]),
            .scan_select_out (scan [40]),
            .latch_enable_out(latch[40])
            );
        
        // https://github.com/andars/universal-turing-machine-w5s8
        scan_wrapper_341174563322724948 #(.NUM_IOS(8)) scan_wrapper_341174563322724948_40 (
            .clk_in          (clk  [40]),
            .data_in         (data [40]),
            .scan_select_in  (scan [40]),
            .latch_enable_in (latch[40]),
            .clk_out         (clk  [41]),
            .data_out        (data [41]),
            .scan_select_out (scan [41]),
            .latch_enable_out(latch[41])
            );
        
        // https://github.com/vmunoz82/tinytapeout_euler1
        scan_wrapper_341271902949474898 #(.NUM_IOS(8)) scan_wrapper_341271902949474898_41 (
            .clk_in          (clk  [41]),
            .data_in         (data [41]),
            .scan_select_in  (scan [41]),
            .latch_enable_in (latch[41]),
            .clk_out         (clk  [42]),
            .data_out        (data [42]),
            .scan_select_out (scan [42]),
            .latch_enable_out(latch[42])
            );
        
        // https://github.com/mikenet213/mikenet213-tt1-verilog
        scan_wrapper_bc4d7220e4fdbf20a574d56ea112a8e1 #(.NUM_IOS(8)) scan_wrapper_bc4d7220e4fdbf20a574d56ea112a8e1_42 (
            .clk_in          (clk  [42]),
            .data_in         (data [42]),
            .scan_select_in  (scan [42]),
            .latch_enable_in (latch[42]),
            .clk_out         (clk  [43]),
            .data_out        (data [43]),
            .scan_select_out (scan [43]),
            .latch_enable_out(latch[43])
            );
        
        // https://github.com/veremenko-y/tinytapeout-ue14500
        scan_wrapper_341178296293130834 #(.NUM_IOS(8)) scan_wrapper_341178296293130834_43 (
            .clk_in          (clk  [43]),
            .data_in         (data [43]),
            .scan_select_in  (scan [43]),
            .latch_enable_in (latch[43]),
            .clk_out         (clk  [44]),
            .data_out        (data [44]),
            .scan_select_out (scan [44]),
            .latch_enable_out(latch[44])
            );
        
        // https://github.com/mikenet213/mikenet213-tt2-verilog
        scan_wrapper_1f985e14df1ed789231bb6e0189d6e39 #(.NUM_IOS(8)) scan_wrapper_1f985e14df1ed789231bb6e0189d6e39_44 (
            .clk_in          (clk  [44]),
            .data_in         (data [44]),
            .scan_select_in  (scan [44]),
            .latch_enable_in (latch[44]),
            .clk_out         (clk  [45]),
            .data_out        (data [45]),
            .scan_select_out (scan [45]),
            .latch_enable_out(latch[45])
            );
        
        // https://github.com/aiunderstand/tinytapeout_asyncbinterconvcomp.git
        scan_wrapper_341277789473735250 #(.NUM_IOS(8)) scan_wrapper_341277789473735250_45 (
            .clk_in          (clk  [45]),
            .data_in         (data [45]),
            .scan_select_in  (scan [45]),
            .latch_enable_in (latch[45]),
            .clk_out         (clk  [46]),
            .data_out        (data [46]),
            .scan_select_out (scan [46]),
            .latch_enable_out(latch[46])
            );
        
        // https://github.com/smunaut/tinytapeout-fifo
        scan_wrapper_341263346544149074 #(.NUM_IOS(8)) scan_wrapper_341263346544149074_46 (
            .clk_in          (clk  [46]),
            .data_in         (data [46]),
            .scan_select_in  (scan [46]),
            .latch_enable_in (latch[46]),
            .clk_out         (clk  [47]),
            .data_out        (data [47]),
            .scan_select_out (scan [47]),
            .latch_enable_out(latch[47])
            );
        
        // https://github.com/nwtechguy/tinytapeout_BCD_counter
        scan_wrapper_341296149788885588 #(.NUM_IOS(8)) scan_wrapper_341296149788885588_47 (
            .clk_in          (clk  [47]),
            .data_in         (data [47]),
            .scan_select_in  (scan [47]),
            .latch_enable_in (latch[47]),
            .clk_out         (clk  [48]),
            .data_out        (data [48]),
            .scan_select_out (scan [48]),
            .latch_enable_out(latch[48])
            );
        
        // https://github.com/kambadur/bcd_to_7seg
        scan_wrapper_341332847867462227 #(.NUM_IOS(8)) scan_wrapper_341332847867462227_48 (
            .clk_in          (clk  [48]),
            .data_in         (data [48]),
            .scan_select_in  (scan [48]),
            .latch_enable_in (latch[48]),
            .clk_out         (clk  [49]),
            .data_out        (data [49]),
            .scan_select_out (scan [49]),
            .latch_enable_out(latch[49])
            );
        
        // https://github.com/bieganski/tinytapeout_bieganski
        scan_wrapper_341337976625693266 #(.NUM_IOS(8)) scan_wrapper_341337976625693266_49 (
            .clk_in          (clk  [49]),
            .data_in         (data [49]),
            .scan_select_in  (scan [49]),
            .latch_enable_in (latch[49]),
            .clk_out         (clk  [50]),
            .data_out        (data [50]),
            .scan_select_out (scan [50]),
            .latch_enable_out(latch[50])
            );
        
        // https://github.com/TomKeddie/tinytapeout-2022-1
        scan_wrapper_341339883600609876 #(.NUM_IOS(8)) scan_wrapper_341339883600609876_50 (
            .clk_in          (clk  [50]),
            .data_in         (data [50]),
            .scan_select_in  (scan [50]),
            .latch_enable_in (latch[50]),
            .clk_out         (clk  [51]),
            .data_out        (data [51]),
            .scan_select_out (scan [51]),
            .latch_enable_out(latch[51])
            );
        
        // https://github.com/r-a-hoggarth/tinytapeGaloisLFSR
        scan_wrapper_341344337258349139 #(.NUM_IOS(8)) scan_wrapper_341344337258349139_51 (
            .clk_in          (clk  [51]),
            .data_in         (data [51]),
            .scan_select_in  (scan [51]),
            .latch_enable_in (latch[51]),
            .clk_out         (clk  [52]),
            .data_out        (data [52]),
            .scan_select_out (scan [52]),
            .latch_enable_out(latch[52])
            );
        
        // https://github.com/adamgreig/tinytapeout-prn
        scan_wrapper_341342096033055316 #(.NUM_IOS(8)) scan_wrapper_341342096033055316_52 (
            .clk_in          (clk  [52]),
            .data_in         (data [52]),
            .scan_select_in  (scan [52]),
            .latch_enable_in (latch[52]),
            .clk_out         (clk  [53]),
            .data_out        (data [53]),
            .scan_select_out (scan [53]),
            .latch_enable_out(latch[53])
            );
        
        // https://github.com/ianloic/tinytapeout-1
        scan_wrapper_341259651269001812 #(.NUM_IOS(8)) scan_wrapper_341259651269001812_53 (
            .clk_in          (clk  [53]),
            .data_in         (data [53]),
            .scan_select_in  (scan [53]),
            .latch_enable_in (latch[53]),
            .clk_out         (clk  [54]),
            .data_out        (data [54]),
            .scan_select_out (scan [54]),
            .latch_enable_out(latch[54])
            );
        
        // https://github.com/sad-electronics/tinytapeout-clock-divider-asic
        scan_wrapper_341353928049295956 #(.NUM_IOS(8)) scan_wrapper_341353928049295956_54 (
            .clk_in          (clk  [54]),
            .data_in         (data [54]),
            .scan_select_in  (scan [54]),
            .latch_enable_in (latch[54]),
            .clk_out         (clk  [55]),
            .data_out        (data [55]),
            .scan_select_out (scan [55]),
            .latch_enable_out(latch[55])
            );
        
        // https://github.com/gatecat/tinytapeout-lutram-test
        scan_wrapper_341353780122485332 #(.NUM_IOS(8)) scan_wrapper_341353780122485332_55 (
            .clk_in          (clk  [55]),
            .data_in         (data [55]),
            .scan_select_in  (scan [55]),
            .latch_enable_in (latch[55]),
            .clk_out         (clk  [56]),
            .data_out        (data [56]),
            .scan_select_out (scan [56]),
            .latch_enable_out(latch[56])
            );
        
        // https://github.com/tommythorn/tinytapeout-4-bit-cpu
        scan_wrapper_341193419111006803 #(.NUM_IOS(8)) scan_wrapper_341193419111006803_56 (
            .clk_in          (clk  [56]),
            .data_in         (data [56]),
            .scan_select_in  (scan [56]),
            .latch_enable_in (latch[56]),
            .clk_out         (clk  [57]),
            .data_out        (data [57]),
            .scan_select_out (scan [57]),
            .latch_enable_out(latch[57])
            );
        
        // https://github.com/wokwi/tt-game-of-life-cell-popcnt
        scan_wrapper_341266732010177108 #(.NUM_IOS(8)) scan_wrapper_341266732010177108_57 (
            .clk_in          (clk  [57]),
            .data_in         (data [57]),
            .scan_select_in  (scan [57]),
            .latch_enable_in (latch[57]),
            .clk_out         (clk  [58]),
            .data_out        (data [58]),
            .scan_select_out (scan [58]),
            .latch_enable_out(latch[58])
            );
        
        // https://github.com/gatecat/tinytapeout-srlut-test
        scan_wrapper_341353777861755476 #(.NUM_IOS(8)) scan_wrapper_341353777861755476_58 (
            .clk_in          (clk  [58]),
            .data_in         (data [58]),
            .scan_select_in  (scan [58]),
            .latch_enable_in (latch[58]),
            .clk_out         (clk  [59]),
            .data_out        (data [59]),
            .scan_select_out (scan [59]),
            .latch_enable_out(latch[59])
            );
        
        // https://github.com/AdDraw/tinytapeout_demo
        scan_wrapper_341359404107432531 #(.NUM_IOS(8)) scan_wrapper_341359404107432531_59 (
            .clk_in          (clk  [59]),
            .data_in         (data [59]),
            .scan_select_in  (scan [59]),
            .latch_enable_in (latch[59]),
            .clk_out         (clk  [60]),
            .data_out        (data [60]),
            .scan_select_out (scan [60]),
            .latch_enable_out(latch[60])
            );
        
        // https://github.com/cpldcpu/tinydice
        scan_wrapper_341315210433266259 #(.NUM_IOS(8)) scan_wrapper_341315210433266259_60 (
            .clk_in          (clk  [60]),
            .data_in         (data [60]),
            .scan_select_in  (scan [60]),
            .latch_enable_in (latch[60]),
            .clk_out         (clk  [61]),
            .data_out        (data [61]),
            .scan_select_out (scan [61]),
            .latch_enable_out(latch[61])
            );
        
        // https://github.com/cpldcpu/tinytapeout_mcpu6bit
        scan_wrapper_341364381657858642 #(.NUM_IOS(8)) scan_wrapper_341364381657858642_61 (
            .clk_in          (clk  [61]),
            .data_in         (data [61]),
            .scan_select_in  (scan [61]),
            .latch_enable_in (latch[61]),
            .clk_out         (clk  [62]),
            .data_out        (data [62]),
            .scan_select_out (scan [62]),
            .latch_enable_out(latch[62])
            );
        
        // https://github.com/azzeloof/tinytapeout-counter
        scan_wrapper_341279123277087315 #(.NUM_IOS(8)) scan_wrapper_341279123277087315_62 (
            .clk_in          (clk  [62]),
            .data_in         (data [62]),
            .scan_select_in  (scan [62]),
            .latch_enable_in (latch[62]),
            .clk_out         (clk  [63]),
            .data_out        (data [63]),
            .scan_select_out (scan [63]),
            .latch_enable_out(latch[63])
            );
        
        // https://github.com/mattvenn/tinytapeout-341802655228625490
        scan_wrapper_341802655228625490 #(.NUM_IOS(8)) scan_wrapper_341802655228625490_63 (
            .clk_in          (clk  [63]),
            .data_in         (data [63]),
            .scan_select_in  (scan [63]),
            .latch_enable_in (latch[63]),
            .clk_out         (clk  [64]),
            .data_out        (data [64]),
            .scan_select_out (scan [64]),
            .latch_enable_out(latch[64])
            );
        
        // https://github.com/mwelling/led-blaster
        scan_wrapper_341382703379120723 #(.NUM_IOS(8)) scan_wrapper_341382703379120723_64 (
            .clk_in          (clk  [64]),
            .data_in         (data [64]),
            .scan_select_in  (scan [64]),
            .latch_enable_in (latch[64]),
            .clk_out         (clk  [65]),
            .data_out        (data [65]),
            .scan_select_out (scan [65]),
            .latch_enable_out(latch[65])
            );
        
        // https://github.com/mwelling/figure-8
        scan_wrapper_341389786199622227 #(.NUM_IOS(8)) scan_wrapper_341389786199622227_65 (
            .clk_in          (clk  [65]),
            .data_in         (data [65]),
            .scan_select_in  (scan [65]),
            .latch_enable_in (latch[65]),
            .clk_out         (clk  [66]),
            .data_out        (data [66]),
            .scan_select_out (scan [66]),
            .latch_enable_out(latch[66])
            );
        
        // https://github.com/gatecat/tinytapeout-fpga-test
        scan_wrapper_341404507891040852 #(.NUM_IOS(8)) scan_wrapper_341404507891040852_66 (
            .clk_in          (clk  [66]),
            .data_in         (data [66]),
            .scan_select_in  (scan [66]),
            .latch_enable_in (latch[66]),
            .clk_out         (clk  [67]),
            .data_out        (data [67]),
            .scan_select_out (scan [67]),
            .latch_enable_out(latch[67])
            );
        
        // https://github.com/cfib/trafficlight-fsm
        scan_wrapper_341410909669818963 #(.NUM_IOS(8)) scan_wrapper_341410909669818963_67 (
            .clk_in          (clk  [67]),
            .data_in         (data [67]),
            .scan_select_in  (scan [67]),
            .latch_enable_in (latch[67]),
            .clk_out         (clk  [68]),
            .data_out        (data [68]),
            .scan_select_out (scan [68]),
            .latch_enable_out(latch[68])
            );
        
        // https://github.com/clj/tinytapeout-verilog-7seg-figure-eight
        scan_wrapper_341063825089364563 #(.NUM_IOS(8)) scan_wrapper_341063825089364563_68 (
            .clk_in          (clk  [68]),
            .data_in         (data [68]),
            .scan_select_in  (scan [68]),
            .latch_enable_in (latch[68]),
            .clk_out         (clk  [69]),
            .data_out        (data [69]),
            .scan_select_out (scan [69]),
            .latch_enable_out(latch[69])
            );
        
        // https://github.com/smunaut/tinytapeout-misc-1
        scan_wrapper_341174480471589458 #(.NUM_IOS(8)) scan_wrapper_341174480471589458_69 (
            .clk_in          (clk  [69]),
            .data_in         (data [69]),
            .scan_select_in  (scan [69]),
            .latch_enable_in (latch[69]),
            .clk_out         (clk  [70]),
            .data_out        (data [70]),
            .scan_select_out (scan [70]),
            .latch_enable_out(latch[70])
            );
        
        // https://github.com/regymm/tinytapeout-funnyblinky
        scan_wrapper_341419328215712339 #(.NUM_IOS(8)) scan_wrapper_341419328215712339_70 (
            .clk_in          (clk  [70]),
            .data_in         (data [70]),
            .scan_select_in  (scan [70]),
            .latch_enable_in (latch[70]),
            .clk_out         (clk  [71]),
            .data_out        (data [71]),
            .scan_select_out (scan [71]),
            .latch_enable_out(latch[71])
            );
        
        // https://github.com/Sirawit7205/tinytapeout-2G57-2G58
        scan_wrapper_341431339142087251 #(.NUM_IOS(8)) scan_wrapper_341431339142087251_71 (
            .clk_in          (clk  [71]),
            .data_in         (data [71]),
            .scan_select_in  (scan [71]),
            .latch_enable_in (latch[71]),
            .clk_out         (clk  [72]),
            .data_out        (data [72]),
            .scan_select_out (scan [72]),
            .latch_enable_out(latch[72])
            );
        
        // https://github.com/Sirawit7205/tinytapeout-2G97-2G98
        scan_wrapper_341432030163108435 #(.NUM_IOS(8)) scan_wrapper_341432030163108435_72 (
            .clk_in          (clk  [72]),
            .data_in         (data [72]),
            .scan_select_in  (scan [72]),
            .latch_enable_in (latch[72]),
            .clk_out         (clk  [73]),
            .data_out        (data [73]),
            .scan_select_out (scan [73]),
            .latch_enable_out(latch[73])
            );
        
        // https://github.com/hosein-mokarian/tinytapeout_counter_3to8_decoder
        scan_wrapper_341440114308678227 #(.NUM_IOS(8)) scan_wrapper_341440114308678227_73 (
            .clk_in          (clk  [73]),
            .data_in         (data [73]),
            .scan_select_in  (scan [73]),
            .latch_enable_in (latch[73]),
            .clk_out         (clk  [74]),
            .data_out        (data [74]),
            .scan_select_out (scan [74]),
            .latch_enable_out(latch[74])
            );
        
        // https://github.com/burtyb/srld
        scan_wrapper_341496918381167187 #(.NUM_IOS(8)) scan_wrapper_341496918381167187_74 (
            .clk_in          (clk  [74]),
            .data_in         (data [74]),
            .scan_select_in  (scan [74]),
            .latch_enable_in (latch[74]),
            .clk_out         (clk  [75]),
            .data_out        (data [75]),
            .scan_select_out (scan [75]),
            .latch_enable_out(latch[75])
            );
        
        // https://github.com/Mahnoor-ismail01/tinytapeout-chromatic-3-to-8-Decoder
        scan_wrapper_341440781874102868 #(.NUM_IOS(8)) scan_wrapper_341440781874102868_75 (
            .clk_in          (clk  [75]),
            .data_in         (data [75]),
            .scan_select_in  (scan [75]),
            .latch_enable_in (latch[75]),
            .clk_out         (clk  [76]),
            .data_out        (data [76]),
            .scan_select_out (scan [76]),
            .latch_enable_out(latch[76])
            );
        
        // https://github.com/Shahzaib2028/tinytapeout-4to2Encoder-2to4Decoder
        scan_wrapper_341444501414347346 #(.NUM_IOS(8)) scan_wrapper_341444501414347346_76 (
            .clk_in          (clk  [76]),
            .data_in         (data [76]),
            .scan_select_in  (scan [76]),
            .latch_enable_in (latch[76]),
            .clk_out         (clk  [77]),
            .data_out        (data [77]),
            .scan_select_out (scan [77]),
            .latch_enable_out(latch[77])
            );
        
        // https://github.com/sfmth/tinytapeout-tinycordic
        scan_wrapper_019235602376235615 #(.NUM_IOS(8)) scan_wrapper_019235602376235615_77 (
            .clk_in          (clk  [77]),
            .data_in         (data [77]),
            .scan_select_in  (scan [77]),
            .latch_enable_in (latch[77]),
            .clk_out         (clk  [78]),
            .data_out        (data [78]),
            .scan_select_out (scan [78]),
            .latch_enable_out(latch[78])
            );
        
        // https://github.com/mm21/tinytapeout-led-matrix
        scan_wrapper_341450853309219412 #(.NUM_IOS(8)) scan_wrapper_341450853309219412_78 (
            .clk_in          (clk  [78]),
            .data_in         (data [78]),
            .scan_select_in  (scan [78]),
            .latch_enable_in (latch[78]),
            .clk_out         (clk  [79]),
            .data_out        (data [79]),
            .scan_select_out (scan [79]),
            .latch_enable_out(latch[79])
            );
        
        // https://github.com/jeanthom/tinytapout-lock
        scan_wrapper_341438392303616596 #(.NUM_IOS(8)) scan_wrapper_341438392303616596_79 (
            .clk_in          (clk  [79]),
            .data_in         (data [79]),
            .scan_select_in  (scan [79]),
            .latch_enable_in (latch[79]),
            .clk_out         (clk  [80]),
            .data_out        (data [80]),
            .scan_select_out (scan [80]),
            .latch_enable_out(latch[80])
            );
        
        // https://github.com/AidanMedcalf/tinytapeout-tinyio
        scan_wrapper_341432284947153491 #(.NUM_IOS(8)) scan_wrapper_341432284947153491_80 (
            .clk_in          (clk  [80]),
            .data_in         (data [80]),
            .scan_select_in  (scan [80]),
            .latch_enable_in (latch[80]),
            .clk_out         (clk  [81]),
            .data_out        (data [81]),
            .scan_select_out (scan [81]),
            .latch_enable_out(latch[81])
            );
        
        // https://github.com/ElectricPotato/tinytapeout-hello-world-uart
        scan_wrapper_341457971277988435 #(.NUM_IOS(8)) scan_wrapper_341457971277988435_81 (
            .clk_in          (clk  [81]),
            .data_in         (data [81]),
            .scan_select_in  (scan [81]),
            .latch_enable_in (latch[81]),
            .clk_out         (clk  [82]),
            .data_out        (data [82]),
            .scan_select_out (scan [82]),
            .latch_enable_out(latch[82])
            );
        
        // https://github.com/abdullahkhalids/TinyTapeout-hamming-code
        scan_wrapper_341399568412312147 #(.NUM_IOS(8)) scan_wrapper_341399568412312147_82 (
            .clk_in          (clk  [82]),
            .data_in         (data [82]),
            .scan_select_in  (scan [82]),
            .latch_enable_in (latch[82]),
            .clk_out         (clk  [83]),
            .data_out        (data [83]),
            .scan_select_out (scan [83]),
            .latch_enable_out(latch[83])
            );
        
        // https://github.com/hossein1387/tinytapeout-verilog-test
        scan_wrapper_341464767397888596 #(.NUM_IOS(8)) scan_wrapper_341464767397888596_83 (
            .clk_in          (clk  [83]),
            .data_in         (data [83]),
            .scan_select_in  (scan [83]),
            .latch_enable_in (latch[83]),
            .clk_out         (clk  [84]),
            .data_out        (data [84]),
            .scan_select_out (scan [84]),
            .latch_enable_out(latch[84])
            );
        
        // https://github.com/ChrisPVille/tinytapeout-FROG4bitCPU
        scan_wrapper_341476989274686036 #(.NUM_IOS(8)) scan_wrapper_341476989274686036_84 (
            .clk_in          (clk  [84]),
            .data_in         (data [84]),
            .scan_select_in  (scan [84]),
            .latch_enable_in (latch[84]),
            .clk_out         (clk  [85]),
            .data_out        (data [85]),
            .scan_select_out (scan [85]),
            .latch_enable_out(latch[85])
            );
        
        // https://github.com/Talha-Ahmed-1/tinytapeout_flop_regfile
        scan_wrapper_341482086419399252 #(.NUM_IOS(8)) scan_wrapper_341482086419399252_85 (
            .clk_in          (clk  [85]),
            .data_in         (data [85]),
            .scan_select_in  (scan [85]),
            .latch_enable_in (latch[85]),
            .clk_out         (clk  [86]),
            .data_out        (data [86]),
            .scan_select_out (scan [86]),
            .latch_enable_out(latch[86])
            );
        
        // https://github.com/skylersaleh/tinytapeout-hello
        scan_wrapper_341452019534398035 #(.NUM_IOS(8)) scan_wrapper_341452019534398035_86 (
            .clk_in          (clk  [86]),
            .data_in         (data [86]),
            .scan_select_in  (scan [86]),
            .latch_enable_in (latch[86]),
            .clk_out         (clk  [87]),
            .data_out        (data [87]),
            .scan_select_out (scan [87]),
            .latch_enable_out(latch[87])
            );
        
        // https://github.com/proppy/tinytapeout-xls-popcount
        scan_wrapper_341497971083313748 #(.NUM_IOS(8)) scan_wrapper_341497971083313748_87 (
            .clk_in          (clk  [87]),
            .data_in         (data [87]),
            .scan_select_in  (scan [87]),
            .latch_enable_in (latch[87]),
            .clk_out         (clk  [88]),
            .data_out        (data [88]),
            .scan_select_out (scan [88]),
            .latch_enable_out(latch[88])
            );
        
        // https://github.com/proppy/tinytapeout-xls-popcount-bithacks
        scan_wrapper_341497964482527828 #(.NUM_IOS(8)) scan_wrapper_341497964482527828_88 (
            .clk_in          (clk  [88]),
            .data_in         (data [88]),
            .scan_select_in  (scan [88]),
            .latch_enable_in (latch[88]),
            .clk_out         (clk  [89]),
            .data_out        (data [89]),
            .scan_select_out (scan [89]),
            .latch_enable_out(latch[89])
            );
        
        // https://github.com/proppy/tinytapeout-xls-inverter
        scan_wrapper_341497938559631956 #(.NUM_IOS(8)) scan_wrapper_341497938559631956_89 (
            .clk_in          (clk  [89]),
            .data_in         (data [89]),
            .scan_select_in  (scan [89]),
            .latch_enable_in (latch[89]),
            .clk_out         (clk  [90]),
            .data_out        (data [90]),
            .scan_select_out (scan [90]),
            .latch_enable_out(latch[90])
            );
        
        // https://github.com/mark64/tinytapeout
        scan_wrapper_341499976001520211 #(.NUM_IOS(8)) scan_wrapper_341499976001520211_90 (
            .clk_in          (clk  [90]),
            .data_in         (data [90]),
            .scan_select_in  (scan [90]),
            .latch_enable_in (latch[90]),
            .clk_out         (clk  [91]),
            .data_out        (data [91]),
            .scan_select_out (scan [91]),
            .latch_enable_out(latch[91])
            );
        
        // https://github.com/dave-roo/ddcomparatorandro
        scan_wrapper_341500800901579348 #(.NUM_IOS(8)) scan_wrapper_341500800901579348_91 (
            .clk_in          (clk  [91]),
            .data_in         (data [91]),
            .scan_select_in  (scan [91]),
            .latch_enable_in (latch[91]),
            .clk_out         (clk  [92]),
            .data_out        (data [92]),
            .scan_select_out (scan [92]),
            .latch_enable_out(latch[92])
            );
        
        // https://github.com/splinedrive/tinytapeout-verilog-4x4-multiplier
        scan_wrapper_341493393195532884 #(.NUM_IOS(8)) scan_wrapper_341493393195532884_92 (
            .clk_in          (clk  [92]),
            .data_in         (data [92]),
            .scan_select_in  (scan [92]),
            .latch_enable_in (latch[92]),
            .clk_out         (clk  [93]),
            .data_out        (data [93]),
            .scan_select_out (scan [93]),
            .latch_enable_out(latch[93])
            );
        
        // https://github.com/ThorKn/tinytapeout_shiftregister_8bit
        scan_wrapper_341506274933867090 #(.NUM_IOS(8)) scan_wrapper_341506274933867090_93 (
            .clk_in          (clk  [93]),
            .data_in         (data [93]),
            .scan_select_in  (scan [93]),
            .latch_enable_in (latch[93]),
            .clk_out         (clk  [94]),
            .data_out        (data [94]),
            .scan_select_out (scan [94]),
            .latch_enable_out(latch[94])
            );
        
        // https://github.com/UDXS/tinytapeout-sqrt
        scan_wrapper_341449297858921043 #(.NUM_IOS(8)) scan_wrapper_341449297858921043_94 (
            .clk_in          (clk  [94]),
            .data_in         (data [94]),
            .scan_select_in  (scan [94]),
            .latch_enable_in (latch[94]),
            .clk_out         (clk  [95]),
            .data_out        (data [95]),
            .scan_select_out (scan [95]),
            .latch_enable_out(latch[95])
            );
        
        // https://github.com/coralmw/tinytapeout-css-feedback
        scan_wrapper_341710255833481812 #(.NUM_IOS(8)) scan_wrapper_341710255833481812_95 (
            .clk_in          (clk  [95]),
            .data_in         (data [95]),
            .scan_select_in  (scan [95]),
            .latch_enable_in (latch[95]),
            .clk_out         (clk  [96]),
            .data_out        (data [96]),
            .scan_select_out (scan [96]),
            .latch_enable_out(latch[96])
            );
        
        // https://github.com/ericsmi/tinytapeout-verilog-div3
        scan_wrapper_340067262721426004 #(.NUM_IOS(8)) scan_wrapper_340067262721426004_96 (
            .clk_in          (clk  [96]),
            .data_in         (data [96]),
            .scan_select_in  (scan [96]),
            .latch_enable_in (latch[96]),
            .clk_out         (clk  [97]),
            .data_out        (data [97]),
            .scan_select_out (scan [97]),
            .latch_enable_out(latch[97])
            );
        
        // https://github.com/fluxfocus/jdtt-logic1.git
        scan_wrapper_341462925422101075 #(.NUM_IOS(8)) scan_wrapper_341462925422101075_97 (
            .clk_in          (clk  [97]),
            .data_in         (data [97]),
            .scan_select_in  (scan [97]),
            .latch_enable_in (latch[97]),
            .clk_out         (clk  [98]),
            .data_out        (data [98]),
            .scan_select_out (scan [98]),
            .latch_enable_out(latch[98])
            );
        
        // https://github.com/anm/nyasic
        scan_wrapper_341520747710120530 #(.NUM_IOS(8)) scan_wrapper_341520747710120530_98 (
            .clk_in          (clk  [98]),
            .data_in         (data [98]),
            .scan_select_in  (scan [98]),
            .latch_enable_in (latch[98]),
            .clk_out         (clk  [99]),
            .data_out        (data [99]),
            .scan_select_out (scan [99]),
            .latch_enable_out(latch[99])
            );
        
        // https://github.com/aiunderstand/tinytapeout_bintristateloadablecounter
        scan_wrapper_341423712597181012 #(.NUM_IOS(8)) scan_wrapper_341423712597181012_99 (
            .clk_in          (clk  [99]),
            .data_in         (data [99]),
            .scan_select_in  (scan [99]),
            .latch_enable_in (latch[99]),
            .clk_out         (clk  [100]),
            .data_out        (data [100]),
            .scan_select_out (scan [100]),
            .latch_enable_out(latch[100])
            );
        
        // https://github.com/ThorKn/tinytapeout_shiftregister_challenge
        scan_wrapper_341516949939814994 #(.NUM_IOS(8)) scan_wrapper_341516949939814994_100 (
            .clk_in          (clk  [100]),
            .data_in         (data [100]),
            .scan_select_in  (scan [100]),
            .latch_enable_in (latch[100]),
            .clk_out         (clk  [101]),
            .data_out        (data [101]),
            .scan_select_out (scan [101]),
            .latch_enable_out(latch[101])
            );
        
        // https://github.com/regymm/tinytapeout-mcpi
        scan_wrapper_341521390605697619 #(.NUM_IOS(8)) scan_wrapper_341521390605697619_101 (
            .clk_in          (clk  [101]),
            .data_in         (data [101]),
            .scan_select_in  (scan [101]),
            .latch_enable_in (latch[101]),
            .clk_out         (clk  [102]),
            .data_out        (data [102]),
            .scan_select_out (scan [102]),
            .latch_enable_out(latch[102])
            );
        
        // https://github.com/todd1251/tinytapeout-figure8
        scan_wrapper_341243232292700755 #(.NUM_IOS(8)) scan_wrapper_341243232292700755_102 (
            .clk_in          (clk  [102]),
            .data_in         (data [102]),
            .scan_select_in  (scan [102]),
            .latch_enable_in (latch[102]),
            .clk_out         (clk  [103]),
            .data_out        (data [103]),
            .scan_select_out (scan [103]),
            .latch_enable_out(latch[103])
            );
        
        // https://github.com/CyberGai/tinytapeout-bcd-counter
        scan_wrapper_341519170869920338 #(.NUM_IOS(8)) scan_wrapper_341519170869920338_103 (
            .clk_in          (clk  [103]),
            .data_in         (data [103]),
            .scan_select_in  (scan [103]),
            .latch_enable_in (latch[103]),
            .clk_out         (clk  [104]),
            .data_out        (data [104]),
            .scan_select_out (scan [104]),
            .latch_enable_out(latch[104])
            );
        
        // https://github.com/georgeyhere/tinytapeout-dice-roller
        scan_wrapper_341446083683025490 #(.NUM_IOS(8)) scan_wrapper_341446083683025490_104 (
            .clk_in          (clk  [104]),
            .data_in         (data [104]),
            .scan_select_in  (scan [104]),
            .latch_enable_in (latch[104]),
            .clk_out         (clk  [105]),
            .data_out        (data [105]),
            .scan_select_out (scan [105]),
            .latch_enable_out(latch[105])
            );
        
        // https://github.com/nayanesh-reddy/2-Bit_Add_Mul_Comp
        scan_wrapper_341524192738411090 #(.NUM_IOS(8)) scan_wrapper_341524192738411090_105 (
            .clk_in          (clk  [105]),
            .data_in         (data [105]),
            .scan_select_in  (scan [105]),
            .latch_enable_in (latch[105]),
            .clk_out         (clk  [106]),
            .data_out        (data [106]),
            .scan_select_out (scan [106]),
            .latch_enable_out(latch[106])
            );
        
        // https://github.com/ryancor/half_addr_asic
        scan_wrapper_341533740987581011 #(.NUM_IOS(8)) scan_wrapper_341533740987581011_106 (
            .clk_in          (clk  [106]),
            .data_in         (data [106]),
            .scan_select_in  (scan [106]),
            .latch_enable_in (latch[106]),
            .clk_out         (clk  [107]),
            .data_out        (data [107]),
            .scan_select_out (scan [107]),
            .latch_enable_out(latch[107])
            );
        
        // https://github.com/hovind/tinytapeout-verilog-test
        scan_wrapper_341431502448362067 #(.NUM_IOS(8)) scan_wrapper_341431502448362067_107 (
            .clk_in          (clk  [107]),
            .data_in         (data [107]),
            .scan_select_in  (scan [107]),
            .latch_enable_in (latch[107]),
            .clk_out         (clk  [108]),
            .data_out        (data [108]),
            .scan_select_out (scan [108]),
            .latch_enable_out(latch[108])
            );
        
        // https://github.com/siriusm46/tinytapeout_bcd_decimal
        scan_wrapper_341473139924927058 #(.NUM_IOS(8)) scan_wrapper_341473139924927058_108 (
            .clk_in          (clk  [108]),
            .data_in         (data [108]),
            .scan_select_in  (scan [108]),
            .latch_enable_in (latch[108]),
            .clk_out         (clk  [109]),
            .data_out        (data [109]),
            .scan_select_out (scan [109]),
            .latch_enable_out(latch[109])
            );
        
        // https://github.com/cpldcpu/tinytapeout_mcpu5
        scan_wrapper_341528610027340372 #(.NUM_IOS(8)) scan_wrapper_341528610027340372_109 (
            .clk_in          (clk  [109]),
            .data_in         (data [109]),
            .scan_select_in  (scan [109]),
            .latch_enable_in (latch[109]),
            .clk_out         (clk  [110]),
            .data_out        (data [110]),
            .scan_select_out (scan [110]),
            .latch_enable_out(latch[110])
            );
        
        // https://github.com/goran-mahovlic/tinytapeout-verilog-piano
        scan_wrapper_341424636358034002 #(.NUM_IOS(8)) scan_wrapper_341424636358034002_110 (
            .clk_in          (clk  [110]),
            .data_in         (data [110]),
            .scan_select_in  (scan [110]),
            .latch_enable_in (latch[110]),
            .clk_out         (clk  [111]),
            .data_out        (data [111]),
            .scan_select_out (scan [111]),
            .latch_enable_out(latch[111])
            );
        
        // https://github.com/andars/universal-turing-machine-aw7s8
        scan_wrapper_341717091617866324 #(.NUM_IOS(8)) scan_wrapper_341717091617866324_111 (
            .clk_in          (clk  [111]),
            .data_in         (data [111]),
            .scan_select_in  (scan [111]),
            .latch_enable_in (latch[111]),
            .clk_out         (clk  [112]),
            .data_out        (data [112]),
            .scan_select_out (scan [112]),
            .latch_enable_out(latch[112])
            );
        
        // https://github.com/marcusmueller/hamming74-tapeout
        scan_wrapper_hamming74 #(.NUM_IOS(8)) scan_wrapper_hamming74_112 (
            .clk_in          (clk  [112]),
            .data_in         (data [112]),
            .scan_select_in  (scan [112]),
            .latch_enable_in (latch[112]),
            .clk_out         (clk  [113]),
            .data_out        (data [113]),
            .scan_select_out (scan [113]),
            .latch_enable_out(latch[113])
            );
        
        // https://github.com/13arn/tinytapeout_counter_steamdeck
        scan_wrapper_341541108650607187 #(.NUM_IOS(8)) scan_wrapper_341541108650607187_113 (
            .clk_in          (clk  [113]),
            .data_in         (data [113]),
            .scan_select_in  (scan [113]),
            .latch_enable_in (latch[113]),
            .clk_out         (clk  [114]),
            .data_out        (data [114]),
            .scan_select_out (scan [114]),
            .latch_enable_out(latch[114])
            );
        
        // https://github.com/johshoff/tinytapeout-verilog
        scan_wrapper_341360223723717202 #(.NUM_IOS(8)) scan_wrapper_341360223723717202_114 (
            .clk_in          (clk  [114]),
            .data_in         (data [114]),
            .scan_select_in  (scan [114]),
            .latch_enable_in (latch[114]),
            .clk_out         (clk  [115]),
            .data_out        (data [115]),
            .scan_select_out (scan [115]),
            .latch_enable_out(latch[115])
            );
        
        // https://github.com/cy384/seven-segment-with-adder
        scan_wrapper_341546888233747026 #(.NUM_IOS(8)) scan_wrapper_341546888233747026_115 (
            .clk_in          (clk  [115]),
            .data_in         (data [115]),
            .scan_select_in  (scan [115]),
            .latch_enable_in (latch[115]),
            .clk_out         (clk  [116]),
            .data_out        (data [116]),
            .scan_select_out (scan [116]),
            .latch_enable_out(latch[116])
            );
        
        // https://github.com/georgerennie/tinytapeout-wokwi-cd4518
        scan_wrapper_340979268609638995 #(.NUM_IOS(8)) scan_wrapper_340979268609638995_116 (
            .clk_in          (clk  [116]),
            .data_in         (data [116]),
            .scan_select_in  (scan [116]),
            .latch_enable_in (latch[116]),
            .clk_out         (clk  [117]),
            .data_out        (data [117]),
            .scan_select_out (scan [117]),
            .latch_enable_out(latch[117])
            );
        
        // https://github.com/ElectricPotato/tinytapeout-picture-printer-b
        scan_wrapper_341542971476279892 #(.NUM_IOS(8)) scan_wrapper_341542971476279892_117 (
            .clk_in          (clk  [117]),
            .data_in         (data [117]),
            .scan_select_in  (scan [117]),
            .latch_enable_in (latch[117]),
            .clk_out         (clk  [118]),
            .data_out        (data [118]),
            .scan_select_out (scan [118]),
            .latch_enable_out(latch[118])
            );
        
        // https://github.com/theFestest/tinytapeout-simple-invert8
        scan_wrapper_341556236196512338 #(.NUM_IOS(8)) scan_wrapper_341556236196512338_118 (
            .clk_in          (clk  [118]),
            .data_in         (data [118]),
            .scan_select_in  (scan [118]),
            .latch_enable_in (latch[118]),
            .clk_out         (clk  [119]),
            .data_out        (data [119]),
            .scan_select_out (scan [119]),
            .latch_enable_out(latch[119])
            );
        
        // https://github.com/ArsenioDev/CustomSiliconTest
        scan_wrapper_341558189536313940 #(.NUM_IOS(8)) scan_wrapper_341558189536313940_119 (
            .clk_in          (clk  [119]),
            .data_in         (data [119]),
            .scan_select_in  (scan [119]),
            .latch_enable_in (latch[119]),
            .clk_out         (clk  [120]),
            .data_out        (data [120]),
            .scan_select_out (scan [120]),
            .latch_enable_out(latch[120])
            );
        
        // https://github.com/mgargano/tinytapeout_alu_with_4bit_7segmetdisplay_decoder
        scan_wrapper_341538994733974098 #(.NUM_IOS(8)) scan_wrapper_341538994733974098_120 (
            .clk_in          (clk  [120]),
            .data_in         (data [120]),
            .scan_select_in  (scan [120]),
            .latch_enable_in (latch[120]),
            .clk_out         (clk  [121]),
            .data_out        (data [121]),
            .scan_select_out (scan [121]),
            .latch_enable_out(latch[121])
            );
        
        // https://github.com/theFestest/tinytapeout-4x4-ram
        scan_wrapper_341557831870186068 #(.NUM_IOS(8)) scan_wrapper_341557831870186068_121 (
            .clk_in          (clk  [121]),
            .data_in         (data [121]),
            .scan_select_in  (scan [121]),
            .latch_enable_in (latch[121]),
            .clk_out         (clk  [122]),
            .data_out        (data [122]),
            .scan_select_out (scan [122]),
            .latch_enable_out(latch[122])
            );
        
        // https://github.com/michael-christen/wokwi-verilog-asic-experiment
        scan_wrapper_341569483755749970 #(.NUM_IOS(8)) scan_wrapper_341569483755749970_122 (
            .clk_in          (clk  [122]),
            .data_in         (data [122]),
            .scan_select_in  (scan [122]),
            .latch_enable_in (latch[122]),
            .clk_out         (clk  [123]),
            .data_out        (data [123]),
            .scan_select_out (scan [123]),
            .latch_enable_out(latch[123])
            );
        
        // https://github.com/craigcc-frii/tinytapeout_craig
        scan_wrapper_341573751072096850 #(.NUM_IOS(8)) scan_wrapper_341573751072096850_123 (
            .clk_in          (clk  [123]),
            .data_in         (data [123]),
            .scan_select_in  (scan [123]),
            .latch_enable_in (latch[123]),
            .clk_out         (clk  [124]),
            .data_out        (data [124]),
            .scan_select_out (scan [124]),
            .latch_enable_out(latch[124])
            );
        
        // https://github.com/youngpines/r2rdac_tinytapeout_demo
        scan_wrapper_341571228858843732 #(.NUM_IOS(8)) scan_wrapper_341571228858843732_124 (
            .clk_in          (clk  [124]),
            .data_in         (data [124]),
            .scan_select_in  (scan [124]),
            .latch_enable_in (latch[124]),
            .clk_out         (clk  [125]),
            .data_out        (data [125]),
            .scan_select_out (scan [125]),
            .latch_enable_out(latch[125])
            );
        
        // https://github.com/toybuilder/learn-tinytapeout
        scan_wrapper_341490465660469844 #(.NUM_IOS(8)) scan_wrapper_341490465660469844_125 (
            .clk_in          (clk  [125]),
            .data_in         (data [125]),
            .scan_select_in  (scan [125]),
            .latch_enable_in (latch[125]),
            .clk_out         (clk  [126]),
            .data_out        (data [126]),
            .scan_select_out (scan [126]),
            .latch_enable_out(latch[126])
            );
        
        // https://github.com/eggsactly/tinytapeout_demo
        scan_wrapper_341581732833657427 #(.NUM_IOS(8)) scan_wrapper_341581732833657427_126 (
            .clk_in          (clk  [126]),
            .data_in         (data [126]),
            .scan_select_in  (scan [126]),
            .latch_enable_in (latch[126]),
            .clk_out         (clk  [127]),
            .data_out        (data [127]),
            .scan_select_out (scan [127]),
            .latch_enable_out(latch[127])
            );
        
        // https://github.com/gsegura96/tinytapeout-chisel
        scan_wrapper_341457494561784402 #(.NUM_IOS(8)) scan_wrapper_341457494561784402_127 (
            .clk_in          (clk  [127]),
            .data_in         (data [127]),
            .scan_select_in  (scan [127]),
            .latch_enable_in (latch[127]),
            .clk_out         (clk  [128]),
            .data_out        (data [128]),
            .scan_select_out (scan [128]),
            .latch_enable_out(latch[128])
            );
        
        // https://github.com/abf149/fbna_like_verilog_abf149
        scan_wrapper_341590933015364178 #(.NUM_IOS(8)) scan_wrapper_341590933015364178_128 (
            .clk_in          (clk  [128]),
            .data_in         (data [128]),
            .scan_select_in  (scan [128]),
            .latch_enable_in (latch[128]),
            .clk_out         (clk  [129]),
            .data_out        (data [129]),
            .scan_select_out (scan [129]),
            .latch_enable_out(latch[129])
            );
        
        // https://github.com/MC-SecPat/tinytapeout_chi2shares
        scan_wrapper_341589685194195540 #(.NUM_IOS(8)) scan_wrapper_341589685194195540_129 (
            .clk_in          (clk  [129]),
            .data_in         (data [129]),
            .scan_select_in  (scan [129]),
            .latch_enable_in (latch[129]),
            .clk_out         (clk  [130]),
            .data_out        (data [130]),
            .scan_select_out (scan [130]),
            .latch_enable_out(latch[130])
            );
        
        // https://github.com/MC-SecPat/tinytapeout_chi3shares
        scan_wrapper_341608574336631379 #(.NUM_IOS(8)) scan_wrapper_341608574336631379_130 (
            .clk_in          (clk  [130]),
            .data_in         (data [130]),
            .scan_select_in  (scan [130]),
            .latch_enable_in (latch[130]),
            .clk_out         (clk  [131]),
            .data_out        (data [131]),
            .scan_select_out (scan [131]),
            .latch_enable_out(latch[131])
            );
        
        // https://github.com/Adil8442/tiny_tapeout_test
        scan_wrapper_341608297106768466 #(.NUM_IOS(8)) scan_wrapper_341608297106768466_131 (
            .clk_in          (clk  [131]),
            .data_in         (data [131]),
            .scan_select_in  (scan [131]),
            .latch_enable_in (latch[131]),
            .clk_out         (clk  [132]),
            .data_out        (data [132]),
            .scan_select_out (scan [132]),
            .latch_enable_out(latch[132])
            );
        
        // https://github.com/mattvenn/tinytapeout-341802448429515346
        scan_wrapper_341802448429515346 #(.NUM_IOS(8)) scan_wrapper_341802448429515346_132 (
            .clk_in          (clk  [132]),
            .data_in         (data [132]),
            .scan_select_in  (scan [132]),
            .latch_enable_in (latch[132]),
            .clk_out         (clk  [133]),
            .data_out        (data [133]),
            .scan_select_out (scan [133]),
            .latch_enable_out(latch[133])
            );
        
        // https://github.com/r4d10n/tinytapeout-HELLo-3orLd-7seg
        scan_wrapper_341609034095264340 #(.NUM_IOS(8)) scan_wrapper_341609034095264340_133 (
            .clk_in          (clk  [133]),
            .data_in         (data [133]),
            .scan_select_in  (scan [133]),
            .latch_enable_in (latch[133]),
            .clk_out         (clk  [134]),
            .data_out        (data [134]),
            .scan_select_out (scan [134]),
            .latch_enable_out(latch[134])
            );
        
        // https://github.com/proppy/tinytapeout-xls-graydec
        scan_wrapper_341617722294010450 #(.NUM_IOS(8)) scan_wrapper_341617722294010450_134 (
            .clk_in          (clk  [134]),
            .data_in         (data [134]),
            .scan_select_in  (scan [134]),
            .latch_enable_in (latch[134]),
            .clk_out         (clk  [135]),
            .data_out        (data [135]),
            .scan_select_out (scan [135]),
            .latch_enable_out(latch[135])
            );
        
        // https://github.com/prabaldutta/tinytapeout_adi
        scan_wrapper_341613097060926036 #(.NUM_IOS(8)) scan_wrapper_341613097060926036_135 (
            .clk_in          (clk  [135]),
            .data_in         (data [135]),
            .scan_select_in  (scan [135]),
            .latch_enable_in (latch[135]),
            .clk_out         (clk  [136]),
            .data_out        (data [136]),
            .scan_select_out (scan [136]),
            .latch_enable_out(latch[136])
            );
        
        // https://github.com/maehw/wokwi-verilog-gds-wolf-goat-cabbage
        scan_wrapper_341614346808328788 #(.NUM_IOS(8)) scan_wrapper_341614346808328788_136 (
            .clk_in          (clk  [136]),
            .data_in         (data [136]),
            .scan_select_in  (scan [136]),
            .latch_enable_in (latch[136]),
            .clk_out         (clk  [137]),
            .data_out        (data [137]),
            .scan_select_out (scan [137]),
            .latch_enable_out(latch[137])
            );
        
        // https://github.com/ThorKn/tinytapeout_pattern_player
        scan_wrapper_341620484740219475 #(.NUM_IOS(8)) scan_wrapper_341620484740219475_137 (
            .clk_in          (clk  [137]),
            .data_in         (data [137]),
            .scan_select_in  (scan [137]),
            .latch_enable_in (latch[137]),
            .clk_out         (clk  [138]),
            .data_out        (data [138]),
            .scan_select_out (scan [138]),
            .latch_enable_out(latch[138])
            );
        
        // https://github.com/rigobertoruiz98/cts_fsm
        scan_wrapper_341624400621077076 #(.NUM_IOS(8)) scan_wrapper_341624400621077076_138 (
            .clk_in          (clk  [138]),
            .data_in         (data [138]),
            .scan_select_in  (scan [138]),
            .latch_enable_in (latch[138]),
            .clk_out         (clk  [139]),
            .data_out        (data [139]),
            .scan_select_out (scan [139]),
            .latch_enable_out(latch[139])
            );
        
        // https://github.com/rajarshiroy/tinytapout0_rajarshi
        scan_wrapper_341614536664547922 #(.NUM_IOS(8)) scan_wrapper_341614536664547922_139 (
            .clk_in          (clk  [139]),
            .data_in         (data [139]),
            .scan_select_in  (scan [139]),
            .latch_enable_in (latch[139]),
            .clk_out         (clk  [140]),
            .data_out        (data [140]),
            .scan_select_out (scan [140]),
            .latch_enable_out(latch[140])
            );
        
        // https://github.com/BarsMonster/MicroASIC
        scan_wrapper_341567111632519764 #(.NUM_IOS(8)) scan_wrapper_341567111632519764_140 (
            .clk_in          (clk  [140]),
            .data_in         (data [140]),
            .scan_select_in  (scan [140]),
            .latch_enable_in (latch[140]),
            .clk_out         (clk  [141]),
            .data_out        (data [141]),
            .scan_select_out (scan [141]),
            .latch_enable_out(latch[141])
            );
        
        // https://github.com/kammoh/tinytapeout-chisel
        scan_wrapper_3398002391929329472 #(.NUM_IOS(8)) scan_wrapper_3398002391929329472_141 (
            .clk_in          (clk  [141]),
            .data_in         (data [141]),
            .scan_select_in  (scan [141]),
            .latch_enable_in (latch[141]),
            .clk_out         (clk  [142]),
            .data_out        (data [142]),
            .scan_select_out (scan [142]),
            .latch_enable_out(latch[142])
            );
        
        // https://github.com/cpldcpu/TinyTapeout_TrainLED
        scan_wrapper_341631485498884690 #(.NUM_IOS(8)) scan_wrapper_341631485498884690_142 (
            .clk_in          (clk  [142]),
            .data_in         (data [142]),
            .scan_select_in  (scan [142]),
            .latch_enable_in (latch[142]),
            .clk_out         (clk  [143]),
            .data_out        (data [143]),
            .scan_select_out (scan [143]),
            .latch_enable_out(latch[143])
            );
        
        // https://github.com/malkam03/tinytapeout-game-of-life
        scan_wrapper_341632596577354323 #(.NUM_IOS(8)) scan_wrapper_341632596577354323_143 (
            .clk_in          (clk  [143]),
            .data_in         (data [143]),
            .scan_select_in  (scan [143]),
            .latch_enable_in (latch[143]),
            .clk_out         (clk  [144]),
            .data_out        (data [144]),
            .scan_select_out (scan [144]),
            .latch_enable_out(latch[144])
            );
        
        // https://github.com/BarsMonster/MicroAsicV
        scan_wrapper_341628725785264722 #(.NUM_IOS(8)) scan_wrapper_341628725785264722_144 (
            .clk_in          (clk  [144]),
            .data_in         (data [144]),
            .scan_select_in  (scan [144]),
            .latch_enable_in (latch[144]),
            .clk_out         (clk  [145]),
            .data_out        (data [145]),
            .scan_select_out (scan [145]),
            .latch_enable_out(latch[145])
            );
        
        // https://github.com/maehw/wokwi-verilog-gds-lowspeed-tiny-uart
        scan_wrapper_341631511790879314 #(.NUM_IOS(8)) scan_wrapper_341631511790879314_145 (
            .clk_in          (clk  [145]),
            .data_in         (data [145]),
            .scan_select_in  (scan [145]),
            .latch_enable_in (latch[145]),
            .clk_out         (clk  [146]),
            .data_out        (data [146]),
            .scan_select_out (scan [146]),
            .latch_enable_out(latch[146])
            );
        
        // https://github.com/smunaut/tinytapeout-smolram
        scan_wrapper_341426151397261906 #(.NUM_IOS(8)) scan_wrapper_341426151397261906_146 (
            .clk_in          (clk  [146]),
            .data_in         (data [146]),
            .scan_select_in  (scan [146]),
            .latch_enable_in (latch[146]),
            .clk_out         (clk  [147]),
            .data_out        (data [147]),
            .scan_select_out (scan [147]),
            .latch_enable_out(latch[147])
            );
        
        // https://github.com/sirejdua/6bit-cellular-automata-tinytapeout
        scan_wrapper_341629415144292948 #(.NUM_IOS(8)) scan_wrapper_341629415144292948_147 (
            .clk_in          (clk  [147]),
            .data_in         (data [147]),
            .scan_select_in  (scan [147]),
            .latch_enable_in (latch[147]),
            .clk_out         (clk  [148]),
            .data_out        (data [148]),
            .scan_select_out (scan [148]),
            .latch_enable_out(latch[148])
            );
        
        // https://github.com/DuaneSand/TinyTapeout-Hello
        scan_wrapper_341637831098106450 #(.NUM_IOS(8)) scan_wrapper_341637831098106450_148 (
            .clk_in          (clk  [148]),
            .data_in         (data [148]),
            .scan_select_in  (scan [148]),
            .latch_enable_in (latch[148]),
            .clk_out         (clk  [149]),
            .data_out        (data [149]),
            .scan_select_out (scan [149]),
            .latch_enable_out(latch[149])
            );
        
        // https://github.com/tzachari/tinytapeout-lab11
        scan_wrapper_341631644820570706 #(.NUM_IOS(8)) scan_wrapper_341631644820570706_149 (
            .clk_in          (clk  [149]),
            .data_in         (data [149]),
            .scan_select_in  (scan [149]),
            .latch_enable_in (latch[149]),
            .clk_out         (clk  [150]),
            .data_out        (data [150]),
            .scan_select_out (scan [150]),
            .latch_enable_out(latch[150])
            );
        
        // https://github.com/mattvenn/tinytapeout-marc
        scan_wrapper_340596276030603858 #(.NUM_IOS(8)) scan_wrapper_340596276030603858_150 (
            .clk_in          (clk  [150]),
            .data_in         (data [150]),
            .scan_select_in  (scan [150]),
            .latch_enable_in (latch[150]),
            .clk_out         (clk  [151]),
            .data_out        (data [151]),
            .scan_select_out (scan [151]),
            .latch_enable_out(latch[151])
            );
        
        // https://github.com/mattvenn/tinytapeout-laura
        scan_wrapper_341678527574180436 #(.NUM_IOS(8)) scan_wrapper_341678527574180436_151 (
            .clk_in          (clk  [151]),
            .data_in         (data [151]),
            .scan_select_in  (scan [151]),
            .latch_enable_in (latch[151]),
            .clk_out         (clk  [152]),
            .data_out        (data [152]),
            .scan_select_out (scan [152]),
            .latch_enable_out(latch[152])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_152 (
            .clk_in          (clk  [152]),
            .data_in         (data [152]),
            .scan_select_in  (scan [152]),
            .latch_enable_in (latch[152]),
            .clk_out         (clk  [153]),
            .data_out        (data [153]),
            .scan_select_out (scan [153]),
            .latch_enable_out(latch[153])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_153 (
            .clk_in          (clk  [153]),
            .data_in         (data [153]),
            .scan_select_in  (scan [153]),
            .latch_enable_in (latch[153]),
            .clk_out         (clk  [154]),
            .data_out        (data [154]),
            .scan_select_out (scan [154]),
            .latch_enable_out(latch[154])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_154 (
            .clk_in          (clk  [154]),
            .data_in         (data [154]),
            .scan_select_in  (scan [154]),
            .latch_enable_in (latch[154]),
            .clk_out         (clk  [155]),
            .data_out        (data [155]),
            .scan_select_out (scan [155]),
            .latch_enable_out(latch[155])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_155 (
            .clk_in          (clk  [155]),
            .data_in         (data [155]),
            .scan_select_in  (scan [155]),
            .latch_enable_in (latch[155]),
            .clk_out         (clk  [156]),
            .data_out        (data [156]),
            .scan_select_out (scan [156]),
            .latch_enable_out(latch[156])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_156 (
            .clk_in          (clk  [156]),
            .data_in         (data [156]),
            .scan_select_in  (scan [156]),
            .latch_enable_in (latch[156]),
            .clk_out         (clk  [157]),
            .data_out        (data [157]),
            .scan_select_out (scan [157]),
            .latch_enable_out(latch[157])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_157 (
            .clk_in          (clk  [157]),
            .data_in         (data [157]),
            .scan_select_in  (scan [157]),
            .latch_enable_in (latch[157]),
            .clk_out         (clk  [158]),
            .data_out        (data [158]),
            .scan_select_out (scan [158]),
            .latch_enable_out(latch[158])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_158 (
            .clk_in          (clk  [158]),
            .data_in         (data [158]),
            .scan_select_in  (scan [158]),
            .latch_enable_in (latch[158]),
            .clk_out         (clk  [159]),
            .data_out        (data [159]),
            .scan_select_out (scan [159]),
            .latch_enable_out(latch[159])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_159 (
            .clk_in          (clk  [159]),
            .data_in         (data [159]),
            .scan_select_in  (scan [159]),
            .latch_enable_in (latch[159]),
            .clk_out         (clk  [160]),
            .data_out        (data [160]),
            .scan_select_out (scan [160]),
            .latch_enable_out(latch[160])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_160 (
            .clk_in          (clk  [160]),
            .data_in         (data [160]),
            .scan_select_in  (scan [160]),
            .latch_enable_in (latch[160]),
            .clk_out         (clk  [161]),
            .data_out        (data [161]),
            .scan_select_out (scan [161]),
            .latch_enable_out(latch[161])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_161 (
            .clk_in          (clk  [161]),
            .data_in         (data [161]),
            .scan_select_in  (scan [161]),
            .latch_enable_in (latch[161]),
            .clk_out         (clk  [162]),
            .data_out        (data [162]),
            .scan_select_out (scan [162]),
            .latch_enable_out(latch[162])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_162 (
            .clk_in          (clk  [162]),
            .data_in         (data [162]),
            .scan_select_in  (scan [162]),
            .latch_enable_in (latch[162]),
            .clk_out         (clk  [163]),
            .data_out        (data [163]),
            .scan_select_out (scan [163]),
            .latch_enable_out(latch[163])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_163 (
            .clk_in          (clk  [163]),
            .data_in         (data [163]),
            .scan_select_in  (scan [163]),
            .latch_enable_in (latch[163]),
            .clk_out         (clk  [164]),
            .data_out        (data [164]),
            .scan_select_out (scan [164]),
            .latch_enable_out(latch[164])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_164 (
            .clk_in          (clk  [164]),
            .data_in         (data [164]),
            .scan_select_in  (scan [164]),
            .latch_enable_in (latch[164]),
            .clk_out         (clk  [165]),
            .data_out        (data [165]),
            .scan_select_out (scan [165]),
            .latch_enable_out(latch[165])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_165 (
            .clk_in          (clk  [165]),
            .data_in         (data [165]),
            .scan_select_in  (scan [165]),
            .latch_enable_in (latch[165]),
            .clk_out         (clk  [166]),
            .data_out        (data [166]),
            .scan_select_out (scan [166]),
            .latch_enable_out(latch[166])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_166 (
            .clk_in          (clk  [166]),
            .data_in         (data [166]),
            .scan_select_in  (scan [166]),
            .latch_enable_in (latch[166]),
            .clk_out         (clk  [167]),
            .data_out        (data [167]),
            .scan_select_out (scan [167]),
            .latch_enable_out(latch[167])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_167 (
            .clk_in          (clk  [167]),
            .data_in         (data [167]),
            .scan_select_in  (scan [167]),
            .latch_enable_in (latch[167]),
            .clk_out         (clk  [168]),
            .data_out        (data [168]),
            .scan_select_out (scan [168]),
            .latch_enable_out(latch[168])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_168 (
            .clk_in          (clk  [168]),
            .data_in         (data [168]),
            .scan_select_in  (scan [168]),
            .latch_enable_in (latch[168]),
            .clk_out         (clk  [169]),
            .data_out        (data [169]),
            .scan_select_out (scan [169]),
            .latch_enable_out(latch[169])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_169 (
            .clk_in          (clk  [169]),
            .data_in         (data [169]),
            .scan_select_in  (scan [169]),
            .latch_enable_in (latch[169]),
            .clk_out         (clk  [170]),
            .data_out        (data [170]),
            .scan_select_out (scan [170]),
            .latch_enable_out(latch[170])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_170 (
            .clk_in          (clk  [170]),
            .data_in         (data [170]),
            .scan_select_in  (scan [170]),
            .latch_enable_in (latch[170]),
            .clk_out         (clk  [171]),
            .data_out        (data [171]),
            .scan_select_out (scan [171]),
            .latch_enable_out(latch[171])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_171 (
            .clk_in          (clk  [171]),
            .data_in         (data [171]),
            .scan_select_in  (scan [171]),
            .latch_enable_in (latch[171]),
            .clk_out         (clk  [172]),
            .data_out        (data [172]),
            .scan_select_out (scan [172]),
            .latch_enable_out(latch[172])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_172 (
            .clk_in          (clk  [172]),
            .data_in         (data [172]),
            .scan_select_in  (scan [172]),
            .latch_enable_in (latch[172]),
            .clk_out         (clk  [173]),
            .data_out        (data [173]),
            .scan_select_out (scan [173]),
            .latch_enable_out(latch[173])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_173 (
            .clk_in          (clk  [173]),
            .data_in         (data [173]),
            .scan_select_in  (scan [173]),
            .latch_enable_in (latch[173]),
            .clk_out         (clk  [174]),
            .data_out        (data [174]),
            .scan_select_out (scan [174]),
            .latch_enable_out(latch[174])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_174 (
            .clk_in          (clk  [174]),
            .data_in         (data [174]),
            .scan_select_in  (scan [174]),
            .latch_enable_in (latch[174]),
            .clk_out         (clk  [175]),
            .data_out        (data [175]),
            .scan_select_out (scan [175]),
            .latch_enable_out(latch[175])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_175 (
            .clk_in          (clk  [175]),
            .data_in         (data [175]),
            .scan_select_in  (scan [175]),
            .latch_enable_in (latch[175]),
            .clk_out         (clk  [176]),
            .data_out        (data [176]),
            .scan_select_out (scan [176]),
            .latch_enable_out(latch[176])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_176 (
            .clk_in          (clk  [176]),
            .data_in         (data [176]),
            .scan_select_in  (scan [176]),
            .latch_enable_in (latch[176]),
            .clk_out         (clk  [177]),
            .data_out        (data [177]),
            .scan_select_out (scan [177]),
            .latch_enable_out(latch[177])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_177 (
            .clk_in          (clk  [177]),
            .data_in         (data [177]),
            .scan_select_in  (scan [177]),
            .latch_enable_in (latch[177]),
            .clk_out         (clk  [178]),
            .data_out        (data [178]),
            .scan_select_out (scan [178]),
            .latch_enable_out(latch[178])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_178 (
            .clk_in          (clk  [178]),
            .data_in         (data [178]),
            .scan_select_in  (scan [178]),
            .latch_enable_in (latch[178]),
            .clk_out         (clk  [179]),
            .data_out        (data [179]),
            .scan_select_out (scan [179]),
            .latch_enable_out(latch[179])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_179 (
            .clk_in          (clk  [179]),
            .data_in         (data [179]),
            .scan_select_in  (scan [179]),
            .latch_enable_in (latch[179]),
            .clk_out         (clk  [180]),
            .data_out        (data [180]),
            .scan_select_out (scan [180]),
            .latch_enable_out(latch[180])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_180 (
            .clk_in          (clk  [180]),
            .data_in         (data [180]),
            .scan_select_in  (scan [180]),
            .latch_enable_in (latch[180]),
            .clk_out         (clk  [181]),
            .data_out        (data [181]),
            .scan_select_out (scan [181]),
            .latch_enable_out(latch[181])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_181 (
            .clk_in          (clk  [181]),
            .data_in         (data [181]),
            .scan_select_in  (scan [181]),
            .latch_enable_in (latch[181]),
            .clk_out         (clk  [182]),
            .data_out        (data [182]),
            .scan_select_out (scan [182]),
            .latch_enable_out(latch[182])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_182 (
            .clk_in          (clk  [182]),
            .data_in         (data [182]),
            .scan_select_in  (scan [182]),
            .latch_enable_in (latch[182]),
            .clk_out         (clk  [183]),
            .data_out        (data [183]),
            .scan_select_out (scan [183]),
            .latch_enable_out(latch[183])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_183 (
            .clk_in          (clk  [183]),
            .data_in         (data [183]),
            .scan_select_in  (scan [183]),
            .latch_enable_in (latch[183]),
            .clk_out         (clk  [184]),
            .data_out        (data [184]),
            .scan_select_out (scan [184]),
            .latch_enable_out(latch[184])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_184 (
            .clk_in          (clk  [184]),
            .data_in         (data [184]),
            .scan_select_in  (scan [184]),
            .latch_enable_in (latch[184]),
            .clk_out         (clk  [185]),
            .data_out        (data [185]),
            .scan_select_out (scan [185]),
            .latch_enable_out(latch[185])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_185 (
            .clk_in          (clk  [185]),
            .data_in         (data [185]),
            .scan_select_in  (scan [185]),
            .latch_enable_in (latch[185]),
            .clk_out         (clk  [186]),
            .data_out        (data [186]),
            .scan_select_out (scan [186]),
            .latch_enable_out(latch[186])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_186 (
            .clk_in          (clk  [186]),
            .data_in         (data [186]),
            .scan_select_in  (scan [186]),
            .latch_enable_in (latch[186]),
            .clk_out         (clk  [187]),
            .data_out        (data [187]),
            .scan_select_out (scan [187]),
            .latch_enable_out(latch[187])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_187 (
            .clk_in          (clk  [187]),
            .data_in         (data [187]),
            .scan_select_in  (scan [187]),
            .latch_enable_in (latch[187]),
            .clk_out         (clk  [188]),
            .data_out        (data [188]),
            .scan_select_out (scan [188]),
            .latch_enable_out(latch[188])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_188 (
            .clk_in          (clk  [188]),
            .data_in         (data [188]),
            .scan_select_in  (scan [188]),
            .latch_enable_in (latch[188]),
            .clk_out         (clk  [189]),
            .data_out        (data [189]),
            .scan_select_out (scan [189]),
            .latch_enable_out(latch[189])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_189 (
            .clk_in          (clk  [189]),
            .data_in         (data [189]),
            .scan_select_in  (scan [189]),
            .latch_enable_in (latch[189]),
            .clk_out         (clk  [190]),
            .data_out        (data [190]),
            .scan_select_out (scan [190]),
            .latch_enable_out(latch[190])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_190 (
            .clk_in          (clk  [190]),
            .data_in         (data [190]),
            .scan_select_in  (scan [190]),
            .latch_enable_in (latch[190]),
            .clk_out         (clk  [191]),
            .data_out        (data [191]),
            .scan_select_out (scan [191]),
            .latch_enable_out(latch[191])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_191 (
            .clk_in          (clk  [191]),
            .data_in         (data [191]),
            .scan_select_in  (scan [191]),
            .latch_enable_in (latch[191]),
            .clk_out         (clk  [192]),
            .data_out        (data [192]),
            .scan_select_out (scan [192]),
            .latch_enable_out(latch[192])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_192 (
            .clk_in          (clk  [192]),
            .data_in         (data [192]),
            .scan_select_in  (scan [192]),
            .latch_enable_in (latch[192]),
            .clk_out         (clk  [193]),
            .data_out        (data [193]),
            .scan_select_out (scan [193]),
            .latch_enable_out(latch[193])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_193 (
            .clk_in          (clk  [193]),
            .data_in         (data [193]),
            .scan_select_in  (scan [193]),
            .latch_enable_in (latch[193]),
            .clk_out         (clk  [194]),
            .data_out        (data [194]),
            .scan_select_out (scan [194]),
            .latch_enable_out(latch[194])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_194 (
            .clk_in          (clk  [194]),
            .data_in         (data [194]),
            .scan_select_in  (scan [194]),
            .latch_enable_in (latch[194]),
            .clk_out         (clk  [195]),
            .data_out        (data [195]),
            .scan_select_out (scan [195]),
            .latch_enable_out(latch[195])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_195 (
            .clk_in          (clk  [195]),
            .data_in         (data [195]),
            .scan_select_in  (scan [195]),
            .latch_enable_in (latch[195]),
            .clk_out         (clk  [196]),
            .data_out        (data [196]),
            .scan_select_out (scan [196]),
            .latch_enable_out(latch[196])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_196 (
            .clk_in          (clk  [196]),
            .data_in         (data [196]),
            .scan_select_in  (scan [196]),
            .latch_enable_in (latch[196]),
            .clk_out         (clk  [197]),
            .data_out        (data [197]),
            .scan_select_out (scan [197]),
            .latch_enable_out(latch[197])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_197 (
            .clk_in          (clk  [197]),
            .data_in         (data [197]),
            .scan_select_in  (scan [197]),
            .latch_enable_in (latch[197]),
            .clk_out         (clk  [198]),
            .data_out        (data [198]),
            .scan_select_out (scan [198]),
            .latch_enable_out(latch[198])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_198 (
            .clk_in          (clk  [198]),
            .data_in         (data [198]),
            .scan_select_in  (scan [198]),
            .latch_enable_in (latch[198]),
            .clk_out         (clk  [199]),
            .data_out        (data [199]),
            .scan_select_out (scan [199]),
            .latch_enable_out(latch[199])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_199 (
            .clk_in          (clk  [199]),
            .data_in         (data [199]),
            .scan_select_in  (scan [199]),
            .latch_enable_in (latch[199]),
            .clk_out         (clk  [200]),
            .data_out        (data [200]),
            .scan_select_out (scan [200]),
            .latch_enable_out(latch[200])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_200 (
            .clk_in          (clk  [200]),
            .data_in         (data [200]),
            .scan_select_in  (scan [200]),
            .latch_enable_in (latch[200]),
            .clk_out         (clk  [201]),
            .data_out        (data [201]),
            .scan_select_out (scan [201]),
            .latch_enable_out(latch[201])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_201 (
            .clk_in          (clk  [201]),
            .data_in         (data [201]),
            .scan_select_in  (scan [201]),
            .latch_enable_in (latch[201]),
            .clk_out         (clk  [202]),
            .data_out        (data [202]),
            .scan_select_out (scan [202]),
            .latch_enable_out(latch[202])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_202 (
            .clk_in          (clk  [202]),
            .data_in         (data [202]),
            .scan_select_in  (scan [202]),
            .latch_enable_in (latch[202]),
            .clk_out         (clk  [203]),
            .data_out        (data [203]),
            .scan_select_out (scan [203]),
            .latch_enable_out(latch[203])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_203 (
            .clk_in          (clk  [203]),
            .data_in         (data [203]),
            .scan_select_in  (scan [203]),
            .latch_enable_in (latch[203]),
            .clk_out         (clk  [204]),
            .data_out        (data [204]),
            .scan_select_out (scan [204]),
            .latch_enable_out(latch[204])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_204 (
            .clk_in          (clk  [204]),
            .data_in         (data [204]),
            .scan_select_in  (scan [204]),
            .latch_enable_in (latch[204]),
            .clk_out         (clk  [205]),
            .data_out        (data [205]),
            .scan_select_out (scan [205]),
            .latch_enable_out(latch[205])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_205 (
            .clk_in          (clk  [205]),
            .data_in         (data [205]),
            .scan_select_in  (scan [205]),
            .latch_enable_in (latch[205]),
            .clk_out         (clk  [206]),
            .data_out        (data [206]),
            .scan_select_out (scan [206]),
            .latch_enable_out(latch[206])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_206 (
            .clk_in          (clk  [206]),
            .data_in         (data [206]),
            .scan_select_in  (scan [206]),
            .latch_enable_in (latch[206]),
            .clk_out         (clk  [207]),
            .data_out        (data [207]),
            .scan_select_out (scan [207]),
            .latch_enable_out(latch[207])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_207 (
            .clk_in          (clk  [207]),
            .data_in         (data [207]),
            .scan_select_in  (scan [207]),
            .latch_enable_in (latch[207]),
            .clk_out         (clk  [208]),
            .data_out        (data [208]),
            .scan_select_out (scan [208]),
            .latch_enable_out(latch[208])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_208 (
            .clk_in          (clk  [208]),
            .data_in         (data [208]),
            .scan_select_in  (scan [208]),
            .latch_enable_in (latch[208]),
            .clk_out         (clk  [209]),
            .data_out        (data [209]),
            .scan_select_out (scan [209]),
            .latch_enable_out(latch[209])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_209 (
            .clk_in          (clk  [209]),
            .data_in         (data [209]),
            .scan_select_in  (scan [209]),
            .latch_enable_in (latch[209]),
            .clk_out         (clk  [210]),
            .data_out        (data [210]),
            .scan_select_out (scan [210]),
            .latch_enable_out(latch[210])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_210 (
            .clk_in          (clk  [210]),
            .data_in         (data [210]),
            .scan_select_in  (scan [210]),
            .latch_enable_in (latch[210]),
            .clk_out         (clk  [211]),
            .data_out        (data [211]),
            .scan_select_out (scan [211]),
            .latch_enable_out(latch[211])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_211 (
            .clk_in          (clk  [211]),
            .data_in         (data [211]),
            .scan_select_in  (scan [211]),
            .latch_enable_in (latch[211]),
            .clk_out         (clk  [212]),
            .data_out        (data [212]),
            .scan_select_out (scan [212]),
            .latch_enable_out(latch[212])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_212 (
            .clk_in          (clk  [212]),
            .data_in         (data [212]),
            .scan_select_in  (scan [212]),
            .latch_enable_in (latch[212]),
            .clk_out         (clk  [213]),
            .data_out        (data [213]),
            .scan_select_out (scan [213]),
            .latch_enable_out(latch[213])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_213 (
            .clk_in          (clk  [213]),
            .data_in         (data [213]),
            .scan_select_in  (scan [213]),
            .latch_enable_in (latch[213]),
            .clk_out         (clk  [214]),
            .data_out        (data [214]),
            .scan_select_out (scan [214]),
            .latch_enable_out(latch[214])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_214 (
            .clk_in          (clk  [214]),
            .data_in         (data [214]),
            .scan_select_in  (scan [214]),
            .latch_enable_in (latch[214]),
            .clk_out         (clk  [215]),
            .data_out        (data [215]),
            .scan_select_out (scan [215]),
            .latch_enable_out(latch[215])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_215 (
            .clk_in          (clk  [215]),
            .data_in         (data [215]),
            .scan_select_in  (scan [215]),
            .latch_enable_in (latch[215]),
            .clk_out         (clk  [216]),
            .data_out        (data [216]),
            .scan_select_out (scan [216]),
            .latch_enable_out(latch[216])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_216 (
            .clk_in          (clk  [216]),
            .data_in         (data [216]),
            .scan_select_in  (scan [216]),
            .latch_enable_in (latch[216]),
            .clk_out         (clk  [217]),
            .data_out        (data [217]),
            .scan_select_out (scan [217]),
            .latch_enable_out(latch[217])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_217 (
            .clk_in          (clk  [217]),
            .data_in         (data [217]),
            .scan_select_in  (scan [217]),
            .latch_enable_in (latch[217]),
            .clk_out         (clk  [218]),
            .data_out        (data [218]),
            .scan_select_out (scan [218]),
            .latch_enable_out(latch[218])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_218 (
            .clk_in          (clk  [218]),
            .data_in         (data [218]),
            .scan_select_in  (scan [218]),
            .latch_enable_in (latch[218]),
            .clk_out         (clk  [219]),
            .data_out        (data [219]),
            .scan_select_out (scan [219]),
            .latch_enable_out(latch[219])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_219 (
            .clk_in          (clk  [219]),
            .data_in         (data [219]),
            .scan_select_in  (scan [219]),
            .latch_enable_in (latch[219]),
            .clk_out         (clk  [220]),
            .data_out        (data [220]),
            .scan_select_out (scan [220]),
            .latch_enable_out(latch[220])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_220 (
            .clk_in          (clk  [220]),
            .data_in         (data [220]),
            .scan_select_in  (scan [220]),
            .latch_enable_in (latch[220]),
            .clk_out         (clk  [221]),
            .data_out        (data [221]),
            .scan_select_out (scan [221]),
            .latch_enable_out(latch[221])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_221 (
            .clk_in          (clk  [221]),
            .data_in         (data [221]),
            .scan_select_in  (scan [221]),
            .latch_enable_in (latch[221]),
            .clk_out         (clk  [222]),
            .data_out        (data [222]),
            .scan_select_out (scan [222]),
            .latch_enable_out(latch[222])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_222 (
            .clk_in          (clk  [222]),
            .data_in         (data [222]),
            .scan_select_in  (scan [222]),
            .latch_enable_in (latch[222]),
            .clk_out         (clk  [223]),
            .data_out        (data [223]),
            .scan_select_out (scan [223]),
            .latch_enable_out(latch[223])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_223 (
            .clk_in          (clk  [223]),
            .data_in         (data [223]),
            .scan_select_in  (scan [223]),
            .latch_enable_in (latch[223]),
            .clk_out         (clk  [224]),
            .data_out        (data [224]),
            .scan_select_out (scan [224]),
            .latch_enable_out(latch[224])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_224 (
            .clk_in          (clk  [224]),
            .data_in         (data [224]),
            .scan_select_in  (scan [224]),
            .latch_enable_in (latch[224]),
            .clk_out         (clk  [225]),
            .data_out        (data [225]),
            .scan_select_out (scan [225]),
            .latch_enable_out(latch[225])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_225 (
            .clk_in          (clk  [225]),
            .data_in         (data [225]),
            .scan_select_in  (scan [225]),
            .latch_enable_in (latch[225]),
            .clk_out         (clk  [226]),
            .data_out        (data [226]),
            .scan_select_out (scan [226]),
            .latch_enable_out(latch[226])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_226 (
            .clk_in          (clk  [226]),
            .data_in         (data [226]),
            .scan_select_in  (scan [226]),
            .latch_enable_in (latch[226]),
            .clk_out         (clk  [227]),
            .data_out        (data [227]),
            .scan_select_out (scan [227]),
            .latch_enable_out(latch[227])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_227 (
            .clk_in          (clk  [227]),
            .data_in         (data [227]),
            .scan_select_in  (scan [227]),
            .latch_enable_in (latch[227]),
            .clk_out         (clk  [228]),
            .data_out        (data [228]),
            .scan_select_out (scan [228]),
            .latch_enable_out(latch[228])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_228 (
            .clk_in          (clk  [228]),
            .data_in         (data [228]),
            .scan_select_in  (scan [228]),
            .latch_enable_in (latch[228]),
            .clk_out         (clk  [229]),
            .data_out        (data [229]),
            .scan_select_out (scan [229]),
            .latch_enable_out(latch[229])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_229 (
            .clk_in          (clk  [229]),
            .data_in         (data [229]),
            .scan_select_in  (scan [229]),
            .latch_enable_in (latch[229]),
            .clk_out         (clk  [230]),
            .data_out        (data [230]),
            .scan_select_out (scan [230]),
            .latch_enable_out(latch[230])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_230 (
            .clk_in          (clk  [230]),
            .data_in         (data [230]),
            .scan_select_in  (scan [230]),
            .latch_enable_in (latch[230]),
            .clk_out         (clk  [231]),
            .data_out        (data [231]),
            .scan_select_out (scan [231]),
            .latch_enable_out(latch[231])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_231 (
            .clk_in          (clk  [231]),
            .data_in         (data [231]),
            .scan_select_in  (scan [231]),
            .latch_enable_in (latch[231]),
            .clk_out         (clk  [232]),
            .data_out        (data [232]),
            .scan_select_out (scan [232]),
            .latch_enable_out(latch[232])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_232 (
            .clk_in          (clk  [232]),
            .data_in         (data [232]),
            .scan_select_in  (scan [232]),
            .latch_enable_in (latch[232]),
            .clk_out         (clk  [233]),
            .data_out        (data [233]),
            .scan_select_out (scan [233]),
            .latch_enable_out(latch[233])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_233 (
            .clk_in          (clk  [233]),
            .data_in         (data [233]),
            .scan_select_in  (scan [233]),
            .latch_enable_in (latch[233]),
            .clk_out         (clk  [234]),
            .data_out        (data [234]),
            .scan_select_out (scan [234]),
            .latch_enable_out(latch[234])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_234 (
            .clk_in          (clk  [234]),
            .data_in         (data [234]),
            .scan_select_in  (scan [234]),
            .latch_enable_in (latch[234]),
            .clk_out         (clk  [235]),
            .data_out        (data [235]),
            .scan_select_out (scan [235]),
            .latch_enable_out(latch[235])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_235 (
            .clk_in          (clk  [235]),
            .data_in         (data [235]),
            .scan_select_in  (scan [235]),
            .latch_enable_in (latch[235]),
            .clk_out         (clk  [236]),
            .data_out        (data [236]),
            .scan_select_out (scan [236]),
            .latch_enable_out(latch[236])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_236 (
            .clk_in          (clk  [236]),
            .data_in         (data [236]),
            .scan_select_in  (scan [236]),
            .latch_enable_in (latch[236]),
            .clk_out         (clk  [237]),
            .data_out        (data [237]),
            .scan_select_out (scan [237]),
            .latch_enable_out(latch[237])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_237 (
            .clk_in          (clk  [237]),
            .data_in         (data [237]),
            .scan_select_in  (scan [237]),
            .latch_enable_in (latch[237]),
            .clk_out         (clk  [238]),
            .data_out        (data [238]),
            .scan_select_out (scan [238]),
            .latch_enable_out(latch[238])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_238 (
            .clk_in          (clk  [238]),
            .data_in         (data [238]),
            .scan_select_in  (scan [238]),
            .latch_enable_in (latch[238]),
            .clk_out         (clk  [239]),
            .data_out        (data [239]),
            .scan_select_out (scan [239]),
            .latch_enable_out(latch[239])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_239 (
            .clk_in          (clk  [239]),
            .data_in         (data [239]),
            .scan_select_in  (scan [239]),
            .latch_enable_in (latch[239]),
            .clk_out         (clk  [240]),
            .data_out        (data [240]),
            .scan_select_out (scan [240]),
            .latch_enable_out(latch[240])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_240 (
            .clk_in          (clk  [240]),
            .data_in         (data [240]),
            .scan_select_in  (scan [240]),
            .latch_enable_in (latch[240]),
            .clk_out         (clk  [241]),
            .data_out        (data [241]),
            .scan_select_out (scan [241]),
            .latch_enable_out(latch[241])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_241 (
            .clk_in          (clk  [241]),
            .data_in         (data [241]),
            .scan_select_in  (scan [241]),
            .latch_enable_in (latch[241]),
            .clk_out         (clk  [242]),
            .data_out        (data [242]),
            .scan_select_out (scan [242]),
            .latch_enable_out(latch[242])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_242 (
            .clk_in          (clk  [242]),
            .data_in         (data [242]),
            .scan_select_in  (scan [242]),
            .latch_enable_in (latch[242]),
            .clk_out         (clk  [243]),
            .data_out        (data [243]),
            .scan_select_out (scan [243]),
            .latch_enable_out(latch[243])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_243 (
            .clk_in          (clk  [243]),
            .data_in         (data [243]),
            .scan_select_in  (scan [243]),
            .latch_enable_in (latch[243]),
            .clk_out         (clk  [244]),
            .data_out        (data [244]),
            .scan_select_out (scan [244]),
            .latch_enable_out(latch[244])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_244 (
            .clk_in          (clk  [244]),
            .data_in         (data [244]),
            .scan_select_in  (scan [244]),
            .latch_enable_in (latch[244]),
            .clk_out         (clk  [245]),
            .data_out        (data [245]),
            .scan_select_out (scan [245]),
            .latch_enable_out(latch[245])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_245 (
            .clk_in          (clk  [245]),
            .data_in         (data [245]),
            .scan_select_in  (scan [245]),
            .latch_enable_in (latch[245]),
            .clk_out         (clk  [246]),
            .data_out        (data [246]),
            .scan_select_out (scan [246]),
            .latch_enable_out(latch[246])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_246 (
            .clk_in          (clk  [246]),
            .data_in         (data [246]),
            .scan_select_in  (scan [246]),
            .latch_enable_in (latch[246]),
            .clk_out         (clk  [247]),
            .data_out        (data [247]),
            .scan_select_out (scan [247]),
            .latch_enable_out(latch[247])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_247 (
            .clk_in          (clk  [247]),
            .data_in         (data [247]),
            .scan_select_in  (scan [247]),
            .latch_enable_in (latch[247]),
            .clk_out         (clk  [248]),
            .data_out        (data [248]),
            .scan_select_out (scan [248]),
            .latch_enable_out(latch[248])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_248 (
            .clk_in          (clk  [248]),
            .data_in         (data [248]),
            .scan_select_in  (scan [248]),
            .latch_enable_in (latch[248]),
            .clk_out         (clk  [249]),
            .data_out        (data [249]),
            .scan_select_out (scan [249]),
            .latch_enable_out(latch[249])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_249 (
            .clk_in          (clk  [249]),
            .data_in         (data [249]),
            .scan_select_in  (scan [249]),
            .latch_enable_in (latch[249]),
            .clk_out         (clk  [250]),
            .data_out        (data [250]),
            .scan_select_out (scan [250]),
            .latch_enable_out(latch[250])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_250 (
            .clk_in          (clk  [250]),
            .data_in         (data [250]),
            .scan_select_in  (scan [250]),
            .latch_enable_in (latch[250]),
            .clk_out         (clk  [251]),
            .data_out        (data [251]),
            .scan_select_out (scan [251]),
            .latch_enable_out(latch[251])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_251 (
            .clk_in          (clk  [251]),
            .data_in         (data [251]),
            .scan_select_in  (scan [251]),
            .latch_enable_in (latch[251]),
            .clk_out         (clk  [252]),
            .data_out        (data [252]),
            .scan_select_out (scan [252]),
            .latch_enable_out(latch[252])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_252 (
            .clk_in          (clk  [252]),
            .data_in         (data [252]),
            .scan_select_in  (scan [252]),
            .latch_enable_in (latch[252]),
            .clk_out         (clk  [253]),
            .data_out        (data [253]),
            .scan_select_out (scan [253]),
            .latch_enable_out(latch[253])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_253 (
            .clk_in          (clk  [253]),
            .data_in         (data [253]),
            .scan_select_in  (scan [253]),
            .latch_enable_in (latch[253]),
            .clk_out         (clk  [254]),
            .data_out        (data [254]),
            .scan_select_out (scan [254]),
            .latch_enable_out(latch[254])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_254 (
            .clk_in          (clk  [254]),
            .data_in         (data [254]),
            .scan_select_in  (scan [254]),
            .latch_enable_in (latch[254]),
            .clk_out         (clk  [255]),
            .data_out        (data [255]),
            .scan_select_out (scan [255]),
            .latch_enable_out(latch[255])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_255 (
            .clk_in          (clk  [255]),
            .data_in         (data [255]),
            .scan_select_in  (scan [255]),
            .latch_enable_in (latch[255]),
            .clk_out         (clk  [256]),
            .data_out        (data [256]),
            .scan_select_out (scan [256]),
            .latch_enable_out(latch[256])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_256 (
            .clk_in          (clk  [256]),
            .data_in         (data [256]),
            .scan_select_in  (scan [256]),
            .latch_enable_in (latch[256]),
            .clk_out         (clk  [257]),
            .data_out        (data [257]),
            .scan_select_out (scan [257]),
            .latch_enable_out(latch[257])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_257 (
            .clk_in          (clk  [257]),
            .data_in         (data [257]),
            .scan_select_in  (scan [257]),
            .latch_enable_in (latch[257]),
            .clk_out         (clk  [258]),
            .data_out        (data [258]),
            .scan_select_out (scan [258]),
            .latch_enable_out(latch[258])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_258 (
            .clk_in          (clk  [258]),
            .data_in         (data [258]),
            .scan_select_in  (scan [258]),
            .latch_enable_in (latch[258]),
            .clk_out         (clk  [259]),
            .data_out        (data [259]),
            .scan_select_out (scan [259]),
            .latch_enable_out(latch[259])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_259 (
            .clk_in          (clk  [259]),
            .data_in         (data [259]),
            .scan_select_in  (scan [259]),
            .latch_enable_in (latch[259]),
            .clk_out         (clk  [260]),
            .data_out        (data [260]),
            .scan_select_out (scan [260]),
            .latch_enable_out(latch[260])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_260 (
            .clk_in          (clk  [260]),
            .data_in         (data [260]),
            .scan_select_in  (scan [260]),
            .latch_enable_in (latch[260]),
            .clk_out         (clk  [261]),
            .data_out        (data [261]),
            .scan_select_out (scan [261]),
            .latch_enable_out(latch[261])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_261 (
            .clk_in          (clk  [261]),
            .data_in         (data [261]),
            .scan_select_in  (scan [261]),
            .latch_enable_in (latch[261]),
            .clk_out         (clk  [262]),
            .data_out        (data [262]),
            .scan_select_out (scan [262]),
            .latch_enable_out(latch[262])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_262 (
            .clk_in          (clk  [262]),
            .data_in         (data [262]),
            .scan_select_in  (scan [262]),
            .latch_enable_in (latch[262]),
            .clk_out         (clk  [263]),
            .data_out        (data [263]),
            .scan_select_out (scan [263]),
            .latch_enable_out(latch[263])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_263 (
            .clk_in          (clk  [263]),
            .data_in         (data [263]),
            .scan_select_in  (scan [263]),
            .latch_enable_in (latch[263]),
            .clk_out         (clk  [264]),
            .data_out        (data [264]),
            .scan_select_out (scan [264]),
            .latch_enable_out(latch[264])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_264 (
            .clk_in          (clk  [264]),
            .data_in         (data [264]),
            .scan_select_in  (scan [264]),
            .latch_enable_in (latch[264]),
            .clk_out         (clk  [265]),
            .data_out        (data [265]),
            .scan_select_out (scan [265]),
            .latch_enable_out(latch[265])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_265 (
            .clk_in          (clk  [265]),
            .data_in         (data [265]),
            .scan_select_in  (scan [265]),
            .latch_enable_in (latch[265]),
            .clk_out         (clk  [266]),
            .data_out        (data [266]),
            .scan_select_out (scan [266]),
            .latch_enable_out(latch[266])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_266 (
            .clk_in          (clk  [266]),
            .data_in         (data [266]),
            .scan_select_in  (scan [266]),
            .latch_enable_in (latch[266]),
            .clk_out         (clk  [267]),
            .data_out        (data [267]),
            .scan_select_out (scan [267]),
            .latch_enable_out(latch[267])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_267 (
            .clk_in          (clk  [267]),
            .data_in         (data [267]),
            .scan_select_in  (scan [267]),
            .latch_enable_in (latch[267]),
            .clk_out         (clk  [268]),
            .data_out        (data [268]),
            .scan_select_out (scan [268]),
            .latch_enable_out(latch[268])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_268 (
            .clk_in          (clk  [268]),
            .data_in         (data [268]),
            .scan_select_in  (scan [268]),
            .latch_enable_in (latch[268]),
            .clk_out         (clk  [269]),
            .data_out        (data [269]),
            .scan_select_out (scan [269]),
            .latch_enable_out(latch[269])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_269 (
            .clk_in          (clk  [269]),
            .data_in         (data [269]),
            .scan_select_in  (scan [269]),
            .latch_enable_in (latch[269]),
            .clk_out         (clk  [270]),
            .data_out        (data [270]),
            .scan_select_out (scan [270]),
            .latch_enable_out(latch[270])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_270 (
            .clk_in          (clk  [270]),
            .data_in         (data [270]),
            .scan_select_in  (scan [270]),
            .latch_enable_in (latch[270]),
            .clk_out         (clk  [271]),
            .data_out        (data [271]),
            .scan_select_out (scan [271]),
            .latch_enable_out(latch[271])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_271 (
            .clk_in          (clk  [271]),
            .data_in         (data [271]),
            .scan_select_in  (scan [271]),
            .latch_enable_in (latch[271]),
            .clk_out         (clk  [272]),
            .data_out        (data [272]),
            .scan_select_out (scan [272]),
            .latch_enable_out(latch[272])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_272 (
            .clk_in          (clk  [272]),
            .data_in         (data [272]),
            .scan_select_in  (scan [272]),
            .latch_enable_in (latch[272]),
            .clk_out         (clk  [273]),
            .data_out        (data [273]),
            .scan_select_out (scan [273]),
            .latch_enable_out(latch[273])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_273 (
            .clk_in          (clk  [273]),
            .data_in         (data [273]),
            .scan_select_in  (scan [273]),
            .latch_enable_in (latch[273]),
            .clk_out         (clk  [274]),
            .data_out        (data [274]),
            .scan_select_out (scan [274]),
            .latch_enable_out(latch[274])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_274 (
            .clk_in          (clk  [274]),
            .data_in         (data [274]),
            .scan_select_in  (scan [274]),
            .latch_enable_in (latch[274]),
            .clk_out         (clk  [275]),
            .data_out        (data [275]),
            .scan_select_out (scan [275]),
            .latch_enable_out(latch[275])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_275 (
            .clk_in          (clk  [275]),
            .data_in         (data [275]),
            .scan_select_in  (scan [275]),
            .latch_enable_in (latch[275]),
            .clk_out         (clk  [276]),
            .data_out        (data [276]),
            .scan_select_out (scan [276]),
            .latch_enable_out(latch[276])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_276 (
            .clk_in          (clk  [276]),
            .data_in         (data [276]),
            .scan_select_in  (scan [276]),
            .latch_enable_in (latch[276]),
            .clk_out         (clk  [277]),
            .data_out        (data [277]),
            .scan_select_out (scan [277]),
            .latch_enable_out(latch[277])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_277 (
            .clk_in          (clk  [277]),
            .data_in         (data [277]),
            .scan_select_in  (scan [277]),
            .latch_enable_in (latch[277]),
            .clk_out         (clk  [278]),
            .data_out        (data [278]),
            .scan_select_out (scan [278]),
            .latch_enable_out(latch[278])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_278 (
            .clk_in          (clk  [278]),
            .data_in         (data [278]),
            .scan_select_in  (scan [278]),
            .latch_enable_in (latch[278]),
            .clk_out         (clk  [279]),
            .data_out        (data [279]),
            .scan_select_out (scan [279]),
            .latch_enable_out(latch[279])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_279 (
            .clk_in          (clk  [279]),
            .data_in         (data [279]),
            .scan_select_in  (scan [279]),
            .latch_enable_in (latch[279]),
            .clk_out         (clk  [280]),
            .data_out        (data [280]),
            .scan_select_out (scan [280]),
            .latch_enable_out(latch[280])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_280 (
            .clk_in          (clk  [280]),
            .data_in         (data [280]),
            .scan_select_in  (scan [280]),
            .latch_enable_in (latch[280]),
            .clk_out         (clk  [281]),
            .data_out        (data [281]),
            .scan_select_out (scan [281]),
            .latch_enable_out(latch[281])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_281 (
            .clk_in          (clk  [281]),
            .data_in         (data [281]),
            .scan_select_in  (scan [281]),
            .latch_enable_in (latch[281]),
            .clk_out         (clk  [282]),
            .data_out        (data [282]),
            .scan_select_out (scan [282]),
            .latch_enable_out(latch[282])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_282 (
            .clk_in          (clk  [282]),
            .data_in         (data [282]),
            .scan_select_in  (scan [282]),
            .latch_enable_in (latch[282]),
            .clk_out         (clk  [283]),
            .data_out        (data [283]),
            .scan_select_out (scan [283]),
            .latch_enable_out(latch[283])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_283 (
            .clk_in          (clk  [283]),
            .data_in         (data [283]),
            .scan_select_in  (scan [283]),
            .latch_enable_in (latch[283]),
            .clk_out         (clk  [284]),
            .data_out        (data [284]),
            .scan_select_out (scan [284]),
            .latch_enable_out(latch[284])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_284 (
            .clk_in          (clk  [284]),
            .data_in         (data [284]),
            .scan_select_in  (scan [284]),
            .latch_enable_in (latch[284]),
            .clk_out         (clk  [285]),
            .data_out        (data [285]),
            .scan_select_out (scan [285]),
            .latch_enable_out(latch[285])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_285 (
            .clk_in          (clk  [285]),
            .data_in         (data [285]),
            .scan_select_in  (scan [285]),
            .latch_enable_in (latch[285]),
            .clk_out         (clk  [286]),
            .data_out        (data [286]),
            .scan_select_out (scan [286]),
            .latch_enable_out(latch[286])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_286 (
            .clk_in          (clk  [286]),
            .data_in         (data [286]),
            .scan_select_in  (scan [286]),
            .latch_enable_in (latch[286]),
            .clk_out         (clk  [287]),
            .data_out        (data [287]),
            .scan_select_out (scan [287]),
            .latch_enable_out(latch[287])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_287 (
            .clk_in          (clk  [287]),
            .data_in         (data [287]),
            .scan_select_in  (scan [287]),
            .latch_enable_in (latch[287]),
            .clk_out         (clk  [288]),
            .data_out        (data [288]),
            .scan_select_out (scan [288]),
            .latch_enable_out(latch[288])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_288 (
            .clk_in          (clk  [288]),
            .data_in         (data [288]),
            .scan_select_in  (scan [288]),
            .latch_enable_in (latch[288]),
            .clk_out         (clk  [289]),
            .data_out        (data [289]),
            .scan_select_out (scan [289]),
            .latch_enable_out(latch[289])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_289 (
            .clk_in          (clk  [289]),
            .data_in         (data [289]),
            .scan_select_in  (scan [289]),
            .latch_enable_in (latch[289]),
            .clk_out         (clk  [290]),
            .data_out        (data [290]),
            .scan_select_out (scan [290]),
            .latch_enable_out(latch[290])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_290 (
            .clk_in          (clk  [290]),
            .data_in         (data [290]),
            .scan_select_in  (scan [290]),
            .latch_enable_in (latch[290]),
            .clk_out         (clk  [291]),
            .data_out        (data [291]),
            .scan_select_out (scan [291]),
            .latch_enable_out(latch[291])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_291 (
            .clk_in          (clk  [291]),
            .data_in         (data [291]),
            .scan_select_in  (scan [291]),
            .latch_enable_in (latch[291]),
            .clk_out         (clk  [292]),
            .data_out        (data [292]),
            .scan_select_out (scan [292]),
            .latch_enable_out(latch[292])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_292 (
            .clk_in          (clk  [292]),
            .data_in         (data [292]),
            .scan_select_in  (scan [292]),
            .latch_enable_in (latch[292]),
            .clk_out         (clk  [293]),
            .data_out        (data [293]),
            .scan_select_out (scan [293]),
            .latch_enable_out(latch[293])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_293 (
            .clk_in          (clk  [293]),
            .data_in         (data [293]),
            .scan_select_in  (scan [293]),
            .latch_enable_in (latch[293]),
            .clk_out         (clk  [294]),
            .data_out        (data [294]),
            .scan_select_out (scan [294]),
            .latch_enable_out(latch[294])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_294 (
            .clk_in          (clk  [294]),
            .data_in         (data [294]),
            .scan_select_in  (scan [294]),
            .latch_enable_in (latch[294]),
            .clk_out         (clk  [295]),
            .data_out        (data [295]),
            .scan_select_out (scan [295]),
            .latch_enable_out(latch[295])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_295 (
            .clk_in          (clk  [295]),
            .data_in         (data [295]),
            .scan_select_in  (scan [295]),
            .latch_enable_in (latch[295]),
            .clk_out         (clk  [296]),
            .data_out        (data [296]),
            .scan_select_out (scan [296]),
            .latch_enable_out(latch[296])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_296 (
            .clk_in          (clk  [296]),
            .data_in         (data [296]),
            .scan_select_in  (scan [296]),
            .latch_enable_in (latch[296]),
            .clk_out         (clk  [297]),
            .data_out        (data [297]),
            .scan_select_out (scan [297]),
            .latch_enable_out(latch[297])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_297 (
            .clk_in          (clk  [297]),
            .data_in         (data [297]),
            .scan_select_in  (scan [297]),
            .latch_enable_in (latch[297]),
            .clk_out         (clk  [298]),
            .data_out        (data [298]),
            .scan_select_out (scan [298]),
            .latch_enable_out(latch[298])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_298 (
            .clk_in          (clk  [298]),
            .data_in         (data [298]),
            .scan_select_in  (scan [298]),
            .latch_enable_in (latch[298]),
            .clk_out         (clk  [299]),
            .data_out        (data [299]),
            .scan_select_out (scan [299]),
            .latch_enable_out(latch[299])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_299 (
            .clk_in          (clk  [299]),
            .data_in         (data [299]),
            .scan_select_in  (scan [299]),
            .latch_enable_in (latch[299]),
            .clk_out         (clk  [300]),
            .data_out        (data [300]),
            .scan_select_out (scan [300]),
            .latch_enable_out(latch[300])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_300 (
            .clk_in          (clk  [300]),
            .data_in         (data [300]),
            .scan_select_in  (scan [300]),
            .latch_enable_in (latch[300]),
            .clk_out         (clk  [301]),
            .data_out        (data [301]),
            .scan_select_out (scan [301]),
            .latch_enable_out(latch[301])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_301 (
            .clk_in          (clk  [301]),
            .data_in         (data [301]),
            .scan_select_in  (scan [301]),
            .latch_enable_in (latch[301]),
            .clk_out         (clk  [302]),
            .data_out        (data [302]),
            .scan_select_out (scan [302]),
            .latch_enable_out(latch[302])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_302 (
            .clk_in          (clk  [302]),
            .data_in         (data [302]),
            .scan_select_in  (scan [302]),
            .latch_enable_in (latch[302]),
            .clk_out         (clk  [303]),
            .data_out        (data [303]),
            .scan_select_out (scan [303]),
            .latch_enable_out(latch[303])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_303 (
            .clk_in          (clk  [303]),
            .data_in         (data [303]),
            .scan_select_in  (scan [303]),
            .latch_enable_in (latch[303]),
            .clk_out         (clk  [304]),
            .data_out        (data [304]),
            .scan_select_out (scan [304]),
            .latch_enable_out(latch[304])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_304 (
            .clk_in          (clk  [304]),
            .data_in         (data [304]),
            .scan_select_in  (scan [304]),
            .latch_enable_in (latch[304]),
            .clk_out         (clk  [305]),
            .data_out        (data [305]),
            .scan_select_out (scan [305]),
            .latch_enable_out(latch[305])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_305 (
            .clk_in          (clk  [305]),
            .data_in         (data [305]),
            .scan_select_in  (scan [305]),
            .latch_enable_in (latch[305]),
            .clk_out         (clk  [306]),
            .data_out        (data [306]),
            .scan_select_out (scan [306]),
            .latch_enable_out(latch[306])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_306 (
            .clk_in          (clk  [306]),
            .data_in         (data [306]),
            .scan_select_in  (scan [306]),
            .latch_enable_in (latch[306]),
            .clk_out         (clk  [307]),
            .data_out        (data [307]),
            .scan_select_out (scan [307]),
            .latch_enable_out(latch[307])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_307 (
            .clk_in          (clk  [307]),
            .data_in         (data [307]),
            .scan_select_in  (scan [307]),
            .latch_enable_in (latch[307]),
            .clk_out         (clk  [308]),
            .data_out        (data [308]),
            .scan_select_out (scan [308]),
            .latch_enable_out(latch[308])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_308 (
            .clk_in          (clk  [308]),
            .data_in         (data [308]),
            .scan_select_in  (scan [308]),
            .latch_enable_in (latch[308]),
            .clk_out         (clk  [309]),
            .data_out        (data [309]),
            .scan_select_out (scan [309]),
            .latch_enable_out(latch[309])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_309 (
            .clk_in          (clk  [309]),
            .data_in         (data [309]),
            .scan_select_in  (scan [309]),
            .latch_enable_in (latch[309]),
            .clk_out         (clk  [310]),
            .data_out        (data [310]),
            .scan_select_out (scan [310]),
            .latch_enable_out(latch[310])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_310 (
            .clk_in          (clk  [310]),
            .data_in         (data [310]),
            .scan_select_in  (scan [310]),
            .latch_enable_in (latch[310]),
            .clk_out         (clk  [311]),
            .data_out        (data [311]),
            .scan_select_out (scan [311]),
            .latch_enable_out(latch[311])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_311 (
            .clk_in          (clk  [311]),
            .data_in         (data [311]),
            .scan_select_in  (scan [311]),
            .latch_enable_in (latch[311]),
            .clk_out         (clk  [312]),
            .data_out        (data [312]),
            .scan_select_out (scan [312]),
            .latch_enable_out(latch[312])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_312 (
            .clk_in          (clk  [312]),
            .data_in         (data [312]),
            .scan_select_in  (scan [312]),
            .latch_enable_in (latch[312]),
            .clk_out         (clk  [313]),
            .data_out        (data [313]),
            .scan_select_out (scan [313]),
            .latch_enable_out(latch[313])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_313 (
            .clk_in          (clk  [313]),
            .data_in         (data [313]),
            .scan_select_in  (scan [313]),
            .latch_enable_in (latch[313]),
            .clk_out         (clk  [314]),
            .data_out        (data [314]),
            .scan_select_out (scan [314]),
            .latch_enable_out(latch[314])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_314 (
            .clk_in          (clk  [314]),
            .data_in         (data [314]),
            .scan_select_in  (scan [314]),
            .latch_enable_in (latch[314]),
            .clk_out         (clk  [315]),
            .data_out        (data [315]),
            .scan_select_out (scan [315]),
            .latch_enable_out(latch[315])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_315 (
            .clk_in          (clk  [315]),
            .data_in         (data [315]),
            .scan_select_in  (scan [315]),
            .latch_enable_in (latch[315]),
            .clk_out         (clk  [316]),
            .data_out        (data [316]),
            .scan_select_out (scan [316]),
            .latch_enable_out(latch[316])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_316 (
            .clk_in          (clk  [316]),
            .data_in         (data [316]),
            .scan_select_in  (scan [316]),
            .latch_enable_in (latch[316]),
            .clk_out         (clk  [317]),
            .data_out        (data [317]),
            .scan_select_out (scan [317]),
            .latch_enable_out(latch[317])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_317 (
            .clk_in          (clk  [317]),
            .data_in         (data [317]),
            .scan_select_in  (scan [317]),
            .latch_enable_in (latch[317]),
            .clk_out         (clk  [318]),
            .data_out        (data [318]),
            .scan_select_out (scan [318]),
            .latch_enable_out(latch[318])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_318 (
            .clk_in          (clk  [318]),
            .data_in         (data [318]),
            .scan_select_in  (scan [318]),
            .latch_enable_in (latch[318]),
            .clk_out         (clk  [319]),
            .data_out        (data [319]),
            .scan_select_out (scan [319]),
            .latch_enable_out(latch[319])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_319 (
            .clk_in          (clk  [319]),
            .data_in         (data [319]),
            .scan_select_in  (scan [319]),
            .latch_enable_in (latch[319]),
            .clk_out         (clk  [320]),
            .data_out        (data [320]),
            .scan_select_out (scan [320]),
            .latch_enable_out(latch[320])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_320 (
            .clk_in          (clk  [320]),
            .data_in         (data [320]),
            .scan_select_in  (scan [320]),
            .latch_enable_in (latch[320]),
            .clk_out         (clk  [321]),
            .data_out        (data [321]),
            .scan_select_out (scan [321]),
            .latch_enable_out(latch[321])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_321 (
            .clk_in          (clk  [321]),
            .data_in         (data [321]),
            .scan_select_in  (scan [321]),
            .latch_enable_in (latch[321]),
            .clk_out         (clk  [322]),
            .data_out        (data [322]),
            .scan_select_out (scan [322]),
            .latch_enable_out(latch[322])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_322 (
            .clk_in          (clk  [322]),
            .data_in         (data [322]),
            .scan_select_in  (scan [322]),
            .latch_enable_in (latch[322]),
            .clk_out         (clk  [323]),
            .data_out        (data [323]),
            .scan_select_out (scan [323]),
            .latch_enable_out(latch[323])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_323 (
            .clk_in          (clk  [323]),
            .data_in         (data [323]),
            .scan_select_in  (scan [323]),
            .latch_enable_in (latch[323]),
            .clk_out         (clk  [324]),
            .data_out        (data [324]),
            .scan_select_out (scan [324]),
            .latch_enable_out(latch[324])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_324 (
            .clk_in          (clk  [324]),
            .data_in         (data [324]),
            .scan_select_in  (scan [324]),
            .latch_enable_in (latch[324]),
            .clk_out         (clk  [325]),
            .data_out        (data [325]),
            .scan_select_out (scan [325]),
            .latch_enable_out(latch[325])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_325 (
            .clk_in          (clk  [325]),
            .data_in         (data [325]),
            .scan_select_in  (scan [325]),
            .latch_enable_in (latch[325]),
            .clk_out         (clk  [326]),
            .data_out        (data [326]),
            .scan_select_out (scan [326]),
            .latch_enable_out(latch[326])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_326 (
            .clk_in          (clk  [326]),
            .data_in         (data [326]),
            .scan_select_in  (scan [326]),
            .latch_enable_in (latch[326]),
            .clk_out         (clk  [327]),
            .data_out        (data [327]),
            .scan_select_out (scan [327]),
            .latch_enable_out(latch[327])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_327 (
            .clk_in          (clk  [327]),
            .data_in         (data [327]),
            .scan_select_in  (scan [327]),
            .latch_enable_in (latch[327]),
            .clk_out         (clk  [328]),
            .data_out        (data [328]),
            .scan_select_out (scan [328]),
            .latch_enable_out(latch[328])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_328 (
            .clk_in          (clk  [328]),
            .data_in         (data [328]),
            .scan_select_in  (scan [328]),
            .latch_enable_in (latch[328]),
            .clk_out         (clk  [329]),
            .data_out        (data [329]),
            .scan_select_out (scan [329]),
            .latch_enable_out(latch[329])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_329 (
            .clk_in          (clk  [329]),
            .data_in         (data [329]),
            .scan_select_in  (scan [329]),
            .latch_enable_in (latch[329]),
            .clk_out         (clk  [330]),
            .data_out        (data [330]),
            .scan_select_out (scan [330]),
            .latch_enable_out(latch[330])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_330 (
            .clk_in          (clk  [330]),
            .data_in         (data [330]),
            .scan_select_in  (scan [330]),
            .latch_enable_in (latch[330]),
            .clk_out         (clk  [331]),
            .data_out        (data [331]),
            .scan_select_out (scan [331]),
            .latch_enable_out(latch[331])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_331 (
            .clk_in          (clk  [331]),
            .data_in         (data [331]),
            .scan_select_in  (scan [331]),
            .latch_enable_in (latch[331]),
            .clk_out         (clk  [332]),
            .data_out        (data [332]),
            .scan_select_out (scan [332]),
            .latch_enable_out(latch[332])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_332 (
            .clk_in          (clk  [332]),
            .data_in         (data [332]),
            .scan_select_in  (scan [332]),
            .latch_enable_in (latch[332]),
            .clk_out         (clk  [333]),
            .data_out        (data [333]),
            .scan_select_out (scan [333]),
            .latch_enable_out(latch[333])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_333 (
            .clk_in          (clk  [333]),
            .data_in         (data [333]),
            .scan_select_in  (scan [333]),
            .latch_enable_in (latch[333]),
            .clk_out         (clk  [334]),
            .data_out        (data [334]),
            .scan_select_out (scan [334]),
            .latch_enable_out(latch[334])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_334 (
            .clk_in          (clk  [334]),
            .data_in         (data [334]),
            .scan_select_in  (scan [334]),
            .latch_enable_in (latch[334]),
            .clk_out         (clk  [335]),
            .data_out        (data [335]),
            .scan_select_out (scan [335]),
            .latch_enable_out(latch[335])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_335 (
            .clk_in          (clk  [335]),
            .data_in         (data [335]),
            .scan_select_in  (scan [335]),
            .latch_enable_in (latch[335]),
            .clk_out         (clk  [336]),
            .data_out        (data [336]),
            .scan_select_out (scan [336]),
            .latch_enable_out(latch[336])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_336 (
            .clk_in          (clk  [336]),
            .data_in         (data [336]),
            .scan_select_in  (scan [336]),
            .latch_enable_in (latch[336]),
            .clk_out         (clk  [337]),
            .data_out        (data [337]),
            .scan_select_out (scan [337]),
            .latch_enable_out(latch[337])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_337 (
            .clk_in          (clk  [337]),
            .data_in         (data [337]),
            .scan_select_in  (scan [337]),
            .latch_enable_in (latch[337]),
            .clk_out         (clk  [338]),
            .data_out        (data [338]),
            .scan_select_out (scan [338]),
            .latch_enable_out(latch[338])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_338 (
            .clk_in          (clk  [338]),
            .data_in         (data [338]),
            .scan_select_in  (scan [338]),
            .latch_enable_in (latch[338]),
            .clk_out         (clk  [339]),
            .data_out        (data [339]),
            .scan_select_out (scan [339]),
            .latch_enable_out(latch[339])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_339 (
            .clk_in          (clk  [339]),
            .data_in         (data [339]),
            .scan_select_in  (scan [339]),
            .latch_enable_in (latch[339]),
            .clk_out         (clk  [340]),
            .data_out        (data [340]),
            .scan_select_out (scan [340]),
            .latch_enable_out(latch[340])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_340 (
            .clk_in          (clk  [340]),
            .data_in         (data [340]),
            .scan_select_in  (scan [340]),
            .latch_enable_in (latch[340]),
            .clk_out         (clk  [341]),
            .data_out        (data [341]),
            .scan_select_out (scan [341]),
            .latch_enable_out(latch[341])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_341 (
            .clk_in          (clk  [341]),
            .data_in         (data [341]),
            .scan_select_in  (scan [341]),
            .latch_enable_in (latch[341]),
            .clk_out         (clk  [342]),
            .data_out        (data [342]),
            .scan_select_out (scan [342]),
            .latch_enable_out(latch[342])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_342 (
            .clk_in          (clk  [342]),
            .data_in         (data [342]),
            .scan_select_in  (scan [342]),
            .latch_enable_in (latch[342]),
            .clk_out         (clk  [343]),
            .data_out        (data [343]),
            .scan_select_out (scan [343]),
            .latch_enable_out(latch[343])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_343 (
            .clk_in          (clk  [343]),
            .data_in         (data [343]),
            .scan_select_in  (scan [343]),
            .latch_enable_in (latch[343]),
            .clk_out         (clk  [344]),
            .data_out        (data [344]),
            .scan_select_out (scan [344]),
            .latch_enable_out(latch[344])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_344 (
            .clk_in          (clk  [344]),
            .data_in         (data [344]),
            .scan_select_in  (scan [344]),
            .latch_enable_in (latch[344]),
            .clk_out         (clk  [345]),
            .data_out        (data [345]),
            .scan_select_out (scan [345]),
            .latch_enable_out(latch[345])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_345 (
            .clk_in          (clk  [345]),
            .data_in         (data [345]),
            .scan_select_in  (scan [345]),
            .latch_enable_in (latch[345]),
            .clk_out         (clk  [346]),
            .data_out        (data [346]),
            .scan_select_out (scan [346]),
            .latch_enable_out(latch[346])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_346 (
            .clk_in          (clk  [346]),
            .data_in         (data [346]),
            .scan_select_in  (scan [346]),
            .latch_enable_in (latch[346]),
            .clk_out         (clk  [347]),
            .data_out        (data [347]),
            .scan_select_out (scan [347]),
            .latch_enable_out(latch[347])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_347 (
            .clk_in          (clk  [347]),
            .data_in         (data [347]),
            .scan_select_in  (scan [347]),
            .latch_enable_in (latch[347]),
            .clk_out         (clk  [348]),
            .data_out        (data [348]),
            .scan_select_out (scan [348]),
            .latch_enable_out(latch[348])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_348 (
            .clk_in          (clk  [348]),
            .data_in         (data [348]),
            .scan_select_in  (scan [348]),
            .latch_enable_in (latch[348]),
            .clk_out         (clk  [349]),
            .data_out        (data [349]),
            .scan_select_out (scan [349]),
            .latch_enable_out(latch[349])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_349 (
            .clk_in          (clk  [349]),
            .data_in         (data [349]),
            .scan_select_in  (scan [349]),
            .latch_enable_in (latch[349]),
            .clk_out         (clk  [350]),
            .data_out        (data [350]),
            .scan_select_out (scan [350]),
            .latch_enable_out(latch[350])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_350 (
            .clk_in          (clk  [350]),
            .data_in         (data [350]),
            .scan_select_in  (scan [350]),
            .latch_enable_in (latch[350]),
            .clk_out         (clk  [351]),
            .data_out        (data [351]),
            .scan_select_out (scan [351]),
            .latch_enable_out(latch[351])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_351 (
            .clk_in          (clk  [351]),
            .data_in         (data [351]),
            .scan_select_in  (scan [351]),
            .latch_enable_in (latch[351]),
            .clk_out         (clk  [352]),
            .data_out        (data [352]),
            .scan_select_out (scan [352]),
            .latch_enable_out(latch[352])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_352 (
            .clk_in          (clk  [352]),
            .data_in         (data [352]),
            .scan_select_in  (scan [352]),
            .latch_enable_in (latch[352]),
            .clk_out         (clk  [353]),
            .data_out        (data [353]),
            .scan_select_out (scan [353]),
            .latch_enable_out(latch[353])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_353 (
            .clk_in          (clk  [353]),
            .data_in         (data [353]),
            .scan_select_in  (scan [353]),
            .latch_enable_in (latch[353]),
            .clk_out         (clk  [354]),
            .data_out        (data [354]),
            .scan_select_out (scan [354]),
            .latch_enable_out(latch[354])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_354 (
            .clk_in          (clk  [354]),
            .data_in         (data [354]),
            .scan_select_in  (scan [354]),
            .latch_enable_in (latch[354]),
            .clk_out         (clk  [355]),
            .data_out        (data [355]),
            .scan_select_out (scan [355]),
            .latch_enable_out(latch[355])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_355 (
            .clk_in          (clk  [355]),
            .data_in         (data [355]),
            .scan_select_in  (scan [355]),
            .latch_enable_in (latch[355]),
            .clk_out         (clk  [356]),
            .data_out        (data [356]),
            .scan_select_out (scan [356]),
            .latch_enable_out(latch[356])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_356 (
            .clk_in          (clk  [356]),
            .data_in         (data [356]),
            .scan_select_in  (scan [356]),
            .latch_enable_in (latch[356]),
            .clk_out         (clk  [357]),
            .data_out        (data [357]),
            .scan_select_out (scan [357]),
            .latch_enable_out(latch[357])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_357 (
            .clk_in          (clk  [357]),
            .data_in         (data [357]),
            .scan_select_in  (scan [357]),
            .latch_enable_in (latch[357]),
            .clk_out         (clk  [358]),
            .data_out        (data [358]),
            .scan_select_out (scan [358]),
            .latch_enable_out(latch[358])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_358 (
            .clk_in          (clk  [358]),
            .data_in         (data [358]),
            .scan_select_in  (scan [358]),
            .latch_enable_in (latch[358]),
            .clk_out         (clk  [359]),
            .data_out        (data [359]),
            .scan_select_out (scan [359]),
            .latch_enable_out(latch[359])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_359 (
            .clk_in          (clk  [359]),
            .data_in         (data [359]),
            .scan_select_in  (scan [359]),
            .latch_enable_in (latch[359]),
            .clk_out         (clk  [360]),
            .data_out        (data [360]),
            .scan_select_out (scan [360]),
            .latch_enable_out(latch[360])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_360 (
            .clk_in          (clk  [360]),
            .data_in         (data [360]),
            .scan_select_in  (scan [360]),
            .latch_enable_in (latch[360]),
            .clk_out         (clk  [361]),
            .data_out        (data [361]),
            .scan_select_out (scan [361]),
            .latch_enable_out(latch[361])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_361 (
            .clk_in          (clk  [361]),
            .data_in         (data [361]),
            .scan_select_in  (scan [361]),
            .latch_enable_in (latch[361]),
            .clk_out         (clk  [362]),
            .data_out        (data [362]),
            .scan_select_out (scan [362]),
            .latch_enable_out(latch[362])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_362 (
            .clk_in          (clk  [362]),
            .data_in         (data [362]),
            .scan_select_in  (scan [362]),
            .latch_enable_in (latch[362]),
            .clk_out         (clk  [363]),
            .data_out        (data [363]),
            .scan_select_out (scan [363]),
            .latch_enable_out(latch[363])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_363 (
            .clk_in          (clk  [363]),
            .data_in         (data [363]),
            .scan_select_in  (scan [363]),
            .latch_enable_in (latch[363]),
            .clk_out         (clk  [364]),
            .data_out        (data [364]),
            .scan_select_out (scan [364]),
            .latch_enable_out(latch[364])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_364 (
            .clk_in          (clk  [364]),
            .data_in         (data [364]),
            .scan_select_in  (scan [364]),
            .latch_enable_in (latch[364]),
            .clk_out         (clk  [365]),
            .data_out        (data [365]),
            .scan_select_out (scan [365]),
            .latch_enable_out(latch[365])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_365 (
            .clk_in          (clk  [365]),
            .data_in         (data [365]),
            .scan_select_in  (scan [365]),
            .latch_enable_in (latch[365]),
            .clk_out         (clk  [366]),
            .data_out        (data [366]),
            .scan_select_out (scan [366]),
            .latch_enable_out(latch[366])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_366 (
            .clk_in          (clk  [366]),
            .data_in         (data [366]),
            .scan_select_in  (scan [366]),
            .latch_enable_in (latch[366]),
            .clk_out         (clk  [367]),
            .data_out        (data [367]),
            .scan_select_out (scan [367]),
            .latch_enable_out(latch[367])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_367 (
            .clk_in          (clk  [367]),
            .data_in         (data [367]),
            .scan_select_in  (scan [367]),
            .latch_enable_in (latch[367]),
            .clk_out         (clk  [368]),
            .data_out        (data [368]),
            .scan_select_out (scan [368]),
            .latch_enable_out(latch[368])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_368 (
            .clk_in          (clk  [368]),
            .data_in         (data [368]),
            .scan_select_in  (scan [368]),
            .latch_enable_in (latch[368]),
            .clk_out         (clk  [369]),
            .data_out        (data [369]),
            .scan_select_out (scan [369]),
            .latch_enable_out(latch[369])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_369 (
            .clk_in          (clk  [369]),
            .data_in         (data [369]),
            .scan_select_in  (scan [369]),
            .latch_enable_in (latch[369]),
            .clk_out         (clk  [370]),
            .data_out        (data [370]),
            .scan_select_out (scan [370]),
            .latch_enable_out(latch[370])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_370 (
            .clk_in          (clk  [370]),
            .data_in         (data [370]),
            .scan_select_in  (scan [370]),
            .latch_enable_in (latch[370]),
            .clk_out         (clk  [371]),
            .data_out        (data [371]),
            .scan_select_out (scan [371]),
            .latch_enable_out(latch[371])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_371 (
            .clk_in          (clk  [371]),
            .data_in         (data [371]),
            .scan_select_in  (scan [371]),
            .latch_enable_in (latch[371]),
            .clk_out         (clk  [372]),
            .data_out        (data [372]),
            .scan_select_out (scan [372]),
            .latch_enable_out(latch[372])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_372 (
            .clk_in          (clk  [372]),
            .data_in         (data [372]),
            .scan_select_in  (scan [372]),
            .latch_enable_in (latch[372]),
            .clk_out         (clk  [373]),
            .data_out        (data [373]),
            .scan_select_out (scan [373]),
            .latch_enable_out(latch[373])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_373 (
            .clk_in          (clk  [373]),
            .data_in         (data [373]),
            .scan_select_in  (scan [373]),
            .latch_enable_in (latch[373]),
            .clk_out         (clk  [374]),
            .data_out        (data [374]),
            .scan_select_out (scan [374]),
            .latch_enable_out(latch[374])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_374 (
            .clk_in          (clk  [374]),
            .data_in         (data [374]),
            .scan_select_in  (scan [374]),
            .latch_enable_in (latch[374]),
            .clk_out         (clk  [375]),
            .data_out        (data [375]),
            .scan_select_out (scan [375]),
            .latch_enable_out(latch[375])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_375 (
            .clk_in          (clk  [375]),
            .data_in         (data [375]),
            .scan_select_in  (scan [375]),
            .latch_enable_in (latch[375]),
            .clk_out         (clk  [376]),
            .data_out        (data [376]),
            .scan_select_out (scan [376]),
            .latch_enable_out(latch[376])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_376 (
            .clk_in          (clk  [376]),
            .data_in         (data [376]),
            .scan_select_in  (scan [376]),
            .latch_enable_in (latch[376]),
            .clk_out         (clk  [377]),
            .data_out        (data [377]),
            .scan_select_out (scan [377]),
            .latch_enable_out(latch[377])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_377 (
            .clk_in          (clk  [377]),
            .data_in         (data [377]),
            .scan_select_in  (scan [377]),
            .latch_enable_in (latch[377]),
            .clk_out         (clk  [378]),
            .data_out        (data [378]),
            .scan_select_out (scan [378]),
            .latch_enable_out(latch[378])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_378 (
            .clk_in          (clk  [378]),
            .data_in         (data [378]),
            .scan_select_in  (scan [378]),
            .latch_enable_in (latch[378]),
            .clk_out         (clk  [379]),
            .data_out        (data [379]),
            .scan_select_out (scan [379]),
            .latch_enable_out(latch[379])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_379 (
            .clk_in          (clk  [379]),
            .data_in         (data [379]),
            .scan_select_in  (scan [379]),
            .latch_enable_in (latch[379]),
            .clk_out         (clk  [380]),
            .data_out        (data [380]),
            .scan_select_out (scan [380]),
            .latch_enable_out(latch[380])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_380 (
            .clk_in          (clk  [380]),
            .data_in         (data [380]),
            .scan_select_in  (scan [380]),
            .latch_enable_in (latch[380]),
            .clk_out         (clk  [381]),
            .data_out        (data [381]),
            .scan_select_out (scan [381]),
            .latch_enable_out(latch[381])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_381 (
            .clk_in          (clk  [381]),
            .data_in         (data [381]),
            .scan_select_in  (scan [381]),
            .latch_enable_in (latch[381]),
            .clk_out         (clk  [382]),
            .data_out        (data [382]),
            .scan_select_out (scan [382]),
            .latch_enable_out(latch[382])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_382 (
            .clk_in          (clk  [382]),
            .data_in         (data [382]),
            .scan_select_in  (scan [382]),
            .latch_enable_in (latch[382]),
            .clk_out         (clk  [383]),
            .data_out        (data [383]),
            .scan_select_out (scan [383]),
            .latch_enable_out(latch[383])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_383 (
            .clk_in          (clk  [383]),
            .data_in         (data [383]),
            .scan_select_in  (scan [383]),
            .latch_enable_in (latch[383]),
            .clk_out         (clk  [384]),
            .data_out        (data [384]),
            .scan_select_out (scan [384]),
            .latch_enable_out(latch[384])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_384 (
            .clk_in          (clk  [384]),
            .data_in         (data [384]),
            .scan_select_in  (scan [384]),
            .latch_enable_in (latch[384]),
            .clk_out         (clk  [385]),
            .data_out        (data [385]),
            .scan_select_out (scan [385]),
            .latch_enable_out(latch[385])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_385 (
            .clk_in          (clk  [385]),
            .data_in         (data [385]),
            .scan_select_in  (scan [385]),
            .latch_enable_in (latch[385]),
            .clk_out         (clk  [386]),
            .data_out        (data [386]),
            .scan_select_out (scan [386]),
            .latch_enable_out(latch[386])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_386 (
            .clk_in          (clk  [386]),
            .data_in         (data [386]),
            .scan_select_in  (scan [386]),
            .latch_enable_in (latch[386]),
            .clk_out         (clk  [387]),
            .data_out        (data [387]),
            .scan_select_out (scan [387]),
            .latch_enable_out(latch[387])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_387 (
            .clk_in          (clk  [387]),
            .data_in         (data [387]),
            .scan_select_in  (scan [387]),
            .latch_enable_in (latch[387]),
            .clk_out         (clk  [388]),
            .data_out        (data [388]),
            .scan_select_out (scan [388]),
            .latch_enable_out(latch[388])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_388 (
            .clk_in          (clk  [388]),
            .data_in         (data [388]),
            .scan_select_in  (scan [388]),
            .latch_enable_in (latch[388]),
            .clk_out         (clk  [389]),
            .data_out        (data [389]),
            .scan_select_out (scan [389]),
            .latch_enable_out(latch[389])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_389 (
            .clk_in          (clk  [389]),
            .data_in         (data [389]),
            .scan_select_in  (scan [389]),
            .latch_enable_in (latch[389]),
            .clk_out         (clk  [390]),
            .data_out        (data [390]),
            .scan_select_out (scan [390]),
            .latch_enable_out(latch[390])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_390 (
            .clk_in          (clk  [390]),
            .data_in         (data [390]),
            .scan_select_in  (scan [390]),
            .latch_enable_in (latch[390]),
            .clk_out         (clk  [391]),
            .data_out        (data [391]),
            .scan_select_out (scan [391]),
            .latch_enable_out(latch[391])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_391 (
            .clk_in          (clk  [391]),
            .data_in         (data [391]),
            .scan_select_in  (scan [391]),
            .latch_enable_in (latch[391]),
            .clk_out         (clk  [392]),
            .data_out        (data [392]),
            .scan_select_out (scan [392]),
            .latch_enable_out(latch[392])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_392 (
            .clk_in          (clk  [392]),
            .data_in         (data [392]),
            .scan_select_in  (scan [392]),
            .latch_enable_in (latch[392]),
            .clk_out         (clk  [393]),
            .data_out        (data [393]),
            .scan_select_out (scan [393]),
            .latch_enable_out(latch[393])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_393 (
            .clk_in          (clk  [393]),
            .data_in         (data [393]),
            .scan_select_in  (scan [393]),
            .latch_enable_in (latch[393]),
            .clk_out         (clk  [394]),
            .data_out        (data [394]),
            .scan_select_out (scan [394]),
            .latch_enable_out(latch[394])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_394 (
            .clk_in          (clk  [394]),
            .data_in         (data [394]),
            .scan_select_in  (scan [394]),
            .latch_enable_in (latch[394]),
            .clk_out         (clk  [395]),
            .data_out        (data [395]),
            .scan_select_out (scan [395]),
            .latch_enable_out(latch[395])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_395 (
            .clk_in          (clk  [395]),
            .data_in         (data [395]),
            .scan_select_in  (scan [395]),
            .latch_enable_in (latch[395]),
            .clk_out         (clk  [396]),
            .data_out        (data [396]),
            .scan_select_out (scan [396]),
            .latch_enable_out(latch[396])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_396 (
            .clk_in          (clk  [396]),
            .data_in         (data [396]),
            .scan_select_in  (scan [396]),
            .latch_enable_in (latch[396]),
            .clk_out         (clk  [397]),
            .data_out        (data [397]),
            .scan_select_out (scan [397]),
            .latch_enable_out(latch[397])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_397 (
            .clk_in          (clk  [397]),
            .data_in         (data [397]),
            .scan_select_in  (scan [397]),
            .latch_enable_in (latch[397]),
            .clk_out         (clk  [398]),
            .data_out        (data [398]),
            .scan_select_out (scan [398]),
            .latch_enable_out(latch[398])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_398 (
            .clk_in          (clk  [398]),
            .data_in         (data [398]),
            .scan_select_in  (scan [398]),
            .latch_enable_in (latch[398]),
            .clk_out         (clk  [399]),
            .data_out        (data [399]),
            .scan_select_out (scan [399]),
            .latch_enable_out(latch[399])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_399 (
            .clk_in          (clk  [399]),
            .data_in         (data [399]),
            .scan_select_in  (scan [399]),
            .latch_enable_in (latch[399]),
            .clk_out         (clk  [400]),
            .data_out        (data [400]),
            .scan_select_out (scan [400]),
            .latch_enable_out(latch[400])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_400 (
            .clk_in          (clk  [400]),
            .data_in         (data [400]),
            .scan_select_in  (scan [400]),
            .latch_enable_in (latch[400]),
            .clk_out         (clk  [401]),
            .data_out        (data [401]),
            .scan_select_out (scan [401]),
            .latch_enable_out(latch[401])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_401 (
            .clk_in          (clk  [401]),
            .data_in         (data [401]),
            .scan_select_in  (scan [401]),
            .latch_enable_in (latch[401]),
            .clk_out         (clk  [402]),
            .data_out        (data [402]),
            .scan_select_out (scan [402]),
            .latch_enable_out(latch[402])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_402 (
            .clk_in          (clk  [402]),
            .data_in         (data [402]),
            .scan_select_in  (scan [402]),
            .latch_enable_in (latch[402]),
            .clk_out         (clk  [403]),
            .data_out        (data [403]),
            .scan_select_out (scan [403]),
            .latch_enable_out(latch[403])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_403 (
            .clk_in          (clk  [403]),
            .data_in         (data [403]),
            .scan_select_in  (scan [403]),
            .latch_enable_in (latch[403]),
            .clk_out         (clk  [404]),
            .data_out        (data [404]),
            .scan_select_out (scan [404]),
            .latch_enable_out(latch[404])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_404 (
            .clk_in          (clk  [404]),
            .data_in         (data [404]),
            .scan_select_in  (scan [404]),
            .latch_enable_in (latch[404]),
            .clk_out         (clk  [405]),
            .data_out        (data [405]),
            .scan_select_out (scan [405]),
            .latch_enable_out(latch[405])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_405 (
            .clk_in          (clk  [405]),
            .data_in         (data [405]),
            .scan_select_in  (scan [405]),
            .latch_enable_in (latch[405]),
            .clk_out         (clk  [406]),
            .data_out        (data [406]),
            .scan_select_out (scan [406]),
            .latch_enable_out(latch[406])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_406 (
            .clk_in          (clk  [406]),
            .data_in         (data [406]),
            .scan_select_in  (scan [406]),
            .latch_enable_in (latch[406]),
            .clk_out         (clk  [407]),
            .data_out        (data [407]),
            .scan_select_out (scan [407]),
            .latch_enable_out(latch[407])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_407 (
            .clk_in          (clk  [407]),
            .data_in         (data [407]),
            .scan_select_in  (scan [407]),
            .latch_enable_in (latch[407]),
            .clk_out         (clk  [408]),
            .data_out        (data [408]),
            .scan_select_out (scan [408]),
            .latch_enable_out(latch[408])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_408 (
            .clk_in          (clk  [408]),
            .data_in         (data [408]),
            .scan_select_in  (scan [408]),
            .latch_enable_in (latch[408]),
            .clk_out         (clk  [409]),
            .data_out        (data [409]),
            .scan_select_out (scan [409]),
            .latch_enable_out(latch[409])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_409 (
            .clk_in          (clk  [409]),
            .data_in         (data [409]),
            .scan_select_in  (scan [409]),
            .latch_enable_in (latch[409]),
            .clk_out         (clk  [410]),
            .data_out        (data [410]),
            .scan_select_out (scan [410]),
            .latch_enable_out(latch[410])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_410 (
            .clk_in          (clk  [410]),
            .data_in         (data [410]),
            .scan_select_in  (scan [410]),
            .latch_enable_in (latch[410]),
            .clk_out         (clk  [411]),
            .data_out        (data [411]),
            .scan_select_out (scan [411]),
            .latch_enable_out(latch[411])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_411 (
            .clk_in          (clk  [411]),
            .data_in         (data [411]),
            .scan_select_in  (scan [411]),
            .latch_enable_in (latch[411]),
            .clk_out         (clk  [412]),
            .data_out        (data [412]),
            .scan_select_out (scan [412]),
            .latch_enable_out(latch[412])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_412 (
            .clk_in          (clk  [412]),
            .data_in         (data [412]),
            .scan_select_in  (scan [412]),
            .latch_enable_in (latch[412]),
            .clk_out         (clk  [413]),
            .data_out        (data [413]),
            .scan_select_out (scan [413]),
            .latch_enable_out(latch[413])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_413 (
            .clk_in          (clk  [413]),
            .data_in         (data [413]),
            .scan_select_in  (scan [413]),
            .latch_enable_in (latch[413]),
            .clk_out         (clk  [414]),
            .data_out        (data [414]),
            .scan_select_out (scan [414]),
            .latch_enable_out(latch[414])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_414 (
            .clk_in          (clk  [414]),
            .data_in         (data [414]),
            .scan_select_in  (scan [414]),
            .latch_enable_in (latch[414]),
            .clk_out         (clk  [415]),
            .data_out        (data [415]),
            .scan_select_out (scan [415]),
            .latch_enable_out(latch[415])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_415 (
            .clk_in          (clk  [415]),
            .data_in         (data [415]),
            .scan_select_in  (scan [415]),
            .latch_enable_in (latch[415]),
            .clk_out         (clk  [416]),
            .data_out        (data [416]),
            .scan_select_out (scan [416]),
            .latch_enable_out(latch[416])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_416 (
            .clk_in          (clk  [416]),
            .data_in         (data [416]),
            .scan_select_in  (scan [416]),
            .latch_enable_in (latch[416]),
            .clk_out         (clk  [417]),
            .data_out        (data [417]),
            .scan_select_out (scan [417]),
            .latch_enable_out(latch[417])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_417 (
            .clk_in          (clk  [417]),
            .data_in         (data [417]),
            .scan_select_in  (scan [417]),
            .latch_enable_in (latch[417]),
            .clk_out         (clk  [418]),
            .data_out        (data [418]),
            .scan_select_out (scan [418]),
            .latch_enable_out(latch[418])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_418 (
            .clk_in          (clk  [418]),
            .data_in         (data [418]),
            .scan_select_in  (scan [418]),
            .latch_enable_in (latch[418]),
            .clk_out         (clk  [419]),
            .data_out        (data [419]),
            .scan_select_out (scan [419]),
            .latch_enable_out(latch[419])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_419 (
            .clk_in          (clk  [419]),
            .data_in         (data [419]),
            .scan_select_in  (scan [419]),
            .latch_enable_in (latch[419]),
            .clk_out         (clk  [420]),
            .data_out        (data [420]),
            .scan_select_out (scan [420]),
            .latch_enable_out(latch[420])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_420 (
            .clk_in          (clk  [420]),
            .data_in         (data [420]),
            .scan_select_in  (scan [420]),
            .latch_enable_in (latch[420]),
            .clk_out         (clk  [421]),
            .data_out        (data [421]),
            .scan_select_out (scan [421]),
            .latch_enable_out(latch[421])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_421 (
            .clk_in          (clk  [421]),
            .data_in         (data [421]),
            .scan_select_in  (scan [421]),
            .latch_enable_in (latch[421]),
            .clk_out         (clk  [422]),
            .data_out        (data [422]),
            .scan_select_out (scan [422]),
            .latch_enable_out(latch[422])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_422 (
            .clk_in          (clk  [422]),
            .data_in         (data [422]),
            .scan_select_in  (scan [422]),
            .latch_enable_in (latch[422]),
            .clk_out         (clk  [423]),
            .data_out        (data [423]),
            .scan_select_out (scan [423]),
            .latch_enable_out(latch[423])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_423 (
            .clk_in          (clk  [423]),
            .data_in         (data [423]),
            .scan_select_in  (scan [423]),
            .latch_enable_in (latch[423]),
            .clk_out         (clk  [424]),
            .data_out        (data [424]),
            .scan_select_out (scan [424]),
            .latch_enable_out(latch[424])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_424 (
            .clk_in          (clk  [424]),
            .data_in         (data [424]),
            .scan_select_in  (scan [424]),
            .latch_enable_in (latch[424]),
            .clk_out         (clk  [425]),
            .data_out        (data [425]),
            .scan_select_out (scan [425]),
            .latch_enable_out(latch[425])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_425 (
            .clk_in          (clk  [425]),
            .data_in         (data [425]),
            .scan_select_in  (scan [425]),
            .latch_enable_in (latch[425]),
            .clk_out         (clk  [426]),
            .data_out        (data [426]),
            .scan_select_out (scan [426]),
            .latch_enable_out(latch[426])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_426 (
            .clk_in          (clk  [426]),
            .data_in         (data [426]),
            .scan_select_in  (scan [426]),
            .latch_enable_in (latch[426]),
            .clk_out         (clk  [427]),
            .data_out        (data [427]),
            .scan_select_out (scan [427]),
            .latch_enable_out(latch[427])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_427 (
            .clk_in          (clk  [427]),
            .data_in         (data [427]),
            .scan_select_in  (scan [427]),
            .latch_enable_in (latch[427]),
            .clk_out         (clk  [428]),
            .data_out        (data [428]),
            .scan_select_out (scan [428]),
            .latch_enable_out(latch[428])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_428 (
            .clk_in          (clk  [428]),
            .data_in         (data [428]),
            .scan_select_in  (scan [428]),
            .latch_enable_in (latch[428]),
            .clk_out         (clk  [429]),
            .data_out        (data [429]),
            .scan_select_out (scan [429]),
            .latch_enable_out(latch[429])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_429 (
            .clk_in          (clk  [429]),
            .data_in         (data [429]),
            .scan_select_in  (scan [429]),
            .latch_enable_in (latch[429]),
            .clk_out         (clk  [430]),
            .data_out        (data [430]),
            .scan_select_out (scan [430]),
            .latch_enable_out(latch[430])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_430 (
            .clk_in          (clk  [430]),
            .data_in         (data [430]),
            .scan_select_in  (scan [430]),
            .latch_enable_in (latch[430]),
            .clk_out         (clk  [431]),
            .data_out        (data [431]),
            .scan_select_out (scan [431]),
            .latch_enable_out(latch[431])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_431 (
            .clk_in          (clk  [431]),
            .data_in         (data [431]),
            .scan_select_in  (scan [431]),
            .latch_enable_in (latch[431]),
            .clk_out         (clk  [432]),
            .data_out        (data [432]),
            .scan_select_out (scan [432]),
            .latch_enable_out(latch[432])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_432 (
            .clk_in          (clk  [432]),
            .data_in         (data [432]),
            .scan_select_in  (scan [432]),
            .latch_enable_in (latch[432]),
            .clk_out         (clk  [433]),
            .data_out        (data [433]),
            .scan_select_out (scan [433]),
            .latch_enable_out(latch[433])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_433 (
            .clk_in          (clk  [433]),
            .data_in         (data [433]),
            .scan_select_in  (scan [433]),
            .latch_enable_in (latch[433]),
            .clk_out         (clk  [434]),
            .data_out        (data [434]),
            .scan_select_out (scan [434]),
            .latch_enable_out(latch[434])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_434 (
            .clk_in          (clk  [434]),
            .data_in         (data [434]),
            .scan_select_in  (scan [434]),
            .latch_enable_in (latch[434]),
            .clk_out         (clk  [435]),
            .data_out        (data [435]),
            .scan_select_out (scan [435]),
            .latch_enable_out(latch[435])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_435 (
            .clk_in          (clk  [435]),
            .data_in         (data [435]),
            .scan_select_in  (scan [435]),
            .latch_enable_in (latch[435]),
            .clk_out         (clk  [436]),
            .data_out        (data [436]),
            .scan_select_out (scan [436]),
            .latch_enable_out(latch[436])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_436 (
            .clk_in          (clk  [436]),
            .data_in         (data [436]),
            .scan_select_in  (scan [436]),
            .latch_enable_in (latch[436]),
            .clk_out         (clk  [437]),
            .data_out        (data [437]),
            .scan_select_out (scan [437]),
            .latch_enable_out(latch[437])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_437 (
            .clk_in          (clk  [437]),
            .data_in         (data [437]),
            .scan_select_in  (scan [437]),
            .latch_enable_in (latch[437]),
            .clk_out         (clk  [438]),
            .data_out        (data [438]),
            .scan_select_out (scan [438]),
            .latch_enable_out(latch[438])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_438 (
            .clk_in          (clk  [438]),
            .data_in         (data [438]),
            .scan_select_in  (scan [438]),
            .latch_enable_in (latch[438]),
            .clk_out         (clk  [439]),
            .data_out        (data [439]),
            .scan_select_out (scan [439]),
            .latch_enable_out(latch[439])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_439 (
            .clk_in          (clk  [439]),
            .data_in         (data [439]),
            .scan_select_in  (scan [439]),
            .latch_enable_in (latch[439]),
            .clk_out         (clk  [440]),
            .data_out        (data [440]),
            .scan_select_out (scan [440]),
            .latch_enable_out(latch[440])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_440 (
            .clk_in          (clk  [440]),
            .data_in         (data [440]),
            .scan_select_in  (scan [440]),
            .latch_enable_in (latch[440]),
            .clk_out         (clk  [441]),
            .data_out        (data [441]),
            .scan_select_out (scan [441]),
            .latch_enable_out(latch[441])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_441 (
            .clk_in          (clk  [441]),
            .data_in         (data [441]),
            .scan_select_in  (scan [441]),
            .latch_enable_in (latch[441]),
            .clk_out         (clk  [442]),
            .data_out        (data [442]),
            .scan_select_out (scan [442]),
            .latch_enable_out(latch[442])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_442 (
            .clk_in          (clk  [442]),
            .data_in         (data [442]),
            .scan_select_in  (scan [442]),
            .latch_enable_in (latch[442]),
            .clk_out         (clk  [443]),
            .data_out        (data [443]),
            .scan_select_out (scan [443]),
            .latch_enable_out(latch[443])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_443 (
            .clk_in          (clk  [443]),
            .data_in         (data [443]),
            .scan_select_in  (scan [443]),
            .latch_enable_in (latch[443]),
            .clk_out         (clk  [444]),
            .data_out        (data [444]),
            .scan_select_out (scan [444]),
            .latch_enable_out(latch[444])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_444 (
            .clk_in          (clk  [444]),
            .data_in         (data [444]),
            .scan_select_in  (scan [444]),
            .latch_enable_in (latch[444]),
            .clk_out         (clk  [445]),
            .data_out        (data [445]),
            .scan_select_out (scan [445]),
            .latch_enable_out(latch[445])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_445 (
            .clk_in          (clk  [445]),
            .data_in         (data [445]),
            .scan_select_in  (scan [445]),
            .latch_enable_in (latch[445]),
            .clk_out         (clk  [446]),
            .data_out        (data [446]),
            .scan_select_out (scan [446]),
            .latch_enable_out(latch[446])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_446 (
            .clk_in          (clk  [446]),
            .data_in         (data [446]),
            .scan_select_in  (scan [446]),
            .latch_enable_in (latch[446]),
            .clk_out         (clk  [447]),
            .data_out        (data [447]),
            .scan_select_out (scan [447]),
            .latch_enable_out(latch[447])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_447 (
            .clk_in          (clk  [447]),
            .data_in         (data [447]),
            .scan_select_in  (scan [447]),
            .latch_enable_in (latch[447]),
            .clk_out         (clk  [448]),
            .data_out        (data [448]),
            .scan_select_out (scan [448]),
            .latch_enable_out(latch[448])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_448 (
            .clk_in          (clk  [448]),
            .data_in         (data [448]),
            .scan_select_in  (scan [448]),
            .latch_enable_in (latch[448]),
            .clk_out         (clk  [449]),
            .data_out        (data [449]),
            .scan_select_out (scan [449]),
            .latch_enable_out(latch[449])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_449 (
            .clk_in          (clk  [449]),
            .data_in         (data [449]),
            .scan_select_in  (scan [449]),
            .latch_enable_in (latch[449]),
            .clk_out         (clk  [450]),
            .data_out        (data [450]),
            .scan_select_out (scan [450]),
            .latch_enable_out(latch[450])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_450 (
            .clk_in          (clk  [450]),
            .data_in         (data [450]),
            .scan_select_in  (scan [450]),
            .latch_enable_in (latch[450]),
            .clk_out         (clk  [451]),
            .data_out        (data [451]),
            .scan_select_out (scan [451]),
            .latch_enable_out(latch[451])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_451 (
            .clk_in          (clk  [451]),
            .data_in         (data [451]),
            .scan_select_in  (scan [451]),
            .latch_enable_in (latch[451]),
            .clk_out         (clk  [452]),
            .data_out        (data [452]),
            .scan_select_out (scan [452]),
            .latch_enable_out(latch[452])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_452 (
            .clk_in          (clk  [452]),
            .data_in         (data [452]),
            .scan_select_in  (scan [452]),
            .latch_enable_in (latch[452]),
            .clk_out         (clk  [453]),
            .data_out        (data [453]),
            .scan_select_out (scan [453]),
            .latch_enable_out(latch[453])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_453 (
            .clk_in          (clk  [453]),
            .data_in         (data [453]),
            .scan_select_in  (scan [453]),
            .latch_enable_in (latch[453]),
            .clk_out         (clk  [454]),
            .data_out        (data [454]),
            .scan_select_out (scan [454]),
            .latch_enable_out(latch[454])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_454 (
            .clk_in          (clk  [454]),
            .data_in         (data [454]),
            .scan_select_in  (scan [454]),
            .latch_enable_in (latch[454]),
            .clk_out         (clk  [455]),
            .data_out        (data [455]),
            .scan_select_out (scan [455]),
            .latch_enable_out(latch[455])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_455 (
            .clk_in          (clk  [455]),
            .data_in         (data [455]),
            .scan_select_in  (scan [455]),
            .latch_enable_in (latch[455]),
            .clk_out         (clk  [456]),
            .data_out        (data [456]),
            .scan_select_out (scan [456]),
            .latch_enable_out(latch[456])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_456 (
            .clk_in          (clk  [456]),
            .data_in         (data [456]),
            .scan_select_in  (scan [456]),
            .latch_enable_in (latch[456]),
            .clk_out         (clk  [457]),
            .data_out        (data [457]),
            .scan_select_out (scan [457]),
            .latch_enable_out(latch[457])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_457 (
            .clk_in          (clk  [457]),
            .data_in         (data [457]),
            .scan_select_in  (scan [457]),
            .latch_enable_in (latch[457]),
            .clk_out         (clk  [458]),
            .data_out        (data [458]),
            .scan_select_out (scan [458]),
            .latch_enable_out(latch[458])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_458 (
            .clk_in          (clk  [458]),
            .data_in         (data [458]),
            .scan_select_in  (scan [458]),
            .latch_enable_in (latch[458]),
            .clk_out         (clk  [459]),
            .data_out        (data [459]),
            .scan_select_out (scan [459]),
            .latch_enable_out(latch[459])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_459 (
            .clk_in          (clk  [459]),
            .data_in         (data [459]),
            .scan_select_in  (scan [459]),
            .latch_enable_in (latch[459]),
            .clk_out         (clk  [460]),
            .data_out        (data [460]),
            .scan_select_out (scan [460]),
            .latch_enable_out(latch[460])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_460 (
            .clk_in          (clk  [460]),
            .data_in         (data [460]),
            .scan_select_in  (scan [460]),
            .latch_enable_in (latch[460]),
            .clk_out         (clk  [461]),
            .data_out        (data [461]),
            .scan_select_out (scan [461]),
            .latch_enable_out(latch[461])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_461 (
            .clk_in          (clk  [461]),
            .data_in         (data [461]),
            .scan_select_in  (scan [461]),
            .latch_enable_in (latch[461]),
            .clk_out         (clk  [462]),
            .data_out        (data [462]),
            .scan_select_out (scan [462]),
            .latch_enable_out(latch[462])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_462 (
            .clk_in          (clk  [462]),
            .data_in         (data [462]),
            .scan_select_in  (scan [462]),
            .latch_enable_in (latch[462]),
            .clk_out         (clk  [463]),
            .data_out        (data [463]),
            .scan_select_out (scan [463]),
            .latch_enable_out(latch[463])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_463 (
            .clk_in          (clk  [463]),
            .data_in         (data [463]),
            .scan_select_in  (scan [463]),
            .latch_enable_in (latch[463]),
            .clk_out         (clk  [464]),
            .data_out        (data [464]),
            .scan_select_out (scan [464]),
            .latch_enable_out(latch[464])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_464 (
            .clk_in          (clk  [464]),
            .data_in         (data [464]),
            .scan_select_in  (scan [464]),
            .latch_enable_in (latch[464]),
            .clk_out         (clk  [465]),
            .data_out        (data [465]),
            .scan_select_out (scan [465]),
            .latch_enable_out(latch[465])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_465 (
            .clk_in          (clk  [465]),
            .data_in         (data [465]),
            .scan_select_in  (scan [465]),
            .latch_enable_in (latch[465]),
            .clk_out         (clk  [466]),
            .data_out        (data [466]),
            .scan_select_out (scan [466]),
            .latch_enable_out(latch[466])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_466 (
            .clk_in          (clk  [466]),
            .data_in         (data [466]),
            .scan_select_in  (scan [466]),
            .latch_enable_in (latch[466]),
            .clk_out         (clk  [467]),
            .data_out        (data [467]),
            .scan_select_out (scan [467]),
            .latch_enable_out(latch[467])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_467 (
            .clk_in          (clk  [467]),
            .data_in         (data [467]),
            .scan_select_in  (scan [467]),
            .latch_enable_in (latch[467]),
            .clk_out         (clk  [468]),
            .data_out        (data [468]),
            .scan_select_out (scan [468]),
            .latch_enable_out(latch[468])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_468 (
            .clk_in          (clk  [468]),
            .data_in         (data [468]),
            .scan_select_in  (scan [468]),
            .latch_enable_in (latch[468]),
            .clk_out         (clk  [469]),
            .data_out        (data [469]),
            .scan_select_out (scan [469]),
            .latch_enable_out(latch[469])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_469 (
            .clk_in          (clk  [469]),
            .data_in         (data [469]),
            .scan_select_in  (scan [469]),
            .latch_enable_in (latch[469]),
            .clk_out         (clk  [470]),
            .data_out        (data [470]),
            .scan_select_out (scan [470]),
            .latch_enable_out(latch[470])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_470 (
            .clk_in          (clk  [470]),
            .data_in         (data [470]),
            .scan_select_in  (scan [470]),
            .latch_enable_in (latch[470]),
            .clk_out         (clk  [471]),
            .data_out        (data [471]),
            .scan_select_out (scan [471]),
            .latch_enable_out(latch[471])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_471 (
            .clk_in          (clk  [471]),
            .data_in         (data [471]),
            .scan_select_in  (scan [471]),
            .latch_enable_in (latch[471]),
            .clk_out         (clk  [472]),
            .data_out        (data [472]),
            .scan_select_out (scan [472]),
            .latch_enable_out(latch[472])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_472 (
            .clk_in          (clk  [472]),
            .data_in         (data [472]),
            .scan_select_in  (scan [472]),
            .latch_enable_in (latch[472]),
            .clk_out         (clk  [473]),
            .data_out        (data [473]),
            .scan_select_out (scan [473]),
            .latch_enable_out(latch[473])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_473 (
            .clk_in          (clk  [473]),
            .data_in         (data [473]),
            .scan_select_in  (scan [473]),
            .latch_enable_in (latch[473]),
            .clk_out         (clk  [474]),
            .data_out        (data [474]),
            .scan_select_out (scan [474]),
            .latch_enable_out(latch[474])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_474 (
            .clk_in          (clk  [474]),
            .data_in         (data [474]),
            .scan_select_in  (scan [474]),
            .latch_enable_in (latch[474]),
            .clk_out         (clk  [475]),
            .data_out        (data [475]),
            .scan_select_out (scan [475]),
            .latch_enable_out(latch[475])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_475 (
            .clk_in          (clk  [475]),
            .data_in         (data [475]),
            .scan_select_in  (scan [475]),
            .latch_enable_in (latch[475]),
            .clk_out         (clk  [476]),
            .data_out        (data [476]),
            .scan_select_out (scan [476]),
            .latch_enable_out(latch[476])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_476 (
            .clk_in          (clk  [476]),
            .data_in         (data [476]),
            .scan_select_in  (scan [476]),
            .latch_enable_in (latch[476]),
            .clk_out         (clk  [477]),
            .data_out        (data [477]),
            .scan_select_out (scan [477]),
            .latch_enable_out(latch[477])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_477 (
            .clk_in          (clk  [477]),
            .data_in         (data [477]),
            .scan_select_in  (scan [477]),
            .latch_enable_in (latch[477]),
            .clk_out         (clk  [478]),
            .data_out        (data [478]),
            .scan_select_out (scan [478]),
            .latch_enable_out(latch[478])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_478 (
            .clk_in          (clk  [478]),
            .data_in         (data [478]),
            .scan_select_in  (scan [478]),
            .latch_enable_in (latch[478]),
            .clk_out         (clk  [479]),
            .data_out        (data [479]),
            .scan_select_out (scan [479]),
            .latch_enable_out(latch[479])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_479 (
            .clk_in          (clk  [479]),
            .data_in         (data [479]),
            .scan_select_in  (scan [479]),
            .latch_enable_in (latch[479]),
            .clk_out         (clk  [480]),
            .data_out        (data [480]),
            .scan_select_out (scan [480]),
            .latch_enable_out(latch[480])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_480 (
            .clk_in          (clk  [480]),
            .data_in         (data [480]),
            .scan_select_in  (scan [480]),
            .latch_enable_in (latch[480]),
            .clk_out         (clk  [481]),
            .data_out        (data [481]),
            .scan_select_out (scan [481]),
            .latch_enable_out(latch[481])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_481 (
            .clk_in          (clk  [481]),
            .data_in         (data [481]),
            .scan_select_in  (scan [481]),
            .latch_enable_in (latch[481]),
            .clk_out         (clk  [482]),
            .data_out        (data [482]),
            .scan_select_out (scan [482]),
            .latch_enable_out(latch[482])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_482 (
            .clk_in          (clk  [482]),
            .data_in         (data [482]),
            .scan_select_in  (scan [482]),
            .latch_enable_in (latch[482]),
            .clk_out         (clk  [483]),
            .data_out        (data [483]),
            .scan_select_out (scan [483]),
            .latch_enable_out(latch[483])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_483 (
            .clk_in          (clk  [483]),
            .data_in         (data [483]),
            .scan_select_in  (scan [483]),
            .latch_enable_in (latch[483]),
            .clk_out         (clk  [484]),
            .data_out        (data [484]),
            .scan_select_out (scan [484]),
            .latch_enable_out(latch[484])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_484 (
            .clk_in          (clk  [484]),
            .data_in         (data [484]),
            .scan_select_in  (scan [484]),
            .latch_enable_in (latch[484]),
            .clk_out         (clk  [485]),
            .data_out        (data [485]),
            .scan_select_out (scan [485]),
            .latch_enable_out(latch[485])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_485 (
            .clk_in          (clk  [485]),
            .data_in         (data [485]),
            .scan_select_in  (scan [485]),
            .latch_enable_in (latch[485]),
            .clk_out         (clk  [486]),
            .data_out        (data [486]),
            .scan_select_out (scan [486]),
            .latch_enable_out(latch[486])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_486 (
            .clk_in          (clk  [486]),
            .data_in         (data [486]),
            .scan_select_in  (scan [486]),
            .latch_enable_in (latch[486]),
            .clk_out         (clk  [487]),
            .data_out        (data [487]),
            .scan_select_out (scan [487]),
            .latch_enable_out(latch[487])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_487 (
            .clk_in          (clk  [487]),
            .data_in         (data [487]),
            .scan_select_in  (scan [487]),
            .latch_enable_in (latch[487]),
            .clk_out         (clk  [488]),
            .data_out        (data [488]),
            .scan_select_out (scan [488]),
            .latch_enable_out(latch[488])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_488 (
            .clk_in          (clk  [488]),
            .data_in         (data [488]),
            .scan_select_in  (scan [488]),
            .latch_enable_in (latch[488]),
            .clk_out         (clk  [489]),
            .data_out        (data [489]),
            .scan_select_out (scan [489]),
            .latch_enable_out(latch[489])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_489 (
            .clk_in          (clk  [489]),
            .data_in         (data [489]),
            .scan_select_in  (scan [489]),
            .latch_enable_in (latch[489]),
            .clk_out         (clk  [490]),
            .data_out        (data [490]),
            .scan_select_out (scan [490]),
            .latch_enable_out(latch[490])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_490 (
            .clk_in          (clk  [490]),
            .data_in         (data [490]),
            .scan_select_in  (scan [490]),
            .latch_enable_in (latch[490]),
            .clk_out         (clk  [491]),
            .data_out        (data [491]),
            .scan_select_out (scan [491]),
            .latch_enable_out(latch[491])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_491 (
            .clk_in          (clk  [491]),
            .data_in         (data [491]),
            .scan_select_in  (scan [491]),
            .latch_enable_in (latch[491]),
            .clk_out         (clk  [492]),
            .data_out        (data [492]),
            .scan_select_out (scan [492]),
            .latch_enable_out(latch[492])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_492 (
            .clk_in          (clk  [492]),
            .data_in         (data [492]),
            .scan_select_in  (scan [492]),
            .latch_enable_in (latch[492]),
            .clk_out         (clk  [493]),
            .data_out        (data [493]),
            .scan_select_out (scan [493]),
            .latch_enable_out(latch[493])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_493 (
            .clk_in          (clk  [493]),
            .data_in         (data [493]),
            .scan_select_in  (scan [493]),
            .latch_enable_in (latch[493]),
            .clk_out         (clk  [494]),
            .data_out        (data [494]),
            .scan_select_out (scan [494]),
            .latch_enable_out(latch[494])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_494 (
            .clk_in          (clk  [494]),
            .data_in         (data [494]),
            .scan_select_in  (scan [494]),
            .latch_enable_in (latch[494]),
            .clk_out         (clk  [495]),
            .data_out        (data [495]),
            .scan_select_out (scan [495]),
            .latch_enable_out(latch[495])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_495 (
            .clk_in          (clk  [495]),
            .data_in         (data [495]),
            .scan_select_in  (scan [495]),
            .latch_enable_in (latch[495]),
            .clk_out         (clk  [496]),
            .data_out        (data [496]),
            .scan_select_out (scan [496]),
            .latch_enable_out(latch[496])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_496 (
            .clk_in          (clk  [496]),
            .data_in         (data [496]),
            .scan_select_in  (scan [496]),
            .latch_enable_in (latch[496]),
            .clk_out         (clk  [497]),
            .data_out        (data [497]),
            .scan_select_out (scan [497]),
            .latch_enable_out(latch[497])
            );
        
        // https://github.com/mattvenn/wokwi_filler
        scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_497 (
            .clk_in          (clk  [497]),
            .data_in         (data [497]),
            .scan_select_in  (scan [497]),
            .latch_enable_in (latch[497]),
            .clk_out         (clk  [498]),
            .data_out        (data [498]),
            .scan_select_out (scan [498]),
            .latch_enable_out(latch[498])
            );
            // end of module instantiation

endmodule	// user_project_wrapper
`default_nettype wire
