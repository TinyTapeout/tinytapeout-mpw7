module scan_wrapper_341426151397261906 (clk_in,
    clk_out,
    data_in,
    data_out,
    latch_enable_in,
    latch_enable_out,
    scan_select_in,
    scan_select_out,
    vccd1,
    vssd1);
 input clk_in;
 output clk_out;
 input data_in;
 output data_out;
 input latch_enable_in;
 output latch_enable_out;
 input scan_select_in;
 output scan_select_out;
 input vccd1;
 input vssd1;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire clk;
 wire data_in_i;
 wire data_out_i;
 wire scan_select_in_i;
 wire \user_module.clk_slow ;
 wire \user_module.eio_in[0] ;
 wire \user_module.eio_in[10] ;
 wire \user_module.eio_in[11] ;
 wire \user_module.eio_in[12] ;
 wire \user_module.eio_in[13] ;
 wire \user_module.eio_in[14] ;
 wire \user_module.eio_in[15] ;
 wire \user_module.eio_in[16] ;
 wire \user_module.eio_in[17] ;
 wire \user_module.eio_in[18] ;
 wire \user_module.eio_in[19] ;
 wire \user_module.eio_in[1] ;
 wire \user_module.eio_in[2] ;
 wire \user_module.eio_in[3] ;
 wire \user_module.eio_in[4] ;
 wire \user_module.eio_in[5] ;
 wire \user_module.eio_in[6] ;
 wire \user_module.eio_in[7] ;
 wire \user_module.eio_in[8] ;
 wire \user_module.eio_in[9] ;
 wire \user_module.eio_latch_n[0] ;
 wire \user_module.eio_latch_n[1] ;
 wire \user_module.eio_latch_n[2] ;
 wire \user_module.eio_latch_n[3] ;
 wire \user_module.eio_latch_n[4] ;
 wire \user_module.eio_out[0] ;
 wire \user_module.eio_out[1] ;
 wire \user_module.eio_out[2] ;
 wire \user_module.eio_out[3] ;
 wire \user_module.eio_out[4] ;
 wire \user_module.eio_out[5] ;
 wire \user_module.eio_out[6] ;
 wire \user_module.eio_out[7] ;
 wire \user_module.io_in[0] ;
 wire \user_module.io_in[1] ;
 wire \user_module.io_in[2] ;
 wire \user_module.io_in[3] ;
 wire \user_module.io_in[4] ;
 wire \user_module.io_in[5] ;
 wire \user_module.io_in[6] ;
 wire \user_module.io_in[7] ;
 wire \user_module.io_out[0] ;
 wire \user_module.io_out[1] ;
 wire \user_module.io_out[2] ;
 wire \user_module.io_out[3] ;
 wire \user_module.io_out[4] ;
 wire \user_module.io_out[5] ;
 wire \user_module.io_out[6] ;
 wire \user_module.io_out[7] ;
 wire \user_module.latch_in ;
 wire \user_module.ram_I.clk_dly ;
 wire \user_module.ram_I.raddr_dec_I.in[0] ;
 wire \user_module.ram_I.raddr_dec_I.in[1] ;
 wire \user_module.ram_I.raddr_dec_I.out[0] ;
 wire \user_module.ram_I.raddr_dec_I.out[1] ;
 wire \user_module.ram_I.raddr_dec_I.out[2] ;
 wire \user_module.ram_I.raddr_dec_I.out[3] ;
 wire \user_module.ram_I.raddr_r[0] ;
 wire \user_module.ram_I.raddr_r[1] ;
 wire \user_module.ram_I.rdata_inv[0] ;
 wire \user_module.ram_I.rdata_inv[1] ;
 wire \user_module.ram_I.rdata_inv[2] ;
 wire \user_module.ram_I.rdata_inv[3] ;
 wire \user_module.ram_I.rdata_inv[4] ;
 wire \user_module.ram_I.rdata_inv[5] ;
 wire \user_module.ram_I.rdata_inv[6] ;
 wire \user_module.ram_I.rdata_inv[7] ;
 wire \user_module.ram_I.rdata_le_n ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in0_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in0_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in0_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in0_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in0_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in0_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in0_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in0_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in1_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in1_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in1_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in1_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in1_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in1_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in1_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in1_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in2_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in2_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in2_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in2_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in2_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in2_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in2_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in2_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in3_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in3_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in3_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in3_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in3_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in3_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in3_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_in3_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_out_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_out_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_out_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_out_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_out_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_out_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_out_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[0].l_out_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in0_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in0_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in0_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in0_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in0_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in0_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in0_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in0_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in1_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in1_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in1_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in1_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in1_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in1_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in1_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in1_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in2_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in2_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in2_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in2_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in2_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in2_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in2_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in2_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in3_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in3_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in3_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in3_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in3_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in3_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in3_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_in3_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_out_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_out_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_out_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_out_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_out_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_out_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_out_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[12].l_out_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in0_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in0_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in0_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in0_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in0_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in0_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in0_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in0_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in1_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in1_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in1_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in1_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in1_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in1_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in1_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in1_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in2_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in2_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in2_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in2_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in2_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in2_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in2_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in2_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in3_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in3_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in3_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in3_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in3_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in3_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in3_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_in3_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_out_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_out_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_out_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_out_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_out_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_out_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_out_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[4].l_out_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in0_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in0_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in0_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in0_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in0_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in0_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in0_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in0_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in1_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in1_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in1_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in1_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in1_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in1_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in1_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in1_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in2_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in2_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in2_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in2_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in2_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in2_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in2_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in2_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in3_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in3_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in3_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in3_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in3_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in3_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in3_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_in3_mux[7] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_out_mux[0] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_out_mux[1] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_out_mux[2] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_out_mux[3] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_out_mux[4] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_out_mux[5] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_out_mux[6] ;
 wire \user_module.ram_I.rdata_sel_loop[8].l_out_mux[7] ;
 wire \user_module.ram_I.rdata_tbuf[0] ;
 wire \user_module.ram_I.rdata_tbuf[1] ;
 wire \user_module.ram_I.rdata_tbuf[2] ;
 wire \user_module.ram_I.rdata_tbuf[3] ;
 wire \user_module.ram_I.rdata_tbuf[4] ;
 wire \user_module.ram_I.rdata_tbuf[5] ;
 wire \user_module.ram_I.rdata_tbuf[6] ;
 wire \user_module.ram_I.rdata_tbuf[7] ;
 wire \user_module.ram_I.re_r ;
 wire \user_module.ram_I.store_gate[0] ;
 wire \user_module.ram_I.store_gate[10] ;
 wire \user_module.ram_I.store_gate[11] ;
 wire \user_module.ram_I.store_gate[12] ;
 wire \user_module.ram_I.store_gate[13] ;
 wire \user_module.ram_I.store_gate[14] ;
 wire \user_module.ram_I.store_gate[15] ;
 wire \user_module.ram_I.store_gate[1] ;
 wire \user_module.ram_I.store_gate[2] ;
 wire \user_module.ram_I.store_gate[3] ;
 wire \user_module.ram_I.store_gate[4] ;
 wire \user_module.ram_I.store_gate[5] ;
 wire \user_module.ram_I.store_gate[6] ;
 wire \user_module.ram_I.store_gate[7] ;
 wire \user_module.ram_I.store_gate[8] ;
 wire \user_module.ram_I.store_gate[9] ;
 wire \user_module.ram_I.store_in[0] ;
 wire \user_module.ram_I.store_in[1] ;
 wire \user_module.ram_I.store_in[2] ;
 wire \user_module.ram_I.store_in[3] ;
 wire \user_module.ram_I.store_in[4] ;
 wire \user_module.ram_I.store_in[5] ;
 wire \user_module.ram_I.store_in[6] ;
 wire \user_module.ram_I.store_in[7] ;
 wire \user_module.ram_I.waddr_dec[0] ;
 wire \user_module.ram_I.waddr_dec[10] ;
 wire \user_module.ram_I.waddr_dec[11] ;
 wire \user_module.ram_I.waddr_dec[12] ;
 wire \user_module.ram_I.waddr_dec[13] ;
 wire \user_module.ram_I.waddr_dec[14] ;
 wire \user_module.ram_I.waddr_dec[15] ;
 wire \user_module.ram_I.waddr_dec[1] ;
 wire \user_module.ram_I.waddr_dec[2] ;
 wire \user_module.ram_I.waddr_dec[3] ;
 wire \user_module.ram_I.waddr_dec[4] ;
 wire \user_module.ram_I.waddr_dec[5] ;
 wire \user_module.ram_I.waddr_dec[6] ;
 wire \user_module.ram_I.waddr_dec[7] ;
 wire \user_module.ram_I.waddr_dec[8] ;
 wire \user_module.ram_I.waddr_dec[9] ;
 wire \user_module.ram_I.waddr_dec_I.in[0] ;
 wire \user_module.ram_I.waddr_dec_I.in[1] ;
 wire \user_module.ram_I.waddr_dec_I.in[2] ;
 wire \user_module.ram_I.waddr_dec_I.in[3] ;
 wire \user_module.ram_I.we_r ;
 wire \user_module.ram_I.wpulse_I.clk_dly ;
 wire \user_module.ram_I.wpulse_I.clk_dly_chain[1] ;
 wire \user_module.ram_I.wpulse_I.clk_dly_chain[2] ;
 wire \user_module.ram_I.wpulse_I.clk_dly_chain[3] ;
 wire \user_module.ram_I.wpulse_I.clk_dly_chain[4] ;
 wire \user_module.ram_I.wpulse_I.clk_dly_chain[5] ;
 wire \user_module.ram_I.wpulse_I.clk_dly_chain[6] ;
 wire \user_module.ram_I.wpulse_I.clk_dly_chain[7] ;
 wire \user_module.ram_I.wpulse_I.pulse ;

 sky130_fd_sc_hd__diode_2 ANTENNA_0 (.DIODE(_03_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_03_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\user_module.ram_I.waddr_dec[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_11_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_12_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_13_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_15_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_16_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_16_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_16_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_16_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_20_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_21_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_21_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_21_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_22_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_22_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_23_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_24_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_24_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_24_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_186 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_25_198 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_170 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_26_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_26_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_27_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_27_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_27_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_172 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_184 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_27_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_27_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_28_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_158 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_170 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_182 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_28_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_29_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_155 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_29_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_29_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_184 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_2_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_2_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_2_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_3_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_4_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_4_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_4_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_6_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_7_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_8_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_9_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _11_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(_06_));
 sky130_fd_sc_hd__conb_1 _12_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(_00_));
 sky130_fd_sc_hd__conb_1 _13_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(_01_));
 sky130_fd_sc_hd__conb_1 _14_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(_02_));
 sky130_fd_sc_hd__conb_1 _15_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(_03_));
 sky130_fd_sc_hd__conb_1 _16_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(_04_));
 sky130_fd_sc_hd__conb_1 _17_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(_05_));
 sky130_fd_sc_hd__conb_1 _18_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(_07_));
 sky130_fd_sc_hd__conb_1 _19_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(_08_));
 sky130_fd_sc_hd__conb_1 _20_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(_09_));
 sky130_fd_sc_hd__conb_1 _21_ (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(_10_));
 sky130_fd_sc_hd__clkbuf_2 input_buf_clk (.A(clk_in),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clk));
 sky130_fd_sc_hd__buf_2 \input_buffers[0]  (.A(latch_enable_in),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.latch_in ));
 sky130_fd_sc_hd__buf_2 \input_buffers[1]  (.A(scan_select_in),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(scan_select_in_i));
 sky130_fd_sc_hd__buf_2 \input_buffers[2]  (.A(data_in),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(data_in_i));
 sky130_fd_sc_hd__dfrtn_1 out_flop (.CLK_N(clk),
    .D(\user_module.io_in[7] ),
    .RESET_B(_00_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(data_out_i));
 sky130_fd_sc_hd__buf_4 \output_buffers[0]  (.A(\user_module.latch_in ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(latch_enable_out));
 sky130_fd_sc_hd__buf_4 \output_buffers[1]  (.A(scan_select_in_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(scan_select_out));
 sky130_fd_sc_hd__buf_4 \output_buffers[2]  (.A(data_out_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(data_out));
 sky130_fd_sc_hd__buf_4 \output_buffers[3]  (.A(clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clk_out));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[0]  (.CLK(clk),
    .D(data_in_i),
    .SCD(\user_module.io_out[0] ),
    .SCE(scan_select_in_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.io_in[0] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[1]  (.CLK(clk),
    .D(\user_module.io_in[0] ),
    .SCD(\user_module.io_out[1] ),
    .SCE(scan_select_in_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.io_in[1] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[2]  (.CLK(clk),
    .D(\user_module.io_in[1] ),
    .SCD(\user_module.io_out[2] ),
    .SCE(scan_select_in_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.io_in[2] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[3]  (.CLK(clk),
    .D(\user_module.io_in[2] ),
    .SCD(\user_module.io_out[3] ),
    .SCE(scan_select_in_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.io_in[3] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[4]  (.CLK(clk),
    .D(\user_module.io_in[3] ),
    .SCD(\user_module.io_out[4] ),
    .SCE(scan_select_in_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.io_in[4] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[5]  (.CLK(clk),
    .D(\user_module.io_in[4] ),
    .SCD(\user_module.io_out[5] ),
    .SCE(scan_select_in_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.io_in[5] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[6]  (.CLK(clk),
    .D(\user_module.io_in[5] ),
    .SCD(\user_module.io_out[6] ),
    .SCE(scan_select_in_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.io_in[6] ));
 sky130_fd_sc_hd__sdfxtp_1 \scan_flop[7]  (.CLK(clk),
    .D(\user_module.io_in[6] ),
    .SCD(\user_module.io_out[7] ),
    .SCE(scan_select_in_i),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.io_in[7] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[0].in_latch_I[0]  (.D(\user_module.io_in[4] ),
    .GATE_N(\user_module.eio_latch_n[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[0] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[0].in_latch_I[1]  (.D(\user_module.io_in[5] ),
    .GATE_N(\user_module.eio_latch_n[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[1] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[0].in_latch_I[2]  (.D(\user_module.io_in[6] ),
    .GATE_N(\user_module.eio_latch_n[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[2] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[0].in_latch_I[3]  (.D(\user_module.io_in[7] ),
    .GATE_N(\user_module.eio_latch_n[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[3] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[1].in_latch_I[0]  (.D(\user_module.io_in[4] ),
    .GATE_N(\user_module.eio_latch_n[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[4] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[1].in_latch_I[1]  (.D(\user_module.io_in[5] ),
    .GATE_N(\user_module.eio_latch_n[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[5] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[1].in_latch_I[2]  (.D(\user_module.io_in[6] ),
    .GATE_N(\user_module.eio_latch_n[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[6] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[1].in_latch_I[3]  (.D(\user_module.io_in[7] ),
    .GATE_N(\user_module.eio_latch_n[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[7] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[2].in_latch_I[0]  (.D(\user_module.io_in[4] ),
    .GATE_N(\user_module.eio_latch_n[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[8] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[2].in_latch_I[1]  (.D(\user_module.io_in[5] ),
    .GATE_N(\user_module.eio_latch_n[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[9] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[2].in_latch_I[2]  (.D(\user_module.io_in[6] ),
    .GATE_N(\user_module.eio_latch_n[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[10] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[2].in_latch_I[3]  (.D(\user_module.io_in[7] ),
    .GATE_N(\user_module.eio_latch_n[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[11] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[3].in_latch_I[0]  (.D(\user_module.io_in[4] ),
    .GATE_N(\user_module.eio_latch_n[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[12] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[3].in_latch_I[1]  (.D(\user_module.io_in[5] ),
    .GATE_N(\user_module.eio_latch_n[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[13] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[3].in_latch_I[2]  (.D(\user_module.io_in[6] ),
    .GATE_N(\user_module.eio_latch_n[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[14] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[3].in_latch_I[3]  (.D(\user_module.io_in[7] ),
    .GATE_N(\user_module.eio_latch_n[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[15] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[4].in_latch_I[0]  (.D(\user_module.io_in[4] ),
    .GATE_N(\user_module.eio_latch_n[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[16] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[4].in_latch_I[1]  (.D(\user_module.io_in[5] ),
    .GATE_N(\user_module.eio_latch_n[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[17] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[4].in_latch_I[2]  (.D(\user_module.io_in[6] ),
    .GATE_N(\user_module.eio_latch_n[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[18] ));
 sky130_fd_sc_hd__dlxtn_1 \user_module.genblk1[4].in_latch_I[3]  (.D(\user_module.io_in[7] ),
    .GATE_N(\user_module.eio_latch_n[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_in[19] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.in_clk_slow_I  (.D(\user_module.io_in[0] ),
    .GATE(\user_module.latch_in ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.clk_slow ));
 sky130_fd_sc_hd__or4b_1 \user_module.in_dec_0_I  (.A(\user_module.io_in[1] ),
    .B(\user_module.io_in[2] ),
    .C(\user_module.io_in[3] ),
    .D_N(\user_module.latch_in ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.eio_latch_n[0] ));
 sky130_fd_sc_hd__nand4bb_1 \user_module.in_dec_1_I  (.A_N(\user_module.io_in[3] ),
    .B_N(\user_module.io_in[2] ),
    .C(\user_module.io_in[1] ),
    .D(\user_module.latch_in ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.eio_latch_n[1] ));
 sky130_fd_sc_hd__nand4bb_1 \user_module.in_dec_2_I  (.A_N(\user_module.io_in[3] ),
    .B_N(\user_module.io_in[1] ),
    .C(\user_module.io_in[2] ),
    .D(\user_module.latch_in ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.eio_latch_n[2] ));
 sky130_fd_sc_hd__nand4b_1 \user_module.in_dec_3_I  (.A_N(\user_module.io_in[3] ),
    .B(\user_module.io_in[2] ),
    .C(\user_module.io_in[1] ),
    .D(\user_module.latch_in ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.eio_latch_n[3] ));
 sky130_fd_sc_hd__nand4bb_1 \user_module.in_dec_4_I  (.A_N(\user_module.io_in[1] ),
    .B_N(\user_module.io_in[2] ),
    .C(\user_module.io_in[3] ),
    .D(\user_module.latch_in ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.eio_latch_n[4] ));
 sky130_fd_sc_hd__mux4_1 \user_module.out_mux_I[0]  (.A0(\user_module.eio_out[0] ),
    .A1(\user_module.eio_in[12] ),
    .A2(\user_module.eio_in[4] ),
    .A3(_01_),
    .S0(\user_module.eio_in[0] ),
    .S1(\user_module.eio_in[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.io_out[0] ));
 sky130_fd_sc_hd__mux4_1 \user_module.out_mux_I[1]  (.A0(\user_module.eio_out[1] ),
    .A1(\user_module.eio_in[13] ),
    .A2(\user_module.eio_in[5] ),
    .A3(_07_),
    .S0(\user_module.eio_in[0] ),
    .S1(\user_module.eio_in[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.io_out[1] ));
 sky130_fd_sc_hd__mux4_1 \user_module.out_mux_I[2]  (.A0(\user_module.eio_out[2] ),
    .A1(\user_module.eio_in[14] ),
    .A2(\user_module.eio_in[6] ),
    .A3(_02_),
    .S0(\user_module.eio_in[0] ),
    .S1(\user_module.eio_in[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.io_out[2] ));
 sky130_fd_sc_hd__mux4_1 \user_module.out_mux_I[3]  (.A0(\user_module.eio_out[3] ),
    .A1(\user_module.eio_in[15] ),
    .A2(\user_module.eio_in[7] ),
    .A3(_08_),
    .S0(\user_module.eio_in[0] ),
    .S1(\user_module.eio_in[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.io_out[3] ));
 sky130_fd_sc_hd__mux4_1 \user_module.out_mux_I[4]  (.A0(\user_module.eio_out[4] ),
    .A1(\user_module.eio_in[16] ),
    .A2(\user_module.eio_in[8] ),
    .A3(_09_),
    .S0(\user_module.eio_in[0] ),
    .S1(\user_module.eio_in[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.io_out[4] ));
 sky130_fd_sc_hd__mux4_1 \user_module.out_mux_I[5]  (.A0(\user_module.eio_out[5] ),
    .A1(\user_module.eio_in[17] ),
    .A2(\user_module.eio_in[9] ),
    .A3(_03_),
    .S0(\user_module.eio_in[0] ),
    .S1(\user_module.eio_in[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.io_out[5] ));
 sky130_fd_sc_hd__mux4_1 \user_module.out_mux_I[6]  (.A0(\user_module.eio_out[6] ),
    .A1(\user_module.eio_in[18] ),
    .A2(\user_module.eio_in[10] ),
    .A3(_10_),
    .S0(\user_module.eio_in[0] ),
    .S1(\user_module.eio_in[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.io_out[6] ));
 sky130_fd_sc_hd__mux4_1 \user_module.out_mux_I[7]  (.A0(\user_module.eio_out[7] ),
    .A1(\user_module.eio_in[19] ),
    .A2(\user_module.eio_in[11] ),
    .A3(_04_),
    .S0(\user_module.eio_in[0] ),
    .S1(\user_module.eio_in[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.io_out[7] ));
 sky130_fd_sc_hd__clkdlybuf4s50_1 \user_module.ram_I.clk_dly_I  (.A(\user_module.clk_slow ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.clk_dly ));
 sky130_fd_sc_hd__nand3_2 \user_module.ram_I.data_le_n_I  (.A(\user_module.clk_slow ),
    .B(\user_module.ram_I.clk_dly ),
    .C(\user_module.ram_I.re_r ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.ram_I.rdata_le_n ));
 sky130_fd_sc_hd__nor2_1 \user_module.ram_I.raddr_dec_I.dec_2_0_I  (.A(\user_module.ram_I.raddr_dec_I.in[0] ),
    .B(\user_module.ram_I.raddr_dec_I.in[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.ram_I.raddr_dec_I.out[0] ));
 sky130_fd_sc_hd__and2b_1 \user_module.ram_I.raddr_dec_I.dec_2_1_I  (.A_N(\user_module.ram_I.raddr_dec_I.in[1] ),
    .B(\user_module.ram_I.raddr_dec_I.in[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.raddr_dec_I.out[1] ));
 sky130_fd_sc_hd__and2b_1 \user_module.ram_I.raddr_dec_I.dec_2_2_I  (.A_N(\user_module.ram_I.raddr_dec_I.in[0] ),
    .B(\user_module.ram_I.raddr_dec_I.in[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.raddr_dec_I.out[2] ));
 sky130_fd_sc_hd__and2_1 \user_module.ram_I.raddr_dec_I.dec_2_3_I  (.A(\user_module.ram_I.raddr_dec_I.in[0] ),
    .B(\user_module.ram_I.raddr_dec_I.in[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.raddr_dec_I.out[3] ));
 sky130_fd_sc_hd__dfxtp_4 \user_module.ram_I.raddr_reg_lsb_I[0]  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.raddr_r[0] ));
 sky130_fd_sc_hd__dfxtp_4 \user_module.ram_I.raddr_reg_lsb_I[1]  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.raddr_r[1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.ram_I.raddr_reg_msb_I[0]  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.raddr_dec_I.in[0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.ram_I.raddr_reg_msb_I[1]  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.raddr_dec_I.in[1] ));
 sky130_fd_sc_hd__inv_1 \user_module.ram_I.rdata_inv_I[0]  (.A(\user_module.ram_I.rdata_tbuf[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.ram_I.rdata_inv[0] ));
 sky130_fd_sc_hd__inv_1 \user_module.ram_I.rdata_inv_I[1]  (.A(\user_module.ram_I.rdata_tbuf[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.ram_I.rdata_inv[1] ));
 sky130_fd_sc_hd__inv_1 \user_module.ram_I.rdata_inv_I[2]  (.A(\user_module.ram_I.rdata_tbuf[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.ram_I.rdata_inv[2] ));
 sky130_fd_sc_hd__inv_1 \user_module.ram_I.rdata_inv_I[3]  (.A(\user_module.ram_I.rdata_tbuf[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.ram_I.rdata_inv[3] ));
 sky130_fd_sc_hd__inv_1 \user_module.ram_I.rdata_inv_I[4]  (.A(\user_module.ram_I.rdata_tbuf[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.ram_I.rdata_inv[4] ));
 sky130_fd_sc_hd__inv_1 \user_module.ram_I.rdata_inv_I[5]  (.A(\user_module.ram_I.rdata_tbuf[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.ram_I.rdata_inv[5] ));
 sky130_fd_sc_hd__inv_1 \user_module.ram_I.rdata_inv_I[6]  (.A(\user_module.ram_I.rdata_tbuf[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.ram_I.rdata_inv[6] ));
 sky130_fd_sc_hd__inv_1 \user_module.ram_I.rdata_inv_I[7]  (.A(\user_module.ram_I.rdata_tbuf[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.ram_I.rdata_inv[7] ));
 sky130_fd_sc_hd__dlxtn_4 \user_module.ram_I.rdata_latch_I[0]  (.D(\user_module.ram_I.rdata_inv[0] ),
    .GATE_N(\user_module.ram_I.rdata_le_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_out[0] ));
 sky130_fd_sc_hd__dlxtn_4 \user_module.ram_I.rdata_latch_I[1]  (.D(\user_module.ram_I.rdata_inv[1] ),
    .GATE_N(\user_module.ram_I.rdata_le_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_out[1] ));
 sky130_fd_sc_hd__dlxtn_4 \user_module.ram_I.rdata_latch_I[2]  (.D(\user_module.ram_I.rdata_inv[2] ),
    .GATE_N(\user_module.ram_I.rdata_le_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_out[2] ));
 sky130_fd_sc_hd__dlxtn_4 \user_module.ram_I.rdata_latch_I[3]  (.D(\user_module.ram_I.rdata_inv[3] ),
    .GATE_N(\user_module.ram_I.rdata_le_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_out[3] ));
 sky130_fd_sc_hd__dlxtn_4 \user_module.ram_I.rdata_latch_I[4]  (.D(\user_module.ram_I.rdata_inv[4] ),
    .GATE_N(\user_module.ram_I.rdata_le_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_out[4] ));
 sky130_fd_sc_hd__dlxtn_4 \user_module.ram_I.rdata_latch_I[5]  (.D(\user_module.ram_I.rdata_inv[5] ),
    .GATE_N(\user_module.ram_I.rdata_le_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_out[5] ));
 sky130_fd_sc_hd__dlxtn_4 \user_module.ram_I.rdata_latch_I[6]  (.D(\user_module.ram_I.rdata_inv[6] ),
    .GATE_N(\user_module.ram_I.rdata_le_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_out[6] ));
 sky130_fd_sc_hd__dlxtn_4 \user_module.ram_I.rdata_latch_I[7]  (.D(\user_module.ram_I.rdata_inv[7] ),
    .GATE_N(\user_module.ram_I.rdata_le_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.eio_out[7] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[0].rdata_mux_I[0]  (.A0(\user_module.ram_I.rdata_sel_loop[0].l_in0_mux[0] ),
    .A1(\user_module.ram_I.rdata_sel_loop[0].l_in1_mux[0] ),
    .A2(\user_module.ram_I.rdata_sel_loop[0].l_in2_mux[0] ),
    .A3(\user_module.ram_I.rdata_sel_loop[0].l_in3_mux[0] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[0].l_out_mux[0] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[0].rdata_mux_I[1]  (.A0(\user_module.ram_I.rdata_sel_loop[0].l_in0_mux[1] ),
    .A1(\user_module.ram_I.rdata_sel_loop[0].l_in1_mux[1] ),
    .A2(\user_module.ram_I.rdata_sel_loop[0].l_in2_mux[1] ),
    .A3(\user_module.ram_I.rdata_sel_loop[0].l_in3_mux[1] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[0].l_out_mux[1] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[0].rdata_mux_I[2]  (.A0(\user_module.ram_I.rdata_sel_loop[0].l_in0_mux[2] ),
    .A1(\user_module.ram_I.rdata_sel_loop[0].l_in1_mux[2] ),
    .A2(\user_module.ram_I.rdata_sel_loop[0].l_in2_mux[2] ),
    .A3(\user_module.ram_I.rdata_sel_loop[0].l_in3_mux[2] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[0].l_out_mux[2] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[0].rdata_mux_I[3]  (.A0(\user_module.ram_I.rdata_sel_loop[0].l_in0_mux[3] ),
    .A1(\user_module.ram_I.rdata_sel_loop[0].l_in1_mux[3] ),
    .A2(\user_module.ram_I.rdata_sel_loop[0].l_in2_mux[3] ),
    .A3(\user_module.ram_I.rdata_sel_loop[0].l_in3_mux[3] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[0].l_out_mux[3] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[0].rdata_mux_I[4]  (.A0(\user_module.ram_I.rdata_sel_loop[0].l_in0_mux[4] ),
    .A1(\user_module.ram_I.rdata_sel_loop[0].l_in1_mux[4] ),
    .A2(\user_module.ram_I.rdata_sel_loop[0].l_in2_mux[4] ),
    .A3(\user_module.ram_I.rdata_sel_loop[0].l_in3_mux[4] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[0].l_out_mux[4] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[0].rdata_mux_I[5]  (.A0(\user_module.ram_I.rdata_sel_loop[0].l_in0_mux[5] ),
    .A1(\user_module.ram_I.rdata_sel_loop[0].l_in1_mux[5] ),
    .A2(\user_module.ram_I.rdata_sel_loop[0].l_in2_mux[5] ),
    .A3(\user_module.ram_I.rdata_sel_loop[0].l_in3_mux[5] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[0].l_out_mux[5] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[0].rdata_mux_I[6]  (.A0(\user_module.ram_I.rdata_sel_loop[0].l_in0_mux[6] ),
    .A1(\user_module.ram_I.rdata_sel_loop[0].l_in1_mux[6] ),
    .A2(\user_module.ram_I.rdata_sel_loop[0].l_in2_mux[6] ),
    .A3(\user_module.ram_I.rdata_sel_loop[0].l_in3_mux[6] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[0].l_out_mux[6] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[0].rdata_mux_I[7]  (.A0(\user_module.ram_I.rdata_sel_loop[0].l_in0_mux[7] ),
    .A1(\user_module.ram_I.rdata_sel_loop[0].l_in1_mux[7] ),
    .A2(\user_module.ram_I.rdata_sel_loop[0].l_in2_mux[7] ),
    .A3(\user_module.ram_I.rdata_sel_loop[0].l_in3_mux[7] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[0].l_out_mux[7] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[0].rdata_tbuf_I[0]  (.A(\user_module.ram_I.rdata_sel_loop[0].l_out_mux[0] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[0] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[0].rdata_tbuf_I[1]  (.A(\user_module.ram_I.rdata_sel_loop[0].l_out_mux[1] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[1] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[0].rdata_tbuf_I[2]  (.A(\user_module.ram_I.rdata_sel_loop[0].l_out_mux[2] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[2] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[0].rdata_tbuf_I[3]  (.A(\user_module.ram_I.rdata_sel_loop[0].l_out_mux[3] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[3] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[0].rdata_tbuf_I[4]  (.A(\user_module.ram_I.rdata_sel_loop[0].l_out_mux[4] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[4] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[0].rdata_tbuf_I[5]  (.A(\user_module.ram_I.rdata_sel_loop[0].l_out_mux[5] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[5] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[0].rdata_tbuf_I[6]  (.A(\user_module.ram_I.rdata_sel_loop[0].l_out_mux[6] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[6] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[0].rdata_tbuf_I[7]  (.A(\user_module.ram_I.rdata_sel_loop[0].l_out_mux[7] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[7] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[12].rdata_mux_I[0]  (.A0(\user_module.ram_I.rdata_sel_loop[12].l_in0_mux[0] ),
    .A1(\user_module.ram_I.rdata_sel_loop[12].l_in1_mux[0] ),
    .A2(\user_module.ram_I.rdata_sel_loop[12].l_in2_mux[0] ),
    .A3(\user_module.ram_I.rdata_sel_loop[12].l_in3_mux[0] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[12].l_out_mux[0] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[12].rdata_mux_I[1]  (.A0(\user_module.ram_I.rdata_sel_loop[12].l_in0_mux[1] ),
    .A1(\user_module.ram_I.rdata_sel_loop[12].l_in1_mux[1] ),
    .A2(\user_module.ram_I.rdata_sel_loop[12].l_in2_mux[1] ),
    .A3(\user_module.ram_I.rdata_sel_loop[12].l_in3_mux[1] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[12].l_out_mux[1] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[12].rdata_mux_I[2]  (.A0(\user_module.ram_I.rdata_sel_loop[12].l_in0_mux[2] ),
    .A1(\user_module.ram_I.rdata_sel_loop[12].l_in1_mux[2] ),
    .A2(\user_module.ram_I.rdata_sel_loop[12].l_in2_mux[2] ),
    .A3(\user_module.ram_I.rdata_sel_loop[12].l_in3_mux[2] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[12].l_out_mux[2] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[12].rdata_mux_I[3]  (.A0(\user_module.ram_I.rdata_sel_loop[12].l_in0_mux[3] ),
    .A1(\user_module.ram_I.rdata_sel_loop[12].l_in1_mux[3] ),
    .A2(\user_module.ram_I.rdata_sel_loop[12].l_in2_mux[3] ),
    .A3(\user_module.ram_I.rdata_sel_loop[12].l_in3_mux[3] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[12].l_out_mux[3] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[12].rdata_mux_I[4]  (.A0(\user_module.ram_I.rdata_sel_loop[12].l_in0_mux[4] ),
    .A1(\user_module.ram_I.rdata_sel_loop[12].l_in1_mux[4] ),
    .A2(\user_module.ram_I.rdata_sel_loop[12].l_in2_mux[4] ),
    .A3(\user_module.ram_I.rdata_sel_loop[12].l_in3_mux[4] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[12].l_out_mux[4] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[12].rdata_mux_I[5]  (.A0(\user_module.ram_I.rdata_sel_loop[12].l_in0_mux[5] ),
    .A1(\user_module.ram_I.rdata_sel_loop[12].l_in1_mux[5] ),
    .A2(\user_module.ram_I.rdata_sel_loop[12].l_in2_mux[5] ),
    .A3(\user_module.ram_I.rdata_sel_loop[12].l_in3_mux[5] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[12].l_out_mux[5] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[12].rdata_mux_I[6]  (.A0(\user_module.ram_I.rdata_sel_loop[12].l_in0_mux[6] ),
    .A1(\user_module.ram_I.rdata_sel_loop[12].l_in1_mux[6] ),
    .A2(\user_module.ram_I.rdata_sel_loop[12].l_in2_mux[6] ),
    .A3(\user_module.ram_I.rdata_sel_loop[12].l_in3_mux[6] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[12].l_out_mux[6] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[12].rdata_mux_I[7]  (.A0(\user_module.ram_I.rdata_sel_loop[12].l_in0_mux[7] ),
    .A1(\user_module.ram_I.rdata_sel_loop[12].l_in1_mux[7] ),
    .A2(\user_module.ram_I.rdata_sel_loop[12].l_in2_mux[7] ),
    .A3(\user_module.ram_I.rdata_sel_loop[12].l_in3_mux[7] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[12].l_out_mux[7] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[12].rdata_tbuf_I[0]  (.A(\user_module.ram_I.rdata_sel_loop[12].l_out_mux[0] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[0] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[12].rdata_tbuf_I[1]  (.A(\user_module.ram_I.rdata_sel_loop[12].l_out_mux[1] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[1] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[12].rdata_tbuf_I[2]  (.A(\user_module.ram_I.rdata_sel_loop[12].l_out_mux[2] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[2] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[12].rdata_tbuf_I[3]  (.A(\user_module.ram_I.rdata_sel_loop[12].l_out_mux[3] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[3] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[12].rdata_tbuf_I[4]  (.A(\user_module.ram_I.rdata_sel_loop[12].l_out_mux[4] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[4] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[12].rdata_tbuf_I[5]  (.A(\user_module.ram_I.rdata_sel_loop[12].l_out_mux[5] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[5] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[12].rdata_tbuf_I[6]  (.A(\user_module.ram_I.rdata_sel_loop[12].l_out_mux[6] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[6] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[12].rdata_tbuf_I[7]  (.A(\user_module.ram_I.rdata_sel_loop[12].l_out_mux[7] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[7] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[4].rdata_mux_I[0]  (.A0(\user_module.ram_I.rdata_sel_loop[4].l_in0_mux[0] ),
    .A1(\user_module.ram_I.rdata_sel_loop[4].l_in1_mux[0] ),
    .A2(\user_module.ram_I.rdata_sel_loop[4].l_in2_mux[0] ),
    .A3(\user_module.ram_I.rdata_sel_loop[4].l_in3_mux[0] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[4].l_out_mux[0] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[4].rdata_mux_I[1]  (.A0(\user_module.ram_I.rdata_sel_loop[4].l_in0_mux[1] ),
    .A1(\user_module.ram_I.rdata_sel_loop[4].l_in1_mux[1] ),
    .A2(\user_module.ram_I.rdata_sel_loop[4].l_in2_mux[1] ),
    .A3(\user_module.ram_I.rdata_sel_loop[4].l_in3_mux[1] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[4].l_out_mux[1] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[4].rdata_mux_I[2]  (.A0(\user_module.ram_I.rdata_sel_loop[4].l_in0_mux[2] ),
    .A1(\user_module.ram_I.rdata_sel_loop[4].l_in1_mux[2] ),
    .A2(\user_module.ram_I.rdata_sel_loop[4].l_in2_mux[2] ),
    .A3(\user_module.ram_I.rdata_sel_loop[4].l_in3_mux[2] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[4].l_out_mux[2] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[4].rdata_mux_I[3]  (.A0(\user_module.ram_I.rdata_sel_loop[4].l_in0_mux[3] ),
    .A1(\user_module.ram_I.rdata_sel_loop[4].l_in1_mux[3] ),
    .A2(\user_module.ram_I.rdata_sel_loop[4].l_in2_mux[3] ),
    .A3(\user_module.ram_I.rdata_sel_loop[4].l_in3_mux[3] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[4].l_out_mux[3] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[4].rdata_mux_I[4]  (.A0(\user_module.ram_I.rdata_sel_loop[4].l_in0_mux[4] ),
    .A1(\user_module.ram_I.rdata_sel_loop[4].l_in1_mux[4] ),
    .A2(\user_module.ram_I.rdata_sel_loop[4].l_in2_mux[4] ),
    .A3(\user_module.ram_I.rdata_sel_loop[4].l_in3_mux[4] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[4].l_out_mux[4] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[4].rdata_mux_I[5]  (.A0(\user_module.ram_I.rdata_sel_loop[4].l_in0_mux[5] ),
    .A1(\user_module.ram_I.rdata_sel_loop[4].l_in1_mux[5] ),
    .A2(\user_module.ram_I.rdata_sel_loop[4].l_in2_mux[5] ),
    .A3(\user_module.ram_I.rdata_sel_loop[4].l_in3_mux[5] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[4].l_out_mux[5] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[4].rdata_mux_I[6]  (.A0(\user_module.ram_I.rdata_sel_loop[4].l_in0_mux[6] ),
    .A1(\user_module.ram_I.rdata_sel_loop[4].l_in1_mux[6] ),
    .A2(\user_module.ram_I.rdata_sel_loop[4].l_in2_mux[6] ),
    .A3(\user_module.ram_I.rdata_sel_loop[4].l_in3_mux[6] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[4].l_out_mux[6] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[4].rdata_mux_I[7]  (.A0(\user_module.ram_I.rdata_sel_loop[4].l_in0_mux[7] ),
    .A1(\user_module.ram_I.rdata_sel_loop[4].l_in1_mux[7] ),
    .A2(\user_module.ram_I.rdata_sel_loop[4].l_in2_mux[7] ),
    .A3(\user_module.ram_I.rdata_sel_loop[4].l_in3_mux[7] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[4].l_out_mux[7] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[4].rdata_tbuf_I[0]  (.A(\user_module.ram_I.rdata_sel_loop[4].l_out_mux[0] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[0] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[4].rdata_tbuf_I[1]  (.A(\user_module.ram_I.rdata_sel_loop[4].l_out_mux[1] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[1] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[4].rdata_tbuf_I[2]  (.A(\user_module.ram_I.rdata_sel_loop[4].l_out_mux[2] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[2] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[4].rdata_tbuf_I[3]  (.A(\user_module.ram_I.rdata_sel_loop[4].l_out_mux[3] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[3] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[4].rdata_tbuf_I[4]  (.A(\user_module.ram_I.rdata_sel_loop[4].l_out_mux[4] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[4] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[4].rdata_tbuf_I[5]  (.A(\user_module.ram_I.rdata_sel_loop[4].l_out_mux[5] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[5] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[4].rdata_tbuf_I[6]  (.A(\user_module.ram_I.rdata_sel_loop[4].l_out_mux[6] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[6] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[4].rdata_tbuf_I[7]  (.A(\user_module.ram_I.rdata_sel_loop[4].l_out_mux[7] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[7] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[8].rdata_mux_I[0]  (.A0(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[0] ),
    .A1(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[0] ),
    .A2(\user_module.ram_I.rdata_sel_loop[8].l_in2_mux[0] ),
    .A3(\user_module.ram_I.rdata_sel_loop[8].l_in3_mux[0] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[8].l_out_mux[0] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[8].rdata_mux_I[1]  (.A0(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[1] ),
    .A1(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[1] ),
    .A2(\user_module.ram_I.rdata_sel_loop[8].l_in2_mux[1] ),
    .A3(\user_module.ram_I.rdata_sel_loop[8].l_in3_mux[1] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[8].l_out_mux[1] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[8].rdata_mux_I[2]  (.A0(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[2] ),
    .A1(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[2] ),
    .A2(\user_module.ram_I.rdata_sel_loop[8].l_in2_mux[2] ),
    .A3(\user_module.ram_I.rdata_sel_loop[8].l_in3_mux[2] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[8].l_out_mux[2] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[8].rdata_mux_I[3]  (.A0(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[3] ),
    .A1(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[3] ),
    .A2(\user_module.ram_I.rdata_sel_loop[8].l_in2_mux[3] ),
    .A3(\user_module.ram_I.rdata_sel_loop[8].l_in3_mux[3] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[8].l_out_mux[3] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[8].rdata_mux_I[4]  (.A0(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[4] ),
    .A1(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[4] ),
    .A2(\user_module.ram_I.rdata_sel_loop[8].l_in2_mux[4] ),
    .A3(\user_module.ram_I.rdata_sel_loop[8].l_in3_mux[4] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[8].l_out_mux[4] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[8].rdata_mux_I[5]  (.A0(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[5] ),
    .A1(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[5] ),
    .A2(\user_module.ram_I.rdata_sel_loop[8].l_in2_mux[5] ),
    .A3(\user_module.ram_I.rdata_sel_loop[8].l_in3_mux[5] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[8].l_out_mux[5] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[8].rdata_mux_I[6]  (.A0(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[6] ),
    .A1(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[6] ),
    .A2(\user_module.ram_I.rdata_sel_loop[8].l_in2_mux[6] ),
    .A3(\user_module.ram_I.rdata_sel_loop[8].l_in3_mux[6] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[8].l_out_mux[6] ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.rdata_sel_loop[8].rdata_mux_I[7]  (.A0(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[7] ),
    .A1(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[7] ),
    .A2(\user_module.ram_I.rdata_sel_loop[8].l_in2_mux[7] ),
    .A3(\user_module.ram_I.rdata_sel_loop[8].l_in3_mux[7] ),
    .S0(\user_module.ram_I.raddr_r[0] ),
    .S1(\user_module.ram_I.raddr_r[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.rdata_sel_loop[8].l_out_mux[7] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[8].rdata_tbuf_I[0]  (.A(\user_module.ram_I.rdata_sel_loop[8].l_out_mux[0] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[0] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[8].rdata_tbuf_I[1]  (.A(\user_module.ram_I.rdata_sel_loop[8].l_out_mux[1] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[1] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[8].rdata_tbuf_I[2]  (.A(\user_module.ram_I.rdata_sel_loop[8].l_out_mux[2] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[2] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[8].rdata_tbuf_I[3]  (.A(\user_module.ram_I.rdata_sel_loop[8].l_out_mux[3] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[3] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[8].rdata_tbuf_I[4]  (.A(\user_module.ram_I.rdata_sel_loop[8].l_out_mux[4] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[4] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[8].rdata_tbuf_I[5]  (.A(\user_module.ram_I.rdata_sel_loop[8].l_out_mux[5] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[5] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[8].rdata_tbuf_I[6]  (.A(\user_module.ram_I.rdata_sel_loop[8].l_out_mux[6] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[6] ));
 sky130_fd_sc_hd__einvp_2 \user_module.ram_I.rdata_sel_loop[8].rdata_tbuf_I[7]  (.A(\user_module.ram_I.rdata_sel_loop[8].l_out_mux[7] ),
    .TE(\user_module.ram_I.raddr_dec_I.out[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Z(\user_module.ram_I.rdata_tbuf[7] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.ram_I.re_reg_I  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.re_r ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[0].store_cell_I[0]  (.D(\user_module.ram_I.store_in[0] ),
    .GATE(\user_module.ram_I.store_gate[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in0_mux[0] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[0].store_cell_I[1]  (.D(\user_module.ram_I.store_in[1] ),
    .GATE(\user_module.ram_I.store_gate[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in0_mux[1] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[0].store_cell_I[2]  (.D(\user_module.ram_I.store_in[2] ),
    .GATE(\user_module.ram_I.store_gate[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in0_mux[2] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[0].store_cell_I[3]  (.D(\user_module.ram_I.store_in[3] ),
    .GATE(\user_module.ram_I.store_gate[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in0_mux[3] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[0].store_cell_I[4]  (.D(\user_module.ram_I.store_in[4] ),
    .GATE(\user_module.ram_I.store_gate[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in0_mux[4] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[0].store_cell_I[5]  (.D(\user_module.ram_I.store_in[5] ),
    .GATE(\user_module.ram_I.store_gate[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in0_mux[5] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[0].store_cell_I[6]  (.D(\user_module.ram_I.store_in[6] ),
    .GATE(\user_module.ram_I.store_gate[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in0_mux[6] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[0].store_cell_I[7]  (.D(\user_module.ram_I.store_in[7] ),
    .GATE(\user_module.ram_I.store_gate[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in0_mux[7] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[10].store_cell_I[0]  (.D(\user_module.ram_I.store_in[0] ),
    .GATE(\user_module.ram_I.store_gate[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in2_mux[0] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[10].store_cell_I[1]  (.D(\user_module.ram_I.store_in[1] ),
    .GATE(\user_module.ram_I.store_gate[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in2_mux[1] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[10].store_cell_I[2]  (.D(\user_module.ram_I.store_in[2] ),
    .GATE(\user_module.ram_I.store_gate[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in2_mux[2] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[10].store_cell_I[3]  (.D(\user_module.ram_I.store_in[3] ),
    .GATE(\user_module.ram_I.store_gate[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in2_mux[3] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[10].store_cell_I[4]  (.D(\user_module.ram_I.store_in[4] ),
    .GATE(\user_module.ram_I.store_gate[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in2_mux[4] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[10].store_cell_I[5]  (.D(\user_module.ram_I.store_in[5] ),
    .GATE(\user_module.ram_I.store_gate[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in2_mux[5] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[10].store_cell_I[6]  (.D(\user_module.ram_I.store_in[6] ),
    .GATE(\user_module.ram_I.store_gate[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in2_mux[6] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[10].store_cell_I[7]  (.D(\user_module.ram_I.store_in[7] ),
    .GATE(\user_module.ram_I.store_gate[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in2_mux[7] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[11].store_cell_I[0]  (.D(\user_module.ram_I.store_in[0] ),
    .GATE(\user_module.ram_I.store_gate[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in3_mux[0] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[11].store_cell_I[1]  (.D(\user_module.ram_I.store_in[1] ),
    .GATE(\user_module.ram_I.store_gate[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in3_mux[1] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[11].store_cell_I[2]  (.D(\user_module.ram_I.store_in[2] ),
    .GATE(\user_module.ram_I.store_gate[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in3_mux[2] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[11].store_cell_I[3]  (.D(\user_module.ram_I.store_in[3] ),
    .GATE(\user_module.ram_I.store_gate[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in3_mux[3] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[11].store_cell_I[4]  (.D(\user_module.ram_I.store_in[4] ),
    .GATE(\user_module.ram_I.store_gate[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in3_mux[4] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[11].store_cell_I[5]  (.D(\user_module.ram_I.store_in[5] ),
    .GATE(\user_module.ram_I.store_gate[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in3_mux[5] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[11].store_cell_I[6]  (.D(\user_module.ram_I.store_in[6] ),
    .GATE(\user_module.ram_I.store_gate[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in3_mux[6] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[11].store_cell_I[7]  (.D(\user_module.ram_I.store_in[7] ),
    .GATE(\user_module.ram_I.store_gate[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in3_mux[7] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[12].store_cell_I[0]  (.D(\user_module.ram_I.store_in[0] ),
    .GATE(\user_module.ram_I.store_gate[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in0_mux[0] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[12].store_cell_I[1]  (.D(\user_module.ram_I.store_in[1] ),
    .GATE(\user_module.ram_I.store_gate[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in0_mux[1] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[12].store_cell_I[2]  (.D(\user_module.ram_I.store_in[2] ),
    .GATE(\user_module.ram_I.store_gate[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in0_mux[2] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[12].store_cell_I[3]  (.D(\user_module.ram_I.store_in[3] ),
    .GATE(\user_module.ram_I.store_gate[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in0_mux[3] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[12].store_cell_I[4]  (.D(\user_module.ram_I.store_in[4] ),
    .GATE(\user_module.ram_I.store_gate[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in0_mux[4] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[12].store_cell_I[5]  (.D(\user_module.ram_I.store_in[5] ),
    .GATE(\user_module.ram_I.store_gate[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in0_mux[5] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[12].store_cell_I[6]  (.D(\user_module.ram_I.store_in[6] ),
    .GATE(\user_module.ram_I.store_gate[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in0_mux[6] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[12].store_cell_I[7]  (.D(\user_module.ram_I.store_in[7] ),
    .GATE(\user_module.ram_I.store_gate[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in0_mux[7] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[13].store_cell_I[0]  (.D(\user_module.ram_I.store_in[0] ),
    .GATE(\user_module.ram_I.store_gate[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in1_mux[0] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[13].store_cell_I[1]  (.D(\user_module.ram_I.store_in[1] ),
    .GATE(\user_module.ram_I.store_gate[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in1_mux[1] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[13].store_cell_I[2]  (.D(\user_module.ram_I.store_in[2] ),
    .GATE(\user_module.ram_I.store_gate[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in1_mux[2] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[13].store_cell_I[3]  (.D(\user_module.ram_I.store_in[3] ),
    .GATE(\user_module.ram_I.store_gate[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in1_mux[3] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[13].store_cell_I[4]  (.D(\user_module.ram_I.store_in[4] ),
    .GATE(\user_module.ram_I.store_gate[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in1_mux[4] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[13].store_cell_I[5]  (.D(\user_module.ram_I.store_in[5] ),
    .GATE(\user_module.ram_I.store_gate[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in1_mux[5] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[13].store_cell_I[6]  (.D(\user_module.ram_I.store_in[6] ),
    .GATE(\user_module.ram_I.store_gate[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in1_mux[6] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[13].store_cell_I[7]  (.D(\user_module.ram_I.store_in[7] ),
    .GATE(\user_module.ram_I.store_gate[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in1_mux[7] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[14].store_cell_I[0]  (.D(\user_module.ram_I.store_in[0] ),
    .GATE(\user_module.ram_I.store_gate[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in2_mux[0] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[14].store_cell_I[1]  (.D(\user_module.ram_I.store_in[1] ),
    .GATE(\user_module.ram_I.store_gate[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in2_mux[1] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[14].store_cell_I[2]  (.D(\user_module.ram_I.store_in[2] ),
    .GATE(\user_module.ram_I.store_gate[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in2_mux[2] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[14].store_cell_I[3]  (.D(\user_module.ram_I.store_in[3] ),
    .GATE(\user_module.ram_I.store_gate[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in2_mux[3] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[14].store_cell_I[4]  (.D(\user_module.ram_I.store_in[4] ),
    .GATE(\user_module.ram_I.store_gate[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in2_mux[4] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[14].store_cell_I[5]  (.D(\user_module.ram_I.store_in[5] ),
    .GATE(\user_module.ram_I.store_gate[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in2_mux[5] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[14].store_cell_I[6]  (.D(\user_module.ram_I.store_in[6] ),
    .GATE(\user_module.ram_I.store_gate[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in2_mux[6] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[14].store_cell_I[7]  (.D(\user_module.ram_I.store_in[7] ),
    .GATE(\user_module.ram_I.store_gate[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in2_mux[7] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[15].store_cell_I[0]  (.D(\user_module.ram_I.store_in[0] ),
    .GATE(\user_module.ram_I.store_gate[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in3_mux[0] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[15].store_cell_I[1]  (.D(\user_module.ram_I.store_in[1] ),
    .GATE(\user_module.ram_I.store_gate[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in3_mux[1] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[15].store_cell_I[2]  (.D(\user_module.ram_I.store_in[2] ),
    .GATE(\user_module.ram_I.store_gate[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in3_mux[2] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[15].store_cell_I[3]  (.D(\user_module.ram_I.store_in[3] ),
    .GATE(\user_module.ram_I.store_gate[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in3_mux[3] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[15].store_cell_I[4]  (.D(\user_module.ram_I.store_in[4] ),
    .GATE(\user_module.ram_I.store_gate[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in3_mux[4] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[15].store_cell_I[5]  (.D(\user_module.ram_I.store_in[5] ),
    .GATE(\user_module.ram_I.store_gate[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in3_mux[5] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[15].store_cell_I[6]  (.D(\user_module.ram_I.store_in[6] ),
    .GATE(\user_module.ram_I.store_gate[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in3_mux[6] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[15].store_cell_I[7]  (.D(\user_module.ram_I.store_in[7] ),
    .GATE(\user_module.ram_I.store_gate[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[12].l_in3_mux[7] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[1].store_cell_I[0]  (.D(\user_module.ram_I.store_in[0] ),
    .GATE(\user_module.ram_I.store_gate[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in1_mux[0] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[1].store_cell_I[1]  (.D(\user_module.ram_I.store_in[1] ),
    .GATE(\user_module.ram_I.store_gate[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in1_mux[1] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[1].store_cell_I[2]  (.D(\user_module.ram_I.store_in[2] ),
    .GATE(\user_module.ram_I.store_gate[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in1_mux[2] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[1].store_cell_I[3]  (.D(\user_module.ram_I.store_in[3] ),
    .GATE(\user_module.ram_I.store_gate[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in1_mux[3] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[1].store_cell_I[4]  (.D(\user_module.ram_I.store_in[4] ),
    .GATE(\user_module.ram_I.store_gate[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in1_mux[4] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[1].store_cell_I[5]  (.D(\user_module.ram_I.store_in[5] ),
    .GATE(\user_module.ram_I.store_gate[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in1_mux[5] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[1].store_cell_I[6]  (.D(\user_module.ram_I.store_in[6] ),
    .GATE(\user_module.ram_I.store_gate[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in1_mux[6] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[1].store_cell_I[7]  (.D(\user_module.ram_I.store_in[7] ),
    .GATE(\user_module.ram_I.store_gate[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in1_mux[7] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[2].store_cell_I[0]  (.D(\user_module.ram_I.store_in[0] ),
    .GATE(\user_module.ram_I.store_gate[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in2_mux[0] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[2].store_cell_I[1]  (.D(\user_module.ram_I.store_in[1] ),
    .GATE(\user_module.ram_I.store_gate[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in2_mux[1] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[2].store_cell_I[2]  (.D(\user_module.ram_I.store_in[2] ),
    .GATE(\user_module.ram_I.store_gate[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in2_mux[2] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[2].store_cell_I[3]  (.D(\user_module.ram_I.store_in[3] ),
    .GATE(\user_module.ram_I.store_gate[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in2_mux[3] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[2].store_cell_I[4]  (.D(\user_module.ram_I.store_in[4] ),
    .GATE(\user_module.ram_I.store_gate[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in2_mux[4] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[2].store_cell_I[5]  (.D(\user_module.ram_I.store_in[5] ),
    .GATE(\user_module.ram_I.store_gate[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in2_mux[5] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[2].store_cell_I[6]  (.D(\user_module.ram_I.store_in[6] ),
    .GATE(\user_module.ram_I.store_gate[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in2_mux[6] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[2].store_cell_I[7]  (.D(\user_module.ram_I.store_in[7] ),
    .GATE(\user_module.ram_I.store_gate[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in2_mux[7] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[3].store_cell_I[0]  (.D(\user_module.ram_I.store_in[0] ),
    .GATE(\user_module.ram_I.store_gate[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in3_mux[0] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[3].store_cell_I[1]  (.D(\user_module.ram_I.store_in[1] ),
    .GATE(\user_module.ram_I.store_gate[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in3_mux[1] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[3].store_cell_I[2]  (.D(\user_module.ram_I.store_in[2] ),
    .GATE(\user_module.ram_I.store_gate[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in3_mux[2] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[3].store_cell_I[3]  (.D(\user_module.ram_I.store_in[3] ),
    .GATE(\user_module.ram_I.store_gate[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in3_mux[3] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[3].store_cell_I[4]  (.D(\user_module.ram_I.store_in[4] ),
    .GATE(\user_module.ram_I.store_gate[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in3_mux[4] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[3].store_cell_I[5]  (.D(\user_module.ram_I.store_in[5] ),
    .GATE(\user_module.ram_I.store_gate[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in3_mux[5] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[3].store_cell_I[6]  (.D(\user_module.ram_I.store_in[6] ),
    .GATE(\user_module.ram_I.store_gate[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in3_mux[6] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[3].store_cell_I[7]  (.D(\user_module.ram_I.store_in[7] ),
    .GATE(\user_module.ram_I.store_gate[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[0].l_in3_mux[7] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[4].store_cell_I[0]  (.D(\user_module.ram_I.store_in[0] ),
    .GATE(\user_module.ram_I.store_gate[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in0_mux[0] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[4].store_cell_I[1]  (.D(\user_module.ram_I.store_in[1] ),
    .GATE(\user_module.ram_I.store_gate[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in0_mux[1] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[4].store_cell_I[2]  (.D(\user_module.ram_I.store_in[2] ),
    .GATE(\user_module.ram_I.store_gate[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in0_mux[2] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[4].store_cell_I[3]  (.D(\user_module.ram_I.store_in[3] ),
    .GATE(\user_module.ram_I.store_gate[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in0_mux[3] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[4].store_cell_I[4]  (.D(\user_module.ram_I.store_in[4] ),
    .GATE(\user_module.ram_I.store_gate[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in0_mux[4] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[4].store_cell_I[5]  (.D(\user_module.ram_I.store_in[5] ),
    .GATE(\user_module.ram_I.store_gate[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in0_mux[5] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[4].store_cell_I[6]  (.D(\user_module.ram_I.store_in[6] ),
    .GATE(\user_module.ram_I.store_gate[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in0_mux[6] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[4].store_cell_I[7]  (.D(\user_module.ram_I.store_in[7] ),
    .GATE(\user_module.ram_I.store_gate[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in0_mux[7] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[5].store_cell_I[0]  (.D(\user_module.ram_I.store_in[0] ),
    .GATE(\user_module.ram_I.store_gate[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in1_mux[0] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[5].store_cell_I[1]  (.D(\user_module.ram_I.store_in[1] ),
    .GATE(\user_module.ram_I.store_gate[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in1_mux[1] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[5].store_cell_I[2]  (.D(\user_module.ram_I.store_in[2] ),
    .GATE(\user_module.ram_I.store_gate[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in1_mux[2] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[5].store_cell_I[3]  (.D(\user_module.ram_I.store_in[3] ),
    .GATE(\user_module.ram_I.store_gate[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in1_mux[3] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[5].store_cell_I[4]  (.D(\user_module.ram_I.store_in[4] ),
    .GATE(\user_module.ram_I.store_gate[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in1_mux[4] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[5].store_cell_I[5]  (.D(\user_module.ram_I.store_in[5] ),
    .GATE(\user_module.ram_I.store_gate[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in1_mux[5] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[5].store_cell_I[6]  (.D(\user_module.ram_I.store_in[6] ),
    .GATE(\user_module.ram_I.store_gate[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in1_mux[6] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[5].store_cell_I[7]  (.D(\user_module.ram_I.store_in[7] ),
    .GATE(\user_module.ram_I.store_gate[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in1_mux[7] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[6].store_cell_I[0]  (.D(\user_module.ram_I.store_in[0] ),
    .GATE(\user_module.ram_I.store_gate[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in2_mux[0] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[6].store_cell_I[1]  (.D(\user_module.ram_I.store_in[1] ),
    .GATE(\user_module.ram_I.store_gate[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in2_mux[1] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[6].store_cell_I[2]  (.D(\user_module.ram_I.store_in[2] ),
    .GATE(\user_module.ram_I.store_gate[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in2_mux[2] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[6].store_cell_I[3]  (.D(\user_module.ram_I.store_in[3] ),
    .GATE(\user_module.ram_I.store_gate[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in2_mux[3] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[6].store_cell_I[4]  (.D(\user_module.ram_I.store_in[4] ),
    .GATE(\user_module.ram_I.store_gate[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in2_mux[4] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[6].store_cell_I[5]  (.D(\user_module.ram_I.store_in[5] ),
    .GATE(\user_module.ram_I.store_gate[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in2_mux[5] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[6].store_cell_I[6]  (.D(\user_module.ram_I.store_in[6] ),
    .GATE(\user_module.ram_I.store_gate[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in2_mux[6] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[6].store_cell_I[7]  (.D(\user_module.ram_I.store_in[7] ),
    .GATE(\user_module.ram_I.store_gate[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in2_mux[7] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[7].store_cell_I[0]  (.D(\user_module.ram_I.store_in[0] ),
    .GATE(\user_module.ram_I.store_gate[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in3_mux[0] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[7].store_cell_I[1]  (.D(\user_module.ram_I.store_in[1] ),
    .GATE(\user_module.ram_I.store_gate[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in3_mux[1] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[7].store_cell_I[2]  (.D(\user_module.ram_I.store_in[2] ),
    .GATE(\user_module.ram_I.store_gate[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in3_mux[2] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[7].store_cell_I[3]  (.D(\user_module.ram_I.store_in[3] ),
    .GATE(\user_module.ram_I.store_gate[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in3_mux[3] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[7].store_cell_I[4]  (.D(\user_module.ram_I.store_in[4] ),
    .GATE(\user_module.ram_I.store_gate[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in3_mux[4] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[7].store_cell_I[5]  (.D(\user_module.ram_I.store_in[5] ),
    .GATE(\user_module.ram_I.store_gate[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in3_mux[5] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[7].store_cell_I[6]  (.D(\user_module.ram_I.store_in[6] ),
    .GATE(\user_module.ram_I.store_gate[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in3_mux[6] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[7].store_cell_I[7]  (.D(\user_module.ram_I.store_in[7] ),
    .GATE(\user_module.ram_I.store_gate[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[4].l_in3_mux[7] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[8].store_cell_I[0]  (.D(\user_module.ram_I.store_in[0] ),
    .GATE(\user_module.ram_I.store_gate[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[0] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[8].store_cell_I[1]  (.D(\user_module.ram_I.store_in[1] ),
    .GATE(\user_module.ram_I.store_gate[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[1] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[8].store_cell_I[2]  (.D(\user_module.ram_I.store_in[2] ),
    .GATE(\user_module.ram_I.store_gate[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[2] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[8].store_cell_I[3]  (.D(\user_module.ram_I.store_in[3] ),
    .GATE(\user_module.ram_I.store_gate[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[3] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[8].store_cell_I[4]  (.D(\user_module.ram_I.store_in[4] ),
    .GATE(\user_module.ram_I.store_gate[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[4] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[8].store_cell_I[5]  (.D(\user_module.ram_I.store_in[5] ),
    .GATE(\user_module.ram_I.store_gate[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[5] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[8].store_cell_I[6]  (.D(\user_module.ram_I.store_in[6] ),
    .GATE(\user_module.ram_I.store_gate[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[6] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[8].store_cell_I[7]  (.D(\user_module.ram_I.store_in[7] ),
    .GATE(\user_module.ram_I.store_gate[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in0_mux[7] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[9].store_cell_I[0]  (.D(\user_module.ram_I.store_in[0] ),
    .GATE(\user_module.ram_I.store_gate[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[0] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[9].store_cell_I[1]  (.D(\user_module.ram_I.store_in[1] ),
    .GATE(\user_module.ram_I.store_gate[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[1] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[9].store_cell_I[2]  (.D(\user_module.ram_I.store_in[2] ),
    .GATE(\user_module.ram_I.store_gate[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[2] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[9].store_cell_I[3]  (.D(\user_module.ram_I.store_in[3] ),
    .GATE(\user_module.ram_I.store_gate[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[3] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[9].store_cell_I[4]  (.D(\user_module.ram_I.store_in[4] ),
    .GATE(\user_module.ram_I.store_gate[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[4] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[9].store_cell_I[5]  (.D(\user_module.ram_I.store_in[5] ),
    .GATE(\user_module.ram_I.store_gate[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[5] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[9].store_cell_I[6]  (.D(\user_module.ram_I.store_in[6] ),
    .GATE(\user_module.ram_I.store_gate[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[6] ));
 sky130_fd_sc_hd__dlxtp_1 \user_module.ram_I.store_cell_loop[9].store_cell_I[7]  (.D(\user_module.ram_I.store_in[7] ),
    .GATE(\user_module.ram_I.store_gate[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.rdata_sel_loop[8].l_in1_mux[7] ));
 sky130_fd_sc_hd__nor4_1 \user_module.ram_I.waddr_dec_I.dec_4_0_I  (.A(\user_module.ram_I.waddr_dec_I.in[0] ),
    .B(\user_module.ram_I.waddr_dec_I.in[1] ),
    .C(\user_module.ram_I.waddr_dec_I.in[2] ),
    .D(\user_module.ram_I.waddr_dec_I.in[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.ram_I.waddr_dec[0] ));
 sky130_fd_sc_hd__and4bb_1 \user_module.ram_I.waddr_dec_I.dec_4_10_I  (.A_N(\user_module.ram_I.waddr_dec_I.in[0] ),
    .B_N(\user_module.ram_I.waddr_dec_I.in[2] ),
    .C(\user_module.ram_I.waddr_dec_I.in[1] ),
    .D(\user_module.ram_I.waddr_dec_I.in[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.waddr_dec[10] ));
 sky130_fd_sc_hd__and4b_1 \user_module.ram_I.waddr_dec_I.dec_4_11_I  (.A_N(\user_module.ram_I.waddr_dec_I.in[2] ),
    .B(\user_module.ram_I.waddr_dec_I.in[0] ),
    .C(\user_module.ram_I.waddr_dec_I.in[1] ),
    .D(\user_module.ram_I.waddr_dec_I.in[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.waddr_dec[11] ));
 sky130_fd_sc_hd__and4bb_1 \user_module.ram_I.waddr_dec_I.dec_4_12_I  (.A_N(\user_module.ram_I.waddr_dec_I.in[0] ),
    .B_N(\user_module.ram_I.waddr_dec_I.in[1] ),
    .C(\user_module.ram_I.waddr_dec_I.in[2] ),
    .D(\user_module.ram_I.waddr_dec_I.in[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.waddr_dec[12] ));
 sky130_fd_sc_hd__and4b_1 \user_module.ram_I.waddr_dec_I.dec_4_13_I  (.A_N(\user_module.ram_I.waddr_dec_I.in[1] ),
    .B(\user_module.ram_I.waddr_dec_I.in[0] ),
    .C(\user_module.ram_I.waddr_dec_I.in[2] ),
    .D(\user_module.ram_I.waddr_dec_I.in[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.waddr_dec[13] ));
 sky130_fd_sc_hd__and4b_1 \user_module.ram_I.waddr_dec_I.dec_4_14_I  (.A_N(\user_module.ram_I.waddr_dec_I.in[0] ),
    .B(\user_module.ram_I.waddr_dec_I.in[1] ),
    .C(\user_module.ram_I.waddr_dec_I.in[2] ),
    .D(\user_module.ram_I.waddr_dec_I.in[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.waddr_dec[14] ));
 sky130_fd_sc_hd__and4_1 \user_module.ram_I.waddr_dec_I.dec_4_15_I  (.A(\user_module.ram_I.waddr_dec_I.in[0] ),
    .B(\user_module.ram_I.waddr_dec_I.in[1] ),
    .C(\user_module.ram_I.waddr_dec_I.in[2] ),
    .D(\user_module.ram_I.waddr_dec_I.in[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.waddr_dec[15] ));
 sky130_fd_sc_hd__nor4b_1 \user_module.ram_I.waddr_dec_I.dec_4_1_I  (.A(\user_module.ram_I.waddr_dec_I.in[1] ),
    .B(\user_module.ram_I.waddr_dec_I.in[2] ),
    .C(\user_module.ram_I.waddr_dec_I.in[3] ),
    .D_N(\user_module.ram_I.waddr_dec_I.in[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.ram_I.waddr_dec[1] ));
 sky130_fd_sc_hd__nor4b_1 \user_module.ram_I.waddr_dec_I.dec_4_2_I  (.A(\user_module.ram_I.waddr_dec_I.in[0] ),
    .B(\user_module.ram_I.waddr_dec_I.in[2] ),
    .C(\user_module.ram_I.waddr_dec_I.in[3] ),
    .D_N(\user_module.ram_I.waddr_dec_I.in[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.ram_I.waddr_dec[2] ));
 sky130_fd_sc_hd__and4bb_1 \user_module.ram_I.waddr_dec_I.dec_4_3_I  (.A_N(\user_module.ram_I.waddr_dec_I.in[2] ),
    .B_N(\user_module.ram_I.waddr_dec_I.in[3] ),
    .C(\user_module.ram_I.waddr_dec_I.in[0] ),
    .D(\user_module.ram_I.waddr_dec_I.in[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.waddr_dec[3] ));
 sky130_fd_sc_hd__nor4b_1 \user_module.ram_I.waddr_dec_I.dec_4_4_I  (.A(\user_module.ram_I.waddr_dec_I.in[0] ),
    .B(\user_module.ram_I.waddr_dec_I.in[1] ),
    .C(\user_module.ram_I.waddr_dec_I.in[3] ),
    .D_N(\user_module.ram_I.waddr_dec_I.in[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.ram_I.waddr_dec[4] ));
 sky130_fd_sc_hd__and4bb_1 \user_module.ram_I.waddr_dec_I.dec_4_5_I  (.A_N(\user_module.ram_I.waddr_dec_I.in[1] ),
    .B_N(\user_module.ram_I.waddr_dec_I.in[3] ),
    .C(\user_module.ram_I.waddr_dec_I.in[0] ),
    .D(\user_module.ram_I.waddr_dec_I.in[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.waddr_dec[5] ));
 sky130_fd_sc_hd__and4bb_1 \user_module.ram_I.waddr_dec_I.dec_4_6_I  (.A_N(\user_module.ram_I.waddr_dec_I.in[0] ),
    .B_N(\user_module.ram_I.waddr_dec_I.in[3] ),
    .C(\user_module.ram_I.waddr_dec_I.in[1] ),
    .D(\user_module.ram_I.waddr_dec_I.in[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.waddr_dec[6] ));
 sky130_fd_sc_hd__and4b_1 \user_module.ram_I.waddr_dec_I.dec_4_7_I  (.A_N(\user_module.ram_I.waddr_dec_I.in[3] ),
    .B(\user_module.ram_I.waddr_dec_I.in[0] ),
    .C(\user_module.ram_I.waddr_dec_I.in[1] ),
    .D(\user_module.ram_I.waddr_dec_I.in[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.waddr_dec[7] ));
 sky130_fd_sc_hd__nor4b_1 \user_module.ram_I.waddr_dec_I.dec_4_8_I  (.A(\user_module.ram_I.waddr_dec_I.in[0] ),
    .B(\user_module.ram_I.waddr_dec_I.in[1] ),
    .C(\user_module.ram_I.waddr_dec_I.in[2] ),
    .D_N(\user_module.ram_I.waddr_dec_I.in[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\user_module.ram_I.waddr_dec[8] ));
 sky130_fd_sc_hd__and4bb_1 \user_module.ram_I.waddr_dec_I.dec_4_9_I  (.A_N(\user_module.ram_I.waddr_dec_I.in[1] ),
    .B_N(\user_module.ram_I.waddr_dec_I.in[2] ),
    .C(\user_module.ram_I.waddr_dec_I.in[0] ),
    .D(\user_module.ram_I.waddr_dec_I.in[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.waddr_dec[9] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.ram_I.waddr_reg_I[0]  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.waddr_dec_I.in[0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.ram_I.waddr_reg_I[1]  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.waddr_dec_I.in[1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.ram_I.waddr_reg_I[2]  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.waddr_dec_I.in[2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.ram_I.waddr_reg_I[3]  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.waddr_dec_I.in[3] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.ram_I.wdata_reg_I[0]  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.store_in[0] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.ram_I.wdata_reg_I[1]  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.store_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.ram_I.wdata_reg_I[2]  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.store_in[2] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.ram_I.wdata_reg_I[3]  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.store_in[3] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.ram_I.wdata_reg_I[4]  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.store_in[4] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.ram_I.wdata_reg_I[5]  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.store_in[5] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.ram_I.wdata_reg_I[6]  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.store_in[6] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.ram_I.wdata_reg_I[7]  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.store_in[7] ));
 sky130_fd_sc_hd__dfxtp_1 \user_module.ram_I.we_reg_I  (.CLK(\user_module.clk_slow ),
    .D(\user_module.eio_in[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\user_module.ram_I.we_r ));
 sky130_fd_sc_hd__mux4_1 \user_module.ram_I.wpulse_I.clk_dly_I  (.A0(\user_module.ram_I.wpulse_I.clk_dly_chain[1] ),
    .A1(\user_module.ram_I.wpulse_I.clk_dly_chain[3] ),
    .A2(\user_module.ram_I.wpulse_I.clk_dly_chain[5] ),
    .A3(\user_module.ram_I.wpulse_I.clk_dly_chain[7] ),
    .S0(_05_),
    .S1(_06_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.wpulse_I.clk_dly ));
 sky130_fd_sc_hd__clkdlybuf4s25_1 \user_module.ram_I.wpulse_I.clk_dly_chain_I[0]  (.A(\user_module.clk_slow ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.wpulse_I.clk_dly_chain[1] ));
 sky130_fd_sc_hd__clkdlybuf4s25_1 \user_module.ram_I.wpulse_I.clk_dly_chain_I[1]  (.A(\user_module.ram_I.wpulse_I.clk_dly_chain[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.wpulse_I.clk_dly_chain[2] ));
 sky130_fd_sc_hd__clkdlybuf4s25_1 \user_module.ram_I.wpulse_I.clk_dly_chain_I[2]  (.A(\user_module.ram_I.wpulse_I.clk_dly_chain[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.wpulse_I.clk_dly_chain[3] ));
 sky130_fd_sc_hd__clkdlybuf4s25_1 \user_module.ram_I.wpulse_I.clk_dly_chain_I[3]  (.A(\user_module.ram_I.wpulse_I.clk_dly_chain[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.wpulse_I.clk_dly_chain[4] ));
 sky130_fd_sc_hd__clkdlybuf4s25_1 \user_module.ram_I.wpulse_I.clk_dly_chain_I[4]  (.A(\user_module.ram_I.wpulse_I.clk_dly_chain[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.wpulse_I.clk_dly_chain[5] ));
 sky130_fd_sc_hd__clkdlybuf4s25_1 \user_module.ram_I.wpulse_I.clk_dly_chain_I[5]  (.A(\user_module.ram_I.wpulse_I.clk_dly_chain[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.wpulse_I.clk_dly_chain[6] ));
 sky130_fd_sc_hd__clkdlybuf4s25_1 \user_module.ram_I.wpulse_I.clk_dly_chain_I[6]  (.A(\user_module.ram_I.wpulse_I.clk_dly_chain[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.wpulse_I.clk_dly_chain[7] ));
 sky130_fd_sc_hd__and3b_4 \user_module.ram_I.wpulse_I.pulse_I  (.A_N(\user_module.clk_slow ),
    .B(\user_module.ram_I.wpulse_I.clk_dly ),
    .C(\user_module.ram_I.we_r ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.wpulse_I.pulse ));
 sky130_fd_sc_hd__and2_4 \user_module.ram_I.wpulse_I.wpulse_I[0]  (.A(\user_module.ram_I.wpulse_I.pulse ),
    .B(\user_module.ram_I.waddr_dec[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.store_gate[0] ));
 sky130_fd_sc_hd__and2_4 \user_module.ram_I.wpulse_I.wpulse_I[10]  (.A(\user_module.ram_I.wpulse_I.pulse ),
    .B(\user_module.ram_I.waddr_dec[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.store_gate[10] ));
 sky130_fd_sc_hd__and2_4 \user_module.ram_I.wpulse_I.wpulse_I[11]  (.A(\user_module.ram_I.wpulse_I.pulse ),
    .B(\user_module.ram_I.waddr_dec[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.store_gate[11] ));
 sky130_fd_sc_hd__and2_4 \user_module.ram_I.wpulse_I.wpulse_I[12]  (.A(\user_module.ram_I.wpulse_I.pulse ),
    .B(\user_module.ram_I.waddr_dec[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.store_gate[12] ));
 sky130_fd_sc_hd__and2_4 \user_module.ram_I.wpulse_I.wpulse_I[13]  (.A(\user_module.ram_I.wpulse_I.pulse ),
    .B(\user_module.ram_I.waddr_dec[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.store_gate[13] ));
 sky130_fd_sc_hd__and2_4 \user_module.ram_I.wpulse_I.wpulse_I[14]  (.A(\user_module.ram_I.wpulse_I.pulse ),
    .B(\user_module.ram_I.waddr_dec[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.store_gate[14] ));
 sky130_fd_sc_hd__and2_4 \user_module.ram_I.wpulse_I.wpulse_I[15]  (.A(\user_module.ram_I.wpulse_I.pulse ),
    .B(\user_module.ram_I.waddr_dec[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.store_gate[15] ));
 sky130_fd_sc_hd__and2_4 \user_module.ram_I.wpulse_I.wpulse_I[1]  (.A(\user_module.ram_I.wpulse_I.pulse ),
    .B(\user_module.ram_I.waddr_dec[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.store_gate[1] ));
 sky130_fd_sc_hd__and2_4 \user_module.ram_I.wpulse_I.wpulse_I[2]  (.A(\user_module.ram_I.wpulse_I.pulse ),
    .B(\user_module.ram_I.waddr_dec[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.store_gate[2] ));
 sky130_fd_sc_hd__and2_4 \user_module.ram_I.wpulse_I.wpulse_I[3]  (.A(\user_module.ram_I.wpulse_I.pulse ),
    .B(\user_module.ram_I.waddr_dec[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.store_gate[3] ));
 sky130_fd_sc_hd__and2_4 \user_module.ram_I.wpulse_I.wpulse_I[4]  (.A(\user_module.ram_I.wpulse_I.pulse ),
    .B(\user_module.ram_I.waddr_dec[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.store_gate[4] ));
 sky130_fd_sc_hd__and2_4 \user_module.ram_I.wpulse_I.wpulse_I[5]  (.A(\user_module.ram_I.wpulse_I.pulse ),
    .B(\user_module.ram_I.waddr_dec[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.store_gate[5] ));
 sky130_fd_sc_hd__and2_4 \user_module.ram_I.wpulse_I.wpulse_I[6]  (.A(\user_module.ram_I.wpulse_I.pulse ),
    .B(\user_module.ram_I.waddr_dec[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.store_gate[6] ));
 sky130_fd_sc_hd__and2_4 \user_module.ram_I.wpulse_I.wpulse_I[7]  (.A(\user_module.ram_I.wpulse_I.pulse ),
    .B(\user_module.ram_I.waddr_dec[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.store_gate[7] ));
 sky130_fd_sc_hd__and2_4 \user_module.ram_I.wpulse_I.wpulse_I[8]  (.A(\user_module.ram_I.wpulse_I.pulse ),
    .B(\user_module.ram_I.waddr_dec[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.store_gate[8] ));
 sky130_fd_sc_hd__and2_4 \user_module.ram_I.wpulse_I.wpulse_I[9]  (.A(\user_module.ram_I.wpulse_I.pulse ),
    .B(\user_module.ram_I.waddr_dec[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\user_module.ram_I.store_gate[9] ));
endmodule
