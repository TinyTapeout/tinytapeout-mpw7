VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO scan_controller
  CLASS BLOCK ;
  FOREIGN scan_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 230.000 BY 100.000 ;
  PIN active_select[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.940 4.000 62.140 ;
    END
  END active_select[0]
  PIN active_select[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 0.000 148.630 4.000 ;
    END
  END active_select[1]
  PIN active_select[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 96.000 142.190 100.000 ;
    END
  END active_select[2]
  PIN active_select[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.910 0.000 58.470 4.000 ;
    END
  END active_select[3]
  PIN active_select[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.150 0.000 193.710 4.000 ;
    END
  END active_select[4]
  PIN active_select[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.490 96.000 23.050 100.000 ;
    END
  END active_select[5]
  PIN active_select[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.050 0.000 177.610 4.000 ;
    END
  END active_select[6]
  PIN active_select[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.170 0.000 164.730 4.000 ;
    END
  END active_select[7]
  PIN active_select[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 54.140 230.000 55.340 ;
    END
  END active_select[8]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 96.000 64.910 100.000 ;
    END
  END clk
  PIN inputs[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.890 0.000 87.450 4.000 ;
    END
  END inputs[0]
  PIN inputs[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.940 4.000 45.140 ;
    END
  END inputs[1]
  PIN inputs[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.090 0.000 119.650 4.000 ;
    END
  END inputs[2]
  PIN inputs[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 67.740 230.000 68.940 ;
    END
  END inputs[3]
  PIN inputs[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.540 4.000 92.740 ;
    END
  END inputs[4]
  PIN inputs[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.930 0.000 29.490 4.000 ;
    END
  END inputs[5]
  PIN inputs[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.690 96.000 216.250 100.000 ;
    END
  END inputs[6]
  PIN inputs[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.610 96.000 171.170 100.000 ;
    END
  END inputs[7]
  PIN oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 20.140 230.000 21.340 ;
    END
  END oeb[0]
  PIN oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.590 96.000 200.150 100.000 ;
    END
  END oeb[1]
  PIN oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.340 4.000 31.540 ;
    END
  END oeb[2]
  PIN oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 84.740 230.000 85.940 ;
    END
  END oeb[3]
  PIN oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.550 96.000 97.110 100.000 ;
    END
  END oeb[4]
  PIN oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END oeb[5]
  PIN oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.510 96.000 155.070 100.000 ;
    END
  END oeb[6]
  PIN oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 37.140 230.000 38.340 ;
    END
  END oeb[7]
  PIN oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.450 96.000 81.010 100.000 ;
    END
  END oeb[8]
  PIN outputs[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.340 4.000 14.540 ;
    END
  END outputs[0]
  PIN outputs[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.970 0.000 132.530 4.000 ;
    END
  END outputs[1]
  PIN outputs[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 96.000 187.270 100.000 ;
    END
  END outputs[2]
  PIN outputs[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.030 0.000 206.590 4.000 ;
    END
  END outputs[3]
  PIN outputs[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.830 0.000 13.390 4.000 ;
    END
  END outputs[4]
  PIN outputs[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.810 0.000 42.370 4.000 ;
    END
  END outputs[5]
  PIN outputs[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.370 96.000 35.930 100.000 ;
    END
  END outputs[6]
  PIN outputs[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.130 0.000 222.690 4.000 ;
    END
  END outputs[7]
  PIN ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.010 0.000 74.570 4.000 ;
    END
  END ready
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.390 96.000 6.950 100.000 ;
    END
  END reset
  PIN scan_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.570 96.000 229.130 100.000 ;
    END
  END scan_clk
  PIN scan_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 96.000 109.990 100.000 ;
    END
  END scan_data_in
  PIN scan_data_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.530 96.000 126.090 100.000 ;
    END
  END scan_data_out
  PIN scan_latch_enable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 0.000 103.550 4.000 ;
    END
  END scan_latch_enable
  PIN scan_select
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.940 4.000 79.140 ;
    END
  END scan_select
  PIN set_clk_div
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.470 96.000 52.030 100.000 ;
    END
  END set_clk_div
  PIN slow_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 6.540 230.000 7.740 ;
    END
  END slow_clk
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 32.090 10.640 33.690 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 86.830 10.640 88.430 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.570 10.640 143.170 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.310 10.640 197.910 87.280 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 59.460 10.640 61.060 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.200 10.640 115.800 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 168.940 10.640 170.540 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 223.680 10.640 225.280 87.280 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 224.480 87.125 ;
      LAYER met1 ;
        RECT 0.070 10.240 229.010 87.280 ;
      LAYER met2 ;
        RECT 0.100 95.720 6.110 96.000 ;
        RECT 7.230 95.720 22.210 96.000 ;
        RECT 23.330 95.720 35.090 96.000 ;
        RECT 36.210 95.720 51.190 96.000 ;
        RECT 52.310 95.720 64.070 96.000 ;
        RECT 65.190 95.720 80.170 96.000 ;
        RECT 81.290 95.720 96.270 96.000 ;
        RECT 97.390 95.720 109.150 96.000 ;
        RECT 110.270 95.720 125.250 96.000 ;
        RECT 126.370 95.720 141.350 96.000 ;
        RECT 142.470 95.720 154.230 96.000 ;
        RECT 155.350 95.720 170.330 96.000 ;
        RECT 171.450 95.720 186.430 96.000 ;
        RECT 187.550 95.720 199.310 96.000 ;
        RECT 200.430 95.720 215.410 96.000 ;
        RECT 216.530 95.720 228.290 96.000 ;
        RECT 0.100 4.280 228.980 95.720 ;
        RECT 0.790 4.000 12.550 4.280 ;
        RECT 13.670 4.000 28.650 4.280 ;
        RECT 29.770 4.000 41.530 4.280 ;
        RECT 42.650 4.000 57.630 4.280 ;
        RECT 58.750 4.000 73.730 4.280 ;
        RECT 74.850 4.000 86.610 4.280 ;
        RECT 87.730 4.000 102.710 4.280 ;
        RECT 103.830 4.000 118.810 4.280 ;
        RECT 119.930 4.000 131.690 4.280 ;
        RECT 132.810 4.000 147.790 4.280 ;
        RECT 148.910 4.000 163.890 4.280 ;
        RECT 165.010 4.000 176.770 4.280 ;
        RECT 177.890 4.000 192.870 4.280 ;
        RECT 193.990 4.000 205.750 4.280 ;
        RECT 206.870 4.000 221.850 4.280 ;
        RECT 222.970 4.000 228.980 4.280 ;
      LAYER met3 ;
        RECT 4.400 91.140 226.010 92.305 ;
        RECT 4.000 86.340 226.010 91.140 ;
        RECT 4.000 84.340 225.600 86.340 ;
        RECT 4.000 79.540 226.010 84.340 ;
        RECT 4.400 77.540 226.010 79.540 ;
        RECT 4.000 69.340 226.010 77.540 ;
        RECT 4.000 67.340 225.600 69.340 ;
        RECT 4.000 62.540 226.010 67.340 ;
        RECT 4.400 60.540 226.010 62.540 ;
        RECT 4.000 55.740 226.010 60.540 ;
        RECT 4.000 53.740 225.600 55.740 ;
        RECT 4.000 45.540 226.010 53.740 ;
        RECT 4.400 43.540 226.010 45.540 ;
        RECT 4.000 38.740 226.010 43.540 ;
        RECT 4.000 36.740 225.600 38.740 ;
        RECT 4.000 31.940 226.010 36.740 ;
        RECT 4.400 29.940 226.010 31.940 ;
        RECT 4.000 21.740 226.010 29.940 ;
        RECT 4.000 19.740 225.600 21.740 ;
        RECT 4.000 14.940 226.010 19.740 ;
        RECT 4.400 12.940 226.010 14.940 ;
        RECT 4.000 8.140 226.010 12.940 ;
        RECT 4.000 6.975 225.600 8.140 ;
  END
END scan_controller
END LIBRARY

