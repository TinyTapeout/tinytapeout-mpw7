* NGSPICE file created from user_project_wrapper.ext - technology: sky130B

* Black-box entry subcircuit for scan_wrapper_341802448429515346 abstract view
.subckt scan_wrapper_341802448429515346 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341262321634509394 abstract view
.subckt scan_wrapper_341262321634509394 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341243232292700755 abstract view
.subckt scan_wrapper_341243232292700755 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341631511790879314 abstract view
.subckt scan_wrapper_341631511790879314 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_339501025136214612 abstract view
.subckt scan_wrapper_339501025136214612 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_1f985e14df1ed789231bb6e0189d6e39 abstract view
.subckt scan_wrapper_1f985e14df1ed789231bb6e0189d6e39 clk_in clk_out data_in data_out
+ latch_enable_in latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341524192738411090 abstract view
.subckt scan_wrapper_341524192738411090 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341628725785264722 abstract view
.subckt scan_wrapper_341628725785264722 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341235575572922964 abstract view
.subckt scan_wrapper_341235575572922964 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341191836498395731 abstract view
.subckt scan_wrapper_341191836498395731 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341631485498884690 abstract view
.subckt scan_wrapper_341631485498884690 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_340979268609638995 abstract view
.subckt scan_wrapper_340979268609638995 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341263346544149074 abstract view
.subckt scan_wrapper_341263346544149074 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341271902949474898 abstract view
.subckt scan_wrapper_341271902949474898 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_hamming74 abstract view
.subckt scan_wrapper_hamming74 clk_in clk_out data_in data_out latch_enable_in latch_enable_out
+ scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341178296293130834 abstract view
.subckt scan_wrapper_341178296293130834 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341399568412312147 abstract view
.subckt scan_wrapper_341399568412312147 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341423712597181012 abstract view
.subckt scan_wrapper_341423712597181012 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341233739099013714 abstract view
.subckt scan_wrapper_341233739099013714 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341571228858843732 abstract view
.subckt scan_wrapper_341571228858843732 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341617722294010450 abstract view
.subckt scan_wrapper_341617722294010450 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341193419111006803 abstract view
.subckt scan_wrapper_341193419111006803 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341360223723717202 abstract view
.subckt scan_wrapper_341360223723717202 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341590933015364178 abstract view
.subckt scan_wrapper_341590933015364178 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341277789473735250 abstract view
.subckt scan_wrapper_341277789473735250 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341182944314917460 abstract view
.subckt scan_wrapper_341182944314917460 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341259651269001812 abstract view
.subckt scan_wrapper_341259651269001812 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341155178824598098 abstract view
.subckt scan_wrapper_341155178824598098 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341315210433266259 abstract view
.subckt scan_wrapper_341315210433266259 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341174563322724948 abstract view
.subckt scan_wrapper_341174563322724948 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341192113929585235 abstract view
.subckt scan_wrapper_341192113929585235 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341164228775772755 abstract view
.subckt scan_wrapper_341164228775772755 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341614346808328788 abstract view
.subckt scan_wrapper_341614346808328788 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341637831098106450 abstract view
.subckt scan_wrapper_341637831098106450 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341432030163108435 abstract view
.subckt scan_wrapper_341432030163108435 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_340596276030603858 abstract view
.subckt scan_wrapper_340596276030603858 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341235973870322258 abstract view
.subckt scan_wrapper_341235973870322258 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341163800289870419 abstract view
.subckt scan_wrapper_341163800289870419 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341404507891040852 abstract view
.subckt scan_wrapper_341404507891040852 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341558189536313940 abstract view
.subckt scan_wrapper_341558189536313940 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341473139924927058 abstract view
.subckt scan_wrapper_341473139924927058 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341431339142087251 abstract view
.subckt scan_wrapper_341431339142087251 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341482086419399252 abstract view
.subckt scan_wrapper_341482086419399252 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_340661930553246290 abstract view
.subckt scan_wrapper_340661930553246290 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341154068332282450 abstract view
.subckt scan_wrapper_341154068332282450 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341438392303616596 abstract view
.subckt scan_wrapper_341438392303616596 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341521390605697619 abstract view
.subckt scan_wrapper_341521390605697619 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341440781874102868 abstract view
.subckt scan_wrapper_341440781874102868 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341224613878956628 abstract view
.subckt scan_wrapper_341224613878956628 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341541108650607187 abstract view
.subckt scan_wrapper_341541108650607187 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341344337258349139 abstract view
.subckt scan_wrapper_341344337258349139 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341457494561784402 abstract view
.subckt scan_wrapper_341457494561784402 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341497964482527828 abstract view
.subckt scan_wrapper_341497964482527828 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341493393195532884 abstract view
.subckt scan_wrapper_341493393195532884 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341499976001520211 abstract view
.subckt scan_wrapper_341499976001520211 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341410909669818963 abstract view
.subckt scan_wrapper_341410909669818963 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341620484740219475 abstract view
.subckt scan_wrapper_341620484740219475 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341339883600609876 abstract view
.subckt scan_wrapper_341339883600609876 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341490465660469844 abstract view
.subckt scan_wrapper_341490465660469844 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341608574336631379 abstract view
.subckt scan_wrapper_341608574336631379 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341802655228625490 abstract view
.subckt scan_wrapper_341802655228625490 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341063825089364563 abstract view
.subckt scan_wrapper_341063825089364563 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341332847867462227 abstract view
.subckt scan_wrapper_341332847867462227 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341136771628663380 abstract view
.subckt scan_wrapper_341136771628663380 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341424636358034002 abstract view
.subckt scan_wrapper_341424636358034002 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341440114308678227 abstract view
.subckt scan_wrapper_341440114308678227 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341178154799333971 abstract view
.subckt scan_wrapper_341178154799333971 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341497938559631956 abstract view
.subckt scan_wrapper_341497938559631956 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341452019534398035 abstract view
.subckt scan_wrapper_341452019534398035 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341500800901579348 abstract view
.subckt scan_wrapper_341500800901579348 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341419328215712339 abstract view
.subckt scan_wrapper_341419328215712339 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341160201697624660 abstract view
.subckt scan_wrapper_341160201697624660 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341342096033055316 abstract view
.subckt scan_wrapper_341342096033055316 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341462925422101075 abstract view
.subckt scan_wrapper_341462925422101075 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341364381657858642 abstract view
.subckt scan_wrapper_341364381657858642 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341516949939814994 abstract view
.subckt scan_wrapper_341516949939814994 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341710255833481812 abstract view
.subckt scan_wrapper_341710255833481812 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341538994733974098 abstract view
.subckt scan_wrapper_341538994733974098 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341457971277988435 abstract view
.subckt scan_wrapper_341457971277988435 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341161378978988626 abstract view
.subckt scan_wrapper_341161378978988626 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341629415144292948 abstract view
.subckt scan_wrapper_341629415144292948 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341188777753969234 abstract view
.subckt scan_wrapper_341188777753969234 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341496918381167187 abstract view
.subckt scan_wrapper_341496918381167187 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341717091617866324 abstract view
.subckt scan_wrapper_341717091617866324 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341589685194195540 abstract view
.subckt scan_wrapper_341589685194195540 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341202178192441940 abstract view
.subckt scan_wrapper_341202178192441940 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341337976625693266 abstract view
.subckt scan_wrapper_341337976625693266 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341476989274686036 abstract view
.subckt scan_wrapper_341476989274686036 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_339800239192932947 abstract view
.subckt scan_wrapper_339800239192932947 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_340285391309374034 abstract view
.subckt scan_wrapper_340285391309374034 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_339688086163161683 abstract view
.subckt scan_wrapper_339688086163161683 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341154161238213203 abstract view
.subckt scan_wrapper_341154161238213203 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341160271679586899 abstract view
.subckt scan_wrapper_341160271679586899 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341194143598379604 abstract view
.subckt scan_wrapper_341194143598379604 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341573751072096850 abstract view
.subckt scan_wrapper_341573751072096850 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341450853309219412 abstract view
.subckt scan_wrapper_341450853309219412 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341542971476279892 abstract view
.subckt scan_wrapper_341542971476279892 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341519170869920338 abstract view
.subckt scan_wrapper_341519170869920338 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341240110454407762 abstract view
.subckt scan_wrapper_341240110454407762 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_340318610245288530 abstract view
.subckt scan_wrapper_340318610245288530 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341556236196512338 abstract view
.subckt scan_wrapper_341556236196512338 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341389786199622227 abstract view
.subckt scan_wrapper_341389786199622227 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341162950004834900 abstract view
.subckt scan_wrapper_341162950004834900 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_bc4d7220e4fdbf20a574d56ea112a8e1 abstract view
.subckt scan_wrapper_bc4d7220e4fdbf20a574d56ea112a8e1 clk_in clk_out data_in data_out
+ latch_enable_in latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341382703379120723 abstract view
.subckt scan_wrapper_341382703379120723 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341167691532337747 abstract view
.subckt scan_wrapper_341167691532337747 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341192621088047698 abstract view
.subckt scan_wrapper_341192621088047698 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341431502448362067 abstract view
.subckt scan_wrapper_341431502448362067 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341444501414347346 abstract view
.subckt scan_wrapper_341444501414347346 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341520747710120530 abstract view
.subckt scan_wrapper_341520747710120530 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341296149788885588 abstract view
.subckt scan_wrapper_341296149788885588 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341567111632519764 abstract view
.subckt scan_wrapper_341567111632519764 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341353928049295956 abstract view
.subckt scan_wrapper_341353928049295956 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341432284947153491 abstract view
.subckt scan_wrapper_341432284947153491 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341353777861755476 abstract view
.subckt scan_wrapper_341353777861755476 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341159915403870803 abstract view
.subckt scan_wrapper_341159915403870803 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341449297858921043 abstract view
.subckt scan_wrapper_341449297858921043 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341205508016833108 abstract view
.subckt scan_wrapper_341205508016833108 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341557831870186068 abstract view
.subckt scan_wrapper_341557831870186068 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_340218629792465491 abstract view
.subckt scan_wrapper_340218629792465491 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341631644820570706 abstract view
.subckt scan_wrapper_341631644820570706 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341608297106768466 abstract view
.subckt scan_wrapper_341608297106768466 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341569483755749970 abstract view
.subckt scan_wrapper_341569483755749970 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341279123277087315 abstract view
.subckt scan_wrapper_341279123277087315 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341353780122485332 abstract view
.subckt scan_wrapper_341353780122485332 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341624400621077076 abstract view
.subckt scan_wrapper_341624400621077076 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341632596577354323 abstract view
.subckt scan_wrapper_341632596577354323 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341266732010177108 abstract view
.subckt scan_wrapper_341266732010177108 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341528610027340372 abstract view
.subckt scan_wrapper_341528610027340372 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341464767397888596 abstract view
.subckt scan_wrapper_341464767397888596 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341497971083313748 abstract view
.subckt scan_wrapper_341497971083313748 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341164910646919762 abstract view
.subckt scan_wrapper_341164910646919762 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_340067262721426004 abstract view
.subckt scan_wrapper_340067262721426004 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341174480471589458 abstract view
.subckt scan_wrapper_341174480471589458 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341678527574180436 abstract view
.subckt scan_wrapper_341678527574180436 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_controller abstract view
.subckt scan_controller active_select[0] active_select[1] active_select[2] active_select[3]
+ active_select[4] active_select[5] active_select[6] active_select[7] active_select[8]
+ clk driver_sel[0] driver_sel[1] inputs[0] inputs[1] inputs[2] inputs[3] inputs[4]
+ inputs[5] inputs[6] inputs[7] la_scan_clk_in la_scan_data_in la_scan_data_out la_scan_latch_en
+ la_scan_select oeb[0] oeb[10] oeb[11] oeb[12] oeb[13] oeb[14] oeb[15] oeb[16] oeb[17]
+ oeb[18] oeb[19] oeb[1] oeb[20] oeb[21] oeb[22] oeb[23] oeb[24] oeb[25] oeb[26] oeb[27]
+ oeb[28] oeb[29] oeb[2] oeb[30] oeb[31] oeb[32] oeb[33] oeb[34] oeb[35] oeb[36] oeb[37]
+ oeb[3] oeb[4] oeb[5] oeb[6] oeb[7] oeb[8] oeb[9] outputs[0] outputs[1] outputs[2]
+ outputs[3] outputs[4] outputs[5] outputs[6] outputs[7] ready reset scan_clk_in scan_clk_out
+ scan_data_in scan_data_out scan_latch_en scan_select set_clk_div slow_clk vccd1
+ vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_019235602376235615 abstract view
.subckt scan_wrapper_019235602376235615 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341178481588044372 abstract view
.subckt scan_wrapper_341178481588044372 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341426151397261906 abstract view
.subckt scan_wrapper_341426151397261906 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341152580068442706 abstract view
.subckt scan_wrapper_341152580068442706 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341533740987581011 abstract view
.subckt scan_wrapper_341533740987581011 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341446083683025490 abstract view
.subckt scan_wrapper_341446083683025490 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341609034095264340 abstract view
.subckt scan_wrapper_341609034095264340 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341614536664547922 abstract view
.subckt scan_wrapper_341614536664547922 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341264068701586004 abstract view
.subckt scan_wrapper_341264068701586004 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341546888233747026 abstract view
.subckt scan_wrapper_341546888233747026 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341506274933867090 abstract view
.subckt scan_wrapper_341506274933867090 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341581732833657427 abstract view
.subckt scan_wrapper_341581732833657427 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_340579111348994642 abstract view
.subckt scan_wrapper_340579111348994642 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341613097060926036 abstract view
.subckt scan_wrapper_341613097060926036 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341176884318437971 abstract view
.subckt scan_wrapper_341176884318437971 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_wrapper_341359404107432531 abstract view
.subckt scan_wrapper_341359404107432531 clk_in clk_out data_in data_out latch_enable_in
+ latch_enable_out scan_select_in scan_select_out vccd1 vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xscan_wrapper_341802448429515346_132 scan_wrapper_341802448429515346_132/clk_in scan_wrapper_341609034095264340_133/clk_in
+ scan_wrapper_341802448429515346_132/data_in scan_wrapper_341609034095264340_133/data_in
+ scan_wrapper_341802448429515346_132/latch_enable_in scan_wrapper_341609034095264340_133/latch_enable_in
+ scan_wrapper_341802448429515346_132/scan_select_in scan_wrapper_341609034095264340_133/scan_select_in
+ vccd1 vssd1 scan_wrapper_341802448429515346
Xscan_wrapper_341262321634509394_39 scan_wrapper_341262321634509394_39/clk_in scan_wrapper_341174563322724948_40/clk_in
+ scan_wrapper_341262321634509394_39/data_in scan_wrapper_341174563322724948_40/data_in
+ scan_wrapper_341262321634509394_39/latch_enable_in scan_wrapper_341174563322724948_40/latch_enable_in
+ scan_wrapper_341262321634509394_39/scan_select_in scan_wrapper_341174563322724948_40/scan_select_in
+ vccd1 vssd1 scan_wrapper_341262321634509394
Xscan_wrapper_341243232292700755_102 scan_wrapper_341243232292700755_102/clk_in scan_wrapper_341519170869920338_103/clk_in
+ scan_wrapper_341243232292700755_102/data_in scan_wrapper_341519170869920338_103/data_in
+ scan_wrapper_341243232292700755_102/latch_enable_in scan_wrapper_341519170869920338_103/latch_enable_in
+ scan_wrapper_341243232292700755_102/scan_select_in scan_wrapper_341519170869920338_103/scan_select_in
+ vccd1 vssd1 scan_wrapper_341243232292700755
Xscan_wrapper_341631511790879314_144 scan_wrapper_341631511790879314_144/clk_in scan_wrapper_341426151397261906_145/clk_in
+ scan_wrapper_341631511790879314_144/data_in scan_wrapper_341426151397261906_145/data_in
+ scan_wrapper_341631511790879314_144/latch_enable_in scan_wrapper_341426151397261906_145/latch_enable_in
+ scan_wrapper_341631511790879314_144/scan_select_in scan_wrapper_341426151397261906_145/scan_select_in
+ vccd1 vssd1 scan_wrapper_341631511790879314
Xscan_wrapper_339501025136214612_379 scan_wrapper_339501025136214612_379/clk_in scan_wrapper_339501025136214612_380/clk_in
+ scan_wrapper_339501025136214612_379/data_in scan_wrapper_339501025136214612_380/data_in
+ scan_wrapper_339501025136214612_379/latch_enable_in scan_wrapper_339501025136214612_380/latch_enable_in
+ scan_wrapper_339501025136214612_379/scan_select_in scan_wrapper_339501025136214612_380/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_313 scan_wrapper_339501025136214612_313/clk_in scan_wrapper_339501025136214612_314/clk_in
+ scan_wrapper_339501025136214612_313/data_in scan_wrapper_339501025136214612_314/data_in
+ scan_wrapper_339501025136214612_313/latch_enable_in scan_wrapper_339501025136214612_314/latch_enable_in
+ scan_wrapper_339501025136214612_313/scan_select_in scan_wrapper_339501025136214612_314/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_302 scan_wrapper_339501025136214612_302/clk_in scan_wrapper_339501025136214612_303/clk_in
+ scan_wrapper_339501025136214612_302/data_in scan_wrapper_339501025136214612_303/data_in
+ scan_wrapper_339501025136214612_302/latch_enable_in scan_wrapper_339501025136214612_303/latch_enable_in
+ scan_wrapper_339501025136214612_302/scan_select_in scan_wrapper_339501025136214612_303/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_324 scan_wrapper_339501025136214612_324/clk_in scan_wrapper_339501025136214612_325/clk_in
+ scan_wrapper_339501025136214612_324/data_in scan_wrapper_339501025136214612_325/data_in
+ scan_wrapper_339501025136214612_324/latch_enable_in scan_wrapper_339501025136214612_325/latch_enable_in
+ scan_wrapper_339501025136214612_324/scan_select_in scan_wrapper_339501025136214612_325/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_335 scan_wrapper_339501025136214612_335/clk_in scan_wrapper_339501025136214612_336/clk_in
+ scan_wrapper_339501025136214612_335/data_in scan_wrapper_339501025136214612_336/data_in
+ scan_wrapper_339501025136214612_335/latch_enable_in scan_wrapper_339501025136214612_336/latch_enable_in
+ scan_wrapper_339501025136214612_335/scan_select_in scan_wrapper_339501025136214612_336/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_357 scan_wrapper_339501025136214612_357/clk_in scan_wrapper_339501025136214612_358/clk_in
+ scan_wrapper_339501025136214612_357/data_in scan_wrapper_339501025136214612_358/data_in
+ scan_wrapper_339501025136214612_357/latch_enable_in scan_wrapper_339501025136214612_358/latch_enable_in
+ scan_wrapper_339501025136214612_357/scan_select_in scan_wrapper_339501025136214612_358/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_346 scan_wrapper_339501025136214612_346/clk_in scan_wrapper_339501025136214612_347/clk_in
+ scan_wrapper_339501025136214612_346/data_in scan_wrapper_339501025136214612_347/data_in
+ scan_wrapper_339501025136214612_346/latch_enable_in scan_wrapper_339501025136214612_347/latch_enable_in
+ scan_wrapper_339501025136214612_346/scan_select_in scan_wrapper_339501025136214612_347/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_368 scan_wrapper_339501025136214612_368/clk_in scan_wrapper_339501025136214612_369/clk_in
+ scan_wrapper_339501025136214612_368/data_in scan_wrapper_339501025136214612_369/data_in
+ scan_wrapper_339501025136214612_368/latch_enable_in scan_wrapper_339501025136214612_369/latch_enable_in
+ scan_wrapper_339501025136214612_368/scan_select_in scan_wrapper_339501025136214612_369/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_1f985e14df1ed789231bb6e0189d6e39_44 scan_wrapper_341178296293130834_43/clk_out
+ scan_wrapper_341277789473735250_45/clk_in scan_wrapper_341178296293130834_43/data_out
+ scan_wrapper_341277789473735250_45/data_in scan_wrapper_341178296293130834_43/latch_enable_out
+ scan_wrapper_341277789473735250_45/latch_enable_in scan_wrapper_341178296293130834_43/scan_select_out
+ scan_wrapper_341277789473735250_45/scan_select_in vccd1 vssd1 scan_wrapper_1f985e14df1ed789231bb6e0189d6e39
Xscan_wrapper_341524192738411090_105 scan_wrapper_341524192738411090_105/clk_in scan_wrapper_341533740987581011_106/clk_in
+ scan_wrapper_341524192738411090_105/data_in scan_wrapper_341533740987581011_106/data_in
+ scan_wrapper_341524192738411090_105/latch_enable_in scan_wrapper_341533740987581011_106/latch_enable_in
+ scan_wrapper_341524192738411090_105/scan_select_in scan_wrapper_341533740987581011_106/scan_select_in
+ vccd1 vssd1 scan_wrapper_341524192738411090
Xscan_wrapper_339501025136214612_154 scan_wrapper_339501025136214612_154/clk_in scan_wrapper_339501025136214612_155/clk_in
+ scan_wrapper_339501025136214612_154/data_in scan_wrapper_339501025136214612_155/data_in
+ scan_wrapper_339501025136214612_154/latch_enable_in scan_wrapper_339501025136214612_155/latch_enable_in
+ scan_wrapper_339501025136214612_154/scan_select_in scan_wrapper_339501025136214612_155/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_165 scan_wrapper_339501025136214612_165/clk_in scan_wrapper_339501025136214612_166/clk_in
+ scan_wrapper_339501025136214612_165/data_in scan_wrapper_339501025136214612_166/data_in
+ scan_wrapper_339501025136214612_165/latch_enable_in scan_wrapper_339501025136214612_166/latch_enable_in
+ scan_wrapper_339501025136214612_165/scan_select_in scan_wrapper_339501025136214612_166/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_176 scan_wrapper_339501025136214612_176/clk_in scan_wrapper_339501025136214612_177/clk_in
+ scan_wrapper_339501025136214612_176/data_in scan_wrapper_339501025136214612_177/data_in
+ scan_wrapper_339501025136214612_176/latch_enable_in scan_wrapper_339501025136214612_177/latch_enable_in
+ scan_wrapper_339501025136214612_176/scan_select_in scan_wrapper_339501025136214612_177/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_187 scan_wrapper_339501025136214612_187/clk_in scan_wrapper_339501025136214612_188/clk_in
+ scan_wrapper_339501025136214612_187/data_in scan_wrapper_339501025136214612_188/data_in
+ scan_wrapper_339501025136214612_187/latch_enable_in scan_wrapper_339501025136214612_188/latch_enable_in
+ scan_wrapper_339501025136214612_187/scan_select_in scan_wrapper_339501025136214612_188/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_198 scan_wrapper_339501025136214612_198/clk_in scan_wrapper_339501025136214612_199/clk_in
+ scan_wrapper_339501025136214612_198/data_in scan_wrapper_339501025136214612_199/data_in
+ scan_wrapper_339501025136214612_198/latch_enable_in scan_wrapper_339501025136214612_199/latch_enable_in
+ scan_wrapper_339501025136214612_198/scan_select_in scan_wrapper_339501025136214612_199/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341628725785264722_143 scan_wrapper_341628725785264722_143/clk_in scan_wrapper_341631511790879314_144/clk_in
+ scan_wrapper_341628725785264722_143/data_in scan_wrapper_341631511790879314_144/data_in
+ scan_wrapper_341628725785264722_143/latch_enable_in scan_wrapper_341631511790879314_144/latch_enable_in
+ scan_wrapper_341628725785264722_143/scan_select_in scan_wrapper_341631511790879314_144/scan_select_in
+ vccd1 vssd1 scan_wrapper_341628725785264722
Xscan_wrapper_341235575572922964_33 scan_wrapper_341235575572922964_33/clk_in scan_wrapper_341164910646919762_34/clk_in
+ scan_wrapper_341235575572922964_33/data_in scan_wrapper_341164910646919762_34/data_in
+ scan_wrapper_341235575572922964_33/latch_enable_in scan_wrapper_341164910646919762_34/latch_enable_in
+ scan_wrapper_341235575572922964_33/scan_select_in scan_wrapper_341164910646919762_34/scan_select_in
+ vccd1 vssd1 scan_wrapper_341235575572922964
Xscan_wrapper_341191836498395731_27 scan_wrapper_341191836498395731_27/clk_in scan_wrapper_341192113929585235_28/clk_in
+ scan_wrapper_341191836498395731_27/data_in scan_wrapper_341192113929585235_28/data_in
+ scan_wrapper_341191836498395731_27/latch_enable_in scan_wrapper_341192113929585235_28/latch_enable_in
+ scan_wrapper_341191836498395731_27/scan_select_in scan_wrapper_341192113929585235_28/scan_select_in
+ vccd1 vssd1 scan_wrapper_341191836498395731
Xscan_wrapper_339501025136214612_314 scan_wrapper_339501025136214612_314/clk_in scan_wrapper_339501025136214612_315/clk_in
+ scan_wrapper_339501025136214612_314/data_in scan_wrapper_339501025136214612_315/data_in
+ scan_wrapper_339501025136214612_314/latch_enable_in scan_wrapper_339501025136214612_315/latch_enable_in
+ scan_wrapper_339501025136214612_314/scan_select_in scan_wrapper_339501025136214612_315/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_303 scan_wrapper_339501025136214612_303/clk_in scan_wrapper_339501025136214612_304/clk_in
+ scan_wrapper_339501025136214612_303/data_in scan_wrapper_339501025136214612_304/data_in
+ scan_wrapper_339501025136214612_303/latch_enable_in scan_wrapper_339501025136214612_304/latch_enable_in
+ scan_wrapper_339501025136214612_303/scan_select_in scan_wrapper_339501025136214612_304/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_325 scan_wrapper_339501025136214612_325/clk_in scan_wrapper_339501025136214612_326/clk_in
+ scan_wrapper_339501025136214612_325/data_in scan_wrapper_339501025136214612_326/data_in
+ scan_wrapper_339501025136214612_325/latch_enable_in scan_wrapper_339501025136214612_326/latch_enable_in
+ scan_wrapper_339501025136214612_325/scan_select_in scan_wrapper_339501025136214612_326/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_336 scan_wrapper_339501025136214612_336/clk_in scan_wrapper_339501025136214612_337/clk_in
+ scan_wrapper_339501025136214612_336/data_in scan_wrapper_339501025136214612_337/data_in
+ scan_wrapper_339501025136214612_336/latch_enable_in scan_wrapper_339501025136214612_337/latch_enable_in
+ scan_wrapper_339501025136214612_336/scan_select_in scan_wrapper_339501025136214612_337/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_347 scan_wrapper_339501025136214612_347/clk_in scan_wrapper_339501025136214612_348/clk_in
+ scan_wrapper_339501025136214612_347/data_in scan_wrapper_339501025136214612_348/data_in
+ scan_wrapper_339501025136214612_347/latch_enable_in scan_wrapper_339501025136214612_348/latch_enable_in
+ scan_wrapper_339501025136214612_347/scan_select_in scan_wrapper_339501025136214612_348/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_358 scan_wrapper_339501025136214612_358/clk_in scan_wrapper_339501025136214612_359/clk_in
+ scan_wrapper_339501025136214612_358/data_in scan_wrapper_339501025136214612_359/data_in
+ scan_wrapper_339501025136214612_358/latch_enable_in scan_wrapper_339501025136214612_359/latch_enable_in
+ scan_wrapper_339501025136214612_358/scan_select_in scan_wrapper_339501025136214612_359/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_369 scan_wrapper_339501025136214612_369/clk_in scan_wrapper_339501025136214612_370/clk_in
+ scan_wrapper_339501025136214612_369/data_in scan_wrapper_339501025136214612_370/data_in
+ scan_wrapper_339501025136214612_369/latch_enable_in scan_wrapper_339501025136214612_370/latch_enable_in
+ scan_wrapper_339501025136214612_369/scan_select_in scan_wrapper_339501025136214612_370/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_155 scan_wrapper_339501025136214612_155/clk_in scan_wrapper_339501025136214612_156/clk_in
+ scan_wrapper_339501025136214612_155/data_in scan_wrapper_339501025136214612_156/data_in
+ scan_wrapper_339501025136214612_155/latch_enable_in scan_wrapper_339501025136214612_156/latch_enable_in
+ scan_wrapper_339501025136214612_155/scan_select_in scan_wrapper_339501025136214612_156/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_166 scan_wrapper_339501025136214612_166/clk_in scan_wrapper_339501025136214612_167/clk_in
+ scan_wrapper_339501025136214612_166/data_in scan_wrapper_339501025136214612_167/data_in
+ scan_wrapper_339501025136214612_166/latch_enable_in scan_wrapper_339501025136214612_167/latch_enable_in
+ scan_wrapper_339501025136214612_166/scan_select_in scan_wrapper_339501025136214612_167/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_177 scan_wrapper_339501025136214612_177/clk_in scan_wrapper_339501025136214612_178/clk_in
+ scan_wrapper_339501025136214612_177/data_in scan_wrapper_339501025136214612_178/data_in
+ scan_wrapper_339501025136214612_177/latch_enable_in scan_wrapper_339501025136214612_178/latch_enable_in
+ scan_wrapper_339501025136214612_177/scan_select_in scan_wrapper_339501025136214612_178/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_188 scan_wrapper_339501025136214612_188/clk_in scan_wrapper_339501025136214612_189/clk_in
+ scan_wrapper_339501025136214612_188/data_in scan_wrapper_339501025136214612_189/data_in
+ scan_wrapper_339501025136214612_188/latch_enable_in scan_wrapper_339501025136214612_189/latch_enable_in
+ scan_wrapper_339501025136214612_188/scan_select_in scan_wrapper_339501025136214612_189/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_199 scan_wrapper_339501025136214612_199/clk_in scan_wrapper_339501025136214612_200/clk_in
+ scan_wrapper_339501025136214612_199/data_in scan_wrapper_339501025136214612_200/data_in
+ scan_wrapper_339501025136214612_199/latch_enable_in scan_wrapper_339501025136214612_200/latch_enable_in
+ scan_wrapper_339501025136214612_199/scan_select_in scan_wrapper_339501025136214612_200/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341631485498884690_141 scan_wrapper_341631485498884690_141/clk_in scan_wrapper_341632596577354323_142/clk_in
+ scan_wrapper_341631485498884690_141/data_in scan_wrapper_341632596577354323_142/data_in
+ scan_wrapper_341631485498884690_141/latch_enable_in scan_wrapper_341632596577354323_142/latch_enable_in
+ scan_wrapper_341631485498884690_141/scan_select_in scan_wrapper_341632596577354323_142/scan_select_in
+ vccd1 vssd1 scan_wrapper_341631485498884690
Xscan_wrapper_340979268609638995_116 scan_wrapper_340979268609638995_116/clk_in scan_wrapper_341542971476279892_117/clk_in
+ scan_wrapper_340979268609638995_116/data_in scan_wrapper_341542971476279892_117/data_in
+ scan_wrapper_340979268609638995_116/latch_enable_in scan_wrapper_341542971476279892_117/latch_enable_in
+ scan_wrapper_340979268609638995_116/scan_select_in scan_wrapper_341542971476279892_117/scan_select_in
+ vccd1 vssd1 scan_wrapper_340979268609638995
Xscan_wrapper_341263346544149074_46 scan_wrapper_341263346544149074_46/clk_in scan_wrapper_341296149788885588_47/clk_in
+ scan_wrapper_341263346544149074_46/data_in scan_wrapper_341296149788885588_47/data_in
+ scan_wrapper_341263346544149074_46/latch_enable_in scan_wrapper_341296149788885588_47/latch_enable_in
+ scan_wrapper_341263346544149074_46/scan_select_in scan_wrapper_341296149788885588_47/scan_select_in
+ vccd1 vssd1 scan_wrapper_341263346544149074
Xscan_wrapper_341271902949474898_41 scan_wrapper_341271902949474898_41/clk_in scan_wrapper_341271902949474898_41/clk_out
+ scan_wrapper_341271902949474898_41/data_in scan_wrapper_341271902949474898_41/data_out
+ scan_wrapper_341271902949474898_41/latch_enable_in scan_wrapper_341271902949474898_41/latch_enable_out
+ scan_wrapper_341271902949474898_41/scan_select_in scan_wrapper_341271902949474898_41/scan_select_out
+ vccd1 vssd1 scan_wrapper_341271902949474898
Xscan_wrapper_339501025136214612_0 scan_controller/scan_clk_out scan_wrapper_339688086163161683_1/clk_in
+ scan_controller/scan_data_out scan_wrapper_339688086163161683_1/data_in scan_controller/scan_latch_en
+ scan_wrapper_339688086163161683_1/latch_enable_in scan_controller/scan_select scan_wrapper_339688086163161683_1/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_hamming74_112 scan_wrapper_hamming74_112/clk_in scan_wrapper_hamming74_112/clk_out
+ scan_wrapper_hamming74_112/data_in scan_wrapper_hamming74_112/data_out scan_wrapper_hamming74_112/latch_enable_in
+ scan_wrapper_hamming74_112/latch_enable_out scan_wrapper_hamming74_112/scan_select_in
+ scan_wrapper_hamming74_112/scan_select_out vccd1 vssd1 scan_wrapper_hamming74
Xscan_wrapper_339501025136214612_315 scan_wrapper_339501025136214612_315/clk_in scan_wrapper_339501025136214612_316/clk_in
+ scan_wrapper_339501025136214612_315/data_in scan_wrapper_339501025136214612_316/data_in
+ scan_wrapper_339501025136214612_315/latch_enable_in scan_wrapper_339501025136214612_316/latch_enable_in
+ scan_wrapper_339501025136214612_315/scan_select_in scan_wrapper_339501025136214612_316/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_304 scan_wrapper_339501025136214612_304/clk_in scan_wrapper_339501025136214612_305/clk_in
+ scan_wrapper_339501025136214612_304/data_in scan_wrapper_339501025136214612_305/data_in
+ scan_wrapper_339501025136214612_304/latch_enable_in scan_wrapper_339501025136214612_305/latch_enable_in
+ scan_wrapper_339501025136214612_304/scan_select_in scan_wrapper_339501025136214612_305/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_326 scan_wrapper_339501025136214612_326/clk_in scan_wrapper_339501025136214612_327/clk_in
+ scan_wrapper_339501025136214612_326/data_in scan_wrapper_339501025136214612_327/data_in
+ scan_wrapper_339501025136214612_326/latch_enable_in scan_wrapper_339501025136214612_327/latch_enable_in
+ scan_wrapper_339501025136214612_326/scan_select_in scan_wrapper_339501025136214612_327/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_337 scan_wrapper_339501025136214612_337/clk_in scan_wrapper_339501025136214612_338/clk_in
+ scan_wrapper_339501025136214612_337/data_in scan_wrapper_339501025136214612_338/data_in
+ scan_wrapper_339501025136214612_337/latch_enable_in scan_wrapper_339501025136214612_338/latch_enable_in
+ scan_wrapper_339501025136214612_337/scan_select_in scan_wrapper_339501025136214612_338/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_348 scan_wrapper_339501025136214612_348/clk_in scan_wrapper_339501025136214612_349/clk_in
+ scan_wrapper_339501025136214612_348/data_in scan_wrapper_339501025136214612_349/data_in
+ scan_wrapper_339501025136214612_348/latch_enable_in scan_wrapper_339501025136214612_349/latch_enable_in
+ scan_wrapper_339501025136214612_348/scan_select_in scan_wrapper_339501025136214612_349/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_359 scan_wrapper_339501025136214612_359/clk_in scan_wrapper_339501025136214612_360/clk_in
+ scan_wrapper_339501025136214612_359/data_in scan_wrapper_339501025136214612_360/data_in
+ scan_wrapper_339501025136214612_359/latch_enable_in scan_wrapper_339501025136214612_360/latch_enable_in
+ scan_wrapper_339501025136214612_359/scan_select_in scan_wrapper_339501025136214612_360/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_156 scan_wrapper_339501025136214612_156/clk_in scan_wrapper_339501025136214612_157/clk_in
+ scan_wrapper_339501025136214612_156/data_in scan_wrapper_339501025136214612_157/data_in
+ scan_wrapper_339501025136214612_156/latch_enable_in scan_wrapper_339501025136214612_157/latch_enable_in
+ scan_wrapper_339501025136214612_156/scan_select_in scan_wrapper_339501025136214612_157/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_167 scan_wrapper_339501025136214612_167/clk_in scan_wrapper_339501025136214612_168/clk_in
+ scan_wrapper_339501025136214612_167/data_in scan_wrapper_339501025136214612_168/data_in
+ scan_wrapper_339501025136214612_167/latch_enable_in scan_wrapper_339501025136214612_168/latch_enable_in
+ scan_wrapper_339501025136214612_167/scan_select_in scan_wrapper_339501025136214612_168/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_189 scan_wrapper_339501025136214612_189/clk_in scan_wrapper_339501025136214612_190/clk_in
+ scan_wrapper_339501025136214612_189/data_in scan_wrapper_339501025136214612_190/data_in
+ scan_wrapper_339501025136214612_189/latch_enable_in scan_wrapper_339501025136214612_190/latch_enable_in
+ scan_wrapper_339501025136214612_189/scan_select_in scan_wrapper_339501025136214612_190/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_178 scan_wrapper_339501025136214612_178/clk_in scan_wrapper_339501025136214612_179/clk_in
+ scan_wrapper_339501025136214612_178/data_in scan_wrapper_339501025136214612_179/data_in
+ scan_wrapper_339501025136214612_178/latch_enable_in scan_wrapper_339501025136214612_179/latch_enable_in
+ scan_wrapper_339501025136214612_178/scan_select_in scan_wrapper_339501025136214612_179/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341178296293130834_43 scan_wrapper_341178296293130834_43/clk_in scan_wrapper_341178296293130834_43/clk_out
+ scan_wrapper_341178296293130834_43/data_in scan_wrapper_341178296293130834_43/data_out
+ scan_wrapper_341178296293130834_43/latch_enable_in scan_wrapper_341178296293130834_43/latch_enable_out
+ scan_wrapper_341178296293130834_43/scan_select_in scan_wrapper_341178296293130834_43/scan_select_out
+ vccd1 vssd1 scan_wrapper_341178296293130834
Xscan_wrapper_341399568412312147_82 scan_wrapper_341399568412312147_82/clk_in scan_wrapper_341464767397888596_83/clk_in
+ scan_wrapper_341399568412312147_82/data_in scan_wrapper_341464767397888596_83/data_in
+ scan_wrapper_341399568412312147_82/latch_enable_in scan_wrapper_341464767397888596_83/latch_enable_in
+ scan_wrapper_341399568412312147_82/scan_select_in scan_wrapper_341464767397888596_83/scan_select_in
+ vccd1 vssd1 scan_wrapper_341399568412312147
Xscan_wrapper_341423712597181012_99 scan_wrapper_341423712597181012_99/clk_in scan_wrapper_341516949939814994_100/clk_in
+ scan_wrapper_341423712597181012_99/data_in scan_wrapper_341516949939814994_100/data_in
+ scan_wrapper_341423712597181012_99/latch_enable_in scan_wrapper_341516949939814994_100/latch_enable_in
+ scan_wrapper_341423712597181012_99/scan_select_in scan_wrapper_341516949939814994_100/scan_select_in
+ vccd1 vssd1 scan_wrapper_341423712597181012
Xscan_wrapper_341233739099013714_35 scan_wrapper_341233739099013714_35/clk_in scan_wrapper_341240110454407762_36/clk_in
+ scan_wrapper_341233739099013714_35/data_in scan_wrapper_341240110454407762_36/data_in
+ scan_wrapper_341233739099013714_35/latch_enable_in scan_wrapper_341240110454407762_36/latch_enable_in
+ scan_wrapper_341233739099013714_35/scan_select_in scan_wrapper_341240110454407762_36/scan_select_in
+ vccd1 vssd1 scan_wrapper_341233739099013714
Xscan_wrapper_341571228858843732_124 scan_wrapper_341571228858843732_124/clk_in scan_wrapper_341490465660469844_125/clk_in
+ scan_wrapper_341571228858843732_124/data_in scan_wrapper_341490465660469844_125/data_in
+ scan_wrapper_341571228858843732_124/latch_enable_in scan_wrapper_341490465660469844_125/latch_enable_in
+ scan_wrapper_341571228858843732_124/scan_select_in scan_wrapper_341490465660469844_125/scan_select_in
+ vccd1 vssd1 scan_wrapper_341571228858843732
Xscan_wrapper_339501025136214612_316 scan_wrapper_339501025136214612_316/clk_in scan_wrapper_339501025136214612_317/clk_in
+ scan_wrapper_339501025136214612_316/data_in scan_wrapper_339501025136214612_317/data_in
+ scan_wrapper_339501025136214612_316/latch_enable_in scan_wrapper_339501025136214612_317/latch_enable_in
+ scan_wrapper_339501025136214612_316/scan_select_in scan_wrapper_339501025136214612_317/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_305 scan_wrapper_339501025136214612_305/clk_in scan_wrapper_339501025136214612_306/clk_in
+ scan_wrapper_339501025136214612_305/data_in scan_wrapper_339501025136214612_306/data_in
+ scan_wrapper_339501025136214612_305/latch_enable_in scan_wrapper_339501025136214612_306/latch_enable_in
+ scan_wrapper_339501025136214612_305/scan_select_in scan_wrapper_339501025136214612_306/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_327 scan_wrapper_339501025136214612_327/clk_in scan_wrapper_339501025136214612_328/clk_in
+ scan_wrapper_339501025136214612_327/data_in scan_wrapper_339501025136214612_328/data_in
+ scan_wrapper_339501025136214612_327/latch_enable_in scan_wrapper_339501025136214612_328/latch_enable_in
+ scan_wrapper_339501025136214612_327/scan_select_in scan_wrapper_339501025136214612_328/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_349 scan_wrapper_339501025136214612_349/clk_in scan_wrapper_339501025136214612_350/clk_in
+ scan_wrapper_339501025136214612_349/data_in scan_wrapper_339501025136214612_350/data_in
+ scan_wrapper_339501025136214612_349/latch_enable_in scan_wrapper_339501025136214612_350/latch_enable_in
+ scan_wrapper_339501025136214612_349/scan_select_in scan_wrapper_339501025136214612_350/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_338 scan_wrapper_339501025136214612_338/clk_in scan_wrapper_339501025136214612_339/clk_in
+ scan_wrapper_339501025136214612_338/data_in scan_wrapper_339501025136214612_339/data_in
+ scan_wrapper_339501025136214612_338/latch_enable_in scan_wrapper_339501025136214612_339/latch_enable_in
+ scan_wrapper_339501025136214612_338/scan_select_in scan_wrapper_339501025136214612_339/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341617722294010450_134 scan_wrapper_341617722294010450_134/clk_in scan_wrapper_341613097060926036_135/clk_in
+ scan_wrapper_341617722294010450_134/data_in scan_wrapper_341613097060926036_135/data_in
+ scan_wrapper_341617722294010450_134/latch_enable_in scan_wrapper_341613097060926036_135/latch_enable_in
+ scan_wrapper_341617722294010450_134/scan_select_in scan_wrapper_341613097060926036_135/scan_select_in
+ vccd1 vssd1 scan_wrapper_341617722294010450
Xscan_wrapper_339501025136214612_157 scan_wrapper_339501025136214612_157/clk_in scan_wrapper_339501025136214612_158/clk_in
+ scan_wrapper_339501025136214612_157/data_in scan_wrapper_339501025136214612_158/data_in
+ scan_wrapper_339501025136214612_157/latch_enable_in scan_wrapper_339501025136214612_158/latch_enable_in
+ scan_wrapper_339501025136214612_157/scan_select_in scan_wrapper_339501025136214612_158/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_168 scan_wrapper_339501025136214612_168/clk_in scan_wrapper_339501025136214612_169/clk_in
+ scan_wrapper_339501025136214612_168/data_in scan_wrapper_339501025136214612_169/data_in
+ scan_wrapper_339501025136214612_168/latch_enable_in scan_wrapper_339501025136214612_169/latch_enable_in
+ scan_wrapper_339501025136214612_168/scan_select_in scan_wrapper_339501025136214612_169/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_179 scan_wrapper_339501025136214612_179/clk_in scan_wrapper_339501025136214612_180/clk_in
+ scan_wrapper_339501025136214612_179/data_in scan_wrapper_339501025136214612_180/data_in
+ scan_wrapper_339501025136214612_179/latch_enable_in scan_wrapper_339501025136214612_180/latch_enable_in
+ scan_wrapper_339501025136214612_179/scan_select_in scan_wrapper_339501025136214612_180/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_317 scan_wrapper_339501025136214612_317/clk_in scan_wrapper_339501025136214612_318/clk_in
+ scan_wrapper_339501025136214612_317/data_in scan_wrapper_339501025136214612_318/data_in
+ scan_wrapper_339501025136214612_317/latch_enable_in scan_wrapper_339501025136214612_318/latch_enable_in
+ scan_wrapper_339501025136214612_317/scan_select_in scan_wrapper_339501025136214612_318/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_306 scan_wrapper_339501025136214612_306/clk_in scan_wrapper_339501025136214612_307/clk_in
+ scan_wrapper_339501025136214612_306/data_in scan_wrapper_339501025136214612_307/data_in
+ scan_wrapper_339501025136214612_306/latch_enable_in scan_wrapper_339501025136214612_307/latch_enable_in
+ scan_wrapper_339501025136214612_306/scan_select_in scan_wrapper_339501025136214612_307/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_328 scan_wrapper_339501025136214612_328/clk_in scan_wrapper_339501025136214612_329/clk_in
+ scan_wrapper_339501025136214612_328/data_in scan_wrapper_339501025136214612_329/data_in
+ scan_wrapper_339501025136214612_328/latch_enable_in scan_wrapper_339501025136214612_329/latch_enable_in
+ scan_wrapper_339501025136214612_328/scan_select_in scan_wrapper_339501025136214612_329/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_339 scan_wrapper_339501025136214612_339/clk_in scan_wrapper_339501025136214612_340/clk_in
+ scan_wrapper_339501025136214612_339/data_in scan_wrapper_339501025136214612_340/data_in
+ scan_wrapper_339501025136214612_339/latch_enable_in scan_wrapper_339501025136214612_340/latch_enable_in
+ scan_wrapper_339501025136214612_339/scan_select_in scan_wrapper_339501025136214612_340/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341193419111006803_56 scan_wrapper_341193419111006803_56/clk_in scan_wrapper_341266732010177108_57/clk_in
+ scan_wrapper_341193419111006803_56/data_in scan_wrapper_341266732010177108_57/data_in
+ scan_wrapper_341193419111006803_56/latch_enable_in scan_wrapper_341266732010177108_57/latch_enable_in
+ scan_wrapper_341193419111006803_56/scan_select_in scan_wrapper_341266732010177108_57/scan_select_in
+ vccd1 vssd1 scan_wrapper_341193419111006803
Xscan_wrapper_339501025136214612_158 scan_wrapper_339501025136214612_158/clk_in scan_wrapper_339501025136214612_159/clk_in
+ scan_wrapper_339501025136214612_158/data_in scan_wrapper_339501025136214612_159/data_in
+ scan_wrapper_339501025136214612_158/latch_enable_in scan_wrapper_339501025136214612_159/latch_enable_in
+ scan_wrapper_339501025136214612_158/scan_select_in scan_wrapper_339501025136214612_159/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_169 scan_wrapper_339501025136214612_169/clk_in scan_wrapper_339501025136214612_170/clk_in
+ scan_wrapper_339501025136214612_169/data_in scan_wrapper_339501025136214612_170/data_in
+ scan_wrapper_339501025136214612_169/latch_enable_in scan_wrapper_339501025136214612_170/latch_enable_in
+ scan_wrapper_339501025136214612_169/scan_select_in scan_wrapper_339501025136214612_170/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341360223723717202_114 scan_wrapper_341360223723717202_114/clk_in scan_wrapper_341546888233747026_115/clk_in
+ scan_wrapper_341360223723717202_114/data_in scan_wrapper_341546888233747026_115/data_in
+ scan_wrapper_341360223723717202_114/latch_enable_in scan_wrapper_341546888233747026_115/latch_enable_in
+ scan_wrapper_341360223723717202_114/scan_select_in scan_wrapper_341546888233747026_115/scan_select_in
+ vccd1 vssd1 scan_wrapper_341360223723717202
Xscan_wrapper_341590933015364178_128 scan_wrapper_341590933015364178_128/clk_in scan_wrapper_341589685194195540_129/clk_in
+ scan_wrapper_341590933015364178_128/data_in scan_wrapper_341589685194195540_129/data_in
+ scan_wrapper_341590933015364178_128/latch_enable_in scan_wrapper_341589685194195540_129/latch_enable_in
+ scan_wrapper_341590933015364178_128/scan_select_in scan_wrapper_341589685194195540_129/scan_select_in
+ vccd1 vssd1 scan_wrapper_341590933015364178
Xscan_wrapper_341277789473735250_45 scan_wrapper_341277789473735250_45/clk_in scan_wrapper_341263346544149074_46/clk_in
+ scan_wrapper_341277789473735250_45/data_in scan_wrapper_341263346544149074_46/data_in
+ scan_wrapper_341277789473735250_45/latch_enable_in scan_wrapper_341263346544149074_46/latch_enable_in
+ scan_wrapper_341277789473735250_45/scan_select_in scan_wrapper_341263346544149074_46/scan_select_in
+ vccd1 vssd1 scan_wrapper_341277789473735250
Xscan_wrapper_339501025136214612_307 scan_wrapper_339501025136214612_307/clk_in scan_wrapper_339501025136214612_308/clk_in
+ scan_wrapper_339501025136214612_307/data_in scan_wrapper_339501025136214612_308/data_in
+ scan_wrapper_339501025136214612_307/latch_enable_in scan_wrapper_339501025136214612_308/latch_enable_in
+ scan_wrapper_339501025136214612_307/scan_select_in scan_wrapper_339501025136214612_308/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_318 scan_wrapper_339501025136214612_318/clk_in scan_wrapper_339501025136214612_319/clk_in
+ scan_wrapper_339501025136214612_318/data_in scan_wrapper_339501025136214612_319/data_in
+ scan_wrapper_339501025136214612_318/latch_enable_in scan_wrapper_339501025136214612_319/latch_enable_in
+ scan_wrapper_339501025136214612_318/scan_select_in scan_wrapper_339501025136214612_319/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_329 scan_wrapper_339501025136214612_329/clk_in scan_wrapper_339501025136214612_330/clk_in
+ scan_wrapper_339501025136214612_329/data_in scan_wrapper_339501025136214612_330/data_in
+ scan_wrapper_339501025136214612_329/latch_enable_in scan_wrapper_339501025136214612_330/latch_enable_in
+ scan_wrapper_339501025136214612_329/scan_select_in scan_wrapper_339501025136214612_330/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341182944314917460_21 scan_wrapper_341182944314917460_21/clk_in scan_wrapper_341188777753969234_22/clk_in
+ scan_wrapper_341182944314917460_21/data_in scan_wrapper_341188777753969234_22/data_in
+ scan_wrapper_341182944314917460_21/latch_enable_in scan_wrapper_341188777753969234_22/latch_enable_in
+ scan_wrapper_341182944314917460_21/scan_select_in scan_wrapper_341188777753969234_22/scan_select_in
+ vccd1 vssd1 scan_wrapper_341182944314917460
Xscan_wrapper_339501025136214612_159 scan_wrapper_339501025136214612_159/clk_in scan_wrapper_339501025136214612_160/clk_in
+ scan_wrapper_339501025136214612_159/data_in scan_wrapper_339501025136214612_160/data_in
+ scan_wrapper_339501025136214612_159/latch_enable_in scan_wrapper_339501025136214612_160/latch_enable_in
+ scan_wrapper_339501025136214612_159/scan_select_in scan_wrapper_339501025136214612_160/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_490 scan_wrapper_339501025136214612_490/clk_in scan_wrapper_339501025136214612_491/clk_in
+ scan_wrapper_339501025136214612_490/data_in scan_wrapper_339501025136214612_491/data_in
+ scan_wrapper_339501025136214612_490/latch_enable_in scan_wrapper_339501025136214612_491/latch_enable_in
+ scan_wrapper_339501025136214612_490/scan_select_in scan_wrapper_339501025136214612_491/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341259651269001812_53 scan_wrapper_341259651269001812_53/clk_in scan_wrapper_341353928049295956_54/clk_in
+ scan_wrapper_341259651269001812_53/data_in scan_wrapper_341353928049295956_54/data_in
+ scan_wrapper_341259651269001812_53/latch_enable_in scan_wrapper_341353928049295956_54/latch_enable_in
+ scan_wrapper_341259651269001812_53/scan_select_in scan_wrapper_341353928049295956_54/scan_select_in
+ vccd1 vssd1 scan_wrapper_341259651269001812
Xscan_wrapper_341155178824598098_16 scan_wrapper_341155178824598098_16/clk_in scan_wrapper_341167691532337747_17/clk_in
+ scan_wrapper_341155178824598098_16/data_in scan_wrapper_341167691532337747_17/data_in
+ scan_wrapper_341155178824598098_16/latch_enable_in scan_wrapper_341167691532337747_17/latch_enable_in
+ scan_wrapper_341155178824598098_16/scan_select_in scan_wrapper_341167691532337747_17/scan_select_in
+ vccd1 vssd1 scan_wrapper_341155178824598098
Xscan_wrapper_339501025136214612_308 scan_wrapper_339501025136214612_308/clk_in scan_wrapper_339501025136214612_309/clk_in
+ scan_wrapper_339501025136214612_308/data_in scan_wrapper_339501025136214612_309/data_in
+ scan_wrapper_339501025136214612_308/latch_enable_in scan_wrapper_339501025136214612_309/latch_enable_in
+ scan_wrapper_339501025136214612_308/scan_select_in scan_wrapper_339501025136214612_309/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_319 scan_wrapper_339501025136214612_319/clk_in scan_wrapper_339501025136214612_320/clk_in
+ scan_wrapper_339501025136214612_319/data_in scan_wrapper_339501025136214612_320/data_in
+ scan_wrapper_339501025136214612_319/latch_enable_in scan_wrapper_339501025136214612_320/latch_enable_in
+ scan_wrapper_339501025136214612_319/scan_select_in scan_wrapper_339501025136214612_320/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341315210433266259_60 scan_wrapper_341315210433266259_60/clk_in scan_wrapper_341364381657858642_61/clk_in
+ scan_wrapper_341315210433266259_60/data_in scan_wrapper_341364381657858642_61/data_in
+ scan_wrapper_341315210433266259_60/latch_enable_in scan_wrapper_341364381657858642_61/latch_enable_in
+ scan_wrapper_341315210433266259_60/scan_select_in scan_wrapper_341364381657858642_61/scan_select_in
+ vccd1 vssd1 scan_wrapper_341315210433266259
Xscan_wrapper_339501025136214612_491 scan_wrapper_339501025136214612_491/clk_in scan_wrapper_339501025136214612_492/clk_in
+ scan_wrapper_339501025136214612_491/data_in scan_wrapper_339501025136214612_492/data_in
+ scan_wrapper_339501025136214612_491/latch_enable_in scan_wrapper_339501025136214612_492/latch_enable_in
+ scan_wrapper_339501025136214612_491/scan_select_in scan_wrapper_339501025136214612_492/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_480 scan_wrapper_339501025136214612_480/clk_in scan_wrapper_339501025136214612_481/clk_in
+ scan_wrapper_339501025136214612_480/data_in scan_wrapper_339501025136214612_481/data_in
+ scan_wrapper_339501025136214612_480/latch_enable_in scan_wrapper_339501025136214612_481/latch_enable_in
+ scan_wrapper_339501025136214612_480/scan_select_in scan_wrapper_339501025136214612_481/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341174563322724948_40 scan_wrapper_341174563322724948_40/clk_in scan_wrapper_341271902949474898_41/clk_in
+ scan_wrapper_341174563322724948_40/data_in scan_wrapper_341271902949474898_41/data_in
+ scan_wrapper_341174563322724948_40/latch_enable_in scan_wrapper_341271902949474898_41/latch_enable_in
+ scan_wrapper_341174563322724948_40/scan_select_in scan_wrapper_341271902949474898_41/scan_select_in
+ vccd1 vssd1 scan_wrapper_341174563322724948
Xscan_wrapper_341192113929585235_28 scan_wrapper_341192113929585235_28/clk_in scan_wrapper_341192621088047698_29/clk_in
+ scan_wrapper_341192113929585235_28/data_in scan_wrapper_341192621088047698_29/data_in
+ scan_wrapper_341192113929585235_28/latch_enable_in scan_wrapper_341192621088047698_29/latch_enable_in
+ scan_wrapper_341192113929585235_28/scan_select_in scan_wrapper_341192621088047698_29/scan_select_in
+ vccd1 vssd1 scan_wrapper_341192113929585235
Xscan_wrapper_339501025136214612_309 scan_wrapper_339501025136214612_309/clk_in scan_wrapper_339501025136214612_310/clk_in
+ scan_wrapper_339501025136214612_309/data_in scan_wrapper_339501025136214612_310/data_in
+ scan_wrapper_339501025136214612_309/latch_enable_in scan_wrapper_339501025136214612_310/latch_enable_in
+ scan_wrapper_339501025136214612_309/scan_select_in scan_wrapper_339501025136214612_310/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_492 scan_wrapper_339501025136214612_492/clk_in scan_wrapper_339501025136214612_493/clk_in
+ scan_wrapper_339501025136214612_492/data_in scan_wrapper_339501025136214612_493/data_in
+ scan_wrapper_339501025136214612_492/latch_enable_in scan_wrapper_339501025136214612_493/latch_enable_in
+ scan_wrapper_339501025136214612_492/scan_select_in scan_wrapper_339501025136214612_493/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_481 scan_wrapper_339501025136214612_481/clk_in scan_wrapper_339501025136214612_482/clk_in
+ scan_wrapper_339501025136214612_481/data_in scan_wrapper_339501025136214612_482/data_in
+ scan_wrapper_339501025136214612_481/latch_enable_in scan_wrapper_339501025136214612_482/latch_enable_in
+ scan_wrapper_339501025136214612_481/scan_select_in scan_wrapper_339501025136214612_482/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_470 scan_wrapper_339501025136214612_470/clk_in scan_wrapper_339501025136214612_471/clk_in
+ scan_wrapper_339501025136214612_470/data_in scan_wrapper_339501025136214612_471/data_in
+ scan_wrapper_339501025136214612_470/latch_enable_in scan_wrapper_339501025136214612_471/latch_enable_in
+ scan_wrapper_339501025136214612_470/scan_select_in scan_wrapper_339501025136214612_471/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341164228775772755_38 scan_wrapper_341164228775772755_38/clk_in scan_wrapper_341262321634509394_39/clk_in
+ scan_wrapper_341164228775772755_38/data_in scan_wrapper_341262321634509394_39/data_in
+ scan_wrapper_341164228775772755_38/latch_enable_in scan_wrapper_341262321634509394_39/latch_enable_in
+ scan_wrapper_341164228775772755_38/scan_select_in scan_wrapper_341262321634509394_39/scan_select_in
+ vccd1 vssd1 scan_wrapper_341164228775772755
Xscan_wrapper_341614346808328788_136 scan_wrapper_341614346808328788_136/clk_in scan_wrapper_341620484740219475_137/clk_in
+ scan_wrapper_341614346808328788_136/data_in scan_wrapper_341620484740219475_137/data_in
+ scan_wrapper_341614346808328788_136/latch_enable_in scan_wrapper_341620484740219475_137/latch_enable_in
+ scan_wrapper_341614346808328788_136/scan_select_in scan_wrapper_341620484740219475_137/scan_select_in
+ vccd1 vssd1 scan_wrapper_341614346808328788
Xscan_wrapper_341637831098106450_147 scan_wrapper_341637831098106450_147/clk_in scan_wrapper_341631644820570706_148/clk_in
+ scan_wrapper_341637831098106450_147/data_in scan_wrapper_341631644820570706_148/data_in
+ scan_wrapper_341637831098106450_147/latch_enable_in scan_wrapper_341631644820570706_148/latch_enable_in
+ scan_wrapper_341637831098106450_147/scan_select_in scan_wrapper_341631644820570706_148/scan_select_in
+ vccd1 vssd1 scan_wrapper_341637831098106450
Xscan_wrapper_341432030163108435_72 scan_wrapper_341432030163108435_72/clk_in scan_wrapper_341440114308678227_73/clk_in
+ scan_wrapper_341432030163108435_72/data_in scan_wrapper_341440114308678227_73/data_in
+ scan_wrapper_341432030163108435_72/latch_enable_in scan_wrapper_341440114308678227_73/latch_enable_in
+ scan_wrapper_341432030163108435_72/scan_select_in scan_wrapper_341440114308678227_73/scan_select_in
+ vccd1 vssd1 scan_wrapper_341432030163108435
Xscan_wrapper_339501025136214612_493 scan_wrapper_339501025136214612_493/clk_in scan_wrapper_339501025136214612_494/clk_in
+ scan_wrapper_339501025136214612_493/data_in scan_wrapper_339501025136214612_494/data_in
+ scan_wrapper_339501025136214612_493/latch_enable_in scan_wrapper_339501025136214612_494/latch_enable_in
+ scan_wrapper_339501025136214612_493/scan_select_in scan_wrapper_339501025136214612_494/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_482 scan_wrapper_339501025136214612_482/clk_in scan_wrapper_339501025136214612_483/clk_in
+ scan_wrapper_339501025136214612_482/data_in scan_wrapper_339501025136214612_483/data_in
+ scan_wrapper_339501025136214612_482/latch_enable_in scan_wrapper_339501025136214612_483/latch_enable_in
+ scan_wrapper_339501025136214612_482/scan_select_in scan_wrapper_339501025136214612_483/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_460 scan_wrapper_339501025136214612_460/clk_in scan_wrapper_339501025136214612_461/clk_in
+ scan_wrapper_339501025136214612_460/data_in scan_wrapper_339501025136214612_461/data_in
+ scan_wrapper_339501025136214612_460/latch_enable_in scan_wrapper_339501025136214612_461/latch_enable_in
+ scan_wrapper_339501025136214612_460/scan_select_in scan_wrapper_339501025136214612_461/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_471 scan_wrapper_339501025136214612_471/clk_in scan_wrapper_339501025136214612_472/clk_in
+ scan_wrapper_339501025136214612_471/data_in scan_wrapper_339501025136214612_472/data_in
+ scan_wrapper_339501025136214612_471/latch_enable_in scan_wrapper_339501025136214612_472/latch_enable_in
+ scan_wrapper_339501025136214612_471/scan_select_in scan_wrapper_339501025136214612_472/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_290 scan_wrapper_339501025136214612_290/clk_in scan_wrapper_339501025136214612_291/clk_in
+ scan_wrapper_339501025136214612_290/data_in scan_wrapper_339501025136214612_291/data_in
+ scan_wrapper_339501025136214612_290/latch_enable_in scan_wrapper_339501025136214612_291/latch_enable_in
+ scan_wrapper_339501025136214612_290/scan_select_in scan_wrapper_339501025136214612_291/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_340596276030603858_149 scan_wrapper_340596276030603858_149/clk_in scan_wrapper_341678527574180436_150/clk_in
+ scan_wrapper_340596276030603858_149/data_in scan_wrapper_341678527574180436_150/data_in
+ scan_wrapper_340596276030603858_149/latch_enable_in scan_wrapper_341678527574180436_150/latch_enable_in
+ scan_wrapper_340596276030603858_149/scan_select_in scan_wrapper_341678527574180436_150/scan_select_in
+ vccd1 vssd1 scan_wrapper_340596276030603858
Xscan_wrapper_341235973870322258_32 scan_wrapper_341235973870322258_32/clk_in scan_wrapper_341235575572922964_33/clk_in
+ scan_wrapper_341235973870322258_32/data_in scan_wrapper_341235575572922964_33/data_in
+ scan_wrapper_341235973870322258_32/latch_enable_in scan_wrapper_341235575572922964_33/latch_enable_in
+ scan_wrapper_341235973870322258_32/scan_select_in scan_wrapper_341235575572922964_33/scan_select_in
+ vccd1 vssd1 scan_wrapper_341235973870322258
Xscan_wrapper_341163800289870419_12 scan_wrapper_341163800289870419_12/clk_in scan_wrapper_341160271679586899_13/clk_in
+ scan_wrapper_341163800289870419_12/data_in scan_wrapper_341160271679586899_13/data_in
+ scan_wrapper_341163800289870419_12/latch_enable_in scan_wrapper_341160271679586899_13/latch_enable_in
+ scan_wrapper_341163800289870419_12/scan_select_in scan_wrapper_341160271679586899_13/scan_select_in
+ vccd1 vssd1 scan_wrapper_341163800289870419
Xscan_wrapper_341404507891040852_66 scan_wrapper_341404507891040852_66/clk_in scan_wrapper_341410909669818963_67/clk_in
+ scan_wrapper_341404507891040852_66/data_in scan_wrapper_341410909669818963_67/data_in
+ scan_wrapper_341404507891040852_66/latch_enable_in scan_wrapper_341410909669818963_67/latch_enable_in
+ scan_wrapper_341404507891040852_66/scan_select_in scan_wrapper_341410909669818963_67/scan_select_in
+ vccd1 vssd1 scan_wrapper_341404507891040852
Xscan_wrapper_341558189536313940_119 scan_wrapper_341558189536313940_119/clk_in scan_wrapper_341538994733974098_120/clk_in
+ scan_wrapper_341558189536313940_119/data_in scan_wrapper_341538994733974098_120/data_in
+ scan_wrapper_341558189536313940_119/latch_enable_in scan_wrapper_341538994733974098_120/latch_enable_in
+ scan_wrapper_341558189536313940_119/scan_select_in scan_wrapper_341538994733974098_120/scan_select_in
+ vccd1 vssd1 scan_wrapper_341558189536313940
Xscan_wrapper_339501025136214612_494 scan_wrapper_339501025136214612_494/clk_in scan_wrapper_339501025136214612_495/clk_in
+ scan_wrapper_339501025136214612_494/data_in scan_wrapper_339501025136214612_495/data_in
+ scan_wrapper_339501025136214612_494/latch_enable_in scan_wrapper_339501025136214612_495/latch_enable_in
+ scan_wrapper_339501025136214612_494/scan_select_in scan_wrapper_339501025136214612_495/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_483 scan_wrapper_339501025136214612_483/clk_in scan_wrapper_339501025136214612_484/clk_in
+ scan_wrapper_339501025136214612_483/data_in scan_wrapper_339501025136214612_484/data_in
+ scan_wrapper_339501025136214612_483/latch_enable_in scan_wrapper_339501025136214612_484/latch_enable_in
+ scan_wrapper_339501025136214612_483/scan_select_in scan_wrapper_339501025136214612_484/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_461 scan_wrapper_339501025136214612_461/clk_in scan_wrapper_339501025136214612_462/clk_in
+ scan_wrapper_339501025136214612_461/data_in scan_wrapper_339501025136214612_462/data_in
+ scan_wrapper_339501025136214612_461/latch_enable_in scan_wrapper_339501025136214612_462/latch_enable_in
+ scan_wrapper_339501025136214612_461/scan_select_in scan_wrapper_339501025136214612_462/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_472 scan_wrapper_339501025136214612_472/clk_in scan_wrapper_339501025136214612_473/clk_in
+ scan_wrapper_339501025136214612_472/data_in scan_wrapper_339501025136214612_473/data_in
+ scan_wrapper_339501025136214612_472/latch_enable_in scan_wrapper_339501025136214612_473/latch_enable_in
+ scan_wrapper_339501025136214612_472/scan_select_in scan_wrapper_339501025136214612_473/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_450 scan_wrapper_339501025136214612_450/clk_in scan_wrapper_339501025136214612_451/clk_in
+ scan_wrapper_339501025136214612_450/data_in scan_wrapper_339501025136214612_451/data_in
+ scan_wrapper_339501025136214612_450/latch_enable_in scan_wrapper_339501025136214612_451/latch_enable_in
+ scan_wrapper_339501025136214612_450/scan_select_in scan_wrapper_339501025136214612_451/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_280 scan_wrapper_339501025136214612_280/clk_in scan_wrapper_339501025136214612_281/clk_in
+ scan_wrapper_339501025136214612_280/data_in scan_wrapper_339501025136214612_281/data_in
+ scan_wrapper_339501025136214612_280/latch_enable_in scan_wrapper_339501025136214612_281/latch_enable_in
+ scan_wrapper_339501025136214612_280/scan_select_in scan_wrapper_339501025136214612_281/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_291 scan_wrapper_339501025136214612_291/clk_in scan_wrapper_339501025136214612_292/clk_in
+ scan_wrapper_339501025136214612_291/data_in scan_wrapper_339501025136214612_292/data_in
+ scan_wrapper_339501025136214612_291/latch_enable_in scan_wrapper_339501025136214612_292/latch_enable_in
+ scan_wrapper_339501025136214612_291/scan_select_in scan_wrapper_339501025136214612_292/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341473139924927058_108 scan_wrapper_341473139924927058_108/clk_in scan_wrapper_341528610027340372_109/clk_in
+ scan_wrapper_341473139924927058_108/data_in scan_wrapper_341528610027340372_109/data_in
+ scan_wrapper_341473139924927058_108/latch_enable_in scan_wrapper_341528610027340372_109/latch_enable_in
+ scan_wrapper_341473139924927058_108/scan_select_in scan_wrapper_341528610027340372_109/scan_select_in
+ vccd1 vssd1 scan_wrapper_341473139924927058
Xscan_wrapper_339501025136214612_495 scan_wrapper_339501025136214612_495/clk_in scan_wrapper_339501025136214612_496/clk_in
+ scan_wrapper_339501025136214612_495/data_in scan_wrapper_339501025136214612_496/data_in
+ scan_wrapper_339501025136214612_495/latch_enable_in scan_wrapper_339501025136214612_496/latch_enable_in
+ scan_wrapper_339501025136214612_495/scan_select_in scan_wrapper_339501025136214612_496/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_484 scan_wrapper_339501025136214612_484/clk_in scan_wrapper_339501025136214612_485/clk_in
+ scan_wrapper_339501025136214612_484/data_in scan_wrapper_339501025136214612_485/data_in
+ scan_wrapper_339501025136214612_484/latch_enable_in scan_wrapper_339501025136214612_485/latch_enable_in
+ scan_wrapper_339501025136214612_484/scan_select_in scan_wrapper_339501025136214612_485/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_462 scan_wrapper_339501025136214612_462/clk_in scan_wrapper_339501025136214612_463/clk_in
+ scan_wrapper_339501025136214612_462/data_in scan_wrapper_339501025136214612_463/data_in
+ scan_wrapper_339501025136214612_462/latch_enable_in scan_wrapper_339501025136214612_463/latch_enable_in
+ scan_wrapper_339501025136214612_462/scan_select_in scan_wrapper_339501025136214612_463/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_473 scan_wrapper_339501025136214612_473/clk_in scan_wrapper_339501025136214612_474/clk_in
+ scan_wrapper_339501025136214612_473/data_in scan_wrapper_339501025136214612_474/data_in
+ scan_wrapper_339501025136214612_473/latch_enable_in scan_wrapper_339501025136214612_474/latch_enable_in
+ scan_wrapper_339501025136214612_473/scan_select_in scan_wrapper_339501025136214612_474/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_451 scan_wrapper_339501025136214612_451/clk_in scan_wrapper_339501025136214612_452/clk_in
+ scan_wrapper_339501025136214612_451/data_in scan_wrapper_339501025136214612_452/data_in
+ scan_wrapper_339501025136214612_451/latch_enable_in scan_wrapper_339501025136214612_452/latch_enable_in
+ scan_wrapper_339501025136214612_451/scan_select_in scan_wrapper_339501025136214612_452/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_440 scan_wrapper_339501025136214612_440/clk_in scan_wrapper_339501025136214612_441/clk_in
+ scan_wrapper_339501025136214612_440/data_in scan_wrapper_339501025136214612_441/data_in
+ scan_wrapper_339501025136214612_440/latch_enable_in scan_wrapper_339501025136214612_441/latch_enable_in
+ scan_wrapper_339501025136214612_440/scan_select_in scan_wrapper_339501025136214612_441/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341431339142087251_71 scan_wrapper_341431339142087251_71/clk_in scan_wrapper_341432030163108435_72/clk_in
+ scan_wrapper_341431339142087251_71/data_in scan_wrapper_341432030163108435_72/data_in
+ scan_wrapper_341431339142087251_71/latch_enable_in scan_wrapper_341432030163108435_72/latch_enable_in
+ scan_wrapper_341431339142087251_71/scan_select_in scan_wrapper_341432030163108435_72/scan_select_in
+ vccd1 vssd1 scan_wrapper_341431339142087251
Xscan_wrapper_339501025136214612_270 scan_wrapper_339501025136214612_270/clk_in scan_wrapper_339501025136214612_271/clk_in
+ scan_wrapper_339501025136214612_270/data_in scan_wrapper_339501025136214612_271/data_in
+ scan_wrapper_339501025136214612_270/latch_enable_in scan_wrapper_339501025136214612_271/latch_enable_in
+ scan_wrapper_339501025136214612_270/scan_select_in scan_wrapper_339501025136214612_271/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_281 scan_wrapper_339501025136214612_281/clk_in scan_wrapper_339501025136214612_282/clk_in
+ scan_wrapper_339501025136214612_281/data_in scan_wrapper_339501025136214612_282/data_in
+ scan_wrapper_339501025136214612_281/latch_enable_in scan_wrapper_339501025136214612_282/latch_enable_in
+ scan_wrapper_339501025136214612_281/scan_select_in scan_wrapper_339501025136214612_282/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_292 scan_wrapper_339501025136214612_292/clk_in scan_wrapper_339501025136214612_293/clk_in
+ scan_wrapper_339501025136214612_292/data_in scan_wrapper_339501025136214612_293/data_in
+ scan_wrapper_339501025136214612_292/latch_enable_in scan_wrapper_339501025136214612_293/latch_enable_in
+ scan_wrapper_339501025136214612_292/scan_select_in scan_wrapper_339501025136214612_293/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341482086419399252_85 scan_wrapper_341482086419399252_85/clk_in scan_wrapper_341452019534398035_86/clk_in
+ scan_wrapper_341482086419399252_85/data_in scan_wrapper_341452019534398035_86/data_in
+ scan_wrapper_341482086419399252_85/latch_enable_in scan_wrapper_341452019534398035_86/latch_enable_in
+ scan_wrapper_341482086419399252_85/scan_select_in scan_wrapper_341452019534398035_86/scan_select_in
+ vccd1 vssd1 scan_wrapper_341482086419399252
Xscan_wrapper_340661930553246290_5 scan_wrapper_340661930553246290_5/clk_in scan_wrapper_341136771628663380_6/clk_in
+ scan_wrapper_340661930553246290_5/data_in scan_wrapper_341136771628663380_6/data_in
+ scan_wrapper_340661930553246290_5/latch_enable_in scan_wrapper_341136771628663380_6/latch_enable_in
+ scan_wrapper_340661930553246290_5/scan_select_in scan_wrapper_341136771628663380_6/scan_select_in
+ vccd1 vssd1 scan_wrapper_340661930553246290
Xscan_wrapper_339501025136214612_496 scan_wrapper_339501025136214612_496/clk_in scan_wrapper_339501025136214612_497/clk_in
+ scan_wrapper_339501025136214612_496/data_in scan_wrapper_339501025136214612_497/data_in
+ scan_wrapper_339501025136214612_496/latch_enable_in scan_wrapper_339501025136214612_497/latch_enable_in
+ scan_wrapper_339501025136214612_496/scan_select_in scan_wrapper_339501025136214612_497/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_485 scan_wrapper_339501025136214612_485/clk_in scan_wrapper_339501025136214612_486/clk_in
+ scan_wrapper_339501025136214612_485/data_in scan_wrapper_339501025136214612_486/data_in
+ scan_wrapper_339501025136214612_485/latch_enable_in scan_wrapper_339501025136214612_486/latch_enable_in
+ scan_wrapper_339501025136214612_485/scan_select_in scan_wrapper_339501025136214612_486/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_463 scan_wrapper_339501025136214612_463/clk_in scan_wrapper_339501025136214612_464/clk_in
+ scan_wrapper_339501025136214612_463/data_in scan_wrapper_339501025136214612_464/data_in
+ scan_wrapper_339501025136214612_463/latch_enable_in scan_wrapper_339501025136214612_464/latch_enable_in
+ scan_wrapper_339501025136214612_463/scan_select_in scan_wrapper_339501025136214612_464/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_474 scan_wrapper_339501025136214612_474/clk_in scan_wrapper_339501025136214612_475/clk_in
+ scan_wrapper_339501025136214612_474/data_in scan_wrapper_339501025136214612_475/data_in
+ scan_wrapper_339501025136214612_474/latch_enable_in scan_wrapper_339501025136214612_475/latch_enable_in
+ scan_wrapper_339501025136214612_474/scan_select_in scan_wrapper_339501025136214612_475/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_452 scan_wrapper_339501025136214612_452/clk_in scan_wrapper_339501025136214612_453/clk_in
+ scan_wrapper_339501025136214612_452/data_in scan_wrapper_339501025136214612_453/data_in
+ scan_wrapper_339501025136214612_452/latch_enable_in scan_wrapper_339501025136214612_453/latch_enable_in
+ scan_wrapper_339501025136214612_452/scan_select_in scan_wrapper_339501025136214612_453/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_441 scan_wrapper_339501025136214612_441/clk_in scan_wrapper_339501025136214612_442/clk_in
+ scan_wrapper_339501025136214612_441/data_in scan_wrapper_339501025136214612_442/data_in
+ scan_wrapper_339501025136214612_441/latch_enable_in scan_wrapper_339501025136214612_442/latch_enable_in
+ scan_wrapper_339501025136214612_441/scan_select_in scan_wrapper_339501025136214612_442/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_430 scan_wrapper_339501025136214612_430/clk_in scan_wrapper_339501025136214612_431/clk_in
+ scan_wrapper_339501025136214612_430/data_in scan_wrapper_339501025136214612_431/data_in
+ scan_wrapper_339501025136214612_430/latch_enable_in scan_wrapper_339501025136214612_431/latch_enable_in
+ scan_wrapper_339501025136214612_430/scan_select_in scan_wrapper_339501025136214612_431/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341154068332282450_10 scan_wrapper_341159915403870803_9/clk_out scan_wrapper_341160201697624660_11/clk_in
+ scan_wrapper_341159915403870803_9/data_out scan_wrapper_341160201697624660_11/data_in
+ scan_wrapper_341159915403870803_9/latch_enable_out scan_wrapper_341160201697624660_11/latch_enable_in
+ scan_wrapper_341159915403870803_9/scan_select_out scan_wrapper_341160201697624660_11/scan_select_in
+ vccd1 vssd1 scan_wrapper_341154068332282450
Xscan_wrapper_339501025136214612_271 scan_wrapper_339501025136214612_271/clk_in scan_wrapper_339501025136214612_272/clk_in
+ scan_wrapper_339501025136214612_271/data_in scan_wrapper_339501025136214612_272/data_in
+ scan_wrapper_339501025136214612_271/latch_enable_in scan_wrapper_339501025136214612_272/latch_enable_in
+ scan_wrapper_339501025136214612_271/scan_select_in scan_wrapper_339501025136214612_272/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_260 scan_wrapper_339501025136214612_260/clk_in scan_wrapper_339501025136214612_261/clk_in
+ scan_wrapper_339501025136214612_260/data_in scan_wrapper_339501025136214612_261/data_in
+ scan_wrapper_339501025136214612_260/latch_enable_in scan_wrapper_339501025136214612_261/latch_enable_in
+ scan_wrapper_339501025136214612_260/scan_select_in scan_wrapper_339501025136214612_261/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_282 scan_wrapper_339501025136214612_282/clk_in scan_wrapper_339501025136214612_283/clk_in
+ scan_wrapper_339501025136214612_282/data_in scan_wrapper_339501025136214612_283/data_in
+ scan_wrapper_339501025136214612_282/latch_enable_in scan_wrapper_339501025136214612_283/latch_enable_in
+ scan_wrapper_339501025136214612_282/scan_select_in scan_wrapper_339501025136214612_283/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_293 scan_wrapper_339501025136214612_293/clk_in scan_wrapper_339501025136214612_294/clk_in
+ scan_wrapper_339501025136214612_293/data_in scan_wrapper_339501025136214612_294/data_in
+ scan_wrapper_339501025136214612_293/latch_enable_in scan_wrapper_339501025136214612_294/latch_enable_in
+ scan_wrapper_339501025136214612_293/scan_select_in scan_wrapper_339501025136214612_294/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341438392303616596_79 scan_wrapper_341438392303616596_79/clk_in scan_wrapper_341432284947153491_80/clk_in
+ scan_wrapper_341438392303616596_79/data_in scan_wrapper_341432284947153491_80/data_in
+ scan_wrapper_341438392303616596_79/latch_enable_in scan_wrapper_341432284947153491_80/latch_enable_in
+ scan_wrapper_341438392303616596_79/scan_select_in scan_wrapper_341432284947153491_80/scan_select_in
+ vccd1 vssd1 scan_wrapper_341438392303616596
Xscan_wrapper_341521390605697619_101 scan_wrapper_341521390605697619_101/clk_in scan_wrapper_341243232292700755_102/clk_in
+ scan_wrapper_341521390605697619_101/data_in scan_wrapper_341243232292700755_102/data_in
+ scan_wrapper_341521390605697619_101/latch_enable_in scan_wrapper_341243232292700755_102/latch_enable_in
+ scan_wrapper_341521390605697619_101/scan_select_in scan_wrapper_341243232292700755_102/scan_select_in
+ vccd1 vssd1 scan_wrapper_341521390605697619
Xscan_wrapper_341440781874102868_75 scan_wrapper_341440781874102868_75/clk_in scan_wrapper_341444501414347346_76/clk_in
+ scan_wrapper_341440781874102868_75/data_in scan_wrapper_341444501414347346_76/data_in
+ scan_wrapper_341440781874102868_75/latch_enable_in scan_wrapper_341444501414347346_76/latch_enable_in
+ scan_wrapper_341440781874102868_75/scan_select_in scan_wrapper_341444501414347346_76/scan_select_in
+ vccd1 vssd1 scan_wrapper_341440781874102868
Xscan_wrapper_341224613878956628_31 scan_wrapper_341224613878956628_31/clk_in scan_wrapper_341235973870322258_32/clk_in
+ scan_wrapper_341224613878956628_31/data_in scan_wrapper_341235973870322258_32/data_in
+ scan_wrapper_341224613878956628_31/latch_enable_in scan_wrapper_341235973870322258_32/latch_enable_in
+ scan_wrapper_341224613878956628_31/scan_select_in scan_wrapper_341235973870322258_32/scan_select_in
+ vccd1 vssd1 scan_wrapper_341224613878956628
Xscan_wrapper_341541108650607187_113 scan_wrapper_hamming74_112/clk_out scan_wrapper_341360223723717202_114/clk_in
+ scan_wrapper_hamming74_112/data_out scan_wrapper_341360223723717202_114/data_in
+ scan_wrapper_hamming74_112/latch_enable_out scan_wrapper_341360223723717202_114/latch_enable_in
+ scan_wrapper_hamming74_112/scan_select_out scan_wrapper_341360223723717202_114/scan_select_in
+ vccd1 vssd1 scan_wrapper_341541108650607187
Xscan_wrapper_341344337258349139_51 scan_wrapper_341344337258349139_51/clk_in scan_wrapper_341342096033055316_52/clk_in
+ scan_wrapper_341344337258349139_51/data_in scan_wrapper_341342096033055316_52/data_in
+ scan_wrapper_341344337258349139_51/latch_enable_in scan_wrapper_341342096033055316_52/latch_enable_in
+ scan_wrapper_341344337258349139_51/scan_select_in scan_wrapper_341342096033055316_52/scan_select_in
+ vccd1 vssd1 scan_wrapper_341344337258349139
Xscan_wrapper_339501025136214612_497 scan_wrapper_339501025136214612_497/clk_in scan_controller/scan_clk_in
+ scan_wrapper_339501025136214612_497/data_in scan_controller/scan_data_in scan_wrapper_339501025136214612_497/latch_enable_in
+ scan_wrapper_339501025136214612_497/latch_enable_out scan_wrapper_339501025136214612_497/scan_select_in
+ scan_wrapper_339501025136214612_497/scan_select_out vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_486 scan_wrapper_339501025136214612_486/clk_in scan_wrapper_339501025136214612_487/clk_in
+ scan_wrapper_339501025136214612_486/data_in scan_wrapper_339501025136214612_487/data_in
+ scan_wrapper_339501025136214612_486/latch_enable_in scan_wrapper_339501025136214612_487/latch_enable_in
+ scan_wrapper_339501025136214612_486/scan_select_in scan_wrapper_339501025136214612_487/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_464 scan_wrapper_339501025136214612_464/clk_in scan_wrapper_339501025136214612_465/clk_in
+ scan_wrapper_339501025136214612_464/data_in scan_wrapper_339501025136214612_465/data_in
+ scan_wrapper_339501025136214612_464/latch_enable_in scan_wrapper_339501025136214612_465/latch_enable_in
+ scan_wrapper_339501025136214612_464/scan_select_in scan_wrapper_339501025136214612_465/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_475 scan_wrapper_339501025136214612_475/clk_in scan_wrapper_339501025136214612_476/clk_in
+ scan_wrapper_339501025136214612_475/data_in scan_wrapper_339501025136214612_476/data_in
+ scan_wrapper_339501025136214612_475/latch_enable_in scan_wrapper_339501025136214612_476/latch_enable_in
+ scan_wrapper_339501025136214612_475/scan_select_in scan_wrapper_339501025136214612_476/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_453 scan_wrapper_339501025136214612_453/clk_in scan_wrapper_339501025136214612_454/clk_in
+ scan_wrapper_339501025136214612_453/data_in scan_wrapper_339501025136214612_454/data_in
+ scan_wrapper_339501025136214612_453/latch_enable_in scan_wrapper_339501025136214612_454/latch_enable_in
+ scan_wrapper_339501025136214612_453/scan_select_in scan_wrapper_339501025136214612_454/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_442 scan_wrapper_339501025136214612_442/clk_in scan_wrapper_339501025136214612_443/clk_in
+ scan_wrapper_339501025136214612_442/data_in scan_wrapper_339501025136214612_443/data_in
+ scan_wrapper_339501025136214612_442/latch_enable_in scan_wrapper_339501025136214612_443/latch_enable_in
+ scan_wrapper_339501025136214612_442/scan_select_in scan_wrapper_339501025136214612_443/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_420 scan_wrapper_339501025136214612_420/clk_in scan_wrapper_339501025136214612_421/clk_in
+ scan_wrapper_339501025136214612_420/data_in scan_wrapper_339501025136214612_421/data_in
+ scan_wrapper_339501025136214612_420/latch_enable_in scan_wrapper_339501025136214612_421/latch_enable_in
+ scan_wrapper_339501025136214612_420/scan_select_in scan_wrapper_339501025136214612_421/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_431 scan_wrapper_339501025136214612_431/clk_in scan_wrapper_339501025136214612_432/clk_in
+ scan_wrapper_339501025136214612_431/data_in scan_wrapper_339501025136214612_432/data_in
+ scan_wrapper_339501025136214612_431/latch_enable_in scan_wrapper_339501025136214612_432/latch_enable_in
+ scan_wrapper_339501025136214612_431/scan_select_in scan_wrapper_339501025136214612_432/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_250 scan_wrapper_339501025136214612_250/clk_in scan_wrapper_339501025136214612_251/clk_in
+ scan_wrapper_339501025136214612_250/data_in scan_wrapper_339501025136214612_251/data_in
+ scan_wrapper_339501025136214612_250/latch_enable_in scan_wrapper_339501025136214612_251/latch_enable_in
+ scan_wrapper_339501025136214612_250/scan_select_in scan_wrapper_339501025136214612_251/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_272 scan_wrapper_339501025136214612_272/clk_in scan_wrapper_339501025136214612_273/clk_in
+ scan_wrapper_339501025136214612_272/data_in scan_wrapper_339501025136214612_273/data_in
+ scan_wrapper_339501025136214612_272/latch_enable_in scan_wrapper_339501025136214612_273/latch_enable_in
+ scan_wrapper_339501025136214612_272/scan_select_in scan_wrapper_339501025136214612_273/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_261 scan_wrapper_339501025136214612_261/clk_in scan_wrapper_339501025136214612_262/clk_in
+ scan_wrapper_339501025136214612_261/data_in scan_wrapper_339501025136214612_262/data_in
+ scan_wrapper_339501025136214612_261/latch_enable_in scan_wrapper_339501025136214612_262/latch_enable_in
+ scan_wrapper_339501025136214612_261/scan_select_in scan_wrapper_339501025136214612_262/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_283 scan_wrapper_339501025136214612_283/clk_in scan_wrapper_339501025136214612_284/clk_in
+ scan_wrapper_339501025136214612_283/data_in scan_wrapper_339501025136214612_284/data_in
+ scan_wrapper_339501025136214612_283/latch_enable_in scan_wrapper_339501025136214612_284/latch_enable_in
+ scan_wrapper_339501025136214612_283/scan_select_in scan_wrapper_339501025136214612_284/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_294 scan_wrapper_339501025136214612_294/clk_in scan_wrapper_339501025136214612_295/clk_in
+ scan_wrapper_339501025136214612_294/data_in scan_wrapper_339501025136214612_295/data_in
+ scan_wrapper_339501025136214612_294/latch_enable_in scan_wrapper_339501025136214612_295/latch_enable_in
+ scan_wrapper_339501025136214612_294/scan_select_in scan_wrapper_339501025136214612_295/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341457494561784402_127 scan_wrapper_341457494561784402_127/clk_in scan_wrapper_341590933015364178_128/clk_in
+ scan_wrapper_341457494561784402_127/data_in scan_wrapper_341590933015364178_128/data_in
+ scan_wrapper_341457494561784402_127/latch_enable_in scan_wrapper_341590933015364178_128/latch_enable_in
+ scan_wrapper_341457494561784402_127/scan_select_in scan_wrapper_341590933015364178_128/scan_select_in
+ vccd1 vssd1 scan_wrapper_341457494561784402
Xscan_wrapper_341497964482527828_88 scan_wrapper_341497964482527828_88/clk_in scan_wrapper_341497938559631956_89/clk_in
+ scan_wrapper_341497964482527828_88/data_in scan_wrapper_341497938559631956_89/data_in
+ scan_wrapper_341497964482527828_88/latch_enable_in scan_wrapper_341497938559631956_89/latch_enable_in
+ scan_wrapper_341497964482527828_88/scan_select_in scan_wrapper_341497938559631956_89/scan_select_in
+ vccd1 vssd1 scan_wrapper_341497964482527828
Xscan_wrapper_339501025136214612_487 scan_wrapper_339501025136214612_487/clk_in scan_wrapper_339501025136214612_488/clk_in
+ scan_wrapper_339501025136214612_487/data_in scan_wrapper_339501025136214612_488/data_in
+ scan_wrapper_339501025136214612_487/latch_enable_in scan_wrapper_339501025136214612_488/latch_enable_in
+ scan_wrapper_339501025136214612_487/scan_select_in scan_wrapper_339501025136214612_488/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_465 scan_wrapper_339501025136214612_465/clk_in scan_wrapper_339501025136214612_466/clk_in
+ scan_wrapper_339501025136214612_465/data_in scan_wrapper_339501025136214612_466/data_in
+ scan_wrapper_339501025136214612_465/latch_enable_in scan_wrapper_339501025136214612_466/latch_enable_in
+ scan_wrapper_339501025136214612_465/scan_select_in scan_wrapper_339501025136214612_466/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_476 scan_wrapper_339501025136214612_476/clk_in scan_wrapper_339501025136214612_477/clk_in
+ scan_wrapper_339501025136214612_476/data_in scan_wrapper_339501025136214612_477/data_in
+ scan_wrapper_339501025136214612_476/latch_enable_in scan_wrapper_339501025136214612_477/latch_enable_in
+ scan_wrapper_339501025136214612_476/scan_select_in scan_wrapper_339501025136214612_477/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_454 scan_wrapper_339501025136214612_454/clk_in scan_wrapper_339501025136214612_455/clk_in
+ scan_wrapper_339501025136214612_454/data_in scan_wrapper_339501025136214612_455/data_in
+ scan_wrapper_339501025136214612_454/latch_enable_in scan_wrapper_339501025136214612_455/latch_enable_in
+ scan_wrapper_339501025136214612_454/scan_select_in scan_wrapper_339501025136214612_455/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_443 scan_wrapper_339501025136214612_443/clk_in scan_wrapper_339501025136214612_444/clk_in
+ scan_wrapper_339501025136214612_443/data_in scan_wrapper_339501025136214612_444/data_in
+ scan_wrapper_339501025136214612_443/latch_enable_in scan_wrapper_339501025136214612_444/latch_enable_in
+ scan_wrapper_339501025136214612_443/scan_select_in scan_wrapper_339501025136214612_444/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_421 scan_wrapper_339501025136214612_421/clk_in scan_wrapper_339501025136214612_422/clk_in
+ scan_wrapper_339501025136214612_421/data_in scan_wrapper_339501025136214612_422/data_in
+ scan_wrapper_339501025136214612_421/latch_enable_in scan_wrapper_339501025136214612_422/latch_enable_in
+ scan_wrapper_339501025136214612_421/scan_select_in scan_wrapper_339501025136214612_422/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_432 scan_wrapper_339501025136214612_432/clk_in scan_wrapper_339501025136214612_433/clk_in
+ scan_wrapper_339501025136214612_432/data_in scan_wrapper_339501025136214612_433/data_in
+ scan_wrapper_339501025136214612_432/latch_enable_in scan_wrapper_339501025136214612_433/latch_enable_in
+ scan_wrapper_339501025136214612_432/scan_select_in scan_wrapper_339501025136214612_433/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_410 scan_wrapper_339501025136214612_410/clk_in scan_wrapper_339501025136214612_411/clk_in
+ scan_wrapper_339501025136214612_410/data_in scan_wrapper_339501025136214612_411/data_in
+ scan_wrapper_339501025136214612_410/latch_enable_in scan_wrapper_339501025136214612_411/latch_enable_in
+ scan_wrapper_339501025136214612_410/scan_select_in scan_wrapper_339501025136214612_411/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341493393195532884_92 scan_wrapper_341493393195532884_92/clk_in scan_wrapper_341506274933867090_93/clk_in
+ scan_wrapper_341493393195532884_92/data_in scan_wrapper_341506274933867090_93/data_in
+ scan_wrapper_341493393195532884_92/latch_enable_in scan_wrapper_341506274933867090_93/latch_enable_in
+ scan_wrapper_341493393195532884_92/scan_select_in scan_wrapper_341506274933867090_93/scan_select_in
+ vccd1 vssd1 scan_wrapper_341493393195532884
Xscan_wrapper_339501025136214612_240 scan_wrapper_339501025136214612_240/clk_in scan_wrapper_339501025136214612_241/clk_in
+ scan_wrapper_339501025136214612_240/data_in scan_wrapper_339501025136214612_241/data_in
+ scan_wrapper_339501025136214612_240/latch_enable_in scan_wrapper_339501025136214612_241/latch_enable_in
+ scan_wrapper_339501025136214612_240/scan_select_in scan_wrapper_339501025136214612_241/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_251 scan_wrapper_339501025136214612_251/clk_in scan_wrapper_339501025136214612_252/clk_in
+ scan_wrapper_339501025136214612_251/data_in scan_wrapper_339501025136214612_252/data_in
+ scan_wrapper_339501025136214612_251/latch_enable_in scan_wrapper_339501025136214612_252/latch_enable_in
+ scan_wrapper_339501025136214612_251/scan_select_in scan_wrapper_339501025136214612_252/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_273 scan_wrapper_339501025136214612_273/clk_in scan_wrapper_339501025136214612_274/clk_in
+ scan_wrapper_339501025136214612_273/data_in scan_wrapper_339501025136214612_274/data_in
+ scan_wrapper_339501025136214612_273/latch_enable_in scan_wrapper_339501025136214612_274/latch_enable_in
+ scan_wrapper_339501025136214612_273/scan_select_in scan_wrapper_339501025136214612_274/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_262 scan_wrapper_339501025136214612_262/clk_in scan_wrapper_339501025136214612_263/clk_in
+ scan_wrapper_339501025136214612_262/data_in scan_wrapper_339501025136214612_263/data_in
+ scan_wrapper_339501025136214612_262/latch_enable_in scan_wrapper_339501025136214612_263/latch_enable_in
+ scan_wrapper_339501025136214612_262/scan_select_in scan_wrapper_339501025136214612_263/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_284 scan_wrapper_339501025136214612_284/clk_in scan_wrapper_339501025136214612_285/clk_in
+ scan_wrapper_339501025136214612_284/data_in scan_wrapper_339501025136214612_285/data_in
+ scan_wrapper_339501025136214612_284/latch_enable_in scan_wrapper_339501025136214612_285/latch_enable_in
+ scan_wrapper_339501025136214612_284/scan_select_in scan_wrapper_339501025136214612_285/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_295 scan_wrapper_339501025136214612_295/clk_in scan_wrapper_339501025136214612_296/clk_in
+ scan_wrapper_339501025136214612_295/data_in scan_wrapper_339501025136214612_296/data_in
+ scan_wrapper_339501025136214612_295/latch_enable_in scan_wrapper_339501025136214612_296/latch_enable_in
+ scan_wrapper_339501025136214612_295/scan_select_in scan_wrapper_339501025136214612_296/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341499976001520211_90 scan_wrapper_341499976001520211_90/clk_in scan_wrapper_341500800901579348_91/clk_in
+ scan_wrapper_341499976001520211_90/data_in scan_wrapper_341500800901579348_91/data_in
+ scan_wrapper_341499976001520211_90/latch_enable_in scan_wrapper_341500800901579348_91/latch_enable_in
+ scan_wrapper_341499976001520211_90/scan_select_in scan_wrapper_341500800901579348_91/scan_select_in
+ vccd1 vssd1 scan_wrapper_341499976001520211
Xscan_wrapper_341410909669818963_67 scan_wrapper_341410909669818963_67/clk_in scan_wrapper_341063825089364563_68/clk_in
+ scan_wrapper_341410909669818963_67/data_in scan_wrapper_341063825089364563_68/data_in
+ scan_wrapper_341410909669818963_67/latch_enable_in scan_wrapper_341063825089364563_68/latch_enable_in
+ scan_wrapper_341410909669818963_67/scan_select_in scan_wrapper_341063825089364563_68/scan_select_in
+ vccd1 vssd1 scan_wrapper_341410909669818963
Xscan_wrapper_341620484740219475_137 scan_wrapper_341620484740219475_137/clk_in scan_wrapper_341624400621077076_138/clk_in
+ scan_wrapper_341620484740219475_137/data_in scan_wrapper_341624400621077076_138/data_in
+ scan_wrapper_341620484740219475_137/latch_enable_in scan_wrapper_341624400621077076_138/latch_enable_in
+ scan_wrapper_341620484740219475_137/scan_select_in scan_wrapper_341624400621077076_138/scan_select_in
+ vccd1 vssd1 scan_wrapper_341620484740219475
Xscan_wrapper_339501025136214612_488 scan_wrapper_339501025136214612_488/clk_in scan_wrapper_339501025136214612_489/clk_in
+ scan_wrapper_339501025136214612_488/data_in scan_wrapper_339501025136214612_489/data_in
+ scan_wrapper_339501025136214612_488/latch_enable_in scan_wrapper_339501025136214612_489/latch_enable_in
+ scan_wrapper_339501025136214612_488/scan_select_in scan_wrapper_339501025136214612_489/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_466 scan_wrapper_339501025136214612_466/clk_in scan_wrapper_339501025136214612_467/clk_in
+ scan_wrapper_339501025136214612_466/data_in scan_wrapper_339501025136214612_467/data_in
+ scan_wrapper_339501025136214612_466/latch_enable_in scan_wrapper_339501025136214612_467/latch_enable_in
+ scan_wrapper_339501025136214612_466/scan_select_in scan_wrapper_339501025136214612_467/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_477 scan_wrapper_339501025136214612_477/clk_in scan_wrapper_339501025136214612_478/clk_in
+ scan_wrapper_339501025136214612_477/data_in scan_wrapper_339501025136214612_478/data_in
+ scan_wrapper_339501025136214612_477/latch_enable_in scan_wrapper_339501025136214612_478/latch_enable_in
+ scan_wrapper_339501025136214612_477/scan_select_in scan_wrapper_339501025136214612_478/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_455 scan_wrapper_339501025136214612_455/clk_in scan_wrapper_339501025136214612_456/clk_in
+ scan_wrapper_339501025136214612_455/data_in scan_wrapper_339501025136214612_456/data_in
+ scan_wrapper_339501025136214612_455/latch_enable_in scan_wrapper_339501025136214612_456/latch_enable_in
+ scan_wrapper_339501025136214612_455/scan_select_in scan_wrapper_339501025136214612_456/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_444 scan_wrapper_339501025136214612_444/clk_in scan_wrapper_339501025136214612_445/clk_in
+ scan_wrapper_339501025136214612_444/data_in scan_wrapper_339501025136214612_445/data_in
+ scan_wrapper_339501025136214612_444/latch_enable_in scan_wrapper_339501025136214612_445/latch_enable_in
+ scan_wrapper_339501025136214612_444/scan_select_in scan_wrapper_339501025136214612_445/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_422 scan_wrapper_339501025136214612_422/clk_in scan_wrapper_339501025136214612_423/clk_in
+ scan_wrapper_339501025136214612_422/data_in scan_wrapper_339501025136214612_423/data_in
+ scan_wrapper_339501025136214612_422/latch_enable_in scan_wrapper_339501025136214612_423/latch_enable_in
+ scan_wrapper_339501025136214612_422/scan_select_in scan_wrapper_339501025136214612_423/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_433 scan_wrapper_339501025136214612_433/clk_in scan_wrapper_339501025136214612_434/clk_in
+ scan_wrapper_339501025136214612_433/data_in scan_wrapper_339501025136214612_434/data_in
+ scan_wrapper_339501025136214612_433/latch_enable_in scan_wrapper_339501025136214612_434/latch_enable_in
+ scan_wrapper_339501025136214612_433/scan_select_in scan_wrapper_339501025136214612_434/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_411 scan_wrapper_339501025136214612_411/clk_in scan_wrapper_339501025136214612_412/clk_in
+ scan_wrapper_339501025136214612_411/data_in scan_wrapper_339501025136214612_412/data_in
+ scan_wrapper_339501025136214612_411/latch_enable_in scan_wrapper_339501025136214612_412/latch_enable_in
+ scan_wrapper_339501025136214612_411/scan_select_in scan_wrapper_339501025136214612_412/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_400 scan_wrapper_339501025136214612_400/clk_in scan_wrapper_339501025136214612_401/clk_in
+ scan_wrapper_339501025136214612_400/data_in scan_wrapper_339501025136214612_401/data_in
+ scan_wrapper_339501025136214612_400/latch_enable_in scan_wrapper_339501025136214612_401/latch_enable_in
+ scan_wrapper_339501025136214612_400/scan_select_in scan_wrapper_339501025136214612_401/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_230 scan_wrapper_339501025136214612_230/clk_in scan_wrapper_339501025136214612_231/clk_in
+ scan_wrapper_339501025136214612_230/data_in scan_wrapper_339501025136214612_231/data_in
+ scan_wrapper_339501025136214612_230/latch_enable_in scan_wrapper_339501025136214612_231/latch_enable_in
+ scan_wrapper_339501025136214612_230/scan_select_in scan_wrapper_339501025136214612_231/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_241 scan_wrapper_339501025136214612_241/clk_in scan_wrapper_339501025136214612_242/clk_in
+ scan_wrapper_339501025136214612_241/data_in scan_wrapper_339501025136214612_242/data_in
+ scan_wrapper_339501025136214612_241/latch_enable_in scan_wrapper_339501025136214612_242/latch_enable_in
+ scan_wrapper_339501025136214612_241/scan_select_in scan_wrapper_339501025136214612_242/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_252 scan_wrapper_339501025136214612_252/clk_in scan_wrapper_339501025136214612_253/clk_in
+ scan_wrapper_339501025136214612_252/data_in scan_wrapper_339501025136214612_253/data_in
+ scan_wrapper_339501025136214612_252/latch_enable_in scan_wrapper_339501025136214612_253/latch_enable_in
+ scan_wrapper_339501025136214612_252/scan_select_in scan_wrapper_339501025136214612_253/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_274 scan_wrapper_339501025136214612_274/clk_in scan_wrapper_339501025136214612_275/clk_in
+ scan_wrapper_339501025136214612_274/data_in scan_wrapper_339501025136214612_275/data_in
+ scan_wrapper_339501025136214612_274/latch_enable_in scan_wrapper_339501025136214612_275/latch_enable_in
+ scan_wrapper_339501025136214612_274/scan_select_in scan_wrapper_339501025136214612_275/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_263 scan_wrapper_339501025136214612_263/clk_in scan_wrapper_339501025136214612_264/clk_in
+ scan_wrapper_339501025136214612_263/data_in scan_wrapper_339501025136214612_264/data_in
+ scan_wrapper_339501025136214612_263/latch_enable_in scan_wrapper_339501025136214612_264/latch_enable_in
+ scan_wrapper_339501025136214612_263/scan_select_in scan_wrapper_339501025136214612_264/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_285 scan_wrapper_339501025136214612_285/clk_in scan_wrapper_339501025136214612_286/clk_in
+ scan_wrapper_339501025136214612_285/data_in scan_wrapper_339501025136214612_286/data_in
+ scan_wrapper_339501025136214612_285/latch_enable_in scan_wrapper_339501025136214612_286/latch_enable_in
+ scan_wrapper_339501025136214612_285/scan_select_in scan_wrapper_339501025136214612_286/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_296 scan_wrapper_339501025136214612_296/clk_in scan_wrapper_339501025136214612_297/clk_in
+ scan_wrapper_339501025136214612_296/data_in scan_wrapper_339501025136214612_297/data_in
+ scan_wrapper_339501025136214612_296/latch_enable_in scan_wrapper_339501025136214612_297/latch_enable_in
+ scan_wrapper_339501025136214612_296/scan_select_in scan_wrapper_339501025136214612_297/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341339883600609876_50 scan_wrapper_341339883600609876_50/clk_in scan_wrapper_341344337258349139_51/clk_in
+ scan_wrapper_341339883600609876_50/data_in scan_wrapper_341344337258349139_51/data_in
+ scan_wrapper_341339883600609876_50/latch_enable_in scan_wrapper_341344337258349139_51/latch_enable_in
+ scan_wrapper_341339883600609876_50/scan_select_in scan_wrapper_341344337258349139_51/scan_select_in
+ vccd1 vssd1 scan_wrapper_341339883600609876
Xscan_wrapper_341490465660469844_125 scan_wrapper_341490465660469844_125/clk_in scan_wrapper_341581732833657427_126/clk_in
+ scan_wrapper_341490465660469844_125/data_in scan_wrapper_341581732833657427_126/data_in
+ scan_wrapper_341490465660469844_125/latch_enable_in scan_wrapper_341581732833657427_126/latch_enable_in
+ scan_wrapper_341490465660469844_125/scan_select_in scan_wrapper_341581732833657427_126/scan_select_in
+ vccd1 vssd1 scan_wrapper_341490465660469844
Xscan_wrapper_341608574336631379_130 scan_wrapper_341608574336631379_130/clk_in scan_wrapper_341608297106768466_131/clk_in
+ scan_wrapper_341608574336631379_130/data_in scan_wrapper_341608297106768466_131/data_in
+ scan_wrapper_341608574336631379_130/latch_enable_in scan_wrapper_341608297106768466_131/latch_enable_in
+ scan_wrapper_341608574336631379_130/scan_select_in scan_wrapper_341608297106768466_131/scan_select_in
+ vccd1 vssd1 scan_wrapper_341608574336631379
Xscan_wrapper_341802655228625490_63 scan_wrapper_341802655228625490_63/clk_in scan_wrapper_341382703379120723_64/clk_in
+ scan_wrapper_341802655228625490_63/data_in scan_wrapper_341382703379120723_64/data_in
+ scan_wrapper_341802655228625490_63/latch_enable_in scan_wrapper_341382703379120723_64/latch_enable_in
+ scan_wrapper_341802655228625490_63/scan_select_in scan_wrapper_341382703379120723_64/scan_select_in
+ vccd1 vssd1 scan_wrapper_341802655228625490
Xscan_wrapper_339501025136214612_423 scan_wrapper_339501025136214612_423/clk_in scan_wrapper_339501025136214612_424/clk_in
+ scan_wrapper_339501025136214612_423/data_in scan_wrapper_339501025136214612_424/data_in
+ scan_wrapper_339501025136214612_423/latch_enable_in scan_wrapper_339501025136214612_424/latch_enable_in
+ scan_wrapper_339501025136214612_423/scan_select_in scan_wrapper_339501025136214612_424/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_434 scan_wrapper_339501025136214612_434/clk_in scan_wrapper_339501025136214612_435/clk_in
+ scan_wrapper_339501025136214612_434/data_in scan_wrapper_339501025136214612_435/data_in
+ scan_wrapper_339501025136214612_434/latch_enable_in scan_wrapper_339501025136214612_435/latch_enable_in
+ scan_wrapper_339501025136214612_434/scan_select_in scan_wrapper_339501025136214612_435/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_412 scan_wrapper_339501025136214612_412/clk_in scan_wrapper_339501025136214612_413/clk_in
+ scan_wrapper_339501025136214612_412/data_in scan_wrapper_339501025136214612_413/data_in
+ scan_wrapper_339501025136214612_412/latch_enable_in scan_wrapper_339501025136214612_413/latch_enable_in
+ scan_wrapper_339501025136214612_412/scan_select_in scan_wrapper_339501025136214612_413/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_401 scan_wrapper_339501025136214612_401/clk_in scan_wrapper_339501025136214612_402/clk_in
+ scan_wrapper_339501025136214612_401/data_in scan_wrapper_339501025136214612_402/data_in
+ scan_wrapper_339501025136214612_401/latch_enable_in scan_wrapper_339501025136214612_402/latch_enable_in
+ scan_wrapper_339501025136214612_401/scan_select_in scan_wrapper_339501025136214612_402/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_489 scan_wrapper_339501025136214612_489/clk_in scan_wrapper_339501025136214612_490/clk_in
+ scan_wrapper_339501025136214612_489/data_in scan_wrapper_339501025136214612_490/data_in
+ scan_wrapper_339501025136214612_489/latch_enable_in scan_wrapper_339501025136214612_490/latch_enable_in
+ scan_wrapper_339501025136214612_489/scan_select_in scan_wrapper_339501025136214612_490/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_478 scan_wrapper_339501025136214612_478/clk_in scan_wrapper_339501025136214612_479/clk_in
+ scan_wrapper_339501025136214612_478/data_in scan_wrapper_339501025136214612_479/data_in
+ scan_wrapper_339501025136214612_478/latch_enable_in scan_wrapper_339501025136214612_479/latch_enable_in
+ scan_wrapper_339501025136214612_478/scan_select_in scan_wrapper_339501025136214612_479/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_467 scan_wrapper_339501025136214612_467/clk_in scan_wrapper_339501025136214612_468/clk_in
+ scan_wrapper_339501025136214612_467/data_in scan_wrapper_339501025136214612_468/data_in
+ scan_wrapper_339501025136214612_467/latch_enable_in scan_wrapper_339501025136214612_468/latch_enable_in
+ scan_wrapper_339501025136214612_467/scan_select_in scan_wrapper_339501025136214612_468/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_456 scan_wrapper_339501025136214612_456/clk_in scan_wrapper_339501025136214612_457/clk_in
+ scan_wrapper_339501025136214612_456/data_in scan_wrapper_339501025136214612_457/data_in
+ scan_wrapper_339501025136214612_456/latch_enable_in scan_wrapper_339501025136214612_457/latch_enable_in
+ scan_wrapper_339501025136214612_456/scan_select_in scan_wrapper_339501025136214612_457/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_445 scan_wrapper_339501025136214612_445/clk_in scan_wrapper_339501025136214612_446/clk_in
+ scan_wrapper_339501025136214612_445/data_in scan_wrapper_339501025136214612_446/data_in
+ scan_wrapper_339501025136214612_445/latch_enable_in scan_wrapper_339501025136214612_446/latch_enable_in
+ scan_wrapper_339501025136214612_445/scan_select_in scan_wrapper_339501025136214612_446/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_231 scan_wrapper_339501025136214612_231/clk_in scan_wrapper_339501025136214612_232/clk_in
+ scan_wrapper_339501025136214612_231/data_in scan_wrapper_339501025136214612_232/data_in
+ scan_wrapper_339501025136214612_231/latch_enable_in scan_wrapper_339501025136214612_232/latch_enable_in
+ scan_wrapper_339501025136214612_231/scan_select_in scan_wrapper_339501025136214612_232/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_220 scan_wrapper_339501025136214612_220/clk_in scan_wrapper_339501025136214612_221/clk_in
+ scan_wrapper_339501025136214612_220/data_in scan_wrapper_339501025136214612_221/data_in
+ scan_wrapper_339501025136214612_220/latch_enable_in scan_wrapper_339501025136214612_221/latch_enable_in
+ scan_wrapper_339501025136214612_220/scan_select_in scan_wrapper_339501025136214612_221/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_242 scan_wrapper_339501025136214612_242/clk_in scan_wrapper_339501025136214612_243/clk_in
+ scan_wrapper_339501025136214612_242/data_in scan_wrapper_339501025136214612_243/data_in
+ scan_wrapper_339501025136214612_242/latch_enable_in scan_wrapper_339501025136214612_243/latch_enable_in
+ scan_wrapper_339501025136214612_242/scan_select_in scan_wrapper_339501025136214612_243/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_253 scan_wrapper_339501025136214612_253/clk_in scan_wrapper_339501025136214612_254/clk_in
+ scan_wrapper_339501025136214612_253/data_in scan_wrapper_339501025136214612_254/data_in
+ scan_wrapper_339501025136214612_253/latch_enable_in scan_wrapper_339501025136214612_254/latch_enable_in
+ scan_wrapper_339501025136214612_253/scan_select_in scan_wrapper_339501025136214612_254/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_275 scan_wrapper_339501025136214612_275/clk_in scan_wrapper_339501025136214612_276/clk_in
+ scan_wrapper_339501025136214612_275/data_in scan_wrapper_339501025136214612_276/data_in
+ scan_wrapper_339501025136214612_275/latch_enable_in scan_wrapper_339501025136214612_276/latch_enable_in
+ scan_wrapper_339501025136214612_275/scan_select_in scan_wrapper_339501025136214612_276/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_264 scan_wrapper_339501025136214612_264/clk_in scan_wrapper_339501025136214612_265/clk_in
+ scan_wrapper_339501025136214612_264/data_in scan_wrapper_339501025136214612_265/data_in
+ scan_wrapper_339501025136214612_264/latch_enable_in scan_wrapper_339501025136214612_265/latch_enable_in
+ scan_wrapper_339501025136214612_264/scan_select_in scan_wrapper_339501025136214612_265/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_286 scan_wrapper_339501025136214612_286/clk_in scan_wrapper_339501025136214612_287/clk_in
+ scan_wrapper_339501025136214612_286/data_in scan_wrapper_339501025136214612_287/data_in
+ scan_wrapper_339501025136214612_286/latch_enable_in scan_wrapper_339501025136214612_287/latch_enable_in
+ scan_wrapper_339501025136214612_286/scan_select_in scan_wrapper_339501025136214612_287/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_297 scan_wrapper_339501025136214612_297/clk_in scan_wrapper_339501025136214612_298/clk_in
+ scan_wrapper_339501025136214612_297/data_in scan_wrapper_339501025136214612_298/data_in
+ scan_wrapper_339501025136214612_297/latch_enable_in scan_wrapper_339501025136214612_298/latch_enable_in
+ scan_wrapper_339501025136214612_297/scan_select_in scan_wrapper_339501025136214612_298/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341063825089364563_68 scan_wrapper_341063825089364563_68/clk_in scan_wrapper_341174480471589458_69/clk_in
+ scan_wrapper_341063825089364563_68/data_in scan_wrapper_341174480471589458_69/data_in
+ scan_wrapper_341063825089364563_68/latch_enable_in scan_wrapper_341174480471589458_69/latch_enable_in
+ scan_wrapper_341063825089364563_68/scan_select_in scan_wrapper_341174480471589458_69/scan_select_in
+ vccd1 vssd1 scan_wrapper_341063825089364563
Xscan_wrapper_341332847867462227_48 scan_wrapper_341332847867462227_48/clk_in scan_wrapper_341337976625693266_49/clk_in
+ scan_wrapper_341332847867462227_48/data_in scan_wrapper_341337976625693266_49/data_in
+ scan_wrapper_341332847867462227_48/latch_enable_in scan_wrapper_341337976625693266_49/latch_enable_in
+ scan_wrapper_341332847867462227_48/scan_select_in scan_wrapper_341337976625693266_49/scan_select_in
+ vccd1 vssd1 scan_wrapper_341332847867462227
Xscan_wrapper_341136771628663380_6 scan_wrapper_341136771628663380_6/clk_in scan_wrapper_339800239192932947_7/clk_in
+ scan_wrapper_341136771628663380_6/data_in scan_wrapper_339800239192932947_7/data_in
+ scan_wrapper_341136771628663380_6/latch_enable_in scan_wrapper_339800239192932947_7/latch_enable_in
+ scan_wrapper_341136771628663380_6/scan_select_in scan_wrapper_339800239192932947_7/scan_select_in
+ vccd1 vssd1 scan_wrapper_341136771628663380
Xscan_wrapper_341424636358034002_110 scan_wrapper_341424636358034002_110/clk_in scan_wrapper_341717091617866324_111/clk_in
+ scan_wrapper_341424636358034002_110/data_in scan_wrapper_341717091617866324_111/data_in
+ scan_wrapper_341424636358034002_110/latch_enable_in scan_wrapper_341717091617866324_111/latch_enable_in
+ scan_wrapper_341424636358034002_110/scan_select_in scan_wrapper_341717091617866324_111/scan_select_in
+ vccd1 vssd1 scan_wrapper_341424636358034002
Xscan_wrapper_341440114308678227_73 scan_wrapper_341440114308678227_73/clk_in scan_wrapper_341496918381167187_74/clk_in
+ scan_wrapper_341440114308678227_73/data_in scan_wrapper_341496918381167187_74/data_in
+ scan_wrapper_341440114308678227_73/latch_enable_in scan_wrapper_341496918381167187_74/latch_enable_in
+ scan_wrapper_341440114308678227_73/scan_select_in scan_wrapper_341496918381167187_74/scan_select_in
+ vccd1 vssd1 scan_wrapper_341440114308678227
Xscan_wrapper_339501025136214612_479 scan_wrapper_339501025136214612_479/clk_in scan_wrapper_339501025136214612_480/clk_in
+ scan_wrapper_339501025136214612_479/data_in scan_wrapper_339501025136214612_480/data_in
+ scan_wrapper_339501025136214612_479/latch_enable_in scan_wrapper_339501025136214612_480/latch_enable_in
+ scan_wrapper_339501025136214612_479/scan_select_in scan_wrapper_339501025136214612_480/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_468 scan_wrapper_339501025136214612_468/clk_in scan_wrapper_339501025136214612_469/clk_in
+ scan_wrapper_339501025136214612_468/data_in scan_wrapper_339501025136214612_469/data_in
+ scan_wrapper_339501025136214612_468/latch_enable_in scan_wrapper_339501025136214612_469/latch_enable_in
+ scan_wrapper_339501025136214612_468/scan_select_in scan_wrapper_339501025136214612_469/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_457 scan_wrapper_339501025136214612_457/clk_in scan_wrapper_339501025136214612_458/clk_in
+ scan_wrapper_339501025136214612_457/data_in scan_wrapper_339501025136214612_458/data_in
+ scan_wrapper_339501025136214612_457/latch_enable_in scan_wrapper_339501025136214612_458/latch_enable_in
+ scan_wrapper_339501025136214612_457/scan_select_in scan_wrapper_339501025136214612_458/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_446 scan_wrapper_339501025136214612_446/clk_in scan_wrapper_339501025136214612_447/clk_in
+ scan_wrapper_339501025136214612_446/data_in scan_wrapper_339501025136214612_447/data_in
+ scan_wrapper_339501025136214612_446/latch_enable_in scan_wrapper_339501025136214612_447/latch_enable_in
+ scan_wrapper_339501025136214612_446/scan_select_in scan_wrapper_339501025136214612_447/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_424 scan_wrapper_339501025136214612_424/clk_in scan_wrapper_339501025136214612_425/clk_in
+ scan_wrapper_339501025136214612_424/data_in scan_wrapper_339501025136214612_425/data_in
+ scan_wrapper_339501025136214612_424/latch_enable_in scan_wrapper_339501025136214612_425/latch_enable_in
+ scan_wrapper_339501025136214612_424/scan_select_in scan_wrapper_339501025136214612_425/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_435 scan_wrapper_339501025136214612_435/clk_in scan_wrapper_339501025136214612_436/clk_in
+ scan_wrapper_339501025136214612_435/data_in scan_wrapper_339501025136214612_436/data_in
+ scan_wrapper_339501025136214612_435/latch_enable_in scan_wrapper_339501025136214612_436/latch_enable_in
+ scan_wrapper_339501025136214612_435/scan_select_in scan_wrapper_339501025136214612_436/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_413 scan_wrapper_339501025136214612_413/clk_in scan_wrapper_339501025136214612_414/clk_in
+ scan_wrapper_339501025136214612_413/data_in scan_wrapper_339501025136214612_414/data_in
+ scan_wrapper_339501025136214612_413/latch_enable_in scan_wrapper_339501025136214612_414/latch_enable_in
+ scan_wrapper_339501025136214612_413/scan_select_in scan_wrapper_339501025136214612_414/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_402 scan_wrapper_339501025136214612_402/clk_in scan_wrapper_339501025136214612_403/clk_in
+ scan_wrapper_339501025136214612_402/data_in scan_wrapper_339501025136214612_403/data_in
+ scan_wrapper_339501025136214612_402/latch_enable_in scan_wrapper_339501025136214612_403/latch_enable_in
+ scan_wrapper_339501025136214612_402/scan_select_in scan_wrapper_339501025136214612_403/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_210 scan_wrapper_339501025136214612_210/clk_in scan_wrapper_339501025136214612_211/clk_in
+ scan_wrapper_339501025136214612_210/data_in scan_wrapper_339501025136214612_211/data_in
+ scan_wrapper_339501025136214612_210/latch_enable_in scan_wrapper_339501025136214612_211/latch_enable_in
+ scan_wrapper_339501025136214612_210/scan_select_in scan_wrapper_339501025136214612_211/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_232 scan_wrapper_339501025136214612_232/clk_in scan_wrapper_339501025136214612_233/clk_in
+ scan_wrapper_339501025136214612_232/data_in scan_wrapper_339501025136214612_233/data_in
+ scan_wrapper_339501025136214612_232/latch_enable_in scan_wrapper_339501025136214612_233/latch_enable_in
+ scan_wrapper_339501025136214612_232/scan_select_in scan_wrapper_339501025136214612_233/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_221 scan_wrapper_339501025136214612_221/clk_in scan_wrapper_339501025136214612_222/clk_in
+ scan_wrapper_339501025136214612_221/data_in scan_wrapper_339501025136214612_222/data_in
+ scan_wrapper_339501025136214612_221/latch_enable_in scan_wrapper_339501025136214612_222/latch_enable_in
+ scan_wrapper_339501025136214612_221/scan_select_in scan_wrapper_339501025136214612_222/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_243 scan_wrapper_339501025136214612_243/clk_in scan_wrapper_339501025136214612_244/clk_in
+ scan_wrapper_339501025136214612_243/data_in scan_wrapper_339501025136214612_244/data_in
+ scan_wrapper_339501025136214612_243/latch_enable_in scan_wrapper_339501025136214612_244/latch_enable_in
+ scan_wrapper_339501025136214612_243/scan_select_in scan_wrapper_339501025136214612_244/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_254 scan_wrapper_339501025136214612_254/clk_in scan_wrapper_339501025136214612_255/clk_in
+ scan_wrapper_339501025136214612_254/data_in scan_wrapper_339501025136214612_255/data_in
+ scan_wrapper_339501025136214612_254/latch_enable_in scan_wrapper_339501025136214612_255/latch_enable_in
+ scan_wrapper_339501025136214612_254/scan_select_in scan_wrapper_339501025136214612_255/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_276 scan_wrapper_339501025136214612_276/clk_in scan_wrapper_339501025136214612_277/clk_in
+ scan_wrapper_339501025136214612_276/data_in scan_wrapper_339501025136214612_277/data_in
+ scan_wrapper_339501025136214612_276/latch_enable_in scan_wrapper_339501025136214612_277/latch_enable_in
+ scan_wrapper_339501025136214612_276/scan_select_in scan_wrapper_339501025136214612_277/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_265 scan_wrapper_339501025136214612_265/clk_in scan_wrapper_339501025136214612_266/clk_in
+ scan_wrapper_339501025136214612_265/data_in scan_wrapper_339501025136214612_266/data_in
+ scan_wrapper_339501025136214612_265/latch_enable_in scan_wrapper_339501025136214612_266/latch_enable_in
+ scan_wrapper_339501025136214612_265/scan_select_in scan_wrapper_339501025136214612_266/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_287 scan_wrapper_339501025136214612_287/clk_in scan_wrapper_339501025136214612_288/clk_in
+ scan_wrapper_339501025136214612_287/data_in scan_wrapper_339501025136214612_288/data_in
+ scan_wrapper_339501025136214612_287/latch_enable_in scan_wrapper_339501025136214612_288/latch_enable_in
+ scan_wrapper_339501025136214612_287/scan_select_in scan_wrapper_339501025136214612_288/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_298 scan_wrapper_339501025136214612_298/clk_in scan_wrapper_339501025136214612_299/clk_in
+ scan_wrapper_339501025136214612_298/data_in scan_wrapper_339501025136214612_299/data_in
+ scan_wrapper_339501025136214612_298/latch_enable_in scan_wrapper_339501025136214612_299/latch_enable_in
+ scan_wrapper_339501025136214612_298/scan_select_in scan_wrapper_339501025136214612_299/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341178154799333971_18 scan_wrapper_341178154799333971_18/clk_in scan_wrapper_341178481588044372_19/clk_in
+ scan_wrapper_341178154799333971_18/data_in scan_wrapper_341178481588044372_19/data_in
+ scan_wrapper_341178154799333971_18/latch_enable_in scan_wrapper_341178481588044372_19/latch_enable_in
+ scan_wrapper_341178154799333971_18/scan_select_in scan_wrapper_341178481588044372_19/scan_select_in
+ vccd1 vssd1 scan_wrapper_341178154799333971
Xscan_wrapper_341497938559631956_89 scan_wrapper_341497938559631956_89/clk_in scan_wrapper_341499976001520211_90/clk_in
+ scan_wrapper_341497938559631956_89/data_in scan_wrapper_341499976001520211_90/data_in
+ scan_wrapper_341497938559631956_89/latch_enable_in scan_wrapper_341499976001520211_90/latch_enable_in
+ scan_wrapper_341497938559631956_89/scan_select_in scan_wrapper_341499976001520211_90/scan_select_in
+ vccd1 vssd1 scan_wrapper_341497938559631956
Xscan_wrapper_341452019534398035_86 scan_wrapper_341452019534398035_86/clk_in scan_wrapper_341497971083313748_87/clk_in
+ scan_wrapper_341452019534398035_86/data_in scan_wrapper_341497971083313748_87/data_in
+ scan_wrapper_341452019534398035_86/latch_enable_in scan_wrapper_341497971083313748_87/latch_enable_in
+ scan_wrapper_341452019534398035_86/scan_select_in scan_wrapper_341497971083313748_87/scan_select_in
+ vccd1 vssd1 scan_wrapper_341452019534398035
Xscan_wrapper_341500800901579348_91 scan_wrapper_341500800901579348_91/clk_in scan_wrapper_341493393195532884_92/clk_in
+ scan_wrapper_341500800901579348_91/data_in scan_wrapper_341493393195532884_92/data_in
+ scan_wrapper_341500800901579348_91/latch_enable_in scan_wrapper_341493393195532884_92/latch_enable_in
+ scan_wrapper_341500800901579348_91/scan_select_in scan_wrapper_341493393195532884_92/scan_select_in
+ vccd1 vssd1 scan_wrapper_341500800901579348
Xscan_wrapper_341419328215712339_70 scan_wrapper_341419328215712339_70/clk_in scan_wrapper_341431339142087251_71/clk_in
+ scan_wrapper_341419328215712339_70/data_in scan_wrapper_341431339142087251_71/data_in
+ scan_wrapper_341419328215712339_70/latch_enable_in scan_wrapper_341431339142087251_71/latch_enable_in
+ scan_wrapper_341419328215712339_70/scan_select_in scan_wrapper_341431339142087251_71/scan_select_in
+ vccd1 vssd1 scan_wrapper_341419328215712339
Xscan_wrapper_341160201697624660_11 scan_wrapper_341160201697624660_11/clk_in scan_wrapper_341163800289870419_12/clk_in
+ scan_wrapper_341160201697624660_11/data_in scan_wrapper_341163800289870419_12/data_in
+ scan_wrapper_341160201697624660_11/latch_enable_in scan_wrapper_341163800289870419_12/latch_enable_in
+ scan_wrapper_341160201697624660_11/scan_select_in scan_wrapper_341163800289870419_12/scan_select_in
+ vccd1 vssd1 scan_wrapper_341160201697624660
Xscan_wrapper_339501025136214612_458 scan_wrapper_339501025136214612_458/clk_in scan_wrapper_339501025136214612_459/clk_in
+ scan_wrapper_339501025136214612_458/data_in scan_wrapper_339501025136214612_459/data_in
+ scan_wrapper_339501025136214612_458/latch_enable_in scan_wrapper_339501025136214612_459/latch_enable_in
+ scan_wrapper_339501025136214612_458/scan_select_in scan_wrapper_339501025136214612_459/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_469 scan_wrapper_339501025136214612_469/clk_in scan_wrapper_339501025136214612_470/clk_in
+ scan_wrapper_339501025136214612_469/data_in scan_wrapper_339501025136214612_470/data_in
+ scan_wrapper_339501025136214612_469/latch_enable_in scan_wrapper_339501025136214612_470/latch_enable_in
+ scan_wrapper_339501025136214612_469/scan_select_in scan_wrapper_339501025136214612_470/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_447 scan_wrapper_339501025136214612_447/clk_in scan_wrapper_339501025136214612_448/clk_in
+ scan_wrapper_339501025136214612_447/data_in scan_wrapper_339501025136214612_448/data_in
+ scan_wrapper_339501025136214612_447/latch_enable_in scan_wrapper_339501025136214612_448/latch_enable_in
+ scan_wrapper_339501025136214612_447/scan_select_in scan_wrapper_339501025136214612_448/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_425 scan_wrapper_339501025136214612_425/clk_in scan_wrapper_339501025136214612_426/clk_in
+ scan_wrapper_339501025136214612_425/data_in scan_wrapper_339501025136214612_426/data_in
+ scan_wrapper_339501025136214612_425/latch_enable_in scan_wrapper_339501025136214612_426/latch_enable_in
+ scan_wrapper_339501025136214612_425/scan_select_in scan_wrapper_339501025136214612_426/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_436 scan_wrapper_339501025136214612_436/clk_in scan_wrapper_339501025136214612_437/clk_in
+ scan_wrapper_339501025136214612_436/data_in scan_wrapper_339501025136214612_437/data_in
+ scan_wrapper_339501025136214612_436/latch_enable_in scan_wrapper_339501025136214612_437/latch_enable_in
+ scan_wrapper_339501025136214612_436/scan_select_in scan_wrapper_339501025136214612_437/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_414 scan_wrapper_339501025136214612_414/clk_in scan_wrapper_339501025136214612_415/clk_in
+ scan_wrapper_339501025136214612_414/data_in scan_wrapper_339501025136214612_415/data_in
+ scan_wrapper_339501025136214612_414/latch_enable_in scan_wrapper_339501025136214612_415/latch_enable_in
+ scan_wrapper_339501025136214612_414/scan_select_in scan_wrapper_339501025136214612_415/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_403 scan_wrapper_339501025136214612_403/clk_in scan_wrapper_339501025136214612_404/clk_in
+ scan_wrapper_339501025136214612_403/data_in scan_wrapper_339501025136214612_404/data_in
+ scan_wrapper_339501025136214612_403/latch_enable_in scan_wrapper_339501025136214612_404/latch_enable_in
+ scan_wrapper_339501025136214612_403/scan_select_in scan_wrapper_339501025136214612_404/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341342096033055316_52 scan_wrapper_341342096033055316_52/clk_in scan_wrapper_341259651269001812_53/clk_in
+ scan_wrapper_341342096033055316_52/data_in scan_wrapper_341259651269001812_53/data_in
+ scan_wrapper_341342096033055316_52/latch_enable_in scan_wrapper_341259651269001812_53/latch_enable_in
+ scan_wrapper_341342096033055316_52/scan_select_in scan_wrapper_341259651269001812_53/scan_select_in
+ vccd1 vssd1 scan_wrapper_341342096033055316
Xscan_wrapper_341462925422101075_97 scan_wrapper_341462925422101075_97/clk_in scan_wrapper_341520747710120530_98/clk_in
+ scan_wrapper_341462925422101075_97/data_in scan_wrapper_341520747710120530_98/data_in
+ scan_wrapper_341462925422101075_97/latch_enable_in scan_wrapper_341520747710120530_98/latch_enable_in
+ scan_wrapper_341462925422101075_97/scan_select_in scan_wrapper_341520747710120530_98/scan_select_in
+ vccd1 vssd1 scan_wrapper_341462925422101075
Xscan_wrapper_339501025136214612_200 scan_wrapper_339501025136214612_200/clk_in scan_wrapper_339501025136214612_201/clk_in
+ scan_wrapper_339501025136214612_200/data_in scan_wrapper_339501025136214612_201/data_in
+ scan_wrapper_339501025136214612_200/latch_enable_in scan_wrapper_339501025136214612_201/latch_enable_in
+ scan_wrapper_339501025136214612_200/scan_select_in scan_wrapper_339501025136214612_201/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_211 scan_wrapper_339501025136214612_211/clk_in scan_wrapper_339501025136214612_212/clk_in
+ scan_wrapper_339501025136214612_211/data_in scan_wrapper_339501025136214612_212/data_in
+ scan_wrapper_339501025136214612_211/latch_enable_in scan_wrapper_339501025136214612_212/latch_enable_in
+ scan_wrapper_339501025136214612_211/scan_select_in scan_wrapper_339501025136214612_212/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_233 scan_wrapper_339501025136214612_233/clk_in scan_wrapper_339501025136214612_234/clk_in
+ scan_wrapper_339501025136214612_233/data_in scan_wrapper_339501025136214612_234/data_in
+ scan_wrapper_339501025136214612_233/latch_enable_in scan_wrapper_339501025136214612_234/latch_enable_in
+ scan_wrapper_339501025136214612_233/scan_select_in scan_wrapper_339501025136214612_234/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_222 scan_wrapper_339501025136214612_222/clk_in scan_wrapper_339501025136214612_223/clk_in
+ scan_wrapper_339501025136214612_222/data_in scan_wrapper_339501025136214612_223/data_in
+ scan_wrapper_339501025136214612_222/latch_enable_in scan_wrapper_339501025136214612_223/latch_enable_in
+ scan_wrapper_339501025136214612_222/scan_select_in scan_wrapper_339501025136214612_223/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_244 scan_wrapper_339501025136214612_244/clk_in scan_wrapper_339501025136214612_245/clk_in
+ scan_wrapper_339501025136214612_244/data_in scan_wrapper_339501025136214612_245/data_in
+ scan_wrapper_339501025136214612_244/latch_enable_in scan_wrapper_339501025136214612_245/latch_enable_in
+ scan_wrapper_339501025136214612_244/scan_select_in scan_wrapper_339501025136214612_245/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_255 scan_wrapper_339501025136214612_255/clk_in scan_wrapper_339501025136214612_256/clk_in
+ scan_wrapper_339501025136214612_255/data_in scan_wrapper_339501025136214612_256/data_in
+ scan_wrapper_339501025136214612_255/latch_enable_in scan_wrapper_339501025136214612_256/latch_enable_in
+ scan_wrapper_339501025136214612_255/scan_select_in scan_wrapper_339501025136214612_256/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_277 scan_wrapper_339501025136214612_277/clk_in scan_wrapper_339501025136214612_278/clk_in
+ scan_wrapper_339501025136214612_277/data_in scan_wrapper_339501025136214612_278/data_in
+ scan_wrapper_339501025136214612_277/latch_enable_in scan_wrapper_339501025136214612_278/latch_enable_in
+ scan_wrapper_339501025136214612_277/scan_select_in scan_wrapper_339501025136214612_278/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_266 scan_wrapper_339501025136214612_266/clk_in scan_wrapper_339501025136214612_267/clk_in
+ scan_wrapper_339501025136214612_266/data_in scan_wrapper_339501025136214612_267/data_in
+ scan_wrapper_339501025136214612_266/latch_enable_in scan_wrapper_339501025136214612_267/latch_enable_in
+ scan_wrapper_339501025136214612_266/scan_select_in scan_wrapper_339501025136214612_267/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_288 scan_wrapper_339501025136214612_288/clk_in scan_wrapper_339501025136214612_289/clk_in
+ scan_wrapper_339501025136214612_288/data_in scan_wrapper_339501025136214612_289/data_in
+ scan_wrapper_339501025136214612_288/latch_enable_in scan_wrapper_339501025136214612_289/latch_enable_in
+ scan_wrapper_339501025136214612_288/scan_select_in scan_wrapper_339501025136214612_289/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_299 scan_wrapper_339501025136214612_299/clk_in scan_wrapper_339501025136214612_300/clk_in
+ scan_wrapper_339501025136214612_299/data_in scan_wrapper_339501025136214612_300/data_in
+ scan_wrapper_339501025136214612_299/latch_enable_in scan_wrapper_339501025136214612_300/latch_enable_in
+ scan_wrapper_339501025136214612_299/scan_select_in scan_wrapper_339501025136214612_300/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341364381657858642_61 scan_wrapper_341364381657858642_61/clk_in scan_wrapper_341279123277087315_62/clk_in
+ scan_wrapper_341364381657858642_61/data_in scan_wrapper_341279123277087315_62/data_in
+ scan_wrapper_341364381657858642_61/latch_enable_in scan_wrapper_341279123277087315_62/latch_enable_in
+ scan_wrapper_341364381657858642_61/scan_select_in scan_wrapper_341279123277087315_62/scan_select_in
+ vccd1 vssd1 scan_wrapper_341364381657858642
Xscan_wrapper_341516949939814994_100 scan_wrapper_341516949939814994_100/clk_in scan_wrapper_341521390605697619_101/clk_in
+ scan_wrapper_341516949939814994_100/data_in scan_wrapper_341521390605697619_101/data_in
+ scan_wrapper_341516949939814994_100/latch_enable_in scan_wrapper_341521390605697619_101/latch_enable_in
+ scan_wrapper_341516949939814994_100/scan_select_in scan_wrapper_341521390605697619_101/scan_select_in
+ vccd1 vssd1 scan_wrapper_341516949939814994
Xscan_wrapper_339501025136214612_459 scan_wrapper_339501025136214612_459/clk_in scan_wrapper_339501025136214612_460/clk_in
+ scan_wrapper_339501025136214612_459/data_in scan_wrapper_339501025136214612_460/data_in
+ scan_wrapper_339501025136214612_459/latch_enable_in scan_wrapper_339501025136214612_460/latch_enable_in
+ scan_wrapper_339501025136214612_459/scan_select_in scan_wrapper_339501025136214612_460/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_448 scan_wrapper_339501025136214612_448/clk_in scan_wrapper_339501025136214612_449/clk_in
+ scan_wrapper_339501025136214612_448/data_in scan_wrapper_339501025136214612_449/data_in
+ scan_wrapper_339501025136214612_448/latch_enable_in scan_wrapper_339501025136214612_449/latch_enable_in
+ scan_wrapper_339501025136214612_448/scan_select_in scan_wrapper_339501025136214612_449/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_426 scan_wrapper_339501025136214612_426/clk_in scan_wrapper_339501025136214612_427/clk_in
+ scan_wrapper_339501025136214612_426/data_in scan_wrapper_339501025136214612_427/data_in
+ scan_wrapper_339501025136214612_426/latch_enable_in scan_wrapper_339501025136214612_427/latch_enable_in
+ scan_wrapper_339501025136214612_426/scan_select_in scan_wrapper_339501025136214612_427/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_437 scan_wrapper_339501025136214612_437/clk_in scan_wrapper_339501025136214612_438/clk_in
+ scan_wrapper_339501025136214612_437/data_in scan_wrapper_339501025136214612_438/data_in
+ scan_wrapper_339501025136214612_437/latch_enable_in scan_wrapper_339501025136214612_438/latch_enable_in
+ scan_wrapper_339501025136214612_437/scan_select_in scan_wrapper_339501025136214612_438/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_415 scan_wrapper_339501025136214612_415/clk_in scan_wrapper_339501025136214612_416/clk_in
+ scan_wrapper_339501025136214612_415/data_in scan_wrapper_339501025136214612_416/data_in
+ scan_wrapper_339501025136214612_415/latch_enable_in scan_wrapper_339501025136214612_416/latch_enable_in
+ scan_wrapper_339501025136214612_415/scan_select_in scan_wrapper_339501025136214612_416/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_404 scan_wrapper_339501025136214612_404/clk_in scan_wrapper_339501025136214612_405/clk_in
+ scan_wrapper_339501025136214612_404/data_in scan_wrapper_339501025136214612_405/data_in
+ scan_wrapper_339501025136214612_404/latch_enable_in scan_wrapper_339501025136214612_405/latch_enable_in
+ scan_wrapper_339501025136214612_404/scan_select_in scan_wrapper_339501025136214612_405/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_201 scan_wrapper_339501025136214612_201/clk_in scan_wrapper_339501025136214612_202/clk_in
+ scan_wrapper_339501025136214612_201/data_in scan_wrapper_339501025136214612_202/data_in
+ scan_wrapper_339501025136214612_201/latch_enable_in scan_wrapper_339501025136214612_202/latch_enable_in
+ scan_wrapper_339501025136214612_201/scan_select_in scan_wrapper_339501025136214612_202/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_212 scan_wrapper_339501025136214612_212/clk_in scan_wrapper_339501025136214612_213/clk_in
+ scan_wrapper_339501025136214612_212/data_in scan_wrapper_339501025136214612_213/data_in
+ scan_wrapper_339501025136214612_212/latch_enable_in scan_wrapper_339501025136214612_213/latch_enable_in
+ scan_wrapper_339501025136214612_212/scan_select_in scan_wrapper_339501025136214612_213/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_234 scan_wrapper_339501025136214612_234/clk_in scan_wrapper_339501025136214612_235/clk_in
+ scan_wrapper_339501025136214612_234/data_in scan_wrapper_339501025136214612_235/data_in
+ scan_wrapper_339501025136214612_234/latch_enable_in scan_wrapper_339501025136214612_235/latch_enable_in
+ scan_wrapper_339501025136214612_234/scan_select_in scan_wrapper_339501025136214612_235/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_223 scan_wrapper_339501025136214612_223/clk_in scan_wrapper_339501025136214612_224/clk_in
+ scan_wrapper_339501025136214612_223/data_in scan_wrapper_339501025136214612_224/data_in
+ scan_wrapper_339501025136214612_223/latch_enable_in scan_wrapper_339501025136214612_224/latch_enable_in
+ scan_wrapper_339501025136214612_223/scan_select_in scan_wrapper_339501025136214612_224/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_245 scan_wrapper_339501025136214612_245/clk_in scan_wrapper_339501025136214612_246/clk_in
+ scan_wrapper_339501025136214612_245/data_in scan_wrapper_339501025136214612_246/data_in
+ scan_wrapper_339501025136214612_245/latch_enable_in scan_wrapper_339501025136214612_246/latch_enable_in
+ scan_wrapper_339501025136214612_245/scan_select_in scan_wrapper_339501025136214612_246/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_256 scan_wrapper_339501025136214612_256/clk_in scan_wrapper_339501025136214612_257/clk_in
+ scan_wrapper_339501025136214612_256/data_in scan_wrapper_339501025136214612_257/data_in
+ scan_wrapper_339501025136214612_256/latch_enable_in scan_wrapper_339501025136214612_257/latch_enable_in
+ scan_wrapper_339501025136214612_256/scan_select_in scan_wrapper_339501025136214612_257/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_267 scan_wrapper_339501025136214612_267/clk_in scan_wrapper_339501025136214612_268/clk_in
+ scan_wrapper_339501025136214612_267/data_in scan_wrapper_339501025136214612_268/data_in
+ scan_wrapper_339501025136214612_267/latch_enable_in scan_wrapper_339501025136214612_268/latch_enable_in
+ scan_wrapper_339501025136214612_267/scan_select_in scan_wrapper_339501025136214612_268/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_278 scan_wrapper_339501025136214612_278/clk_in scan_wrapper_339501025136214612_279/clk_in
+ scan_wrapper_339501025136214612_278/data_in scan_wrapper_339501025136214612_279/data_in
+ scan_wrapper_339501025136214612_278/latch_enable_in scan_wrapper_339501025136214612_279/latch_enable_in
+ scan_wrapper_339501025136214612_278/scan_select_in scan_wrapper_339501025136214612_279/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_289 scan_wrapper_339501025136214612_289/clk_in scan_wrapper_339501025136214612_290/clk_in
+ scan_wrapper_339501025136214612_289/data_in scan_wrapper_339501025136214612_290/data_in
+ scan_wrapper_339501025136214612_289/latch_enable_in scan_wrapper_339501025136214612_290/latch_enable_in
+ scan_wrapper_339501025136214612_289/scan_select_in scan_wrapper_339501025136214612_290/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341710255833481812_95 scan_wrapper_341710255833481812_95/clk_in scan_wrapper_340067262721426004_96/clk_in
+ scan_wrapper_341710255833481812_95/data_in scan_wrapper_340067262721426004_96/data_in
+ scan_wrapper_341710255833481812_95/latch_enable_in scan_wrapper_340067262721426004_96/latch_enable_in
+ scan_wrapper_341710255833481812_95/scan_select_in scan_wrapper_340067262721426004_96/scan_select_in
+ vccd1 vssd1 scan_wrapper_341710255833481812
Xscan_wrapper_341538994733974098_120 scan_wrapper_341538994733974098_120/clk_in scan_wrapper_341557831870186068_121/clk_in
+ scan_wrapper_341538994733974098_120/data_in scan_wrapper_341557831870186068_121/data_in
+ scan_wrapper_341538994733974098_120/latch_enable_in scan_wrapper_341557831870186068_121/latch_enable_in
+ scan_wrapper_341538994733974098_120/scan_select_in scan_wrapper_341557831870186068_121/scan_select_in
+ vccd1 vssd1 scan_wrapper_341538994733974098
Xscan_wrapper_341457971277988435_81 scan_wrapper_341457971277988435_81/clk_in scan_wrapper_341399568412312147_82/clk_in
+ scan_wrapper_341457971277988435_81/data_in scan_wrapper_341399568412312147_82/data_in
+ scan_wrapper_341457971277988435_81/latch_enable_in scan_wrapper_341399568412312147_82/latch_enable_in
+ scan_wrapper_341457971277988435_81/scan_select_in scan_wrapper_341399568412312147_82/scan_select_in
+ vccd1 vssd1 scan_wrapper_341457971277988435
Xscan_wrapper_341161378978988626_14 scan_wrapper_341161378978988626_14/clk_in scan_wrapper_341152580068442706_15/clk_in
+ scan_wrapper_341161378978988626_14/data_in scan_wrapper_341152580068442706_15/data_in
+ scan_wrapper_341161378978988626_14/latch_enable_in scan_wrapper_341152580068442706_15/latch_enable_in
+ scan_wrapper_341161378978988626_14/scan_select_in scan_wrapper_341152580068442706_15/scan_select_in
+ vccd1 vssd1 scan_wrapper_341161378978988626
Xscan_wrapper_339501025136214612_449 scan_wrapper_339501025136214612_449/clk_in scan_wrapper_339501025136214612_450/clk_in
+ scan_wrapper_339501025136214612_449/data_in scan_wrapper_339501025136214612_450/data_in
+ scan_wrapper_339501025136214612_449/latch_enable_in scan_wrapper_339501025136214612_450/latch_enable_in
+ scan_wrapper_339501025136214612_449/scan_select_in scan_wrapper_339501025136214612_450/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_438 scan_wrapper_339501025136214612_438/clk_in scan_wrapper_339501025136214612_439/clk_in
+ scan_wrapper_339501025136214612_438/data_in scan_wrapper_339501025136214612_439/data_in
+ scan_wrapper_339501025136214612_438/latch_enable_in scan_wrapper_339501025136214612_439/latch_enable_in
+ scan_wrapper_339501025136214612_438/scan_select_in scan_wrapper_339501025136214612_439/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_427 scan_wrapper_339501025136214612_427/clk_in scan_wrapper_339501025136214612_428/clk_in
+ scan_wrapper_339501025136214612_427/data_in scan_wrapper_339501025136214612_428/data_in
+ scan_wrapper_339501025136214612_427/latch_enable_in scan_wrapper_339501025136214612_428/latch_enable_in
+ scan_wrapper_339501025136214612_427/scan_select_in scan_wrapper_339501025136214612_428/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_416 scan_wrapper_339501025136214612_416/clk_in scan_wrapper_339501025136214612_417/clk_in
+ scan_wrapper_339501025136214612_416/data_in scan_wrapper_339501025136214612_417/data_in
+ scan_wrapper_339501025136214612_416/latch_enable_in scan_wrapper_339501025136214612_417/latch_enable_in
+ scan_wrapper_339501025136214612_416/scan_select_in scan_wrapper_339501025136214612_417/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_405 scan_wrapper_339501025136214612_405/clk_in scan_wrapper_339501025136214612_406/clk_in
+ scan_wrapper_339501025136214612_405/data_in scan_wrapper_339501025136214612_406/data_in
+ scan_wrapper_339501025136214612_405/latch_enable_in scan_wrapper_339501025136214612_406/latch_enable_in
+ scan_wrapper_339501025136214612_405/scan_select_in scan_wrapper_339501025136214612_406/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341629415144292948_146 scan_wrapper_341629415144292948_146/clk_in scan_wrapper_341637831098106450_147/clk_in
+ scan_wrapper_341629415144292948_146/data_in scan_wrapper_341637831098106450_147/data_in
+ scan_wrapper_341629415144292948_146/latch_enable_in scan_wrapper_341637831098106450_147/latch_enable_in
+ scan_wrapper_341629415144292948_146/scan_select_in scan_wrapper_341637831098106450_147/scan_select_in
+ vccd1 vssd1 scan_wrapper_341629415144292948
Xscan_wrapper_341188777753969234_22 scan_wrapper_341188777753969234_22/clk_in scan_wrapper_341194143598379604_23/clk_in
+ scan_wrapper_341188777753969234_22/data_in scan_wrapper_341194143598379604_23/data_in
+ scan_wrapper_341188777753969234_22/latch_enable_in scan_wrapper_341194143598379604_23/latch_enable_in
+ scan_wrapper_341188777753969234_22/scan_select_in scan_wrapper_341194143598379604_23/scan_select_in
+ vccd1 vssd1 scan_wrapper_341188777753969234
Xscan_wrapper_339501025136214612_202 scan_wrapper_339501025136214612_202/clk_in scan_wrapper_339501025136214612_203/clk_in
+ scan_wrapper_339501025136214612_202/data_in scan_wrapper_339501025136214612_203/data_in
+ scan_wrapper_339501025136214612_202/latch_enable_in scan_wrapper_339501025136214612_203/latch_enable_in
+ scan_wrapper_339501025136214612_202/scan_select_in scan_wrapper_339501025136214612_203/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_213 scan_wrapper_339501025136214612_213/clk_in scan_wrapper_339501025136214612_214/clk_in
+ scan_wrapper_339501025136214612_213/data_in scan_wrapper_339501025136214612_214/data_in
+ scan_wrapper_339501025136214612_213/latch_enable_in scan_wrapper_339501025136214612_214/latch_enable_in
+ scan_wrapper_339501025136214612_213/scan_select_in scan_wrapper_339501025136214612_214/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_235 scan_wrapper_339501025136214612_235/clk_in scan_wrapper_339501025136214612_236/clk_in
+ scan_wrapper_339501025136214612_235/data_in scan_wrapper_339501025136214612_236/data_in
+ scan_wrapper_339501025136214612_235/latch_enable_in scan_wrapper_339501025136214612_236/latch_enable_in
+ scan_wrapper_339501025136214612_235/scan_select_in scan_wrapper_339501025136214612_236/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_224 scan_wrapper_339501025136214612_224/clk_in scan_wrapper_339501025136214612_225/clk_in
+ scan_wrapper_339501025136214612_224/data_in scan_wrapper_339501025136214612_225/data_in
+ scan_wrapper_339501025136214612_224/latch_enable_in scan_wrapper_339501025136214612_225/latch_enable_in
+ scan_wrapper_339501025136214612_224/scan_select_in scan_wrapper_339501025136214612_225/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_246 scan_wrapper_339501025136214612_246/clk_in scan_wrapper_339501025136214612_247/clk_in
+ scan_wrapper_339501025136214612_246/data_in scan_wrapper_339501025136214612_247/data_in
+ scan_wrapper_339501025136214612_246/latch_enable_in scan_wrapper_339501025136214612_247/latch_enable_in
+ scan_wrapper_339501025136214612_246/scan_select_in scan_wrapper_339501025136214612_247/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_257 scan_wrapper_339501025136214612_257/clk_in scan_wrapper_339501025136214612_258/clk_in
+ scan_wrapper_339501025136214612_257/data_in scan_wrapper_339501025136214612_258/data_in
+ scan_wrapper_339501025136214612_257/latch_enable_in scan_wrapper_339501025136214612_258/latch_enable_in
+ scan_wrapper_339501025136214612_257/scan_select_in scan_wrapper_339501025136214612_258/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_268 scan_wrapper_339501025136214612_268/clk_in scan_wrapper_339501025136214612_269/clk_in
+ scan_wrapper_339501025136214612_268/data_in scan_wrapper_339501025136214612_269/data_in
+ scan_wrapper_339501025136214612_268/latch_enable_in scan_wrapper_339501025136214612_269/latch_enable_in
+ scan_wrapper_339501025136214612_268/scan_select_in scan_wrapper_339501025136214612_269/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_279 scan_wrapper_339501025136214612_279/clk_in scan_wrapper_339501025136214612_280/clk_in
+ scan_wrapper_339501025136214612_279/data_in scan_wrapper_339501025136214612_280/data_in
+ scan_wrapper_339501025136214612_279/latch_enable_in scan_wrapper_339501025136214612_280/latch_enable_in
+ scan_wrapper_339501025136214612_279/scan_select_in scan_wrapper_339501025136214612_280/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341496918381167187_74 scan_wrapper_341496918381167187_74/clk_in scan_wrapper_341440781874102868_75/clk_in
+ scan_wrapper_341496918381167187_74/data_in scan_wrapper_341440781874102868_75/data_in
+ scan_wrapper_341496918381167187_74/latch_enable_in scan_wrapper_341440781874102868_75/latch_enable_in
+ scan_wrapper_341496918381167187_74/scan_select_in scan_wrapper_341440781874102868_75/scan_select_in
+ vccd1 vssd1 scan_wrapper_341496918381167187
Xscan_wrapper_341717091617866324_111 scan_wrapper_341717091617866324_111/clk_in scan_wrapper_hamming74_112/clk_in
+ scan_wrapper_341717091617866324_111/data_in scan_wrapper_hamming74_112/data_in scan_wrapper_341717091617866324_111/latch_enable_in
+ scan_wrapper_hamming74_112/latch_enable_in scan_wrapper_341717091617866324_111/scan_select_in
+ scan_wrapper_hamming74_112/scan_select_in vccd1 vssd1 scan_wrapper_341717091617866324
Xscan_wrapper_339501025136214612_439 scan_wrapper_339501025136214612_439/clk_in scan_wrapper_339501025136214612_440/clk_in
+ scan_wrapper_339501025136214612_439/data_in scan_wrapper_339501025136214612_440/data_in
+ scan_wrapper_339501025136214612_439/latch_enable_in scan_wrapper_339501025136214612_440/latch_enable_in
+ scan_wrapper_339501025136214612_439/scan_select_in scan_wrapper_339501025136214612_440/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_428 scan_wrapper_339501025136214612_428/clk_in scan_wrapper_339501025136214612_429/clk_in
+ scan_wrapper_339501025136214612_428/data_in scan_wrapper_339501025136214612_429/data_in
+ scan_wrapper_339501025136214612_428/latch_enable_in scan_wrapper_339501025136214612_429/latch_enable_in
+ scan_wrapper_339501025136214612_428/scan_select_in scan_wrapper_339501025136214612_429/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_417 scan_wrapper_339501025136214612_417/clk_in scan_wrapper_339501025136214612_418/clk_in
+ scan_wrapper_339501025136214612_417/data_in scan_wrapper_339501025136214612_418/data_in
+ scan_wrapper_339501025136214612_417/latch_enable_in scan_wrapper_339501025136214612_418/latch_enable_in
+ scan_wrapper_339501025136214612_417/scan_select_in scan_wrapper_339501025136214612_418/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_406 scan_wrapper_339501025136214612_406/clk_in scan_wrapper_339501025136214612_407/clk_in
+ scan_wrapper_339501025136214612_406/data_in scan_wrapper_339501025136214612_407/data_in
+ scan_wrapper_339501025136214612_406/latch_enable_in scan_wrapper_339501025136214612_407/latch_enable_in
+ scan_wrapper_339501025136214612_406/scan_select_in scan_wrapper_339501025136214612_407/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341589685194195540_129 scan_wrapper_341589685194195540_129/clk_in scan_wrapper_341608574336631379_130/clk_in
+ scan_wrapper_341589685194195540_129/data_in scan_wrapper_341608574336631379_130/data_in
+ scan_wrapper_341589685194195540_129/latch_enable_in scan_wrapper_341608574336631379_130/latch_enable_in
+ scan_wrapper_341589685194195540_129/scan_select_in scan_wrapper_341608574336631379_130/scan_select_in
+ vccd1 vssd1 scan_wrapper_341589685194195540
Xscan_wrapper_339501025136214612_203 scan_wrapper_339501025136214612_203/clk_in scan_wrapper_339501025136214612_204/clk_in
+ scan_wrapper_339501025136214612_203/data_in scan_wrapper_339501025136214612_204/data_in
+ scan_wrapper_339501025136214612_203/latch_enable_in scan_wrapper_339501025136214612_204/latch_enable_in
+ scan_wrapper_339501025136214612_203/scan_select_in scan_wrapper_339501025136214612_204/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_214 scan_wrapper_339501025136214612_214/clk_in scan_wrapper_339501025136214612_215/clk_in
+ scan_wrapper_339501025136214612_214/data_in scan_wrapper_339501025136214612_215/data_in
+ scan_wrapper_339501025136214612_214/latch_enable_in scan_wrapper_339501025136214612_215/latch_enable_in
+ scan_wrapper_339501025136214612_214/scan_select_in scan_wrapper_339501025136214612_215/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_236 scan_wrapper_339501025136214612_236/clk_in scan_wrapper_339501025136214612_237/clk_in
+ scan_wrapper_339501025136214612_236/data_in scan_wrapper_339501025136214612_237/data_in
+ scan_wrapper_339501025136214612_236/latch_enable_in scan_wrapper_339501025136214612_237/latch_enable_in
+ scan_wrapper_339501025136214612_236/scan_select_in scan_wrapper_339501025136214612_237/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_225 scan_wrapper_339501025136214612_225/clk_in scan_wrapper_339501025136214612_226/clk_in
+ scan_wrapper_339501025136214612_225/data_in scan_wrapper_339501025136214612_226/data_in
+ scan_wrapper_339501025136214612_225/latch_enable_in scan_wrapper_339501025136214612_226/latch_enable_in
+ scan_wrapper_339501025136214612_225/scan_select_in scan_wrapper_339501025136214612_226/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_247 scan_wrapper_339501025136214612_247/clk_in scan_wrapper_339501025136214612_248/clk_in
+ scan_wrapper_339501025136214612_247/data_in scan_wrapper_339501025136214612_248/data_in
+ scan_wrapper_339501025136214612_247/latch_enable_in scan_wrapper_339501025136214612_248/latch_enable_in
+ scan_wrapper_339501025136214612_247/scan_select_in scan_wrapper_339501025136214612_248/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_269 scan_wrapper_339501025136214612_269/clk_in scan_wrapper_339501025136214612_270/clk_in
+ scan_wrapper_339501025136214612_269/data_in scan_wrapper_339501025136214612_270/data_in
+ scan_wrapper_339501025136214612_269/latch_enable_in scan_wrapper_339501025136214612_270/latch_enable_in
+ scan_wrapper_339501025136214612_269/scan_select_in scan_wrapper_339501025136214612_270/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_258 scan_wrapper_339501025136214612_258/clk_in scan_wrapper_339501025136214612_259/clk_in
+ scan_wrapper_339501025136214612_258/data_in scan_wrapper_339501025136214612_259/data_in
+ scan_wrapper_339501025136214612_258/latch_enable_in scan_wrapper_339501025136214612_259/latch_enable_in
+ scan_wrapper_339501025136214612_258/scan_select_in scan_wrapper_339501025136214612_259/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341202178192441940_26 scan_wrapper_341202178192441940_26/clk_in scan_wrapper_341191836498395731_27/clk_in
+ scan_wrapper_341202178192441940_26/data_in scan_wrapper_341191836498395731_27/data_in
+ scan_wrapper_341202178192441940_26/latch_enable_in scan_wrapper_341191836498395731_27/latch_enable_in
+ scan_wrapper_341202178192441940_26/scan_select_in scan_wrapper_341191836498395731_27/scan_select_in
+ vccd1 vssd1 scan_wrapper_341202178192441940
Xscan_wrapper_341337976625693266_49 scan_wrapper_341337976625693266_49/clk_in scan_wrapper_341339883600609876_50/clk_in
+ scan_wrapper_341337976625693266_49/data_in scan_wrapper_341339883600609876_50/data_in
+ scan_wrapper_341337976625693266_49/latch_enable_in scan_wrapper_341339883600609876_50/latch_enable_in
+ scan_wrapper_341337976625693266_49/scan_select_in scan_wrapper_341339883600609876_50/scan_select_in
+ vccd1 vssd1 scan_wrapper_341337976625693266
Xscan_wrapper_339501025136214612_418 scan_wrapper_339501025136214612_418/clk_in scan_wrapper_339501025136214612_419/clk_in
+ scan_wrapper_339501025136214612_418/data_in scan_wrapper_339501025136214612_419/data_in
+ scan_wrapper_339501025136214612_418/latch_enable_in scan_wrapper_339501025136214612_419/latch_enable_in
+ scan_wrapper_339501025136214612_418/scan_select_in scan_wrapper_339501025136214612_419/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_429 scan_wrapper_339501025136214612_429/clk_in scan_wrapper_339501025136214612_430/clk_in
+ scan_wrapper_339501025136214612_429/data_in scan_wrapper_339501025136214612_430/data_in
+ scan_wrapper_339501025136214612_429/latch_enable_in scan_wrapper_339501025136214612_430/latch_enable_in
+ scan_wrapper_339501025136214612_429/scan_select_in scan_wrapper_339501025136214612_430/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_407 scan_wrapper_339501025136214612_407/clk_in scan_wrapper_339501025136214612_408/clk_in
+ scan_wrapper_339501025136214612_407/data_in scan_wrapper_339501025136214612_408/data_in
+ scan_wrapper_339501025136214612_407/latch_enable_in scan_wrapper_339501025136214612_408/latch_enable_in
+ scan_wrapper_339501025136214612_407/scan_select_in scan_wrapper_339501025136214612_408/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341476989274686036_84 scan_wrapper_341476989274686036_84/clk_in scan_wrapper_341482086419399252_85/clk_in
+ scan_wrapper_341476989274686036_84/data_in scan_wrapper_341482086419399252_85/data_in
+ scan_wrapper_341476989274686036_84/latch_enable_in scan_wrapper_341482086419399252_85/latch_enable_in
+ scan_wrapper_341476989274686036_84/scan_select_in scan_wrapper_341482086419399252_85/scan_select_in
+ vccd1 vssd1 scan_wrapper_341476989274686036
Xscan_wrapper_339800239192932947_7 scan_wrapper_339800239192932947_7/clk_in scan_wrapper_341154161238213203_8/clk_in
+ scan_wrapper_339800239192932947_7/data_in scan_wrapper_341154161238213203_8/data_in
+ scan_wrapper_339800239192932947_7/latch_enable_in scan_wrapper_341154161238213203_8/latch_enable_in
+ scan_wrapper_339800239192932947_7/scan_select_in scan_wrapper_341154161238213203_8/scan_select_in
+ vccd1 vssd1 scan_wrapper_339800239192932947
Xscan_wrapper_340285391309374034_4 scan_wrapper_340285391309374034_4/clk_in scan_wrapper_340661930553246290_5/clk_in
+ scan_wrapper_340285391309374034_4/data_in scan_wrapper_340661930553246290_5/data_in
+ scan_wrapper_340285391309374034_4/latch_enable_in scan_wrapper_340661930553246290_5/latch_enable_in
+ scan_wrapper_340285391309374034_4/scan_select_in scan_wrapper_340661930553246290_5/scan_select_in
+ vccd1 vssd1 scan_wrapper_340285391309374034
Xscan_wrapper_339688086163161683_1 scan_wrapper_339688086163161683_1/clk_in scan_wrapper_340218629792465491_2/clk_in
+ scan_wrapper_339688086163161683_1/data_in scan_wrapper_340218629792465491_2/data_in
+ scan_wrapper_339688086163161683_1/latch_enable_in scan_wrapper_340218629792465491_2/latch_enable_in
+ scan_wrapper_339688086163161683_1/scan_select_in scan_wrapper_340218629792465491_2/scan_select_in
+ vccd1 vssd1 scan_wrapper_339688086163161683
Xscan_wrapper_339501025136214612_204 scan_wrapper_339501025136214612_204/clk_in scan_wrapper_339501025136214612_205/clk_in
+ scan_wrapper_339501025136214612_204/data_in scan_wrapper_339501025136214612_205/data_in
+ scan_wrapper_339501025136214612_204/latch_enable_in scan_wrapper_339501025136214612_205/latch_enable_in
+ scan_wrapper_339501025136214612_204/scan_select_in scan_wrapper_339501025136214612_205/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_215 scan_wrapper_339501025136214612_215/clk_in scan_wrapper_339501025136214612_216/clk_in
+ scan_wrapper_339501025136214612_215/data_in scan_wrapper_339501025136214612_216/data_in
+ scan_wrapper_339501025136214612_215/latch_enable_in scan_wrapper_339501025136214612_216/latch_enable_in
+ scan_wrapper_339501025136214612_215/scan_select_in scan_wrapper_339501025136214612_216/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_237 scan_wrapper_339501025136214612_237/clk_in scan_wrapper_339501025136214612_238/clk_in
+ scan_wrapper_339501025136214612_237/data_in scan_wrapper_339501025136214612_238/data_in
+ scan_wrapper_339501025136214612_237/latch_enable_in scan_wrapper_339501025136214612_238/latch_enable_in
+ scan_wrapper_339501025136214612_237/scan_select_in scan_wrapper_339501025136214612_238/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_226 scan_wrapper_339501025136214612_226/clk_in scan_wrapper_339501025136214612_227/clk_in
+ scan_wrapper_339501025136214612_226/data_in scan_wrapper_339501025136214612_227/data_in
+ scan_wrapper_339501025136214612_226/latch_enable_in scan_wrapper_339501025136214612_227/latch_enable_in
+ scan_wrapper_339501025136214612_226/scan_select_in scan_wrapper_339501025136214612_227/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_248 scan_wrapper_339501025136214612_248/clk_in scan_wrapper_339501025136214612_249/clk_in
+ scan_wrapper_339501025136214612_248/data_in scan_wrapper_339501025136214612_249/data_in
+ scan_wrapper_339501025136214612_248/latch_enable_in scan_wrapper_339501025136214612_249/latch_enable_in
+ scan_wrapper_339501025136214612_248/scan_select_in scan_wrapper_339501025136214612_249/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_259 scan_wrapper_339501025136214612_259/clk_in scan_wrapper_339501025136214612_260/clk_in
+ scan_wrapper_339501025136214612_259/data_in scan_wrapper_339501025136214612_260/data_in
+ scan_wrapper_339501025136214612_259/latch_enable_in scan_wrapper_339501025136214612_260/latch_enable_in
+ scan_wrapper_339501025136214612_259/scan_select_in scan_wrapper_339501025136214612_260/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341154161238213203_8 scan_wrapper_341154161238213203_8/clk_in scan_wrapper_341159915403870803_9/clk_in
+ scan_wrapper_341154161238213203_8/data_in scan_wrapper_341159915403870803_9/data_in
+ scan_wrapper_341154161238213203_8/latch_enable_in scan_wrapper_341159915403870803_9/latch_enable_in
+ scan_wrapper_341154161238213203_8/scan_select_in scan_wrapper_341159915403870803_9/scan_select_in
+ vccd1 vssd1 scan_wrapper_341154161238213203
Xscan_wrapper_339501025136214612_419 scan_wrapper_339501025136214612_419/clk_in scan_wrapper_339501025136214612_420/clk_in
+ scan_wrapper_339501025136214612_419/data_in scan_wrapper_339501025136214612_420/data_in
+ scan_wrapper_339501025136214612_419/latch_enable_in scan_wrapper_339501025136214612_420/latch_enable_in
+ scan_wrapper_339501025136214612_419/scan_select_in scan_wrapper_339501025136214612_420/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_408 scan_wrapper_339501025136214612_408/clk_in scan_wrapper_339501025136214612_409/clk_in
+ scan_wrapper_339501025136214612_408/data_in scan_wrapper_339501025136214612_409/data_in
+ scan_wrapper_339501025136214612_408/latch_enable_in scan_wrapper_339501025136214612_409/latch_enable_in
+ scan_wrapper_339501025136214612_408/scan_select_in scan_wrapper_339501025136214612_409/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341160271679586899_13 scan_wrapper_341160271679586899_13/clk_in scan_wrapper_341161378978988626_14/clk_in
+ scan_wrapper_341160271679586899_13/data_in scan_wrapper_341161378978988626_14/data_in
+ scan_wrapper_341160271679586899_13/latch_enable_in scan_wrapper_341161378978988626_14/latch_enable_in
+ scan_wrapper_341160271679586899_13/scan_select_in scan_wrapper_341161378978988626_14/scan_select_in
+ vccd1 vssd1 scan_wrapper_341160271679586899
Xscan_wrapper_339501025136214612_205 scan_wrapper_339501025136214612_205/clk_in scan_wrapper_339501025136214612_206/clk_in
+ scan_wrapper_339501025136214612_205/data_in scan_wrapper_339501025136214612_206/data_in
+ scan_wrapper_339501025136214612_205/latch_enable_in scan_wrapper_339501025136214612_206/latch_enable_in
+ scan_wrapper_339501025136214612_205/scan_select_in scan_wrapper_339501025136214612_206/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_216 scan_wrapper_339501025136214612_216/clk_in scan_wrapper_339501025136214612_217/clk_in
+ scan_wrapper_339501025136214612_216/data_in scan_wrapper_339501025136214612_217/data_in
+ scan_wrapper_339501025136214612_216/latch_enable_in scan_wrapper_339501025136214612_217/latch_enable_in
+ scan_wrapper_339501025136214612_216/scan_select_in scan_wrapper_339501025136214612_217/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_227 scan_wrapper_339501025136214612_227/clk_in scan_wrapper_339501025136214612_228/clk_in
+ scan_wrapper_339501025136214612_227/data_in scan_wrapper_339501025136214612_228/data_in
+ scan_wrapper_339501025136214612_227/latch_enable_in scan_wrapper_339501025136214612_228/latch_enable_in
+ scan_wrapper_339501025136214612_227/scan_select_in scan_wrapper_339501025136214612_228/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_238 scan_wrapper_339501025136214612_238/clk_in scan_wrapper_339501025136214612_239/clk_in
+ scan_wrapper_339501025136214612_238/data_in scan_wrapper_339501025136214612_239/data_in
+ scan_wrapper_339501025136214612_238/latch_enable_in scan_wrapper_339501025136214612_239/latch_enable_in
+ scan_wrapper_339501025136214612_238/scan_select_in scan_wrapper_339501025136214612_239/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_249 scan_wrapper_339501025136214612_249/clk_in scan_wrapper_339501025136214612_250/clk_in
+ scan_wrapper_339501025136214612_249/data_in scan_wrapper_339501025136214612_250/data_in
+ scan_wrapper_339501025136214612_249/latch_enable_in scan_wrapper_339501025136214612_250/latch_enable_in
+ scan_wrapper_339501025136214612_249/scan_select_in scan_wrapper_339501025136214612_250/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341194143598379604_23 scan_wrapper_341194143598379604_23/clk_in scan_wrapper_341205508016833108_24/clk_in
+ scan_wrapper_341194143598379604_23/data_in scan_wrapper_341205508016833108_24/data_in
+ scan_wrapper_341194143598379604_23/latch_enable_in scan_wrapper_341205508016833108_24/latch_enable_in
+ scan_wrapper_341194143598379604_23/scan_select_in scan_wrapper_341205508016833108_24/scan_select_in
+ vccd1 vssd1 scan_wrapper_341194143598379604
Xscan_wrapper_341573751072096850_123 scan_wrapper_341573751072096850_123/clk_in scan_wrapper_341571228858843732_124/clk_in
+ scan_wrapper_341573751072096850_123/data_in scan_wrapper_341571228858843732_124/data_in
+ scan_wrapper_341573751072096850_123/latch_enable_in scan_wrapper_341571228858843732_124/latch_enable_in
+ scan_wrapper_341573751072096850_123/scan_select_in scan_wrapper_341571228858843732_124/scan_select_in
+ vccd1 vssd1 scan_wrapper_341573751072096850
Xscan_wrapper_341450853309219412_78 scan_wrapper_341450853309219412_78/clk_in scan_wrapper_341438392303616596_79/clk_in
+ scan_wrapper_341450853309219412_78/data_in scan_wrapper_341438392303616596_79/data_in
+ scan_wrapper_341450853309219412_78/latch_enable_in scan_wrapper_341438392303616596_79/latch_enable_in
+ scan_wrapper_341450853309219412_78/scan_select_in scan_wrapper_341438392303616596_79/scan_select_in
+ vccd1 vssd1 scan_wrapper_341450853309219412
Xscan_wrapper_339501025136214612_409 scan_wrapper_339501025136214612_409/clk_in scan_wrapper_339501025136214612_410/clk_in
+ scan_wrapper_339501025136214612_409/data_in scan_wrapper_339501025136214612_410/data_in
+ scan_wrapper_339501025136214612_409/latch_enable_in scan_wrapper_339501025136214612_410/latch_enable_in
+ scan_wrapper_339501025136214612_409/scan_select_in scan_wrapper_339501025136214612_410/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341542971476279892_117 scan_wrapper_341542971476279892_117/clk_in scan_wrapper_341556236196512338_118/clk_in
+ scan_wrapper_341542971476279892_117/data_in scan_wrapper_341556236196512338_118/data_in
+ scan_wrapper_341542971476279892_117/latch_enable_in scan_wrapper_341556236196512338_118/latch_enable_in
+ scan_wrapper_341542971476279892_117/scan_select_in scan_wrapper_341556236196512338_118/scan_select_in
+ vccd1 vssd1 scan_wrapper_341542971476279892
Xscan_wrapper_341519170869920338_103 scan_wrapper_341519170869920338_103/clk_in scan_wrapper_341446083683025490_104/clk_in
+ scan_wrapper_341519170869920338_103/data_in scan_wrapper_341446083683025490_104/data_in
+ scan_wrapper_341519170869920338_103/latch_enable_in scan_wrapper_341446083683025490_104/latch_enable_in
+ scan_wrapper_341519170869920338_103/scan_select_in scan_wrapper_341446083683025490_104/scan_select_in
+ vccd1 vssd1 scan_wrapper_341519170869920338
Xscan_wrapper_341240110454407762_36 scan_wrapper_341240110454407762_36/clk_in scan_wrapper_341264068701586004_37/clk_in
+ scan_wrapper_341240110454407762_36/data_in scan_wrapper_341264068701586004_37/data_in
+ scan_wrapper_341240110454407762_36/latch_enable_in scan_wrapper_341264068701586004_37/latch_enable_in
+ scan_wrapper_341240110454407762_36/scan_select_in scan_wrapper_341264068701586004_37/scan_select_in
+ vccd1 vssd1 scan_wrapper_341240110454407762
Xscan_wrapper_340318610245288530_3 scan_wrapper_340318610245288530_3/clk_in scan_wrapper_340285391309374034_4/clk_in
+ scan_wrapper_340318610245288530_3/data_in scan_wrapper_340285391309374034_4/data_in
+ scan_wrapper_340318610245288530_3/latch_enable_in scan_wrapper_340285391309374034_4/latch_enable_in
+ scan_wrapper_340318610245288530_3/scan_select_in scan_wrapper_340285391309374034_4/scan_select_in
+ vccd1 vssd1 scan_wrapper_340318610245288530
Xscan_wrapper_339501025136214612_206 scan_wrapper_339501025136214612_206/clk_in scan_wrapper_339501025136214612_207/clk_in
+ scan_wrapper_339501025136214612_206/data_in scan_wrapper_339501025136214612_207/data_in
+ scan_wrapper_339501025136214612_206/latch_enable_in scan_wrapper_339501025136214612_207/latch_enable_in
+ scan_wrapper_339501025136214612_206/scan_select_in scan_wrapper_339501025136214612_207/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_217 scan_wrapper_339501025136214612_217/clk_in scan_wrapper_339501025136214612_218/clk_in
+ scan_wrapper_339501025136214612_217/data_in scan_wrapper_339501025136214612_218/data_in
+ scan_wrapper_339501025136214612_217/latch_enable_in scan_wrapper_339501025136214612_218/latch_enable_in
+ scan_wrapper_339501025136214612_217/scan_select_in scan_wrapper_339501025136214612_218/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_228 scan_wrapper_339501025136214612_228/clk_in scan_wrapper_339501025136214612_229/clk_in
+ scan_wrapper_339501025136214612_228/data_in scan_wrapper_339501025136214612_229/data_in
+ scan_wrapper_339501025136214612_228/latch_enable_in scan_wrapper_339501025136214612_229/latch_enable_in
+ scan_wrapper_339501025136214612_228/scan_select_in scan_wrapper_339501025136214612_229/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_239 scan_wrapper_339501025136214612_239/clk_in scan_wrapper_339501025136214612_240/clk_in
+ scan_wrapper_339501025136214612_239/data_in scan_wrapper_339501025136214612_240/data_in
+ scan_wrapper_339501025136214612_239/latch_enable_in scan_wrapper_339501025136214612_240/latch_enable_in
+ scan_wrapper_339501025136214612_239/scan_select_in scan_wrapper_339501025136214612_240/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341556236196512338_118 scan_wrapper_341556236196512338_118/clk_in scan_wrapper_341558189536313940_119/clk_in
+ scan_wrapper_341556236196512338_118/data_in scan_wrapper_341558189536313940_119/data_in
+ scan_wrapper_341556236196512338_118/latch_enable_in scan_wrapper_341558189536313940_119/latch_enable_in
+ scan_wrapper_341556236196512338_118/scan_select_in scan_wrapper_341558189536313940_119/scan_select_in
+ vccd1 vssd1 scan_wrapper_341556236196512338
Xscan_wrapper_339501025136214612_207 scan_wrapper_339501025136214612_207/clk_in scan_wrapper_339501025136214612_208/clk_in
+ scan_wrapper_339501025136214612_207/data_in scan_wrapper_339501025136214612_208/data_in
+ scan_wrapper_339501025136214612_207/latch_enable_in scan_wrapper_339501025136214612_208/latch_enable_in
+ scan_wrapper_339501025136214612_207/scan_select_in scan_wrapper_339501025136214612_208/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_229 scan_wrapper_339501025136214612_229/clk_in scan_wrapper_339501025136214612_230/clk_in
+ scan_wrapper_339501025136214612_229/data_in scan_wrapper_339501025136214612_230/data_in
+ scan_wrapper_339501025136214612_229/latch_enable_in scan_wrapper_339501025136214612_230/latch_enable_in
+ scan_wrapper_339501025136214612_229/scan_select_in scan_wrapper_339501025136214612_230/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_218 scan_wrapper_339501025136214612_218/clk_in scan_wrapper_339501025136214612_219/clk_in
+ scan_wrapper_339501025136214612_218/data_in scan_wrapper_339501025136214612_219/data_in
+ scan_wrapper_339501025136214612_218/latch_enable_in scan_wrapper_339501025136214612_219/latch_enable_in
+ scan_wrapper_339501025136214612_218/scan_select_in scan_wrapper_339501025136214612_219/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341389786199622227_65 scan_wrapper_341389786199622227_65/clk_in scan_wrapper_341404507891040852_66/clk_in
+ scan_wrapper_341389786199622227_65/data_in scan_wrapper_341404507891040852_66/data_in
+ scan_wrapper_341389786199622227_65/latch_enable_in scan_wrapper_341404507891040852_66/latch_enable_in
+ scan_wrapper_341389786199622227_65/scan_select_in scan_wrapper_341404507891040852_66/scan_select_in
+ vccd1 vssd1 scan_wrapper_341389786199622227
Xscan_wrapper_339501025136214612_390 scan_wrapper_339501025136214612_390/clk_in scan_wrapper_339501025136214612_391/clk_in
+ scan_wrapper_339501025136214612_390/data_in scan_wrapper_339501025136214612_391/data_in
+ scan_wrapper_339501025136214612_390/latch_enable_in scan_wrapper_339501025136214612_391/latch_enable_in
+ scan_wrapper_339501025136214612_390/scan_select_in scan_wrapper_339501025136214612_391/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341162950004834900_25 scan_wrapper_341162950004834900_25/clk_in scan_wrapper_341202178192441940_26/clk_in
+ scan_wrapper_341162950004834900_25/data_in scan_wrapper_341202178192441940_26/data_in
+ scan_wrapper_341162950004834900_25/latch_enable_in scan_wrapper_341202178192441940_26/latch_enable_in
+ scan_wrapper_341162950004834900_25/scan_select_in scan_wrapper_341202178192441940_26/scan_select_in
+ vccd1 vssd1 scan_wrapper_341162950004834900
Xscan_wrapper_bc4d7220e4fdbf20a574d56ea112a8e1_42 scan_wrapper_341271902949474898_41/clk_out
+ scan_wrapper_341178296293130834_43/clk_in scan_wrapper_341271902949474898_41/data_out
+ scan_wrapper_341178296293130834_43/data_in scan_wrapper_341271902949474898_41/latch_enable_out
+ scan_wrapper_341178296293130834_43/latch_enable_in scan_wrapper_341271902949474898_41/scan_select_out
+ scan_wrapper_341178296293130834_43/scan_select_in vccd1 vssd1 scan_wrapper_bc4d7220e4fdbf20a574d56ea112a8e1
Xscan_wrapper_341382703379120723_64 scan_wrapper_341382703379120723_64/clk_in scan_wrapper_341389786199622227_65/clk_in
+ scan_wrapper_341382703379120723_64/data_in scan_wrapper_341389786199622227_65/data_in
+ scan_wrapper_341382703379120723_64/latch_enable_in scan_wrapper_341389786199622227_65/latch_enable_in
+ scan_wrapper_341382703379120723_64/scan_select_in scan_wrapper_341389786199622227_65/scan_select_in
+ vccd1 vssd1 scan_wrapper_341382703379120723
Xscan_wrapper_341167691532337747_17 scan_wrapper_341167691532337747_17/clk_in scan_wrapper_341178154799333971_18/clk_in
+ scan_wrapper_341167691532337747_17/data_in scan_wrapper_341178154799333971_18/data_in
+ scan_wrapper_341167691532337747_17/latch_enable_in scan_wrapper_341178154799333971_18/latch_enable_in
+ scan_wrapper_341167691532337747_17/scan_select_in scan_wrapper_341178154799333971_18/scan_select_in
+ vccd1 vssd1 scan_wrapper_341167691532337747
Xscan_wrapper_339501025136214612_208 scan_wrapper_339501025136214612_208/clk_in scan_wrapper_339501025136214612_209/clk_in
+ scan_wrapper_339501025136214612_208/data_in scan_wrapper_339501025136214612_209/data_in
+ scan_wrapper_339501025136214612_208/latch_enable_in scan_wrapper_339501025136214612_209/latch_enable_in
+ scan_wrapper_339501025136214612_208/scan_select_in scan_wrapper_339501025136214612_209/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_219 scan_wrapper_339501025136214612_219/clk_in scan_wrapper_339501025136214612_220/clk_in
+ scan_wrapper_339501025136214612_219/data_in scan_wrapper_339501025136214612_220/data_in
+ scan_wrapper_339501025136214612_219/latch_enable_in scan_wrapper_339501025136214612_220/latch_enable_in
+ scan_wrapper_339501025136214612_219/scan_select_in scan_wrapper_339501025136214612_220/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341192621088047698_29 scan_wrapper_341192621088047698_29/clk_in scan_wrapper_340579111348994642_30/clk_in
+ scan_wrapper_341192621088047698_29/data_in scan_wrapper_340579111348994642_30/data_in
+ scan_wrapper_341192621088047698_29/latch_enable_in scan_wrapper_340579111348994642_30/latch_enable_in
+ scan_wrapper_341192621088047698_29/scan_select_in scan_wrapper_340579111348994642_30/scan_select_in
+ vccd1 vssd1 scan_wrapper_341192621088047698
Xscan_wrapper_339501025136214612_380 scan_wrapper_339501025136214612_380/clk_in scan_wrapper_339501025136214612_381/clk_in
+ scan_wrapper_339501025136214612_380/data_in scan_wrapper_339501025136214612_381/data_in
+ scan_wrapper_339501025136214612_380/latch_enable_in scan_wrapper_339501025136214612_381/latch_enable_in
+ scan_wrapper_339501025136214612_380/scan_select_in scan_wrapper_339501025136214612_381/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_391 scan_wrapper_339501025136214612_391/clk_in scan_wrapper_339501025136214612_392/clk_in
+ scan_wrapper_339501025136214612_391/data_in scan_wrapper_339501025136214612_392/data_in
+ scan_wrapper_339501025136214612_391/latch_enable_in scan_wrapper_339501025136214612_392/latch_enable_in
+ scan_wrapper_339501025136214612_391/scan_select_in scan_wrapper_339501025136214612_392/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341431502448362067_107 scan_wrapper_341431502448362067_107/clk_in scan_wrapper_341473139924927058_108/clk_in
+ scan_wrapper_341431502448362067_107/data_in scan_wrapper_341473139924927058_108/data_in
+ scan_wrapper_341431502448362067_107/latch_enable_in scan_wrapper_341473139924927058_108/latch_enable_in
+ scan_wrapper_341431502448362067_107/scan_select_in scan_wrapper_341473139924927058_108/scan_select_in
+ vccd1 vssd1 scan_wrapper_341431502448362067
Xscan_wrapper_341444501414347346_76 scan_wrapper_341444501414347346_76/clk_in scan_wrapper_019235602376235615_77/clk_in
+ scan_wrapper_341444501414347346_76/data_in scan_wrapper_019235602376235615_77/data_in
+ scan_wrapper_341444501414347346_76/latch_enable_in scan_wrapper_019235602376235615_77/latch_enable_in
+ scan_wrapper_341444501414347346_76/scan_select_in scan_wrapper_019235602376235615_77/scan_select_in
+ vccd1 vssd1 scan_wrapper_341444501414347346
Xscan_wrapper_341520747710120530_98 scan_wrapper_341520747710120530_98/clk_in scan_wrapper_341423712597181012_99/clk_in
+ scan_wrapper_341520747710120530_98/data_in scan_wrapper_341423712597181012_99/data_in
+ scan_wrapper_341520747710120530_98/latch_enable_in scan_wrapper_341423712597181012_99/latch_enable_in
+ scan_wrapper_341520747710120530_98/scan_select_in scan_wrapper_341423712597181012_99/scan_select_in
+ vccd1 vssd1 scan_wrapper_341520747710120530
Xscan_wrapper_341296149788885588_47 scan_wrapper_341296149788885588_47/clk_in scan_wrapper_341332847867462227_48/clk_in
+ scan_wrapper_341296149788885588_47/data_in scan_wrapper_341332847867462227_48/data_in
+ scan_wrapper_341296149788885588_47/latch_enable_in scan_wrapper_341332847867462227_48/latch_enable_in
+ scan_wrapper_341296149788885588_47/scan_select_in scan_wrapper_341332847867462227_48/scan_select_in
+ vccd1 vssd1 scan_wrapper_341296149788885588
Xscan_wrapper_339501025136214612_209 scan_wrapper_339501025136214612_209/clk_in scan_wrapper_339501025136214612_210/clk_in
+ scan_wrapper_339501025136214612_209/data_in scan_wrapper_339501025136214612_210/data_in
+ scan_wrapper_339501025136214612_209/latch_enable_in scan_wrapper_339501025136214612_210/latch_enable_in
+ scan_wrapper_339501025136214612_209/scan_select_in scan_wrapper_339501025136214612_210/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341567111632519764_140 scan_wrapper_341567111632519764_140/clk_in scan_wrapper_341631485498884690_141/clk_in
+ scan_wrapper_341567111632519764_140/data_in scan_wrapper_341631485498884690_141/data_in
+ scan_wrapper_341567111632519764_140/latch_enable_in scan_wrapper_341631485498884690_141/latch_enable_in
+ scan_wrapper_341567111632519764_140/scan_select_in scan_wrapper_341631485498884690_141/scan_select_in
+ vccd1 vssd1 scan_wrapper_341567111632519764
Xscan_wrapper_339501025136214612_381 scan_wrapper_339501025136214612_381/clk_in scan_wrapper_339501025136214612_382/clk_in
+ scan_wrapper_339501025136214612_381/data_in scan_wrapper_339501025136214612_382/data_in
+ scan_wrapper_339501025136214612_381/latch_enable_in scan_wrapper_339501025136214612_382/latch_enable_in
+ scan_wrapper_339501025136214612_381/scan_select_in scan_wrapper_339501025136214612_382/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_392 scan_wrapper_339501025136214612_392/clk_in scan_wrapper_339501025136214612_393/clk_in
+ scan_wrapper_339501025136214612_392/data_in scan_wrapper_339501025136214612_393/data_in
+ scan_wrapper_339501025136214612_392/latch_enable_in scan_wrapper_339501025136214612_393/latch_enable_in
+ scan_wrapper_339501025136214612_392/scan_select_in scan_wrapper_339501025136214612_393/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_370 scan_wrapper_339501025136214612_370/clk_in scan_wrapper_339501025136214612_371/clk_in
+ scan_wrapper_339501025136214612_370/data_in scan_wrapper_339501025136214612_371/data_in
+ scan_wrapper_339501025136214612_370/latch_enable_in scan_wrapper_339501025136214612_371/latch_enable_in
+ scan_wrapper_339501025136214612_370/scan_select_in scan_wrapper_339501025136214612_371/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341353928049295956_54 scan_wrapper_341353928049295956_54/clk_in scan_wrapper_341353780122485332_55/clk_in
+ scan_wrapper_341353928049295956_54/data_in scan_wrapper_341353780122485332_55/data_in
+ scan_wrapper_341353928049295956_54/latch_enable_in scan_wrapper_341353780122485332_55/latch_enable_in
+ scan_wrapper_341353928049295956_54/scan_select_in scan_wrapper_341353780122485332_55/scan_select_in
+ vccd1 vssd1 scan_wrapper_341353928049295956
Xscan_wrapper_341432284947153491_80 scan_wrapper_341432284947153491_80/clk_in scan_wrapper_341457971277988435_81/clk_in
+ scan_wrapper_341432284947153491_80/data_in scan_wrapper_341457971277988435_81/data_in
+ scan_wrapper_341432284947153491_80/latch_enable_in scan_wrapper_341457971277988435_81/latch_enable_in
+ scan_wrapper_341432284947153491_80/scan_select_in scan_wrapper_341457971277988435_81/scan_select_in
+ vccd1 vssd1 scan_wrapper_341432284947153491
Xscan_wrapper_341353777861755476_58 scan_wrapper_341353777861755476_58/clk_in scan_wrapper_341359404107432531_59/clk_in
+ scan_wrapper_341353777861755476_58/data_in scan_wrapper_341359404107432531_59/data_in
+ scan_wrapper_341353777861755476_58/latch_enable_in scan_wrapper_341359404107432531_59/latch_enable_in
+ scan_wrapper_341353777861755476_58/scan_select_in scan_wrapper_341359404107432531_59/scan_select_in
+ vccd1 vssd1 scan_wrapper_341353777861755476
Xscan_wrapper_339501025136214612_382 scan_wrapper_339501025136214612_382/clk_in scan_wrapper_339501025136214612_383/clk_in
+ scan_wrapper_339501025136214612_382/data_in scan_wrapper_339501025136214612_383/data_in
+ scan_wrapper_339501025136214612_382/latch_enable_in scan_wrapper_339501025136214612_383/latch_enable_in
+ scan_wrapper_339501025136214612_382/scan_select_in scan_wrapper_339501025136214612_383/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_360 scan_wrapper_339501025136214612_360/clk_in scan_wrapper_339501025136214612_361/clk_in
+ scan_wrapper_339501025136214612_360/data_in scan_wrapper_339501025136214612_361/data_in
+ scan_wrapper_339501025136214612_360/latch_enable_in scan_wrapper_339501025136214612_361/latch_enable_in
+ scan_wrapper_339501025136214612_360/scan_select_in scan_wrapper_339501025136214612_361/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_371 scan_wrapper_339501025136214612_371/clk_in scan_wrapper_339501025136214612_372/clk_in
+ scan_wrapper_339501025136214612_371/data_in scan_wrapper_339501025136214612_372/data_in
+ scan_wrapper_339501025136214612_371/latch_enable_in scan_wrapper_339501025136214612_372/latch_enable_in
+ scan_wrapper_339501025136214612_371/scan_select_in scan_wrapper_339501025136214612_372/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_393 scan_wrapper_339501025136214612_393/clk_in scan_wrapper_339501025136214612_394/clk_in
+ scan_wrapper_339501025136214612_393/data_in scan_wrapper_339501025136214612_394/data_in
+ scan_wrapper_339501025136214612_393/latch_enable_in scan_wrapper_339501025136214612_394/latch_enable_in
+ scan_wrapper_339501025136214612_393/scan_select_in scan_wrapper_339501025136214612_394/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_190 scan_wrapper_339501025136214612_190/clk_in scan_wrapper_339501025136214612_191/clk_in
+ scan_wrapper_339501025136214612_190/data_in scan_wrapper_339501025136214612_191/data_in
+ scan_wrapper_339501025136214612_190/latch_enable_in scan_wrapper_339501025136214612_191/latch_enable_in
+ scan_wrapper_339501025136214612_190/scan_select_in scan_wrapper_339501025136214612_191/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341159915403870803_9 scan_wrapper_341159915403870803_9/clk_in scan_wrapper_341159915403870803_9/clk_out
+ scan_wrapper_341159915403870803_9/data_in scan_wrapper_341159915403870803_9/data_out
+ scan_wrapper_341159915403870803_9/latch_enable_in scan_wrapper_341159915403870803_9/latch_enable_out
+ scan_wrapper_341159915403870803_9/scan_select_in scan_wrapper_341159915403870803_9/scan_select_out
+ vccd1 vssd1 scan_wrapper_341159915403870803
Xscan_wrapper_341449297858921043_94 scan_wrapper_341449297858921043_94/clk_in scan_wrapper_341710255833481812_95/clk_in
+ scan_wrapper_341449297858921043_94/data_in scan_wrapper_341710255833481812_95/data_in
+ scan_wrapper_341449297858921043_94/latch_enable_in scan_wrapper_341710255833481812_95/latch_enable_in
+ scan_wrapper_341449297858921043_94/scan_select_in scan_wrapper_341710255833481812_95/scan_select_in
+ vccd1 vssd1 scan_wrapper_341449297858921043
Xscan_wrapper_341205508016833108_24 scan_wrapper_341205508016833108_24/clk_in scan_wrapper_341162950004834900_25/clk_in
+ scan_wrapper_341205508016833108_24/data_in scan_wrapper_341162950004834900_25/data_in
+ scan_wrapper_341205508016833108_24/latch_enable_in scan_wrapper_341162950004834900_25/latch_enable_in
+ scan_wrapper_341205508016833108_24/scan_select_in scan_wrapper_341162950004834900_25/scan_select_in
+ vccd1 vssd1 scan_wrapper_341205508016833108
Xscan_wrapper_341557831870186068_121 scan_wrapper_341557831870186068_121/clk_in scan_wrapper_341569483755749970_122/clk_in
+ scan_wrapper_341557831870186068_121/data_in scan_wrapper_341569483755749970_122/data_in
+ scan_wrapper_341557831870186068_121/latch_enable_in scan_wrapper_341569483755749970_122/latch_enable_in
+ scan_wrapper_341557831870186068_121/scan_select_in scan_wrapper_341569483755749970_122/scan_select_in
+ vccd1 vssd1 scan_wrapper_341557831870186068
Xscan_wrapper_340218629792465491_2 scan_wrapper_340218629792465491_2/clk_in scan_wrapper_340318610245288530_3/clk_in
+ scan_wrapper_340218629792465491_2/data_in scan_wrapper_340318610245288530_3/data_in
+ scan_wrapper_340218629792465491_2/latch_enable_in scan_wrapper_340318610245288530_3/latch_enable_in
+ scan_wrapper_340218629792465491_2/scan_select_in scan_wrapper_340318610245288530_3/scan_select_in
+ vccd1 vssd1 scan_wrapper_340218629792465491
Xscan_wrapper_341631644820570706_148 scan_wrapper_341631644820570706_148/clk_in scan_wrapper_340596276030603858_149/clk_in
+ scan_wrapper_341631644820570706_148/data_in scan_wrapper_340596276030603858_149/data_in
+ scan_wrapper_341631644820570706_148/latch_enable_in scan_wrapper_340596276030603858_149/latch_enable_in
+ scan_wrapper_341631644820570706_148/scan_select_in scan_wrapper_340596276030603858_149/scan_select_in
+ vccd1 vssd1 scan_wrapper_341631644820570706
Xscan_wrapper_339501025136214612_383 scan_wrapper_339501025136214612_383/clk_in scan_wrapper_339501025136214612_384/clk_in
+ scan_wrapper_339501025136214612_383/data_in scan_wrapper_339501025136214612_384/data_in
+ scan_wrapper_339501025136214612_383/latch_enable_in scan_wrapper_339501025136214612_384/latch_enable_in
+ scan_wrapper_339501025136214612_383/scan_select_in scan_wrapper_339501025136214612_384/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_350 scan_wrapper_339501025136214612_350/clk_in scan_wrapper_339501025136214612_351/clk_in
+ scan_wrapper_339501025136214612_350/data_in scan_wrapper_339501025136214612_351/data_in
+ scan_wrapper_339501025136214612_350/latch_enable_in scan_wrapper_339501025136214612_351/latch_enable_in
+ scan_wrapper_339501025136214612_350/scan_select_in scan_wrapper_339501025136214612_351/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_361 scan_wrapper_339501025136214612_361/clk_in scan_wrapper_339501025136214612_362/clk_in
+ scan_wrapper_339501025136214612_361/data_in scan_wrapper_339501025136214612_362/data_in
+ scan_wrapper_339501025136214612_361/latch_enable_in scan_wrapper_339501025136214612_362/latch_enable_in
+ scan_wrapper_339501025136214612_361/scan_select_in scan_wrapper_339501025136214612_362/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_372 scan_wrapper_339501025136214612_372/clk_in scan_wrapper_339501025136214612_373/clk_in
+ scan_wrapper_339501025136214612_372/data_in scan_wrapper_339501025136214612_373/data_in
+ scan_wrapper_339501025136214612_372/latch_enable_in scan_wrapper_339501025136214612_373/latch_enable_in
+ scan_wrapper_339501025136214612_372/scan_select_in scan_wrapper_339501025136214612_373/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_394 scan_wrapper_339501025136214612_394/clk_in scan_wrapper_339501025136214612_395/clk_in
+ scan_wrapper_339501025136214612_394/data_in scan_wrapper_339501025136214612_395/data_in
+ scan_wrapper_339501025136214612_394/latch_enable_in scan_wrapper_339501025136214612_395/latch_enable_in
+ scan_wrapper_339501025136214612_394/scan_select_in scan_wrapper_339501025136214612_395/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341608297106768466_131 scan_wrapper_341608297106768466_131/clk_in scan_wrapper_341802448429515346_132/clk_in
+ scan_wrapper_341608297106768466_131/data_in scan_wrapper_341802448429515346_132/data_in
+ scan_wrapper_341608297106768466_131/latch_enable_in scan_wrapper_341802448429515346_132/latch_enable_in
+ scan_wrapper_341608297106768466_131/scan_select_in scan_wrapper_341802448429515346_132/scan_select_in
+ vccd1 vssd1 scan_wrapper_341608297106768466
Xscan_wrapper_341569483755749970_122 scan_wrapper_341569483755749970_122/clk_in scan_wrapper_341573751072096850_123/clk_in
+ scan_wrapper_341569483755749970_122/data_in scan_wrapper_341573751072096850_123/data_in
+ scan_wrapper_341569483755749970_122/latch_enable_in scan_wrapper_341573751072096850_123/latch_enable_in
+ scan_wrapper_341569483755749970_122/scan_select_in scan_wrapper_341573751072096850_123/scan_select_in
+ vccd1 vssd1 scan_wrapper_341569483755749970
Xscan_wrapper_339501025136214612_191 scan_wrapper_339501025136214612_191/clk_in scan_wrapper_339501025136214612_192/clk_in
+ scan_wrapper_339501025136214612_191/data_in scan_wrapper_339501025136214612_192/data_in
+ scan_wrapper_339501025136214612_191/latch_enable_in scan_wrapper_339501025136214612_192/latch_enable_in
+ scan_wrapper_339501025136214612_191/scan_select_in scan_wrapper_339501025136214612_192/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_180 scan_wrapper_339501025136214612_180/clk_in scan_wrapper_339501025136214612_181/clk_in
+ scan_wrapper_339501025136214612_180/data_in scan_wrapper_339501025136214612_181/data_in
+ scan_wrapper_339501025136214612_180/latch_enable_in scan_wrapper_339501025136214612_181/latch_enable_in
+ scan_wrapper_339501025136214612_180/scan_select_in scan_wrapper_339501025136214612_181/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341279123277087315_62 scan_wrapper_341279123277087315_62/clk_in scan_wrapper_341802655228625490_63/clk_in
+ scan_wrapper_341279123277087315_62/data_in scan_wrapper_341802655228625490_63/data_in
+ scan_wrapper_341279123277087315_62/latch_enable_in scan_wrapper_341802655228625490_63/latch_enable_in
+ scan_wrapper_341279123277087315_62/scan_select_in scan_wrapper_341802655228625490_63/scan_select_in
+ vccd1 vssd1 scan_wrapper_341279123277087315
Xscan_wrapper_341353780122485332_55 scan_wrapper_341353780122485332_55/clk_in scan_wrapper_341193419111006803_56/clk_in
+ scan_wrapper_341353780122485332_55/data_in scan_wrapper_341193419111006803_56/data_in
+ scan_wrapper_341353780122485332_55/latch_enable_in scan_wrapper_341193419111006803_56/latch_enable_in
+ scan_wrapper_341353780122485332_55/scan_select_in scan_wrapper_341193419111006803_56/scan_select_in
+ vccd1 vssd1 scan_wrapper_341353780122485332
Xscan_wrapper_341624400621077076_138 scan_wrapper_341624400621077076_138/clk_in scan_wrapper_341614536664547922_139/clk_in
+ scan_wrapper_341624400621077076_138/data_in scan_wrapper_341614536664547922_139/data_in
+ scan_wrapper_341624400621077076_138/latch_enable_in scan_wrapper_341614536664547922_139/latch_enable_in
+ scan_wrapper_341624400621077076_138/scan_select_in scan_wrapper_341614536664547922_139/scan_select_in
+ vccd1 vssd1 scan_wrapper_341624400621077076
Xscan_wrapper_339501025136214612_384 scan_wrapper_339501025136214612_384/clk_in scan_wrapper_339501025136214612_385/clk_in
+ scan_wrapper_339501025136214612_384/data_in scan_wrapper_339501025136214612_385/data_in
+ scan_wrapper_339501025136214612_384/latch_enable_in scan_wrapper_339501025136214612_385/latch_enable_in
+ scan_wrapper_339501025136214612_384/scan_select_in scan_wrapper_339501025136214612_385/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341632596577354323_142 scan_wrapper_341632596577354323_142/clk_in scan_wrapper_341628725785264722_143/clk_in
+ scan_wrapper_341632596577354323_142/data_in scan_wrapper_341628725785264722_143/data_in
+ scan_wrapper_341632596577354323_142/latch_enable_in scan_wrapper_341628725785264722_143/latch_enable_in
+ scan_wrapper_341632596577354323_142/scan_select_in scan_wrapper_341628725785264722_143/scan_select_in
+ vccd1 vssd1 scan_wrapper_341632596577354323
Xscan_wrapper_339501025136214612_351 scan_wrapper_339501025136214612_351/clk_in scan_wrapper_339501025136214612_352/clk_in
+ scan_wrapper_339501025136214612_351/data_in scan_wrapper_339501025136214612_352/data_in
+ scan_wrapper_339501025136214612_351/latch_enable_in scan_wrapper_339501025136214612_352/latch_enable_in
+ scan_wrapper_339501025136214612_351/scan_select_in scan_wrapper_339501025136214612_352/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_340 scan_wrapper_339501025136214612_340/clk_in scan_wrapper_339501025136214612_341/clk_in
+ scan_wrapper_339501025136214612_340/data_in scan_wrapper_339501025136214612_341/data_in
+ scan_wrapper_339501025136214612_340/latch_enable_in scan_wrapper_339501025136214612_341/latch_enable_in
+ scan_wrapper_339501025136214612_340/scan_select_in scan_wrapper_339501025136214612_341/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_362 scan_wrapper_339501025136214612_362/clk_in scan_wrapper_339501025136214612_363/clk_in
+ scan_wrapper_339501025136214612_362/data_in scan_wrapper_339501025136214612_363/data_in
+ scan_wrapper_339501025136214612_362/latch_enable_in scan_wrapper_339501025136214612_363/latch_enable_in
+ scan_wrapper_339501025136214612_362/scan_select_in scan_wrapper_339501025136214612_363/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_373 scan_wrapper_339501025136214612_373/clk_in scan_wrapper_339501025136214612_374/clk_in
+ scan_wrapper_339501025136214612_373/data_in scan_wrapper_339501025136214612_374/data_in
+ scan_wrapper_339501025136214612_373/latch_enable_in scan_wrapper_339501025136214612_374/latch_enable_in
+ scan_wrapper_339501025136214612_373/scan_select_in scan_wrapper_339501025136214612_374/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_395 scan_wrapper_339501025136214612_395/clk_in scan_wrapper_339501025136214612_396/clk_in
+ scan_wrapper_339501025136214612_395/data_in scan_wrapper_339501025136214612_396/data_in
+ scan_wrapper_339501025136214612_395/latch_enable_in scan_wrapper_339501025136214612_396/latch_enable_in
+ scan_wrapper_339501025136214612_395/scan_select_in scan_wrapper_339501025136214612_396/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341266732010177108_57 scan_wrapper_341266732010177108_57/clk_in scan_wrapper_341353777861755476_58/clk_in
+ scan_wrapper_341266732010177108_57/data_in scan_wrapper_341353777861755476_58/data_in
+ scan_wrapper_341266732010177108_57/latch_enable_in scan_wrapper_341353777861755476_58/latch_enable_in
+ scan_wrapper_341266732010177108_57/scan_select_in scan_wrapper_341353777861755476_58/scan_select_in
+ vccd1 vssd1 scan_wrapper_341266732010177108
Xscan_wrapper_341528610027340372_109 scan_wrapper_341528610027340372_109/clk_in scan_wrapper_341424636358034002_110/clk_in
+ scan_wrapper_341528610027340372_109/data_in scan_wrapper_341424636358034002_110/data_in
+ scan_wrapper_341528610027340372_109/latch_enable_in scan_wrapper_341424636358034002_110/latch_enable_in
+ scan_wrapper_341528610027340372_109/scan_select_in scan_wrapper_341424636358034002_110/scan_select_in
+ vccd1 vssd1 scan_wrapper_341528610027340372
Xscan_wrapper_339501025136214612_170 scan_wrapper_339501025136214612_170/clk_in scan_wrapper_339501025136214612_171/clk_in
+ scan_wrapper_339501025136214612_170/data_in scan_wrapper_339501025136214612_171/data_in
+ scan_wrapper_339501025136214612_170/latch_enable_in scan_wrapper_339501025136214612_171/latch_enable_in
+ scan_wrapper_339501025136214612_170/scan_select_in scan_wrapper_339501025136214612_171/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_192 scan_wrapper_339501025136214612_192/clk_in scan_wrapper_339501025136214612_193/clk_in
+ scan_wrapper_339501025136214612_192/data_in scan_wrapper_339501025136214612_193/data_in
+ scan_wrapper_339501025136214612_192/latch_enable_in scan_wrapper_339501025136214612_193/latch_enable_in
+ scan_wrapper_339501025136214612_192/scan_select_in scan_wrapper_339501025136214612_193/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_181 scan_wrapper_339501025136214612_181/clk_in scan_wrapper_339501025136214612_182/clk_in
+ scan_wrapper_339501025136214612_181/data_in scan_wrapper_339501025136214612_182/data_in
+ scan_wrapper_339501025136214612_181/latch_enable_in scan_wrapper_339501025136214612_182/latch_enable_in
+ scan_wrapper_339501025136214612_181/scan_select_in scan_wrapper_339501025136214612_182/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341464767397888596_83 scan_wrapper_341464767397888596_83/clk_in scan_wrapper_341476989274686036_84/clk_in
+ scan_wrapper_341464767397888596_83/data_in scan_wrapper_341476989274686036_84/data_in
+ scan_wrapper_341464767397888596_83/latch_enable_in scan_wrapper_341476989274686036_84/latch_enable_in
+ scan_wrapper_341464767397888596_83/scan_select_in scan_wrapper_341476989274686036_84/scan_select_in
+ vccd1 vssd1 scan_wrapper_341464767397888596
Xscan_wrapper_341497971083313748_87 scan_wrapper_341497971083313748_87/clk_in scan_wrapper_341497964482527828_88/clk_in
+ scan_wrapper_341497971083313748_87/data_in scan_wrapper_341497964482527828_88/data_in
+ scan_wrapper_341497971083313748_87/latch_enable_in scan_wrapper_341497964482527828_88/latch_enable_in
+ scan_wrapper_341497971083313748_87/scan_select_in scan_wrapper_341497964482527828_88/scan_select_in
+ vccd1 vssd1 scan_wrapper_341497971083313748
Xscan_wrapper_341164910646919762_34 scan_wrapper_341164910646919762_34/clk_in scan_wrapper_341233739099013714_35/clk_in
+ scan_wrapper_341164910646919762_34/data_in scan_wrapper_341233739099013714_35/data_in
+ scan_wrapper_341164910646919762_34/latch_enable_in scan_wrapper_341233739099013714_35/latch_enable_in
+ scan_wrapper_341164910646919762_34/scan_select_in scan_wrapper_341233739099013714_35/scan_select_in
+ vccd1 vssd1 scan_wrapper_341164910646919762
Xscan_wrapper_340067262721426004_96 scan_wrapper_340067262721426004_96/clk_in scan_wrapper_341462925422101075_97/clk_in
+ scan_wrapper_340067262721426004_96/data_in scan_wrapper_341462925422101075_97/data_in
+ scan_wrapper_340067262721426004_96/latch_enable_in scan_wrapper_341462925422101075_97/latch_enable_in
+ scan_wrapper_340067262721426004_96/scan_select_in scan_wrapper_341462925422101075_97/scan_select_in
+ vccd1 vssd1 scan_wrapper_340067262721426004
Xscan_wrapper_341174480471589458_69 scan_wrapper_341174480471589458_69/clk_in scan_wrapper_341419328215712339_70/clk_in
+ scan_wrapper_341174480471589458_69/data_in scan_wrapper_341419328215712339_70/data_in
+ scan_wrapper_341174480471589458_69/latch_enable_in scan_wrapper_341419328215712339_70/latch_enable_in
+ scan_wrapper_341174480471589458_69/scan_select_in scan_wrapper_341419328215712339_70/scan_select_in
+ vccd1 vssd1 scan_wrapper_341174480471589458
Xscan_wrapper_339501025136214612_385 scan_wrapper_339501025136214612_385/clk_in scan_wrapper_339501025136214612_386/clk_in
+ scan_wrapper_339501025136214612_385/data_in scan_wrapper_339501025136214612_386/data_in
+ scan_wrapper_339501025136214612_385/latch_enable_in scan_wrapper_339501025136214612_386/latch_enable_in
+ scan_wrapper_339501025136214612_385/scan_select_in scan_wrapper_339501025136214612_386/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_330 scan_wrapper_339501025136214612_330/clk_in scan_wrapper_339501025136214612_331/clk_in
+ scan_wrapper_339501025136214612_330/data_in scan_wrapper_339501025136214612_331/data_in
+ scan_wrapper_339501025136214612_330/latch_enable_in scan_wrapper_339501025136214612_331/latch_enable_in
+ scan_wrapper_339501025136214612_330/scan_select_in scan_wrapper_339501025136214612_331/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_352 scan_wrapper_339501025136214612_352/clk_in scan_wrapper_339501025136214612_353/clk_in
+ scan_wrapper_339501025136214612_352/data_in scan_wrapper_339501025136214612_353/data_in
+ scan_wrapper_339501025136214612_352/latch_enable_in scan_wrapper_339501025136214612_353/latch_enable_in
+ scan_wrapper_339501025136214612_352/scan_select_in scan_wrapper_339501025136214612_353/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_341 scan_wrapper_339501025136214612_341/clk_in scan_wrapper_339501025136214612_342/clk_in
+ scan_wrapper_339501025136214612_341/data_in scan_wrapper_339501025136214612_342/data_in
+ scan_wrapper_339501025136214612_341/latch_enable_in scan_wrapper_339501025136214612_342/latch_enable_in
+ scan_wrapper_339501025136214612_341/scan_select_in scan_wrapper_339501025136214612_342/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_363 scan_wrapper_339501025136214612_363/clk_in scan_wrapper_339501025136214612_364/clk_in
+ scan_wrapper_339501025136214612_363/data_in scan_wrapper_339501025136214612_364/data_in
+ scan_wrapper_339501025136214612_363/latch_enable_in scan_wrapper_339501025136214612_364/latch_enable_in
+ scan_wrapper_339501025136214612_363/scan_select_in scan_wrapper_339501025136214612_364/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_374 scan_wrapper_339501025136214612_374/clk_in scan_wrapper_339501025136214612_375/clk_in
+ scan_wrapper_339501025136214612_374/data_in scan_wrapper_339501025136214612_375/data_in
+ scan_wrapper_339501025136214612_374/latch_enable_in scan_wrapper_339501025136214612_375/latch_enable_in
+ scan_wrapper_339501025136214612_374/scan_select_in scan_wrapper_339501025136214612_375/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_396 scan_wrapper_339501025136214612_396/clk_in scan_wrapper_339501025136214612_397/clk_in
+ scan_wrapper_339501025136214612_396/data_in scan_wrapper_339501025136214612_397/data_in
+ scan_wrapper_339501025136214612_396/latch_enable_in scan_wrapper_339501025136214612_397/latch_enable_in
+ scan_wrapper_339501025136214612_396/scan_select_in scan_wrapper_339501025136214612_397/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_160 scan_wrapper_339501025136214612_160/clk_in scan_wrapper_339501025136214612_161/clk_in
+ scan_wrapper_339501025136214612_160/data_in scan_wrapper_339501025136214612_161/data_in
+ scan_wrapper_339501025136214612_160/latch_enable_in scan_wrapper_339501025136214612_161/latch_enable_in
+ scan_wrapper_339501025136214612_160/scan_select_in scan_wrapper_339501025136214612_161/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_171 scan_wrapper_339501025136214612_171/clk_in scan_wrapper_339501025136214612_172/clk_in
+ scan_wrapper_339501025136214612_171/data_in scan_wrapper_339501025136214612_172/data_in
+ scan_wrapper_339501025136214612_171/latch_enable_in scan_wrapper_339501025136214612_172/latch_enable_in
+ scan_wrapper_339501025136214612_171/scan_select_in scan_wrapper_339501025136214612_172/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_193 scan_wrapper_339501025136214612_193/clk_in scan_wrapper_339501025136214612_194/clk_in
+ scan_wrapper_339501025136214612_193/data_in scan_wrapper_339501025136214612_194/data_in
+ scan_wrapper_339501025136214612_193/latch_enable_in scan_wrapper_339501025136214612_194/latch_enable_in
+ scan_wrapper_339501025136214612_193/scan_select_in scan_wrapper_339501025136214612_194/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_182 scan_wrapper_339501025136214612_182/clk_in scan_wrapper_339501025136214612_183/clk_in
+ scan_wrapper_339501025136214612_182/data_in scan_wrapper_339501025136214612_183/data_in
+ scan_wrapper_339501025136214612_182/latch_enable_in scan_wrapper_339501025136214612_183/latch_enable_in
+ scan_wrapper_339501025136214612_182/scan_select_in scan_wrapper_339501025136214612_183/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341678527574180436_150 scan_wrapper_341678527574180436_150/clk_in scan_wrapper_339501025136214612_151/clk_in
+ scan_wrapper_341678527574180436_150/data_in scan_wrapper_339501025136214612_151/data_in
+ scan_wrapper_341678527574180436_150/latch_enable_in scan_wrapper_339501025136214612_151/latch_enable_in
+ scan_wrapper_341678527574180436_150/scan_select_in scan_wrapper_339501025136214612_151/scan_select_in
+ vccd1 vssd1 scan_wrapper_341678527574180436
Xscan_controller io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18]
+ io_in[19] io_in[20] wb_clk_i io_in[8] io_in[9] io_in[21] io_in[22] io_in[23] io_in[24]
+ io_in[25] io_in[26] io_in[27] io_in[28] la_data_in[0] la_data_in[1] la_data_out[0]
+ la_data_in[3] la_data_in[2] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[29] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35]
+ io_out[36] io_out[37] wb_rst_i scan_controller/scan_clk_in scan_controller/scan_clk_out
+ scan_controller/scan_data_in scan_controller/scan_data_out scan_controller/scan_latch_en
+ scan_controller/scan_select io_in[11] io_out[10] vccd1 vssd1 scan_controller
Xscan_wrapper_019235602376235615_77 scan_wrapper_019235602376235615_77/clk_in scan_wrapper_341450853309219412_78/clk_in
+ scan_wrapper_019235602376235615_77/data_in scan_wrapper_341450853309219412_78/data_in
+ scan_wrapper_019235602376235615_77/latch_enable_in scan_wrapper_341450853309219412_78/latch_enable_in
+ scan_wrapper_019235602376235615_77/scan_select_in scan_wrapper_341450853309219412_78/scan_select_in
+ vccd1 vssd1 scan_wrapper_019235602376235615
Xscan_wrapper_341178481588044372_19 scan_wrapper_341178481588044372_19/clk_in scan_wrapper_341176884318437971_20/clk_in
+ scan_wrapper_341178481588044372_19/data_in scan_wrapper_341176884318437971_20/data_in
+ scan_wrapper_341178481588044372_19/latch_enable_in scan_wrapper_341176884318437971_20/latch_enable_in
+ scan_wrapper_341178481588044372_19/scan_select_in scan_wrapper_341176884318437971_20/scan_select_in
+ vccd1 vssd1 scan_wrapper_341178481588044372
Xscan_wrapper_341426151397261906_145 scan_wrapper_341426151397261906_145/clk_in scan_wrapper_341629415144292948_146/clk_in
+ scan_wrapper_341426151397261906_145/data_in scan_wrapper_341629415144292948_146/data_in
+ scan_wrapper_341426151397261906_145/latch_enable_in scan_wrapper_341629415144292948_146/latch_enable_in
+ scan_wrapper_341426151397261906_145/scan_select_in scan_wrapper_341629415144292948_146/scan_select_in
+ vccd1 vssd1 scan_wrapper_341426151397261906
Xscan_wrapper_339501025136214612_386 scan_wrapper_339501025136214612_386/clk_in scan_wrapper_339501025136214612_387/clk_in
+ scan_wrapper_339501025136214612_386/data_in scan_wrapper_339501025136214612_387/data_in
+ scan_wrapper_339501025136214612_386/latch_enable_in scan_wrapper_339501025136214612_387/latch_enable_in
+ scan_wrapper_339501025136214612_386/scan_select_in scan_wrapper_339501025136214612_387/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_320 scan_wrapper_339501025136214612_320/clk_in scan_wrapper_339501025136214612_321/clk_in
+ scan_wrapper_339501025136214612_320/data_in scan_wrapper_339501025136214612_321/data_in
+ scan_wrapper_339501025136214612_320/latch_enable_in scan_wrapper_339501025136214612_321/latch_enable_in
+ scan_wrapper_339501025136214612_320/scan_select_in scan_wrapper_339501025136214612_321/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_331 scan_wrapper_339501025136214612_331/clk_in scan_wrapper_339501025136214612_332/clk_in
+ scan_wrapper_339501025136214612_331/data_in scan_wrapper_339501025136214612_332/data_in
+ scan_wrapper_339501025136214612_331/latch_enable_in scan_wrapper_339501025136214612_332/latch_enable_in
+ scan_wrapper_339501025136214612_331/scan_select_in scan_wrapper_339501025136214612_332/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_353 scan_wrapper_339501025136214612_353/clk_in scan_wrapper_339501025136214612_354/clk_in
+ scan_wrapper_339501025136214612_353/data_in scan_wrapper_339501025136214612_354/data_in
+ scan_wrapper_339501025136214612_353/latch_enable_in scan_wrapper_339501025136214612_354/latch_enable_in
+ scan_wrapper_339501025136214612_353/scan_select_in scan_wrapper_339501025136214612_354/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_342 scan_wrapper_339501025136214612_342/clk_in scan_wrapper_339501025136214612_343/clk_in
+ scan_wrapper_339501025136214612_342/data_in scan_wrapper_339501025136214612_343/data_in
+ scan_wrapper_339501025136214612_342/latch_enable_in scan_wrapper_339501025136214612_343/latch_enable_in
+ scan_wrapper_339501025136214612_342/scan_select_in scan_wrapper_339501025136214612_343/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_364 scan_wrapper_339501025136214612_364/clk_in scan_wrapper_339501025136214612_365/clk_in
+ scan_wrapper_339501025136214612_364/data_in scan_wrapper_339501025136214612_365/data_in
+ scan_wrapper_339501025136214612_364/latch_enable_in scan_wrapper_339501025136214612_365/latch_enable_in
+ scan_wrapper_339501025136214612_364/scan_select_in scan_wrapper_339501025136214612_365/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_375 scan_wrapper_339501025136214612_375/clk_in scan_wrapper_339501025136214612_376/clk_in
+ scan_wrapper_339501025136214612_375/data_in scan_wrapper_339501025136214612_376/data_in
+ scan_wrapper_339501025136214612_375/latch_enable_in scan_wrapper_339501025136214612_376/latch_enable_in
+ scan_wrapper_339501025136214612_375/scan_select_in scan_wrapper_339501025136214612_376/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_397 scan_wrapper_339501025136214612_397/clk_in scan_wrapper_339501025136214612_398/clk_in
+ scan_wrapper_339501025136214612_397/data_in scan_wrapper_339501025136214612_398/data_in
+ scan_wrapper_339501025136214612_397/latch_enable_in scan_wrapper_339501025136214612_398/latch_enable_in
+ scan_wrapper_339501025136214612_397/scan_select_in scan_wrapper_339501025136214612_398/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_161 scan_wrapper_339501025136214612_161/clk_in scan_wrapper_339501025136214612_162/clk_in
+ scan_wrapper_339501025136214612_161/data_in scan_wrapper_339501025136214612_162/data_in
+ scan_wrapper_339501025136214612_161/latch_enable_in scan_wrapper_339501025136214612_162/latch_enable_in
+ scan_wrapper_339501025136214612_161/scan_select_in scan_wrapper_339501025136214612_162/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_172 scan_wrapper_339501025136214612_172/clk_in scan_wrapper_339501025136214612_173/clk_in
+ scan_wrapper_339501025136214612_172/data_in scan_wrapper_339501025136214612_173/data_in
+ scan_wrapper_339501025136214612_172/latch_enable_in scan_wrapper_339501025136214612_173/latch_enable_in
+ scan_wrapper_339501025136214612_172/scan_select_in scan_wrapper_339501025136214612_173/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_194 scan_wrapper_339501025136214612_194/clk_in scan_wrapper_339501025136214612_195/clk_in
+ scan_wrapper_339501025136214612_194/data_in scan_wrapper_339501025136214612_195/data_in
+ scan_wrapper_339501025136214612_194/latch_enable_in scan_wrapper_339501025136214612_195/latch_enable_in
+ scan_wrapper_339501025136214612_194/scan_select_in scan_wrapper_339501025136214612_195/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_183 scan_wrapper_339501025136214612_183/clk_in scan_wrapper_339501025136214612_184/clk_in
+ scan_wrapper_339501025136214612_183/data_in scan_wrapper_339501025136214612_184/data_in
+ scan_wrapper_339501025136214612_183/latch_enable_in scan_wrapper_339501025136214612_184/latch_enable_in
+ scan_wrapper_339501025136214612_183/scan_select_in scan_wrapper_339501025136214612_184/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341152580068442706_15 scan_wrapper_341152580068442706_15/clk_in scan_wrapper_341155178824598098_16/clk_in
+ scan_wrapper_341152580068442706_15/data_in scan_wrapper_341155178824598098_16/data_in
+ scan_wrapper_341152580068442706_15/latch_enable_in scan_wrapper_341155178824598098_16/latch_enable_in
+ scan_wrapper_341152580068442706_15/scan_select_in scan_wrapper_341155178824598098_16/scan_select_in
+ vccd1 vssd1 scan_wrapper_341152580068442706
Xscan_wrapper_341533740987581011_106 scan_wrapper_341533740987581011_106/clk_in scan_wrapper_341431502448362067_107/clk_in
+ scan_wrapper_341533740987581011_106/data_in scan_wrapper_341431502448362067_107/data_in
+ scan_wrapper_341533740987581011_106/latch_enable_in scan_wrapper_341431502448362067_107/latch_enable_in
+ scan_wrapper_341533740987581011_106/scan_select_in scan_wrapper_341431502448362067_107/scan_select_in
+ vccd1 vssd1 scan_wrapper_341533740987581011
Xscan_wrapper_341446083683025490_104 scan_wrapper_341446083683025490_104/clk_in scan_wrapper_341524192738411090_105/clk_in
+ scan_wrapper_341446083683025490_104/data_in scan_wrapper_341524192738411090_105/data_in
+ scan_wrapper_341446083683025490_104/latch_enable_in scan_wrapper_341524192738411090_105/latch_enable_in
+ scan_wrapper_341446083683025490_104/scan_select_in scan_wrapper_341524192738411090_105/scan_select_in
+ vccd1 vssd1 scan_wrapper_341446083683025490
Xscan_wrapper_341609034095264340_133 scan_wrapper_341609034095264340_133/clk_in scan_wrapper_341617722294010450_134/clk_in
+ scan_wrapper_341609034095264340_133/data_in scan_wrapper_341617722294010450_134/data_in
+ scan_wrapper_341609034095264340_133/latch_enable_in scan_wrapper_341617722294010450_134/latch_enable_in
+ scan_wrapper_341609034095264340_133/scan_select_in scan_wrapper_341617722294010450_134/scan_select_in
+ vccd1 vssd1 scan_wrapper_341609034095264340
Xscan_wrapper_339501025136214612_398 scan_wrapper_339501025136214612_398/clk_in scan_wrapper_339501025136214612_399/clk_in
+ scan_wrapper_339501025136214612_398/data_in scan_wrapper_339501025136214612_399/data_in
+ scan_wrapper_339501025136214612_398/latch_enable_in scan_wrapper_339501025136214612_399/latch_enable_in
+ scan_wrapper_339501025136214612_398/scan_select_in scan_wrapper_339501025136214612_399/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_387 scan_wrapper_339501025136214612_387/clk_in scan_wrapper_339501025136214612_388/clk_in
+ scan_wrapper_339501025136214612_387/data_in scan_wrapper_339501025136214612_388/data_in
+ scan_wrapper_339501025136214612_387/latch_enable_in scan_wrapper_339501025136214612_388/latch_enable_in
+ scan_wrapper_339501025136214612_387/scan_select_in scan_wrapper_339501025136214612_388/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_310 scan_wrapper_339501025136214612_310/clk_in scan_wrapper_339501025136214612_311/clk_in
+ scan_wrapper_339501025136214612_310/data_in scan_wrapper_339501025136214612_311/data_in
+ scan_wrapper_339501025136214612_310/latch_enable_in scan_wrapper_339501025136214612_311/latch_enable_in
+ scan_wrapper_339501025136214612_310/scan_select_in scan_wrapper_339501025136214612_311/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_321 scan_wrapper_339501025136214612_321/clk_in scan_wrapper_339501025136214612_322/clk_in
+ scan_wrapper_339501025136214612_321/data_in scan_wrapper_339501025136214612_322/data_in
+ scan_wrapper_339501025136214612_321/latch_enable_in scan_wrapper_339501025136214612_322/latch_enable_in
+ scan_wrapper_339501025136214612_321/scan_select_in scan_wrapper_339501025136214612_322/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_332 scan_wrapper_339501025136214612_332/clk_in scan_wrapper_339501025136214612_333/clk_in
+ scan_wrapper_339501025136214612_332/data_in scan_wrapper_339501025136214612_333/data_in
+ scan_wrapper_339501025136214612_332/latch_enable_in scan_wrapper_339501025136214612_333/latch_enable_in
+ scan_wrapper_339501025136214612_332/scan_select_in scan_wrapper_339501025136214612_333/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_354 scan_wrapper_339501025136214612_354/clk_in scan_wrapper_339501025136214612_355/clk_in
+ scan_wrapper_339501025136214612_354/data_in scan_wrapper_339501025136214612_355/data_in
+ scan_wrapper_339501025136214612_354/latch_enable_in scan_wrapper_339501025136214612_355/latch_enable_in
+ scan_wrapper_339501025136214612_354/scan_select_in scan_wrapper_339501025136214612_355/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_343 scan_wrapper_339501025136214612_343/clk_in scan_wrapper_339501025136214612_344/clk_in
+ scan_wrapper_339501025136214612_343/data_in scan_wrapper_339501025136214612_344/data_in
+ scan_wrapper_339501025136214612_343/latch_enable_in scan_wrapper_339501025136214612_344/latch_enable_in
+ scan_wrapper_339501025136214612_343/scan_select_in scan_wrapper_339501025136214612_344/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_365 scan_wrapper_339501025136214612_365/clk_in scan_wrapper_339501025136214612_366/clk_in
+ scan_wrapper_339501025136214612_365/data_in scan_wrapper_339501025136214612_366/data_in
+ scan_wrapper_339501025136214612_365/latch_enable_in scan_wrapper_339501025136214612_366/latch_enable_in
+ scan_wrapper_339501025136214612_365/scan_select_in scan_wrapper_339501025136214612_366/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_376 scan_wrapper_339501025136214612_376/clk_in scan_wrapper_339501025136214612_377/clk_in
+ scan_wrapper_339501025136214612_376/data_in scan_wrapper_339501025136214612_377/data_in
+ scan_wrapper_339501025136214612_376/latch_enable_in scan_wrapper_339501025136214612_377/latch_enable_in
+ scan_wrapper_339501025136214612_376/scan_select_in scan_wrapper_339501025136214612_377/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_151 scan_wrapper_339501025136214612_151/clk_in scan_wrapper_339501025136214612_152/clk_in
+ scan_wrapper_339501025136214612_151/data_in scan_wrapper_339501025136214612_152/data_in
+ scan_wrapper_339501025136214612_151/latch_enable_in scan_wrapper_339501025136214612_152/latch_enable_in
+ scan_wrapper_339501025136214612_151/scan_select_in scan_wrapper_339501025136214612_152/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_162 scan_wrapper_339501025136214612_162/clk_in scan_wrapper_339501025136214612_163/clk_in
+ scan_wrapper_339501025136214612_162/data_in scan_wrapper_339501025136214612_163/data_in
+ scan_wrapper_339501025136214612_162/latch_enable_in scan_wrapper_339501025136214612_163/latch_enable_in
+ scan_wrapper_339501025136214612_162/scan_select_in scan_wrapper_339501025136214612_163/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_173 scan_wrapper_339501025136214612_173/clk_in scan_wrapper_339501025136214612_174/clk_in
+ scan_wrapper_339501025136214612_173/data_in scan_wrapper_339501025136214612_174/data_in
+ scan_wrapper_339501025136214612_173/latch_enable_in scan_wrapper_339501025136214612_174/latch_enable_in
+ scan_wrapper_339501025136214612_173/scan_select_in scan_wrapper_339501025136214612_174/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_184 scan_wrapper_339501025136214612_184/clk_in scan_wrapper_339501025136214612_185/clk_in
+ scan_wrapper_339501025136214612_184/data_in scan_wrapper_339501025136214612_185/data_in
+ scan_wrapper_339501025136214612_184/latch_enable_in scan_wrapper_339501025136214612_185/latch_enable_in
+ scan_wrapper_339501025136214612_184/scan_select_in scan_wrapper_339501025136214612_185/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_195 scan_wrapper_339501025136214612_195/clk_in scan_wrapper_339501025136214612_196/clk_in
+ scan_wrapper_339501025136214612_195/data_in scan_wrapper_339501025136214612_196/data_in
+ scan_wrapper_339501025136214612_195/latch_enable_in scan_wrapper_339501025136214612_196/latch_enable_in
+ scan_wrapper_339501025136214612_195/scan_select_in scan_wrapper_339501025136214612_196/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341614536664547922_139 scan_wrapper_341614536664547922_139/clk_in scan_wrapper_341567111632519764_140/clk_in
+ scan_wrapper_341614536664547922_139/data_in scan_wrapper_341567111632519764_140/data_in
+ scan_wrapper_341614536664547922_139/latch_enable_in scan_wrapper_341567111632519764_140/latch_enable_in
+ scan_wrapper_341614536664547922_139/scan_select_in scan_wrapper_341567111632519764_140/scan_select_in
+ vccd1 vssd1 scan_wrapper_341614536664547922
Xscan_wrapper_341264068701586004_37 scan_wrapper_341264068701586004_37/clk_in scan_wrapper_341164228775772755_38/clk_in
+ scan_wrapper_341264068701586004_37/data_in scan_wrapper_341164228775772755_38/data_in
+ scan_wrapper_341264068701586004_37/latch_enable_in scan_wrapper_341164228775772755_38/latch_enable_in
+ scan_wrapper_341264068701586004_37/scan_select_in scan_wrapper_341164228775772755_38/scan_select_in
+ vccd1 vssd1 scan_wrapper_341264068701586004
Xscan_wrapper_339501025136214612_399 scan_wrapper_339501025136214612_399/clk_in scan_wrapper_339501025136214612_400/clk_in
+ scan_wrapper_339501025136214612_399/data_in scan_wrapper_339501025136214612_400/data_in
+ scan_wrapper_339501025136214612_399/latch_enable_in scan_wrapper_339501025136214612_400/latch_enable_in
+ scan_wrapper_339501025136214612_399/scan_select_in scan_wrapper_339501025136214612_400/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_388 scan_wrapper_339501025136214612_388/clk_in scan_wrapper_339501025136214612_389/clk_in
+ scan_wrapper_339501025136214612_388/data_in scan_wrapper_339501025136214612_389/data_in
+ scan_wrapper_339501025136214612_388/latch_enable_in scan_wrapper_339501025136214612_389/latch_enable_in
+ scan_wrapper_339501025136214612_388/scan_select_in scan_wrapper_339501025136214612_389/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_311 scan_wrapper_339501025136214612_311/clk_in scan_wrapper_339501025136214612_312/clk_in
+ scan_wrapper_339501025136214612_311/data_in scan_wrapper_339501025136214612_312/data_in
+ scan_wrapper_339501025136214612_311/latch_enable_in scan_wrapper_339501025136214612_312/latch_enable_in
+ scan_wrapper_339501025136214612_311/scan_select_in scan_wrapper_339501025136214612_312/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_300 scan_wrapper_339501025136214612_300/clk_in scan_wrapper_339501025136214612_301/clk_in
+ scan_wrapper_339501025136214612_300/data_in scan_wrapper_339501025136214612_301/data_in
+ scan_wrapper_339501025136214612_300/latch_enable_in scan_wrapper_339501025136214612_301/latch_enable_in
+ scan_wrapper_339501025136214612_300/scan_select_in scan_wrapper_339501025136214612_301/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_322 scan_wrapper_339501025136214612_322/clk_in scan_wrapper_339501025136214612_323/clk_in
+ scan_wrapper_339501025136214612_322/data_in scan_wrapper_339501025136214612_323/data_in
+ scan_wrapper_339501025136214612_322/latch_enable_in scan_wrapper_339501025136214612_323/latch_enable_in
+ scan_wrapper_339501025136214612_322/scan_select_in scan_wrapper_339501025136214612_323/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_333 scan_wrapper_339501025136214612_333/clk_in scan_wrapper_339501025136214612_334/clk_in
+ scan_wrapper_339501025136214612_333/data_in scan_wrapper_339501025136214612_334/data_in
+ scan_wrapper_339501025136214612_333/latch_enable_in scan_wrapper_339501025136214612_334/latch_enable_in
+ scan_wrapper_339501025136214612_333/scan_select_in scan_wrapper_339501025136214612_334/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_355 scan_wrapper_339501025136214612_355/clk_in scan_wrapper_339501025136214612_356/clk_in
+ scan_wrapper_339501025136214612_355/data_in scan_wrapper_339501025136214612_356/data_in
+ scan_wrapper_339501025136214612_355/latch_enable_in scan_wrapper_339501025136214612_356/latch_enable_in
+ scan_wrapper_339501025136214612_355/scan_select_in scan_wrapper_339501025136214612_356/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_344 scan_wrapper_339501025136214612_344/clk_in scan_wrapper_339501025136214612_345/clk_in
+ scan_wrapper_339501025136214612_344/data_in scan_wrapper_339501025136214612_345/data_in
+ scan_wrapper_339501025136214612_344/latch_enable_in scan_wrapper_339501025136214612_345/latch_enable_in
+ scan_wrapper_339501025136214612_344/scan_select_in scan_wrapper_339501025136214612_345/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_366 scan_wrapper_339501025136214612_366/clk_in scan_wrapper_339501025136214612_367/clk_in
+ scan_wrapper_339501025136214612_366/data_in scan_wrapper_339501025136214612_367/data_in
+ scan_wrapper_339501025136214612_366/latch_enable_in scan_wrapper_339501025136214612_367/latch_enable_in
+ scan_wrapper_339501025136214612_366/scan_select_in scan_wrapper_339501025136214612_367/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_377 scan_wrapper_339501025136214612_377/clk_in scan_wrapper_339501025136214612_378/clk_in
+ scan_wrapper_339501025136214612_377/data_in scan_wrapper_339501025136214612_378/data_in
+ scan_wrapper_339501025136214612_377/latch_enable_in scan_wrapper_339501025136214612_378/latch_enable_in
+ scan_wrapper_339501025136214612_377/scan_select_in scan_wrapper_339501025136214612_378/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341546888233747026_115 scan_wrapper_341546888233747026_115/clk_in scan_wrapper_340979268609638995_116/clk_in
+ scan_wrapper_341546888233747026_115/data_in scan_wrapper_340979268609638995_116/data_in
+ scan_wrapper_341546888233747026_115/latch_enable_in scan_wrapper_340979268609638995_116/latch_enable_in
+ scan_wrapper_341546888233747026_115/scan_select_in scan_wrapper_340979268609638995_116/scan_select_in
+ vccd1 vssd1 scan_wrapper_341546888233747026
Xscan_wrapper_339501025136214612_152 scan_wrapper_339501025136214612_152/clk_in scan_wrapper_339501025136214612_153/clk_in
+ scan_wrapper_339501025136214612_152/data_in scan_wrapper_339501025136214612_153/data_in
+ scan_wrapper_339501025136214612_152/latch_enable_in scan_wrapper_339501025136214612_153/latch_enable_in
+ scan_wrapper_339501025136214612_152/scan_select_in scan_wrapper_339501025136214612_153/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_163 scan_wrapper_339501025136214612_163/clk_in scan_wrapper_339501025136214612_164/clk_in
+ scan_wrapper_339501025136214612_163/data_in scan_wrapper_339501025136214612_164/data_in
+ scan_wrapper_339501025136214612_163/latch_enable_in scan_wrapper_339501025136214612_164/latch_enable_in
+ scan_wrapper_339501025136214612_163/scan_select_in scan_wrapper_339501025136214612_164/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_174 scan_wrapper_339501025136214612_174/clk_in scan_wrapper_339501025136214612_175/clk_in
+ scan_wrapper_339501025136214612_174/data_in scan_wrapper_339501025136214612_175/data_in
+ scan_wrapper_339501025136214612_174/latch_enable_in scan_wrapper_339501025136214612_175/latch_enable_in
+ scan_wrapper_339501025136214612_174/scan_select_in scan_wrapper_339501025136214612_175/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_196 scan_wrapper_339501025136214612_196/clk_in scan_wrapper_339501025136214612_197/clk_in
+ scan_wrapper_339501025136214612_196/data_in scan_wrapper_339501025136214612_197/data_in
+ scan_wrapper_339501025136214612_196/latch_enable_in scan_wrapper_339501025136214612_197/latch_enable_in
+ scan_wrapper_339501025136214612_196/scan_select_in scan_wrapper_339501025136214612_197/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_185 scan_wrapper_339501025136214612_185/clk_in scan_wrapper_339501025136214612_186/clk_in
+ scan_wrapper_339501025136214612_185/data_in scan_wrapper_339501025136214612_186/data_in
+ scan_wrapper_339501025136214612_185/latch_enable_in scan_wrapper_339501025136214612_186/latch_enable_in
+ scan_wrapper_339501025136214612_185/scan_select_in scan_wrapper_339501025136214612_186/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341506274933867090_93 scan_wrapper_341506274933867090_93/clk_in scan_wrapper_341449297858921043_94/clk_in
+ scan_wrapper_341506274933867090_93/data_in scan_wrapper_341449297858921043_94/data_in
+ scan_wrapper_341506274933867090_93/latch_enable_in scan_wrapper_341449297858921043_94/latch_enable_in
+ scan_wrapper_341506274933867090_93/scan_select_in scan_wrapper_341449297858921043_94/scan_select_in
+ vccd1 vssd1 scan_wrapper_341506274933867090
Xscan_wrapper_341581732833657427_126 scan_wrapper_341581732833657427_126/clk_in scan_wrapper_341457494561784402_127/clk_in
+ scan_wrapper_341581732833657427_126/data_in scan_wrapper_341457494561784402_127/data_in
+ scan_wrapper_341581732833657427_126/latch_enable_in scan_wrapper_341457494561784402_127/latch_enable_in
+ scan_wrapper_341581732833657427_126/scan_select_in scan_wrapper_341457494561784402_127/scan_select_in
+ vccd1 vssd1 scan_wrapper_341581732833657427
Xscan_wrapper_340579111348994642_30 scan_wrapper_340579111348994642_30/clk_in scan_wrapper_341224613878956628_31/clk_in
+ scan_wrapper_340579111348994642_30/data_in scan_wrapper_341224613878956628_31/data_in
+ scan_wrapper_340579111348994642_30/latch_enable_in scan_wrapper_341224613878956628_31/latch_enable_in
+ scan_wrapper_340579111348994642_30/scan_select_in scan_wrapper_341224613878956628_31/scan_select_in
+ vccd1 vssd1 scan_wrapper_340579111348994642
Xscan_wrapper_341613097060926036_135 scan_wrapper_341613097060926036_135/clk_in scan_wrapper_341614346808328788_136/clk_in
+ scan_wrapper_341613097060926036_135/data_in scan_wrapper_341614346808328788_136/data_in
+ scan_wrapper_341613097060926036_135/latch_enable_in scan_wrapper_341614346808328788_136/latch_enable_in
+ scan_wrapper_341613097060926036_135/scan_select_in scan_wrapper_341614346808328788_136/scan_select_in
+ vccd1 vssd1 scan_wrapper_341613097060926036
Xscan_wrapper_339501025136214612_378 scan_wrapper_339501025136214612_378/clk_in scan_wrapper_339501025136214612_379/clk_in
+ scan_wrapper_339501025136214612_378/data_in scan_wrapper_339501025136214612_379/data_in
+ scan_wrapper_339501025136214612_378/latch_enable_in scan_wrapper_339501025136214612_379/latch_enable_in
+ scan_wrapper_339501025136214612_378/scan_select_in scan_wrapper_339501025136214612_379/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_389 scan_wrapper_339501025136214612_389/clk_in scan_wrapper_339501025136214612_390/clk_in
+ scan_wrapper_339501025136214612_389/data_in scan_wrapper_339501025136214612_390/data_in
+ scan_wrapper_339501025136214612_389/latch_enable_in scan_wrapper_339501025136214612_390/latch_enable_in
+ scan_wrapper_339501025136214612_389/scan_select_in scan_wrapper_339501025136214612_390/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_312 scan_wrapper_339501025136214612_312/clk_in scan_wrapper_339501025136214612_313/clk_in
+ scan_wrapper_339501025136214612_312/data_in scan_wrapper_339501025136214612_313/data_in
+ scan_wrapper_339501025136214612_312/latch_enable_in scan_wrapper_339501025136214612_313/latch_enable_in
+ scan_wrapper_339501025136214612_312/scan_select_in scan_wrapper_339501025136214612_313/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_301 scan_wrapper_339501025136214612_301/clk_in scan_wrapper_339501025136214612_302/clk_in
+ scan_wrapper_339501025136214612_301/data_in scan_wrapper_339501025136214612_302/data_in
+ scan_wrapper_339501025136214612_301/latch_enable_in scan_wrapper_339501025136214612_302/latch_enable_in
+ scan_wrapper_339501025136214612_301/scan_select_in scan_wrapper_339501025136214612_302/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_323 scan_wrapper_339501025136214612_323/clk_in scan_wrapper_339501025136214612_324/clk_in
+ scan_wrapper_339501025136214612_323/data_in scan_wrapper_339501025136214612_324/data_in
+ scan_wrapper_339501025136214612_323/latch_enable_in scan_wrapper_339501025136214612_324/latch_enable_in
+ scan_wrapper_339501025136214612_323/scan_select_in scan_wrapper_339501025136214612_324/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_334 scan_wrapper_339501025136214612_334/clk_in scan_wrapper_339501025136214612_335/clk_in
+ scan_wrapper_339501025136214612_334/data_in scan_wrapper_339501025136214612_335/data_in
+ scan_wrapper_339501025136214612_334/latch_enable_in scan_wrapper_339501025136214612_335/latch_enable_in
+ scan_wrapper_339501025136214612_334/scan_select_in scan_wrapper_339501025136214612_335/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_356 scan_wrapper_339501025136214612_356/clk_in scan_wrapper_339501025136214612_357/clk_in
+ scan_wrapper_339501025136214612_356/data_in scan_wrapper_339501025136214612_357/data_in
+ scan_wrapper_339501025136214612_356/latch_enable_in scan_wrapper_339501025136214612_357/latch_enable_in
+ scan_wrapper_339501025136214612_356/scan_select_in scan_wrapper_339501025136214612_357/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_345 scan_wrapper_339501025136214612_345/clk_in scan_wrapper_339501025136214612_346/clk_in
+ scan_wrapper_339501025136214612_345/data_in scan_wrapper_339501025136214612_346/data_in
+ scan_wrapper_339501025136214612_345/latch_enable_in scan_wrapper_339501025136214612_346/latch_enable_in
+ scan_wrapper_339501025136214612_345/scan_select_in scan_wrapper_339501025136214612_346/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_367 scan_wrapper_339501025136214612_367/clk_in scan_wrapper_339501025136214612_368/clk_in
+ scan_wrapper_339501025136214612_367/data_in scan_wrapper_339501025136214612_368/data_in
+ scan_wrapper_339501025136214612_367/latch_enable_in scan_wrapper_339501025136214612_368/latch_enable_in
+ scan_wrapper_339501025136214612_367/scan_select_in scan_wrapper_339501025136214612_368/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341176884318437971_20 scan_wrapper_341176884318437971_20/clk_in scan_wrapper_341182944314917460_21/clk_in
+ scan_wrapper_341176884318437971_20/data_in scan_wrapper_341182944314917460_21/data_in
+ scan_wrapper_341176884318437971_20/latch_enable_in scan_wrapper_341182944314917460_21/latch_enable_in
+ scan_wrapper_341176884318437971_20/scan_select_in scan_wrapper_341182944314917460_21/scan_select_in
+ vccd1 vssd1 scan_wrapper_341176884318437971
Xscan_wrapper_339501025136214612_153 scan_wrapper_339501025136214612_153/clk_in scan_wrapper_339501025136214612_154/clk_in
+ scan_wrapper_339501025136214612_153/data_in scan_wrapper_339501025136214612_154/data_in
+ scan_wrapper_339501025136214612_153/latch_enable_in scan_wrapper_339501025136214612_154/latch_enable_in
+ scan_wrapper_339501025136214612_153/scan_select_in scan_wrapper_339501025136214612_154/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_164 scan_wrapper_339501025136214612_164/clk_in scan_wrapper_339501025136214612_165/clk_in
+ scan_wrapper_339501025136214612_164/data_in scan_wrapper_339501025136214612_165/data_in
+ scan_wrapper_339501025136214612_164/latch_enable_in scan_wrapper_339501025136214612_165/latch_enable_in
+ scan_wrapper_339501025136214612_164/scan_select_in scan_wrapper_339501025136214612_165/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_175 scan_wrapper_339501025136214612_175/clk_in scan_wrapper_339501025136214612_176/clk_in
+ scan_wrapper_339501025136214612_175/data_in scan_wrapper_339501025136214612_176/data_in
+ scan_wrapper_339501025136214612_175/latch_enable_in scan_wrapper_339501025136214612_176/latch_enable_in
+ scan_wrapper_339501025136214612_175/scan_select_in scan_wrapper_339501025136214612_176/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_197 scan_wrapper_339501025136214612_197/clk_in scan_wrapper_339501025136214612_198/clk_in
+ scan_wrapper_339501025136214612_197/data_in scan_wrapper_339501025136214612_198/data_in
+ scan_wrapper_339501025136214612_197/latch_enable_in scan_wrapper_339501025136214612_198/latch_enable_in
+ scan_wrapper_339501025136214612_197/scan_select_in scan_wrapper_339501025136214612_198/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_339501025136214612_186 scan_wrapper_339501025136214612_186/clk_in scan_wrapper_339501025136214612_187/clk_in
+ scan_wrapper_339501025136214612_186/data_in scan_wrapper_339501025136214612_187/data_in
+ scan_wrapper_339501025136214612_186/latch_enable_in scan_wrapper_339501025136214612_187/latch_enable_in
+ scan_wrapper_339501025136214612_186/scan_select_in scan_wrapper_339501025136214612_187/scan_select_in
+ vccd1 vssd1 scan_wrapper_339501025136214612
Xscan_wrapper_341359404107432531_59 scan_wrapper_341359404107432531_59/clk_in scan_wrapper_341315210433266259_60/clk_in
+ scan_wrapper_341359404107432531_59/data_in scan_wrapper_341315210433266259_60/data_in
+ scan_wrapper_341359404107432531_59/latch_enable_in scan_wrapper_341315210433266259_60/latch_enable_in
+ scan_wrapper_341359404107432531_59/scan_select_in scan_wrapper_341315210433266259_60/scan_select_in
+ vccd1 vssd1 scan_wrapper_341359404107432531
.ends

