// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_project_wrapper
 *
 * This wrapper enumerates all of the pins available to the
 * user for the user project.
 *
 * An example user project is provided in this wrapper.  The
 * example should be removed and replaced with the actual
 * user project.
 *
 * THIS FILE HAS BEEN GENERATED USING multi_tools_project CODEGEN
 * IF YOU NEED TO MAKE EDITS TO IT, EDIT codegen/caravel_iface_header.txt
 *
 *-------------------------------------------------------------
 */

module user_project_wrapper #(
    parameter BITS = 32
)(
`ifdef USE_POWER_PINS
    inout vdda1,       // User area 1 3.3V supply
    inout vdda2,       // User area 2 3.3V supply
    inout vssa1,       // User area 1 analog ground
    inout vssa2,       // User area 2 analog ground
    inout vccd1,       // User area 1 1.8V supply
    inout vccd2,       // User area 2 1.8v supply
    inout vssd1,       // User area 1 digital ground
    inout vssd2,       // User area 2 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // Analog (direct connection to GPIO pad---use with caution)
    // Note that analog I/O is not available on the 7 lowest-numbered
    // GPIO pads, and so the analog_io indexing is offset from the
    // GPIO indexing by 7 (also upper 2 GPIOs do not have analog_io).
    inout [`MPRJ_IO_PADS-10:0] analog_io,

    // Independent clock (on independent integer divider)
    input   user_clock2,

    // User maskable interrupt signals
    output [2:0] user_irq
);

    // start of module instantiation

    wire sc_clk_out, sc_data_out, sc_latch_out, sc_scan_out;
    wire sc_clk_in,  sc_data_in;

    scan_controller #(.NUM_DESIGNS(498)) scan_controller (
       .clk                    (wb_clk_i),
       .reset                  (wb_rst_i),
       .active_select          (io_in[20:12]),
       .inputs                 (io_in[28:21]),
       .outputs                (io_out[36:29]),
       .ready                  (io_out[37]),
       .slow_clk               (io_out[10]),
       .set_clk_div            (io_in[11]),

       .scan_clk_out           (sc_clk_out),
       .scan_clk_in            (sc_clk_in),
       .scan_data_out          (sc_data_out),
       .scan_data_in           (sc_data_in),
       .scan_select            (sc_scan_out),
       .scan_latch_en          (sc_latch_out),

       .la_scan_clk_in         (la_data_in[0]),
       .la_scan_data_in        (la_data_in[1]),
       .la_scan_data_out       (la_data_out[0]),
       .la_scan_select         (la_data_in[2]),
       .la_scan_latch_en       (la_data_in[3]),

       .driver_sel             (io_in[9:8]),

       .oeb                    (io_oeb)
    );

    // [000] https://github.com/mattvenn/wokwi_filler
    wire sw_000_clk_out, sw_000_data_out, sw_000_scan_out, sw_000_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_0 (
        .clk_in          (sc_clk_out),
        .data_in         (sc_data_out),
        .scan_select_in  (sc_scan_out),
        .latch_enable_in (sc_latch_out),
        .clk_out         (sw_000_clk_out),
        .data_out        (sw_000_data_out),
        .scan_select_out (sw_000_scan_out),
        .latch_enable_out(sw_000_latch_out)
    );

    // [001] https://github.com/mattvenn/tinytapeout_m_segments
    wire sw_001_clk_out, sw_001_data_out, sw_001_scan_out, sw_001_latch_out;
    scan_wrapper_339688086163161683 #(.NUM_IOS(8)) scan_wrapper_339688086163161683_1 (
        .clk_in          (sw_000_clk_out),
        .data_in         (sw_000_data_out),
        .scan_select_in  (sw_000_scan_out),
        .latch_enable_in (sw_000_latch_out),
        .clk_out         (sw_001_clk_out),
        .data_out        (sw_001_data_out),
        .scan_select_out (sw_001_scan_out),
        .latch_enable_out(sw_001_latch_out)
    );

    // [002] https://github.com/gregdavill/tinytapeout_spin0
    wire sw_002_clk_out, sw_002_data_out, sw_002_scan_out, sw_002_latch_out;
    scan_wrapper_340218629792465491 #(.NUM_IOS(8)) scan_wrapper_340218629792465491_2 (
        .clk_in          (sw_001_clk_out),
        .data_in         (sw_001_data_out),
        .scan_select_in  (sw_001_scan_out),
        .latch_enable_in (sw_001_latch_out),
        .clk_out         (sw_002_clk_out),
        .data_out        (sw_002_data_out),
        .scan_select_out (sw_002_scan_out),
        .latch_enable_out(sw_002_latch_out)
    );

    // [003] https://github.com/mole99/wokwi-1bit-alu
    wire sw_003_clk_out, sw_003_data_out, sw_003_scan_out, sw_003_latch_out;
    scan_wrapper_340318610245288530 #(.NUM_IOS(8)) scan_wrapper_340318610245288530_3 (
        .clk_in          (sw_002_clk_out),
        .data_in         (sw_002_data_out),
        .scan_select_in  (sw_002_scan_out),
        .latch_enable_in (sw_002_latch_out),
        .clk_out         (sw_003_clk_out),
        .data_out        (sw_003_data_out),
        .scan_select_out (sw_003_scan_out),
        .latch_enable_out(sw_003_latch_out)
    );

    // [004] https://github.com/ericsmi/tinytapeout_popcnt.git
    wire sw_004_clk_out, sw_004_data_out, sw_004_scan_out, sw_004_latch_out;
    scan_wrapper_340285391309374034 #(.NUM_IOS(8)) scan_wrapper_340285391309374034_4 (
        .clk_in          (sw_003_clk_out),
        .data_in         (sw_003_data_out),
        .scan_select_in  (sw_003_scan_out),
        .latch_enable_in (sw_003_latch_out),
        .clk_out         (sw_004_clk_out),
        .data_out        (sw_004_data_out),
        .scan_select_out (sw_004_scan_out),
        .latch_enable_out(sw_004_latch_out)
    );

    // [005] https://github.com/krasin/wokwi-guess-my-number
    wire sw_005_clk_out, sw_005_data_out, sw_005_scan_out, sw_005_latch_out;
    scan_wrapper_340661930553246290 #(.NUM_IOS(8)) scan_wrapper_340661930553246290_5 (
        .clk_in          (sw_004_clk_out),
        .data_in         (sw_004_data_out),
        .scan_select_in  (sw_004_scan_out),
        .latch_enable_in (sw_004_latch_out),
        .clk_out         (sw_005_clk_out),
        .data_out        (sw_005_data_out),
        .scan_select_out (sw_005_scan_out),
        .latch_enable_out(sw_005_latch_out)
    );

    // [006] https://github.com/johshoff/barrelshifter-wokwi-gds
    wire sw_006_clk_out, sw_006_data_out, sw_006_scan_out, sw_006_latch_out;
    scan_wrapper_341136771628663380 #(.NUM_IOS(8)) scan_wrapper_341136771628663380_6 (
        .clk_in          (sw_005_clk_out),
        .data_in         (sw_005_data_out),
        .scan_select_in  (sw_005_scan_out),
        .latch_enable_in (sw_005_latch_out),
        .clk_out         (sw_006_clk_out),
        .data_out        (sw_006_data_out),
        .scan_select_out (sw_006_scan_out),
        .latch_enable_out(sw_006_latch_out)
    );

    // [007] https://github.com/pretentious7/tinytapeout
    wire sw_007_clk_out, sw_007_data_out, sw_007_scan_out, sw_007_latch_out;
    scan_wrapper_339800239192932947 #(.NUM_IOS(8)) scan_wrapper_339800239192932947_7 (
        .clk_in          (sw_006_clk_out),
        .data_in         (sw_006_data_out),
        .scan_select_in  (sw_006_scan_out),
        .latch_enable_in (sw_006_latch_out),
        .clk_out         (sw_007_clk_out),
        .data_out        (sw_007_data_out),
        .scan_select_out (sw_007_scan_out),
        .latch_enable_out(sw_007_latch_out)
    );

    // [008] https://github.com/GuzTech/wokwi-ripple-carry-adder
    wire sw_008_clk_out, sw_008_data_out, sw_008_scan_out, sw_008_latch_out;
    scan_wrapper_341154161238213203 #(.NUM_IOS(8)) scan_wrapper_341154161238213203_8 (
        .clk_in          (sw_007_clk_out),
        .data_in         (sw_007_data_out),
        .scan_select_in  (sw_007_scan_out),
        .latch_enable_in (sw_007_latch_out),
        .clk_out         (sw_008_clk_out),
        .data_out        (sw_008_data_out),
        .scan_select_out (sw_008_scan_out),
        .latch_enable_out(sw_008_latch_out)
    );

    // [009] https://github.com/kbeckmann/tinytapeout_kbeckmann1
    wire sw_009_clk_out, sw_009_data_out, sw_009_scan_out, sw_009_latch_out;
    scan_wrapper_341159915403870803 #(.NUM_IOS(8)) scan_wrapper_341159915403870803_9 (
        .clk_in          (sw_008_clk_out),
        .data_in         (sw_008_data_out),
        .scan_select_in  (sw_008_scan_out),
        .latch_enable_in (sw_008_latch_out),
        .clk_out         (sw_009_clk_out),
        .data_out        (sw_009_data_out),
        .scan_select_out (sw_009_scan_out),
        .latch_enable_out(sw_009_latch_out)
    );

    // [010] https://github.com/H-S-S-11/tinytapeout-verilog-test
    wire sw_010_clk_out, sw_010_data_out, sw_010_scan_out, sw_010_latch_out;
    scan_wrapper_341154068332282450 #(.NUM_IOS(8)) scan_wrapper_341154068332282450_10 (
        .clk_in          (sw_009_clk_out),
        .data_in         (sw_009_data_out),
        .scan_select_in  (sw_009_scan_out),
        .latch_enable_in (sw_009_latch_out),
        .clk_out         (sw_010_clk_out),
        .data_out        (sw_010_data_out),
        .scan_select_out (sw_010_scan_out),
        .latch_enable_out(sw_010_latch_out)
    );

    // [011] https://github.com/skerr92/tinytapeout_frequency_div
    wire sw_011_clk_out, sw_011_data_out, sw_011_scan_out, sw_011_latch_out;
    scan_wrapper_341160201697624660 #(.NUM_IOS(8)) scan_wrapper_341160201697624660_11 (
        .clk_in          (sw_010_clk_out),
        .data_in         (sw_010_data_out),
        .scan_select_in  (sw_010_scan_out),
        .latch_enable_in (sw_010_latch_out),
        .clk_out         (sw_011_clk_out),
        .data_out        (sw_011_data_out),
        .scan_select_out (sw_011_scan_out),
        .latch_enable_out(sw_011_latch_out)
    );

    // [012] https://github.com/argunda/tinytapeout_dualedgedetector
    wire sw_012_clk_out, sw_012_data_out, sw_012_scan_out, sw_012_latch_out;
    scan_wrapper_341163800289870419 #(.NUM_IOS(8)) scan_wrapper_341163800289870419_12 (
        .clk_in          (sw_011_clk_out),
        .data_in         (sw_011_data_out),
        .scan_select_in  (sw_011_scan_out),
        .latch_enable_in (sw_011_latch_out),
        .clk_out         (sw_012_clk_out),
        .data_out        (sw_012_data_out),
        .scan_select_out (sw_012_scan_out),
        .latch_enable_out(sw_012_latch_out)
    );

    // [013] https://github.com/libokuohai/tinytapeout-2022-08
    wire sw_013_clk_out, sw_013_data_out, sw_013_scan_out, sw_013_latch_out;
    scan_wrapper_341160271679586899 #(.NUM_IOS(8)) scan_wrapper_341160271679586899_13 (
        .clk_in          (sw_012_clk_out),
        .data_in         (sw_012_data_out),
        .scan_select_in  (sw_012_scan_out),
        .latch_enable_in (sw_012_latch_out),
        .clk_out         (sw_013_clk_out),
        .data_out        (sw_013_data_out),
        .scan_select_out (sw_013_scan_out),
        .latch_enable_out(sw_013_latch_out)
    );

    // [014] https://github.com/jglim/tinytapeout_bcd-dec
    wire sw_014_clk_out, sw_014_data_out, sw_014_scan_out, sw_014_latch_out;
    scan_wrapper_341161378978988626 #(.NUM_IOS(8)) scan_wrapper_341161378978988626_14 (
        .clk_in          (sw_013_clk_out),
        .data_in         (sw_013_data_out),
        .scan_select_in  (sw_013_scan_out),
        .latch_enable_in (sw_013_latch_out),
        .clk_out         (sw_014_clk_out),
        .data_out        (sw_014_data_out),
        .scan_select_out (sw_014_scan_out),
        .latch_enable_out(sw_014_latch_out)
    );

    // [015] https://github.com/jglim/tinytapeout_bcd-7seg
    wire sw_015_clk_out, sw_015_data_out, sw_015_scan_out, sw_015_latch_out;
    scan_wrapper_341152580068442706 #(.NUM_IOS(8)) scan_wrapper_341152580068442706_15 (
        .clk_in          (sw_014_clk_out),
        .data_in         (sw_014_data_out),
        .scan_select_in  (sw_014_scan_out),
        .latch_enable_in (sw_014_latch_out),
        .clk_out         (sw_015_clk_out),
        .data_out        (sw_015_data_out),
        .scan_select_out (sw_015_scan_out),
        .latch_enable_out(sw_015_latch_out)
    );

    // [016] https://github.com/tkuester/wokwi-directghost
    wire sw_016_clk_out, sw_016_data_out, sw_016_scan_out, sw_016_latch_out;
    scan_wrapper_341155178824598098 #(.NUM_IOS(8)) scan_wrapper_341155178824598098_16 (
        .clk_in          (sw_015_clk_out),
        .data_in         (sw_015_data_out),
        .scan_select_in  (sw_015_scan_out),
        .latch_enable_in (sw_015_latch_out),
        .clk_out         (sw_016_clk_out),
        .data_out        (sw_016_data_out),
        .scan_select_out (sw_016_scan_out),
        .latch_enable_out(sw_016_latch_out)
    );

    // [017] https://github.com/shahzaibk23/tinytapeout-barrel-shifter
    wire sw_017_clk_out, sw_017_data_out, sw_017_scan_out, sw_017_latch_out;
    scan_wrapper_341167691532337747 #(.NUM_IOS(8)) scan_wrapper_341167691532337747_17 (
        .clk_in          (sw_016_clk_out),
        .data_in         (sw_016_data_out),
        .scan_select_in  (sw_016_scan_out),
        .latch_enable_in (sw_016_latch_out),
        .clk_out         (sw_017_clk_out),
        .data_out        (sw_017_data_out),
        .scan_select_out (sw_017_scan_out),
        .latch_enable_out(sw_017_latch_out)
    );

    // [018] https://github.com/tcptomato/tinytapeout
    wire sw_018_clk_out, sw_018_data_out, sw_018_scan_out, sw_018_latch_out;
    scan_wrapper_341178154799333971 #(.NUM_IOS(8)) scan_wrapper_341178154799333971_18 (
        .clk_in          (sw_017_clk_out),
        .data_in         (sw_017_data_out),
        .scan_select_in  (sw_017_scan_out),
        .latch_enable_in (sw_017_latch_out),
        .clk_out         (sw_018_clk_out),
        .data_out        (sw_018_data_out),
        .scan_select_out (sw_018_scan_out),
        .latch_enable_out(sw_018_latch_out)
    );

    // [019] https://github.com/DaveyPocket/chaser
    wire sw_019_clk_out, sw_019_data_out, sw_019_scan_out, sw_019_latch_out;
    scan_wrapper_341178481588044372 #(.NUM_IOS(8)) scan_wrapper_341178481588044372_19 (
        .clk_in          (sw_018_clk_out),
        .data_in         (sw_018_data_out),
        .scan_select_in  (sw_018_scan_out),
        .latch_enable_in (sw_018_latch_out),
        .clk_out         (sw_019_clk_out),
        .data_out        (sw_019_data_out),
        .scan_select_out (sw_019_scan_out),
        .latch_enable_out(sw_019_latch_out)
    );

    // [020] https://github.com/GuzTech/tinytapeout-4x4-multiplier
    wire sw_020_clk_out, sw_020_data_out, sw_020_scan_out, sw_020_latch_out;
    scan_wrapper_341176884318437971 #(.NUM_IOS(8)) scan_wrapper_341176884318437971_20 (
        .clk_in          (sw_019_clk_out),
        .data_in         (sw_019_data_out),
        .scan_select_in  (sw_019_scan_out),
        .latch_enable_in (sw_019_latch_out),
        .clk_out         (sw_020_clk_out),
        .data_out        (sw_020_data_out),
        .scan_select_out (sw_020_scan_out),
        .latch_enable_out(sw_020_latch_out)
    );

    // [021] https://github.com/derhexenmeister/tinytapeout_nco
    wire sw_021_clk_out, sw_021_data_out, sw_021_scan_out, sw_021_latch_out;
    scan_wrapper_341182944314917460 #(.NUM_IOS(8)) scan_wrapper_341182944314917460_21 (
        .clk_in          (sw_020_clk_out),
        .data_in         (sw_020_data_out),
        .scan_select_in  (sw_020_scan_out),
        .latch_enable_in (sw_020_latch_out),
        .clk_out         (sw_021_clk_out),
        .data_out        (sw_021_data_out),
        .scan_select_out (sw_021_scan_out),
        .latch_enable_out(sw_021_latch_out)
    );

    // [022] https://github.com/mbalestrini/tinytapeout_rgb_lut_test
    wire sw_022_clk_out, sw_022_data_out, sw_022_scan_out, sw_022_latch_out;
    scan_wrapper_341188777753969234 #(.NUM_IOS(8)) scan_wrapper_341188777753969234_22 (
        .clk_in          (sw_021_clk_out),
        .data_in         (sw_021_data_out),
        .scan_select_in  (sw_021_scan_out),
        .latch_enable_in (sw_021_latch_out),
        .clk_out         (sw_022_clk_out),
        .data_out        (sw_022_data_out),
        .scan_select_out (sw_022_scan_out),
        .latch_enable_out(sw_022_latch_out)
    );

    // [023] https://github.com/derhexenmeister/tinytapeout_updwnbcd
    wire sw_023_clk_out, sw_023_data_out, sw_023_scan_out, sw_023_latch_out;
    scan_wrapper_341194143598379604 #(.NUM_IOS(8)) scan_wrapper_341194143598379604_23 (
        .clk_in          (sw_022_clk_out),
        .data_in         (sw_022_data_out),
        .scan_select_in  (sw_022_scan_out),
        .latch_enable_in (sw_022_latch_out),
        .clk_out         (sw_023_clk_out),
        .data_out        (sw_023_data_out),
        .scan_select_out (sw_023_scan_out),
        .latch_enable_out(sw_023_latch_out)
    );

    // [024] https://github.com/bradysalz/pll_tiny_tapeout_demo
    wire sw_024_clk_out, sw_024_data_out, sw_024_scan_out, sw_024_latch_out;
    scan_wrapper_341205508016833108 #(.NUM_IOS(8)) scan_wrapper_341205508016833108_24 (
        .clk_in          (sw_023_clk_out),
        .data_in         (sw_023_data_out),
        .scan_select_in  (sw_023_scan_out),
        .latch_enable_in (sw_023_latch_out),
        .clk_out         (sw_024_clk_out),
        .data_out        (sw_024_data_out),
        .scan_select_out (sw_024_scan_out),
        .latch_enable_out(sw_024_latch_out)
    );

    // [025] https://github.com/pramitpal/tinytapeout_pramit
    wire sw_025_clk_out, sw_025_data_out, sw_025_scan_out, sw_025_latch_out;
    scan_wrapper_341162950004834900 #(.NUM_IOS(8)) scan_wrapper_341162950004834900_25 (
        .clk_in          (sw_024_clk_out),
        .data_in         (sw_024_data_out),
        .scan_select_in  (sw_024_scan_out),
        .latch_enable_in (sw_024_latch_out),
        .clk_out         (sw_025_clk_out),
        .data_out        (sw_025_data_out),
        .scan_select_out (sw_025_scan_out),
        .latch_enable_out(sw_025_latch_out)
    );

    // [026] https://github.com/gregdavill/tinytapeout-verilog-fifo
    wire sw_026_clk_out, sw_026_data_out, sw_026_scan_out, sw_026_latch_out;
    scan_wrapper_341202178192441940 #(.NUM_IOS(8)) scan_wrapper_341202178192441940_26 (
        .clk_in          (sw_025_clk_out),
        .data_in         (sw_025_data_out),
        .scan_select_in  (sw_025_scan_out),
        .latch_enable_in (sw_025_latch_out),
        .clk_out         (sw_026_clk_out),
        .data_out        (sw_026_data_out),
        .scan_select_out (sw_026_scan_out),
        .latch_enable_out(sw_026_latch_out)
    );

    // [027] https://github.com/gregdavill/tinytapeout-wokwi-74x1G00
    wire sw_027_clk_out, sw_027_data_out, sw_027_scan_out, sw_027_latch_out;
    scan_wrapper_341191836498395731 #(.NUM_IOS(8)) scan_wrapper_341191836498395731_27 (
        .clk_in          (sw_026_clk_out),
        .data_in         (sw_026_data_out),
        .scan_select_in  (sw_026_scan_out),
        .latch_enable_in (sw_026_latch_out),
        .clk_out         (sw_027_clk_out),
        .data_out        (sw_027_data_out),
        .scan_select_out (sw_027_scan_out),
        .latch_enable_out(sw_027_latch_out)
    );

    // [028] https://github.com/gregdavill/tinytapeout-wokwi-74x1G02
    wire sw_028_clk_out, sw_028_data_out, sw_028_scan_out, sw_028_latch_out;
    scan_wrapper_341192113929585235 #(.NUM_IOS(8)) scan_wrapper_341192113929585235_28 (
        .clk_in          (sw_027_clk_out),
        .data_in         (sw_027_data_out),
        .scan_select_in  (sw_027_scan_out),
        .latch_enable_in (sw_027_latch_out),
        .clk_out         (sw_028_clk_out),
        .data_out        (sw_028_data_out),
        .scan_select_out (sw_028_scan_out),
        .latch_enable_out(sw_028_latch_out)
    );

    // [029] https://github.com/gregdavill/tinytapeout-wokwi-74xG198
    wire sw_029_clk_out, sw_029_data_out, sw_029_scan_out, sw_029_latch_out;
    scan_wrapper_341192621088047698 #(.NUM_IOS(8)) scan_wrapper_341192621088047698_29 (
        .clk_in          (sw_028_clk_out),
        .data_in         (sw_028_data_out),
        .scan_select_in  (sw_028_scan_out),
        .latch_enable_in (sw_028_latch_out),
        .clk_out         (sw_029_clk_out),
        .data_out        (sw_029_data_out),
        .scan_select_out (sw_029_scan_out),
        .latch_enable_out(sw_029_latch_out)
    );

    // [030] https://github.com/gregdavill/tinytapeout-verilog-7seg-clock
    wire sw_030_clk_out, sw_030_data_out, sw_030_scan_out, sw_030_latch_out;
    scan_wrapper_340579111348994642 #(.NUM_IOS(8)) scan_wrapper_340579111348994642_30 (
        .clk_in          (sw_029_clk_out),
        .data_in         (sw_029_data_out),
        .scan_select_in  (sw_029_scan_out),
        .latch_enable_in (sw_029_latch_out),
        .clk_out         (sw_030_clk_out),
        .data_out        (sw_030_data_out),
        .scan_select_out (sw_030_scan_out),
        .latch_enable_out(sw_030_latch_out)
    );

    // [031] https://github.com/alanvgreen/tinytapeout4bitadder
    wire sw_031_clk_out, sw_031_data_out, sw_031_scan_out, sw_031_latch_out;
    scan_wrapper_341224613878956628 #(.NUM_IOS(8)) scan_wrapper_341224613878956628_31 (
        .clk_in          (sw_030_clk_out),
        .data_in         (sw_030_data_out),
        .scan_select_in  (sw_030_scan_out),
        .latch_enable_in (sw_030_latch_out),
        .clk_out         (sw_031_clk_out),
        .data_out        (sw_031_data_out),
        .scan_select_out (sw_031_scan_out),
        .latch_enable_out(sw_031_latch_out)
    );

    // [032] https://github.com/benlaurie/twistedringcounter
    wire sw_032_clk_out, sw_032_data_out, sw_032_scan_out, sw_032_latch_out;
    scan_wrapper_341235973870322258 #(.NUM_IOS(8)) scan_wrapper_341235973870322258_32 (
        .clk_in          (sw_031_clk_out),
        .data_in         (sw_031_data_out),
        .scan_select_in  (sw_031_scan_out),
        .latch_enable_in (sw_031_latch_out),
        .clk_out         (sw_032_clk_out),
        .data_out        (sw_032_data_out),
        .scan_select_out (sw_032_scan_out),
        .latch_enable_out(sw_032_latch_out)
    );

    // [033] https://github.com/sureshsugumar/tinytapeout_counter
    wire sw_033_clk_out, sw_033_data_out, sw_033_scan_out, sw_033_latch_out;
    scan_wrapper_341235575572922964 #(.NUM_IOS(8)) scan_wrapper_341235575572922964_33 (
        .clk_in          (sw_032_clk_out),
        .data_in         (sw_032_data_out),
        .scan_select_in  (sw_032_scan_out),
        .latch_enable_in (sw_032_latch_out),
        .clk_out         (sw_033_clk_out),
        .data_out        (sw_033_data_out),
        .scan_select_out (sw_033_scan_out),
        .latch_enable_out(sw_033_latch_out)
    );

    // [034] https://github.com/daniestevez/tinytapeout-verilog
    wire sw_034_clk_out, sw_034_data_out, sw_034_scan_out, sw_034_latch_out;
    scan_wrapper_341164910646919762 #(.NUM_IOS(8)) scan_wrapper_341164910646919762_34 (
        .clk_in          (sw_033_clk_out),
        .data_in         (sw_033_data_out),
        .scan_select_in  (sw_033_scan_out),
        .latch_enable_in (sw_033_latch_out),
        .clk_out         (sw_034_clk_out),
        .data_out        (sw_034_data_out),
        .scan_select_out (sw_034_scan_out),
        .latch_enable_out(sw_034_latch_out)
    );

    // [035] https://github.com/pkuligowski/tinytapeout_tmr
    wire sw_035_clk_out, sw_035_data_out, sw_035_scan_out, sw_035_latch_out;
    scan_wrapper_341233739099013714 #(.NUM_IOS(8)) scan_wrapper_341233739099013714_35 (
        .clk_in          (sw_034_clk_out),
        .data_in         (sw_034_data_out),
        .scan_select_in  (sw_034_scan_out),
        .latch_enable_in (sw_034_latch_out),
        .clk_out         (sw_035_clk_out),
        .data_out        (sw_035_data_out),
        .scan_select_out (sw_035_scan_out),
        .latch_enable_out(sw_035_latch_out)
    );

    // [036] https://github.com/chiplet/tinytapeout-snake
    wire sw_036_clk_out, sw_036_data_out, sw_036_scan_out, sw_036_latch_out;
    scan_wrapper_341240110454407762 #(.NUM_IOS(8)) scan_wrapper_341240110454407762_36 (
        .clk_in          (sw_035_clk_out),
        .data_in         (sw_035_data_out),
        .scan_select_in  (sw_035_scan_out),
        .latch_enable_in (sw_035_latch_out),
        .clk_out         (sw_036_clk_out),
        .data_out        (sw_036_data_out),
        .scan_select_out (sw_036_scan_out),
        .latch_enable_out(sw_036_latch_out)
    );

    // [037] https://github.com/derhexenmeister/tinytapeout_pwm
    wire sw_037_clk_out, sw_037_data_out, sw_037_scan_out, sw_037_latch_out;
    scan_wrapper_341264068701586004 #(.NUM_IOS(8)) scan_wrapper_341264068701586004_37 (
        .clk_in          (sw_036_clk_out),
        .data_in         (sw_036_data_out),
        .scan_select_in  (sw_036_scan_out),
        .latch_enable_in (sw_036_latch_out),
        .clk_out         (sw_037_clk_out),
        .data_out        (sw_037_data_out),
        .scan_select_out (sw_037_scan_out),
        .latch_enable_out(sw_037_latch_out)
    );

    // [038] https://github.com/raha96/tinycharacters-locked
    wire sw_038_clk_out, sw_038_data_out, sw_038_scan_out, sw_038_latch_out;
    scan_wrapper_341164228775772755 #(.NUM_IOS(8)) scan_wrapper_341164228775772755_38 (
        .clk_in          (sw_037_clk_out),
        .data_in         (sw_037_data_out),
        .scan_select_in  (sw_037_scan_out),
        .latch_enable_in (sw_037_latch_out),
        .clk_out         (sw_038_clk_out),
        .data_out        (sw_038_data_out),
        .scan_select_out (sw_038_scan_out),
        .latch_enable_out(sw_038_latch_out)
    );

    // [039] https://github.com/nathancheek/tinytapeout-loop
    wire sw_039_clk_out, sw_039_data_out, sw_039_scan_out, sw_039_latch_out;
    scan_wrapper_341262321634509394 #(.NUM_IOS(8)) scan_wrapper_341262321634509394_39 (
        .clk_in          (sw_038_clk_out),
        .data_in         (sw_038_data_out),
        .scan_select_in  (sw_038_scan_out),
        .latch_enable_in (sw_038_latch_out),
        .clk_out         (sw_039_clk_out),
        .data_out        (sw_039_data_out),
        .scan_select_out (sw_039_scan_out),
        .latch_enable_out(sw_039_latch_out)
    );

    // [040] https://github.com/andars/universal-turing-machine-w5s8
    wire sw_040_clk_out, sw_040_data_out, sw_040_scan_out, sw_040_latch_out;
    scan_wrapper_341174563322724948 #(.NUM_IOS(8)) scan_wrapper_341174563322724948_40 (
        .clk_in          (sw_039_clk_out),
        .data_in         (sw_039_data_out),
        .scan_select_in  (sw_039_scan_out),
        .latch_enable_in (sw_039_latch_out),
        .clk_out         (sw_040_clk_out),
        .data_out        (sw_040_data_out),
        .scan_select_out (sw_040_scan_out),
        .latch_enable_out(sw_040_latch_out)
    );

    // [041] https://github.com/vmunoz82/tinytapeout_euler1
    wire sw_041_clk_out, sw_041_data_out, sw_041_scan_out, sw_041_latch_out;
    scan_wrapper_341271902949474898 #(.NUM_IOS(8)) scan_wrapper_341271902949474898_41 (
        .clk_in          (sw_040_clk_out),
        .data_in         (sw_040_data_out),
        .scan_select_in  (sw_040_scan_out),
        .latch_enable_in (sw_040_latch_out),
        .clk_out         (sw_041_clk_out),
        .data_out        (sw_041_data_out),
        .scan_select_out (sw_041_scan_out),
        .latch_enable_out(sw_041_latch_out)
    );

    // [042] https://github.com/mikenet213/mikenet213-tt1-verilog
    wire sw_042_clk_out, sw_042_data_out, sw_042_scan_out, sw_042_latch_out;
    scan_wrapper_bc4d7220e4fdbf20a574d56ea112a8e1 #(.NUM_IOS(8)) scan_wrapper_bc4d7220e4fdbf20a574d56ea112a8e1_42 (
        .clk_in          (sw_041_clk_out),
        .data_in         (sw_041_data_out),
        .scan_select_in  (sw_041_scan_out),
        .latch_enable_in (sw_041_latch_out),
        .clk_out         (sw_042_clk_out),
        .data_out        (sw_042_data_out),
        .scan_select_out (sw_042_scan_out),
        .latch_enable_out(sw_042_latch_out)
    );

    // [043] https://github.com/veremenko-y/tinytapeout-ue14500
    wire sw_043_clk_out, sw_043_data_out, sw_043_scan_out, sw_043_latch_out;
    scan_wrapper_341178296293130834 #(.NUM_IOS(8)) scan_wrapper_341178296293130834_43 (
        .clk_in          (sw_042_clk_out),
        .data_in         (sw_042_data_out),
        .scan_select_in  (sw_042_scan_out),
        .latch_enable_in (sw_042_latch_out),
        .clk_out         (sw_043_clk_out),
        .data_out        (sw_043_data_out),
        .scan_select_out (sw_043_scan_out),
        .latch_enable_out(sw_043_latch_out)
    );

    // [044] https://github.com/mikenet213/mikenet213-tt2-verilog
    wire sw_044_clk_out, sw_044_data_out, sw_044_scan_out, sw_044_latch_out;
    scan_wrapper_1f985e14df1ed789231bb6e0189d6e39 #(.NUM_IOS(8)) scan_wrapper_1f985e14df1ed789231bb6e0189d6e39_44 (
        .clk_in          (sw_043_clk_out),
        .data_in         (sw_043_data_out),
        .scan_select_in  (sw_043_scan_out),
        .latch_enable_in (sw_043_latch_out),
        .clk_out         (sw_044_clk_out),
        .data_out        (sw_044_data_out),
        .scan_select_out (sw_044_scan_out),
        .latch_enable_out(sw_044_latch_out)
    );

    // [045] https://github.com/aiunderstand/tinytapeout_asyncbinterconvcomp.git
    wire sw_045_clk_out, sw_045_data_out, sw_045_scan_out, sw_045_latch_out;
    scan_wrapper_341277789473735250 #(.NUM_IOS(8)) scan_wrapper_341277789473735250_45 (
        .clk_in          (sw_044_clk_out),
        .data_in         (sw_044_data_out),
        .scan_select_in  (sw_044_scan_out),
        .latch_enable_in (sw_044_latch_out),
        .clk_out         (sw_045_clk_out),
        .data_out        (sw_045_data_out),
        .scan_select_out (sw_045_scan_out),
        .latch_enable_out(sw_045_latch_out)
    );

    // [046] https://github.com/smunaut/tinytapeout-fifo
    wire sw_046_clk_out, sw_046_data_out, sw_046_scan_out, sw_046_latch_out;
    scan_wrapper_341263346544149074 #(.NUM_IOS(8)) scan_wrapper_341263346544149074_46 (
        .clk_in          (sw_045_clk_out),
        .data_in         (sw_045_data_out),
        .scan_select_in  (sw_045_scan_out),
        .latch_enable_in (sw_045_latch_out),
        .clk_out         (sw_046_clk_out),
        .data_out        (sw_046_data_out),
        .scan_select_out (sw_046_scan_out),
        .latch_enable_out(sw_046_latch_out)
    );

    // [047] https://github.com/nwtechguy/tinytapeout_BCD_counter
    wire sw_047_clk_out, sw_047_data_out, sw_047_scan_out, sw_047_latch_out;
    scan_wrapper_341296149788885588 #(.NUM_IOS(8)) scan_wrapper_341296149788885588_47 (
        .clk_in          (sw_046_clk_out),
        .data_in         (sw_046_data_out),
        .scan_select_in  (sw_046_scan_out),
        .latch_enable_in (sw_046_latch_out),
        .clk_out         (sw_047_clk_out),
        .data_out        (sw_047_data_out),
        .scan_select_out (sw_047_scan_out),
        .latch_enable_out(sw_047_latch_out)
    );

    // [048] https://github.com/kambadur/bcd_to_7seg
    wire sw_048_clk_out, sw_048_data_out, sw_048_scan_out, sw_048_latch_out;
    scan_wrapper_341332847867462227 #(.NUM_IOS(8)) scan_wrapper_341332847867462227_48 (
        .clk_in          (sw_047_clk_out),
        .data_in         (sw_047_data_out),
        .scan_select_in  (sw_047_scan_out),
        .latch_enable_in (sw_047_latch_out),
        .clk_out         (sw_048_clk_out),
        .data_out        (sw_048_data_out),
        .scan_select_out (sw_048_scan_out),
        .latch_enable_out(sw_048_latch_out)
    );

    // [049] https://github.com/bieganski/tinytapeout_bieganski
    wire sw_049_clk_out, sw_049_data_out, sw_049_scan_out, sw_049_latch_out;
    scan_wrapper_341337976625693266 #(.NUM_IOS(8)) scan_wrapper_341337976625693266_49 (
        .clk_in          (sw_048_clk_out),
        .data_in         (sw_048_data_out),
        .scan_select_in  (sw_048_scan_out),
        .latch_enable_in (sw_048_latch_out),
        .clk_out         (sw_049_clk_out),
        .data_out        (sw_049_data_out),
        .scan_select_out (sw_049_scan_out),
        .latch_enable_out(sw_049_latch_out)
    );

    // [050] https://github.com/TomKeddie/tinytapeout-2022-1
    wire sw_050_clk_out, sw_050_data_out, sw_050_scan_out, sw_050_latch_out;
    scan_wrapper_341339883600609876 #(.NUM_IOS(8)) scan_wrapper_341339883600609876_50 (
        .clk_in          (sw_049_clk_out),
        .data_in         (sw_049_data_out),
        .scan_select_in  (sw_049_scan_out),
        .latch_enable_in (sw_049_latch_out),
        .clk_out         (sw_050_clk_out),
        .data_out        (sw_050_data_out),
        .scan_select_out (sw_050_scan_out),
        .latch_enable_out(sw_050_latch_out)
    );

    // [051] https://github.com/r-a-hoggarth/tinytapeGaloisLFSR
    wire sw_051_clk_out, sw_051_data_out, sw_051_scan_out, sw_051_latch_out;
    scan_wrapper_341344337258349139 #(.NUM_IOS(8)) scan_wrapper_341344337258349139_51 (
        .clk_in          (sw_050_clk_out),
        .data_in         (sw_050_data_out),
        .scan_select_in  (sw_050_scan_out),
        .latch_enable_in (sw_050_latch_out),
        .clk_out         (sw_051_clk_out),
        .data_out        (sw_051_data_out),
        .scan_select_out (sw_051_scan_out),
        .latch_enable_out(sw_051_latch_out)
    );

    // [052] https://github.com/adamgreig/tinytapeout-prn
    wire sw_052_clk_out, sw_052_data_out, sw_052_scan_out, sw_052_latch_out;
    scan_wrapper_341342096033055316 #(.NUM_IOS(8)) scan_wrapper_341342096033055316_52 (
        .clk_in          (sw_051_clk_out),
        .data_in         (sw_051_data_out),
        .scan_select_in  (sw_051_scan_out),
        .latch_enable_in (sw_051_latch_out),
        .clk_out         (sw_052_clk_out),
        .data_out        (sw_052_data_out),
        .scan_select_out (sw_052_scan_out),
        .latch_enable_out(sw_052_latch_out)
    );

    // [053] https://github.com/ianloic/tinytapeout-1
    wire sw_053_clk_out, sw_053_data_out, sw_053_scan_out, sw_053_latch_out;
    scan_wrapper_341259651269001812 #(.NUM_IOS(8)) scan_wrapper_341259651269001812_53 (
        .clk_in          (sw_052_clk_out),
        .data_in         (sw_052_data_out),
        .scan_select_in  (sw_052_scan_out),
        .latch_enable_in (sw_052_latch_out),
        .clk_out         (sw_053_clk_out),
        .data_out        (sw_053_data_out),
        .scan_select_out (sw_053_scan_out),
        .latch_enable_out(sw_053_latch_out)
    );

    // [054] https://github.com/sad-electronics/tinytapeout-clock-divider-asic
    wire sw_054_clk_out, sw_054_data_out, sw_054_scan_out, sw_054_latch_out;
    scan_wrapper_341353928049295956 #(.NUM_IOS(8)) scan_wrapper_341353928049295956_54 (
        .clk_in          (sw_053_clk_out),
        .data_in         (sw_053_data_out),
        .scan_select_in  (sw_053_scan_out),
        .latch_enable_in (sw_053_latch_out),
        .clk_out         (sw_054_clk_out),
        .data_out        (sw_054_data_out),
        .scan_select_out (sw_054_scan_out),
        .latch_enable_out(sw_054_latch_out)
    );

    // [055] https://github.com/gatecat/tinytapeout-lutram-test
    wire sw_055_clk_out, sw_055_data_out, sw_055_scan_out, sw_055_latch_out;
    scan_wrapper_341353780122485332 #(.NUM_IOS(8)) scan_wrapper_341353780122485332_55 (
        .clk_in          (sw_054_clk_out),
        .data_in         (sw_054_data_out),
        .scan_select_in  (sw_054_scan_out),
        .latch_enable_in (sw_054_latch_out),
        .clk_out         (sw_055_clk_out),
        .data_out        (sw_055_data_out),
        .scan_select_out (sw_055_scan_out),
        .latch_enable_out(sw_055_latch_out)
    );

    // [056] https://github.com/tommythorn/tinytapeout-4-bit-cpu
    wire sw_056_clk_out, sw_056_data_out, sw_056_scan_out, sw_056_latch_out;
    scan_wrapper_341193419111006803 #(.NUM_IOS(8)) scan_wrapper_341193419111006803_56 (
        .clk_in          (sw_055_clk_out),
        .data_in         (sw_055_data_out),
        .scan_select_in  (sw_055_scan_out),
        .latch_enable_in (sw_055_latch_out),
        .clk_out         (sw_056_clk_out),
        .data_out        (sw_056_data_out),
        .scan_select_out (sw_056_scan_out),
        .latch_enable_out(sw_056_latch_out)
    );

    // [057] https://github.com/wokwi/tt-game-of-life-cell-popcnt
    wire sw_057_clk_out, sw_057_data_out, sw_057_scan_out, sw_057_latch_out;
    scan_wrapper_341266732010177108 #(.NUM_IOS(8)) scan_wrapper_341266732010177108_57 (
        .clk_in          (sw_056_clk_out),
        .data_in         (sw_056_data_out),
        .scan_select_in  (sw_056_scan_out),
        .latch_enable_in (sw_056_latch_out),
        .clk_out         (sw_057_clk_out),
        .data_out        (sw_057_data_out),
        .scan_select_out (sw_057_scan_out),
        .latch_enable_out(sw_057_latch_out)
    );

    // [058] https://github.com/gatecat/tinytapeout-srlut-test
    wire sw_058_clk_out, sw_058_data_out, sw_058_scan_out, sw_058_latch_out;
    scan_wrapper_341353777861755476 #(.NUM_IOS(8)) scan_wrapper_341353777861755476_58 (
        .clk_in          (sw_057_clk_out),
        .data_in         (sw_057_data_out),
        .scan_select_in  (sw_057_scan_out),
        .latch_enable_in (sw_057_latch_out),
        .clk_out         (sw_058_clk_out),
        .data_out        (sw_058_data_out),
        .scan_select_out (sw_058_scan_out),
        .latch_enable_out(sw_058_latch_out)
    );

    // [059] https://github.com/AdDraw/tinytapeout_demo
    wire sw_059_clk_out, sw_059_data_out, sw_059_scan_out, sw_059_latch_out;
    scan_wrapper_341359404107432531 #(.NUM_IOS(8)) scan_wrapper_341359404107432531_59 (
        .clk_in          (sw_058_clk_out),
        .data_in         (sw_058_data_out),
        .scan_select_in  (sw_058_scan_out),
        .latch_enable_in (sw_058_latch_out),
        .clk_out         (sw_059_clk_out),
        .data_out        (sw_059_data_out),
        .scan_select_out (sw_059_scan_out),
        .latch_enable_out(sw_059_latch_out)
    );

    // [060] https://github.com/cpldcpu/tinydice
    wire sw_060_clk_out, sw_060_data_out, sw_060_scan_out, sw_060_latch_out;
    scan_wrapper_341315210433266259 #(.NUM_IOS(8)) scan_wrapper_341315210433266259_60 (
        .clk_in          (sw_059_clk_out),
        .data_in         (sw_059_data_out),
        .scan_select_in  (sw_059_scan_out),
        .latch_enable_in (sw_059_latch_out),
        .clk_out         (sw_060_clk_out),
        .data_out        (sw_060_data_out),
        .scan_select_out (sw_060_scan_out),
        .latch_enable_out(sw_060_latch_out)
    );

    // [061] https://github.com/cpldcpu/tinytapeout_mcpu6bit
    wire sw_061_clk_out, sw_061_data_out, sw_061_scan_out, sw_061_latch_out;
    scan_wrapper_341364381657858642 #(.NUM_IOS(8)) scan_wrapper_341364381657858642_61 (
        .clk_in          (sw_060_clk_out),
        .data_in         (sw_060_data_out),
        .scan_select_in  (sw_060_scan_out),
        .latch_enable_in (sw_060_latch_out),
        .clk_out         (sw_061_clk_out),
        .data_out        (sw_061_data_out),
        .scan_select_out (sw_061_scan_out),
        .latch_enable_out(sw_061_latch_out)
    );

    // [062] https://github.com/azzeloof/tinytapeout-counter
    wire sw_062_clk_out, sw_062_data_out, sw_062_scan_out, sw_062_latch_out;
    scan_wrapper_341279123277087315 #(.NUM_IOS(8)) scan_wrapper_341279123277087315_62 (
        .clk_in          (sw_061_clk_out),
        .data_in         (sw_061_data_out),
        .scan_select_in  (sw_061_scan_out),
        .latch_enable_in (sw_061_latch_out),
        .clk_out         (sw_062_clk_out),
        .data_out        (sw_062_data_out),
        .scan_select_out (sw_062_scan_out),
        .latch_enable_out(sw_062_latch_out)
    );

    // [063] https://github.com/mattvenn/tinytapeout-341802655228625490
    wire sw_063_clk_out, sw_063_data_out, sw_063_scan_out, sw_063_latch_out;
    scan_wrapper_341802655228625490 #(.NUM_IOS(8)) scan_wrapper_341802655228625490_63 (
        .clk_in          (sw_062_clk_out),
        .data_in         (sw_062_data_out),
        .scan_select_in  (sw_062_scan_out),
        .latch_enable_in (sw_062_latch_out),
        .clk_out         (sw_063_clk_out),
        .data_out        (sw_063_data_out),
        .scan_select_out (sw_063_scan_out),
        .latch_enable_out(sw_063_latch_out)
    );

    // [064] https://github.com/mwelling/led-blaster
    wire sw_064_clk_out, sw_064_data_out, sw_064_scan_out, sw_064_latch_out;
    scan_wrapper_341382703379120723 #(.NUM_IOS(8)) scan_wrapper_341382703379120723_64 (
        .clk_in          (sw_063_clk_out),
        .data_in         (sw_063_data_out),
        .scan_select_in  (sw_063_scan_out),
        .latch_enable_in (sw_063_latch_out),
        .clk_out         (sw_064_clk_out),
        .data_out        (sw_064_data_out),
        .scan_select_out (sw_064_scan_out),
        .latch_enable_out(sw_064_latch_out)
    );

    // [065] https://github.com/mwelling/figure-8
    wire sw_065_clk_out, sw_065_data_out, sw_065_scan_out, sw_065_latch_out;
    scan_wrapper_341389786199622227 #(.NUM_IOS(8)) scan_wrapper_341389786199622227_65 (
        .clk_in          (sw_064_clk_out),
        .data_in         (sw_064_data_out),
        .scan_select_in  (sw_064_scan_out),
        .latch_enable_in (sw_064_latch_out),
        .clk_out         (sw_065_clk_out),
        .data_out        (sw_065_data_out),
        .scan_select_out (sw_065_scan_out),
        .latch_enable_out(sw_065_latch_out)
    );

    // [066] https://github.com/gatecat/tinytapeout-fpga-test
    wire sw_066_clk_out, sw_066_data_out, sw_066_scan_out, sw_066_latch_out;
    scan_wrapper_341404507891040852 #(.NUM_IOS(8)) scan_wrapper_341404507891040852_66 (
        .clk_in          (sw_065_clk_out),
        .data_in         (sw_065_data_out),
        .scan_select_in  (sw_065_scan_out),
        .latch_enable_in (sw_065_latch_out),
        .clk_out         (sw_066_clk_out),
        .data_out        (sw_066_data_out),
        .scan_select_out (sw_066_scan_out),
        .latch_enable_out(sw_066_latch_out)
    );

    // [067] https://github.com/cfib/trafficlight-fsm
    wire sw_067_clk_out, sw_067_data_out, sw_067_scan_out, sw_067_latch_out;
    scan_wrapper_341410909669818963 #(.NUM_IOS(8)) scan_wrapper_341410909669818963_67 (
        .clk_in          (sw_066_clk_out),
        .data_in         (sw_066_data_out),
        .scan_select_in  (sw_066_scan_out),
        .latch_enable_in (sw_066_latch_out),
        .clk_out         (sw_067_clk_out),
        .data_out        (sw_067_data_out),
        .scan_select_out (sw_067_scan_out),
        .latch_enable_out(sw_067_latch_out)
    );

    // [068] https://github.com/clj/tinytapeout-verilog-7seg-figure-eight
    wire sw_068_clk_out, sw_068_data_out, sw_068_scan_out, sw_068_latch_out;
    scan_wrapper_341063825089364563 #(.NUM_IOS(8)) scan_wrapper_341063825089364563_68 (
        .clk_in          (sw_067_clk_out),
        .data_in         (sw_067_data_out),
        .scan_select_in  (sw_067_scan_out),
        .latch_enable_in (sw_067_latch_out),
        .clk_out         (sw_068_clk_out),
        .data_out        (sw_068_data_out),
        .scan_select_out (sw_068_scan_out),
        .latch_enable_out(sw_068_latch_out)
    );

    // [069] https://github.com/smunaut/tinytapeout-misc-1
    wire sw_069_clk_out, sw_069_data_out, sw_069_scan_out, sw_069_latch_out;
    scan_wrapper_341174480471589458 #(.NUM_IOS(8)) scan_wrapper_341174480471589458_69 (
        .clk_in          (sw_068_clk_out),
        .data_in         (sw_068_data_out),
        .scan_select_in  (sw_068_scan_out),
        .latch_enable_in (sw_068_latch_out),
        .clk_out         (sw_069_clk_out),
        .data_out        (sw_069_data_out),
        .scan_select_out (sw_069_scan_out),
        .latch_enable_out(sw_069_latch_out)
    );

    // [070] https://github.com/regymm/tinytapeout-funnyblinky
    wire sw_070_clk_out, sw_070_data_out, sw_070_scan_out, sw_070_latch_out;
    scan_wrapper_341419328215712339 #(.NUM_IOS(8)) scan_wrapper_341419328215712339_70 (
        .clk_in          (sw_069_clk_out),
        .data_in         (sw_069_data_out),
        .scan_select_in  (sw_069_scan_out),
        .latch_enable_in (sw_069_latch_out),
        .clk_out         (sw_070_clk_out),
        .data_out        (sw_070_data_out),
        .scan_select_out (sw_070_scan_out),
        .latch_enable_out(sw_070_latch_out)
    );

    // [071] https://github.com/Sirawit7205/tinytapeout-2G57-2G58
    wire sw_071_clk_out, sw_071_data_out, sw_071_scan_out, sw_071_latch_out;
    scan_wrapper_341431339142087251 #(.NUM_IOS(8)) scan_wrapper_341431339142087251_71 (
        .clk_in          (sw_070_clk_out),
        .data_in         (sw_070_data_out),
        .scan_select_in  (sw_070_scan_out),
        .latch_enable_in (sw_070_latch_out),
        .clk_out         (sw_071_clk_out),
        .data_out        (sw_071_data_out),
        .scan_select_out (sw_071_scan_out),
        .latch_enable_out(sw_071_latch_out)
    );

    // [072] https://github.com/Sirawit7205/tinytapeout-2G97-2G98
    wire sw_072_clk_out, sw_072_data_out, sw_072_scan_out, sw_072_latch_out;
    scan_wrapper_341432030163108435 #(.NUM_IOS(8)) scan_wrapper_341432030163108435_72 (
        .clk_in          (sw_071_clk_out),
        .data_in         (sw_071_data_out),
        .scan_select_in  (sw_071_scan_out),
        .latch_enable_in (sw_071_latch_out),
        .clk_out         (sw_072_clk_out),
        .data_out        (sw_072_data_out),
        .scan_select_out (sw_072_scan_out),
        .latch_enable_out(sw_072_latch_out)
    );

    // [073] https://github.com/hosein-mokarian/tinytapeout_counter_3to8_decoder
    wire sw_073_clk_out, sw_073_data_out, sw_073_scan_out, sw_073_latch_out;
    scan_wrapper_341440114308678227 #(.NUM_IOS(8)) scan_wrapper_341440114308678227_73 (
        .clk_in          (sw_072_clk_out),
        .data_in         (sw_072_data_out),
        .scan_select_in  (sw_072_scan_out),
        .latch_enable_in (sw_072_latch_out),
        .clk_out         (sw_073_clk_out),
        .data_out        (sw_073_data_out),
        .scan_select_out (sw_073_scan_out),
        .latch_enable_out(sw_073_latch_out)
    );

    // [074] https://github.com/burtyb/srld
    wire sw_074_clk_out, sw_074_data_out, sw_074_scan_out, sw_074_latch_out;
    scan_wrapper_341496918381167187 #(.NUM_IOS(8)) scan_wrapper_341496918381167187_74 (
        .clk_in          (sw_073_clk_out),
        .data_in         (sw_073_data_out),
        .scan_select_in  (sw_073_scan_out),
        .latch_enable_in (sw_073_latch_out),
        .clk_out         (sw_074_clk_out),
        .data_out        (sw_074_data_out),
        .scan_select_out (sw_074_scan_out),
        .latch_enable_out(sw_074_latch_out)
    );

    // [075] https://github.com/Mahnoor-ismail01/tinytapeout-chromatic-3-to-8-Decoder
    wire sw_075_clk_out, sw_075_data_out, sw_075_scan_out, sw_075_latch_out;
    scan_wrapper_341440781874102868 #(.NUM_IOS(8)) scan_wrapper_341440781874102868_75 (
        .clk_in          (sw_074_clk_out),
        .data_in         (sw_074_data_out),
        .scan_select_in  (sw_074_scan_out),
        .latch_enable_in (sw_074_latch_out),
        .clk_out         (sw_075_clk_out),
        .data_out        (sw_075_data_out),
        .scan_select_out (sw_075_scan_out),
        .latch_enable_out(sw_075_latch_out)
    );

    // [076] https://github.com/Shahzaib2028/tinytapeout-4to2Encoder-2to4Decoder
    wire sw_076_clk_out, sw_076_data_out, sw_076_scan_out, sw_076_latch_out;
    scan_wrapper_341444501414347346 #(.NUM_IOS(8)) scan_wrapper_341444501414347346_76 (
        .clk_in          (sw_075_clk_out),
        .data_in         (sw_075_data_out),
        .scan_select_in  (sw_075_scan_out),
        .latch_enable_in (sw_075_latch_out),
        .clk_out         (sw_076_clk_out),
        .data_out        (sw_076_data_out),
        .scan_select_out (sw_076_scan_out),
        .latch_enable_out(sw_076_latch_out)
    );

    // [077] https://github.com/sfmth/tinytapeout-tinycordic
    wire sw_077_clk_out, sw_077_data_out, sw_077_scan_out, sw_077_latch_out;
    scan_wrapper_019235602376235615 #(.NUM_IOS(8)) scan_wrapper_019235602376235615_77 (
        .clk_in          (sw_076_clk_out),
        .data_in         (sw_076_data_out),
        .scan_select_in  (sw_076_scan_out),
        .latch_enable_in (sw_076_latch_out),
        .clk_out         (sw_077_clk_out),
        .data_out        (sw_077_data_out),
        .scan_select_out (sw_077_scan_out),
        .latch_enable_out(sw_077_latch_out)
    );

    // [078] https://github.com/mm21/tinytapeout-led-matrix
    wire sw_078_clk_out, sw_078_data_out, sw_078_scan_out, sw_078_latch_out;
    scan_wrapper_341450853309219412 #(.NUM_IOS(8)) scan_wrapper_341450853309219412_78 (
        .clk_in          (sw_077_clk_out),
        .data_in         (sw_077_data_out),
        .scan_select_in  (sw_077_scan_out),
        .latch_enable_in (sw_077_latch_out),
        .clk_out         (sw_078_clk_out),
        .data_out        (sw_078_data_out),
        .scan_select_out (sw_078_scan_out),
        .latch_enable_out(sw_078_latch_out)
    );

    // [079] https://github.com/jeanthom/tinytapout-lock
    wire sw_079_clk_out, sw_079_data_out, sw_079_scan_out, sw_079_latch_out;
    scan_wrapper_341438392303616596 #(.NUM_IOS(8)) scan_wrapper_341438392303616596_79 (
        .clk_in          (sw_078_clk_out),
        .data_in         (sw_078_data_out),
        .scan_select_in  (sw_078_scan_out),
        .latch_enable_in (sw_078_latch_out),
        .clk_out         (sw_079_clk_out),
        .data_out        (sw_079_data_out),
        .scan_select_out (sw_079_scan_out),
        .latch_enable_out(sw_079_latch_out)
    );

    // [080] https://github.com/AidanMedcalf/tinytapeout-tinyio
    wire sw_080_clk_out, sw_080_data_out, sw_080_scan_out, sw_080_latch_out;
    scan_wrapper_341432284947153491 #(.NUM_IOS(8)) scan_wrapper_341432284947153491_80 (
        .clk_in          (sw_079_clk_out),
        .data_in         (sw_079_data_out),
        .scan_select_in  (sw_079_scan_out),
        .latch_enable_in (sw_079_latch_out),
        .clk_out         (sw_080_clk_out),
        .data_out        (sw_080_data_out),
        .scan_select_out (sw_080_scan_out),
        .latch_enable_out(sw_080_latch_out)
    );

    // [081] https://github.com/ElectricPotato/tinytapeout-hello-world-uart
    wire sw_081_clk_out, sw_081_data_out, sw_081_scan_out, sw_081_latch_out;
    scan_wrapper_341457971277988435 #(.NUM_IOS(8)) scan_wrapper_341457971277988435_81 (
        .clk_in          (sw_080_clk_out),
        .data_in         (sw_080_data_out),
        .scan_select_in  (sw_080_scan_out),
        .latch_enable_in (sw_080_latch_out),
        .clk_out         (sw_081_clk_out),
        .data_out        (sw_081_data_out),
        .scan_select_out (sw_081_scan_out),
        .latch_enable_out(sw_081_latch_out)
    );

    // [082] https://github.com/abdullahkhalids/TinyTapeout-hamming-code
    wire sw_082_clk_out, sw_082_data_out, sw_082_scan_out, sw_082_latch_out;
    scan_wrapper_341399568412312147 #(.NUM_IOS(8)) scan_wrapper_341399568412312147_82 (
        .clk_in          (sw_081_clk_out),
        .data_in         (sw_081_data_out),
        .scan_select_in  (sw_081_scan_out),
        .latch_enable_in (sw_081_latch_out),
        .clk_out         (sw_082_clk_out),
        .data_out        (sw_082_data_out),
        .scan_select_out (sw_082_scan_out),
        .latch_enable_out(sw_082_latch_out)
    );

    // [083] https://github.com/hossein1387/tinytapeout-verilog-test
    wire sw_083_clk_out, sw_083_data_out, sw_083_scan_out, sw_083_latch_out;
    scan_wrapper_341464767397888596 #(.NUM_IOS(8)) scan_wrapper_341464767397888596_83 (
        .clk_in          (sw_082_clk_out),
        .data_in         (sw_082_data_out),
        .scan_select_in  (sw_082_scan_out),
        .latch_enable_in (sw_082_latch_out),
        .clk_out         (sw_083_clk_out),
        .data_out        (sw_083_data_out),
        .scan_select_out (sw_083_scan_out),
        .latch_enable_out(sw_083_latch_out)
    );

    // [084] https://github.com/ChrisPVille/tinytapeout-FROG4bitCPU
    wire sw_084_clk_out, sw_084_data_out, sw_084_scan_out, sw_084_latch_out;
    scan_wrapper_341476989274686036 #(.NUM_IOS(8)) scan_wrapper_341476989274686036_84 (
        .clk_in          (sw_083_clk_out),
        .data_in         (sw_083_data_out),
        .scan_select_in  (sw_083_scan_out),
        .latch_enable_in (sw_083_latch_out),
        .clk_out         (sw_084_clk_out),
        .data_out        (sw_084_data_out),
        .scan_select_out (sw_084_scan_out),
        .latch_enable_out(sw_084_latch_out)
    );

    // [085] https://github.com/Talha-Ahmed-1/tinytapeout_flop_regfile
    wire sw_085_clk_out, sw_085_data_out, sw_085_scan_out, sw_085_latch_out;
    scan_wrapper_341482086419399252 #(.NUM_IOS(8)) scan_wrapper_341482086419399252_85 (
        .clk_in          (sw_084_clk_out),
        .data_in         (sw_084_data_out),
        .scan_select_in  (sw_084_scan_out),
        .latch_enable_in (sw_084_latch_out),
        .clk_out         (sw_085_clk_out),
        .data_out        (sw_085_data_out),
        .scan_select_out (sw_085_scan_out),
        .latch_enable_out(sw_085_latch_out)
    );

    // [086] https://github.com/skylersaleh/tinytapeout-hello
    wire sw_086_clk_out, sw_086_data_out, sw_086_scan_out, sw_086_latch_out;
    scan_wrapper_341452019534398035 #(.NUM_IOS(8)) scan_wrapper_341452019534398035_86 (
        .clk_in          (sw_085_clk_out),
        .data_in         (sw_085_data_out),
        .scan_select_in  (sw_085_scan_out),
        .latch_enable_in (sw_085_latch_out),
        .clk_out         (sw_086_clk_out),
        .data_out        (sw_086_data_out),
        .scan_select_out (sw_086_scan_out),
        .latch_enable_out(sw_086_latch_out)
    );

    // [087] https://github.com/proppy/tinytapeout-xls-popcount
    wire sw_087_clk_out, sw_087_data_out, sw_087_scan_out, sw_087_latch_out;
    scan_wrapper_341497971083313748 #(.NUM_IOS(8)) scan_wrapper_341497971083313748_87 (
        .clk_in          (sw_086_clk_out),
        .data_in         (sw_086_data_out),
        .scan_select_in  (sw_086_scan_out),
        .latch_enable_in (sw_086_latch_out),
        .clk_out         (sw_087_clk_out),
        .data_out        (sw_087_data_out),
        .scan_select_out (sw_087_scan_out),
        .latch_enable_out(sw_087_latch_out)
    );

    // [088] https://github.com/proppy/tinytapeout-xls-popcount-bithacks
    wire sw_088_clk_out, sw_088_data_out, sw_088_scan_out, sw_088_latch_out;
    scan_wrapper_341497964482527828 #(.NUM_IOS(8)) scan_wrapper_341497964482527828_88 (
        .clk_in          (sw_087_clk_out),
        .data_in         (sw_087_data_out),
        .scan_select_in  (sw_087_scan_out),
        .latch_enable_in (sw_087_latch_out),
        .clk_out         (sw_088_clk_out),
        .data_out        (sw_088_data_out),
        .scan_select_out (sw_088_scan_out),
        .latch_enable_out(sw_088_latch_out)
    );

    // [089] https://github.com/proppy/tinytapeout-xls-inverter
    wire sw_089_clk_out, sw_089_data_out, sw_089_scan_out, sw_089_latch_out;
    scan_wrapper_341497938559631956 #(.NUM_IOS(8)) scan_wrapper_341497938559631956_89 (
        .clk_in          (sw_088_clk_out),
        .data_in         (sw_088_data_out),
        .scan_select_in  (sw_088_scan_out),
        .latch_enable_in (sw_088_latch_out),
        .clk_out         (sw_089_clk_out),
        .data_out        (sw_089_data_out),
        .scan_select_out (sw_089_scan_out),
        .latch_enable_out(sw_089_latch_out)
    );

    // [090] https://github.com/mark64/tinytapeout
    wire sw_090_clk_out, sw_090_data_out, sw_090_scan_out, sw_090_latch_out;
    scan_wrapper_341499976001520211 #(.NUM_IOS(8)) scan_wrapper_341499976001520211_90 (
        .clk_in          (sw_089_clk_out),
        .data_in         (sw_089_data_out),
        .scan_select_in  (sw_089_scan_out),
        .latch_enable_in (sw_089_latch_out),
        .clk_out         (sw_090_clk_out),
        .data_out        (sw_090_data_out),
        .scan_select_out (sw_090_scan_out),
        .latch_enable_out(sw_090_latch_out)
    );

    // [091] https://github.com/dave-roo/ddcomparatorandro
    wire sw_091_clk_out, sw_091_data_out, sw_091_scan_out, sw_091_latch_out;
    scan_wrapper_341500800901579348 #(.NUM_IOS(8)) scan_wrapper_341500800901579348_91 (
        .clk_in          (sw_090_clk_out),
        .data_in         (sw_090_data_out),
        .scan_select_in  (sw_090_scan_out),
        .latch_enable_in (sw_090_latch_out),
        .clk_out         (sw_091_clk_out),
        .data_out        (sw_091_data_out),
        .scan_select_out (sw_091_scan_out),
        .latch_enable_out(sw_091_latch_out)
    );

    // [092] https://github.com/splinedrive/tinytapeout-verilog-4x4-multiplier
    wire sw_092_clk_out, sw_092_data_out, sw_092_scan_out, sw_092_latch_out;
    scan_wrapper_341493393195532884 #(.NUM_IOS(8)) scan_wrapper_341493393195532884_92 (
        .clk_in          (sw_091_clk_out),
        .data_in         (sw_091_data_out),
        .scan_select_in  (sw_091_scan_out),
        .latch_enable_in (sw_091_latch_out),
        .clk_out         (sw_092_clk_out),
        .data_out        (sw_092_data_out),
        .scan_select_out (sw_092_scan_out),
        .latch_enable_out(sw_092_latch_out)
    );

    // [093] https://github.com/ThorKn/tinytapeout_shiftregister_8bit
    wire sw_093_clk_out, sw_093_data_out, sw_093_scan_out, sw_093_latch_out;
    scan_wrapper_341506274933867090 #(.NUM_IOS(8)) scan_wrapper_341506274933867090_93 (
        .clk_in          (sw_092_clk_out),
        .data_in         (sw_092_data_out),
        .scan_select_in  (sw_092_scan_out),
        .latch_enable_in (sw_092_latch_out),
        .clk_out         (sw_093_clk_out),
        .data_out        (sw_093_data_out),
        .scan_select_out (sw_093_scan_out),
        .latch_enable_out(sw_093_latch_out)
    );

    // [094] https://github.com/UDXS/tinytapeout-sqrt
    wire sw_094_clk_out, sw_094_data_out, sw_094_scan_out, sw_094_latch_out;
    scan_wrapper_341449297858921043 #(.NUM_IOS(8)) scan_wrapper_341449297858921043_94 (
        .clk_in          (sw_093_clk_out),
        .data_in         (sw_093_data_out),
        .scan_select_in  (sw_093_scan_out),
        .latch_enable_in (sw_093_latch_out),
        .clk_out         (sw_094_clk_out),
        .data_out        (sw_094_data_out),
        .scan_select_out (sw_094_scan_out),
        .latch_enable_out(sw_094_latch_out)
    );

    // [095] https://github.com/coralmw/tinytapeout-css-feedback
    wire sw_095_clk_out, sw_095_data_out, sw_095_scan_out, sw_095_latch_out;
    scan_wrapper_341710255833481812 #(.NUM_IOS(8)) scan_wrapper_341710255833481812_95 (
        .clk_in          (sw_094_clk_out),
        .data_in         (sw_094_data_out),
        .scan_select_in  (sw_094_scan_out),
        .latch_enable_in (sw_094_latch_out),
        .clk_out         (sw_095_clk_out),
        .data_out        (sw_095_data_out),
        .scan_select_out (sw_095_scan_out),
        .latch_enable_out(sw_095_latch_out)
    );

    // [096] https://github.com/ericsmi/tinytapeout-verilog-div3
    wire sw_096_clk_out, sw_096_data_out, sw_096_scan_out, sw_096_latch_out;
    scan_wrapper_340067262721426004 #(.NUM_IOS(8)) scan_wrapper_340067262721426004_96 (
        .clk_in          (sw_095_clk_out),
        .data_in         (sw_095_data_out),
        .scan_select_in  (sw_095_scan_out),
        .latch_enable_in (sw_095_latch_out),
        .clk_out         (sw_096_clk_out),
        .data_out        (sw_096_data_out),
        .scan_select_out (sw_096_scan_out),
        .latch_enable_out(sw_096_latch_out)
    );

    // [097] https://github.com/fluxfocus/jdtt-logic1.git
    wire sw_097_clk_out, sw_097_data_out, sw_097_scan_out, sw_097_latch_out;
    scan_wrapper_341462925422101075 #(.NUM_IOS(8)) scan_wrapper_341462925422101075_97 (
        .clk_in          (sw_096_clk_out),
        .data_in         (sw_096_data_out),
        .scan_select_in  (sw_096_scan_out),
        .latch_enable_in (sw_096_latch_out),
        .clk_out         (sw_097_clk_out),
        .data_out        (sw_097_data_out),
        .scan_select_out (sw_097_scan_out),
        .latch_enable_out(sw_097_latch_out)
    );

    // [098] https://github.com/anm/nyasic
    wire sw_098_clk_out, sw_098_data_out, sw_098_scan_out, sw_098_latch_out;
    scan_wrapper_341520747710120530 #(.NUM_IOS(8)) scan_wrapper_341520747710120530_98 (
        .clk_in          (sw_097_clk_out),
        .data_in         (sw_097_data_out),
        .scan_select_in  (sw_097_scan_out),
        .latch_enable_in (sw_097_latch_out),
        .clk_out         (sw_098_clk_out),
        .data_out        (sw_098_data_out),
        .scan_select_out (sw_098_scan_out),
        .latch_enable_out(sw_098_latch_out)
    );

    // [099] https://github.com/aiunderstand/tinytapeout_bintristateloadablecounter
    wire sw_099_clk_out, sw_099_data_out, sw_099_scan_out, sw_099_latch_out;
    scan_wrapper_341423712597181012 #(.NUM_IOS(8)) scan_wrapper_341423712597181012_99 (
        .clk_in          (sw_098_clk_out),
        .data_in         (sw_098_data_out),
        .scan_select_in  (sw_098_scan_out),
        .latch_enable_in (sw_098_latch_out),
        .clk_out         (sw_099_clk_out),
        .data_out        (sw_099_data_out),
        .scan_select_out (sw_099_scan_out),
        .latch_enable_out(sw_099_latch_out)
    );

    // [100] https://github.com/ThorKn/tinytapeout_shiftregister_challenge
    wire sw_100_clk_out, sw_100_data_out, sw_100_scan_out, sw_100_latch_out;
    scan_wrapper_341516949939814994 #(.NUM_IOS(8)) scan_wrapper_341516949939814994_100 (
        .clk_in          (sw_099_clk_out),
        .data_in         (sw_099_data_out),
        .scan_select_in  (sw_099_scan_out),
        .latch_enable_in (sw_099_latch_out),
        .clk_out         (sw_100_clk_out),
        .data_out        (sw_100_data_out),
        .scan_select_out (sw_100_scan_out),
        .latch_enable_out(sw_100_latch_out)
    );

    // [101] https://github.com/regymm/tinytapeout-mcpi
    wire sw_101_clk_out, sw_101_data_out, sw_101_scan_out, sw_101_latch_out;
    scan_wrapper_341521390605697619 #(.NUM_IOS(8)) scan_wrapper_341521390605697619_101 (
        .clk_in          (sw_100_clk_out),
        .data_in         (sw_100_data_out),
        .scan_select_in  (sw_100_scan_out),
        .latch_enable_in (sw_100_latch_out),
        .clk_out         (sw_101_clk_out),
        .data_out        (sw_101_data_out),
        .scan_select_out (sw_101_scan_out),
        .latch_enable_out(sw_101_latch_out)
    );

    // [102] https://github.com/todd1251/tinytapeout-figure8
    wire sw_102_clk_out, sw_102_data_out, sw_102_scan_out, sw_102_latch_out;
    scan_wrapper_341243232292700755 #(.NUM_IOS(8)) scan_wrapper_341243232292700755_102 (
        .clk_in          (sw_101_clk_out),
        .data_in         (sw_101_data_out),
        .scan_select_in  (sw_101_scan_out),
        .latch_enable_in (sw_101_latch_out),
        .clk_out         (sw_102_clk_out),
        .data_out        (sw_102_data_out),
        .scan_select_out (sw_102_scan_out),
        .latch_enable_out(sw_102_latch_out)
    );

    // [103] https://github.com/CyberGai/tinytapeout-bcd-counter
    wire sw_103_clk_out, sw_103_data_out, sw_103_scan_out, sw_103_latch_out;
    scan_wrapper_341519170869920338 #(.NUM_IOS(8)) scan_wrapper_341519170869920338_103 (
        .clk_in          (sw_102_clk_out),
        .data_in         (sw_102_data_out),
        .scan_select_in  (sw_102_scan_out),
        .latch_enable_in (sw_102_latch_out),
        .clk_out         (sw_103_clk_out),
        .data_out        (sw_103_data_out),
        .scan_select_out (sw_103_scan_out),
        .latch_enable_out(sw_103_latch_out)
    );

    // [104] https://github.com/georgeyhere/tinytapeout-dice-roller
    wire sw_104_clk_out, sw_104_data_out, sw_104_scan_out, sw_104_latch_out;
    scan_wrapper_341446083683025490 #(.NUM_IOS(8)) scan_wrapper_341446083683025490_104 (
        .clk_in          (sw_103_clk_out),
        .data_in         (sw_103_data_out),
        .scan_select_in  (sw_103_scan_out),
        .latch_enable_in (sw_103_latch_out),
        .clk_out         (sw_104_clk_out),
        .data_out        (sw_104_data_out),
        .scan_select_out (sw_104_scan_out),
        .latch_enable_out(sw_104_latch_out)
    );

    // [105] https://github.com/nayanesh-reddy/2-Bit_Add_Mul_Comp
    wire sw_105_clk_out, sw_105_data_out, sw_105_scan_out, sw_105_latch_out;
    scan_wrapper_341524192738411090 #(.NUM_IOS(8)) scan_wrapper_341524192738411090_105 (
        .clk_in          (sw_104_clk_out),
        .data_in         (sw_104_data_out),
        .scan_select_in  (sw_104_scan_out),
        .latch_enable_in (sw_104_latch_out),
        .clk_out         (sw_105_clk_out),
        .data_out        (sw_105_data_out),
        .scan_select_out (sw_105_scan_out),
        .latch_enable_out(sw_105_latch_out)
    );

    // [106] https://github.com/ryancor/half_addr_asic
    wire sw_106_clk_out, sw_106_data_out, sw_106_scan_out, sw_106_latch_out;
    scan_wrapper_341533740987581011 #(.NUM_IOS(8)) scan_wrapper_341533740987581011_106 (
        .clk_in          (sw_105_clk_out),
        .data_in         (sw_105_data_out),
        .scan_select_in  (sw_105_scan_out),
        .latch_enable_in (sw_105_latch_out),
        .clk_out         (sw_106_clk_out),
        .data_out        (sw_106_data_out),
        .scan_select_out (sw_106_scan_out),
        .latch_enable_out(sw_106_latch_out)
    );

    // [107] https://github.com/hovind/tinytapeout-verilog-test
    wire sw_107_clk_out, sw_107_data_out, sw_107_scan_out, sw_107_latch_out;
    scan_wrapper_341431502448362067 #(.NUM_IOS(8)) scan_wrapper_341431502448362067_107 (
        .clk_in          (sw_106_clk_out),
        .data_in         (sw_106_data_out),
        .scan_select_in  (sw_106_scan_out),
        .latch_enable_in (sw_106_latch_out),
        .clk_out         (sw_107_clk_out),
        .data_out        (sw_107_data_out),
        .scan_select_out (sw_107_scan_out),
        .latch_enable_out(sw_107_latch_out)
    );

    // [108] https://github.com/siriusm46/tinytapeout_bcd_decimal
    wire sw_108_clk_out, sw_108_data_out, sw_108_scan_out, sw_108_latch_out;
    scan_wrapper_341473139924927058 #(.NUM_IOS(8)) scan_wrapper_341473139924927058_108 (
        .clk_in          (sw_107_clk_out),
        .data_in         (sw_107_data_out),
        .scan_select_in  (sw_107_scan_out),
        .latch_enable_in (sw_107_latch_out),
        .clk_out         (sw_108_clk_out),
        .data_out        (sw_108_data_out),
        .scan_select_out (sw_108_scan_out),
        .latch_enable_out(sw_108_latch_out)
    );

    // [109] https://github.com/cpldcpu/tinytapeout_mcpu5
    wire sw_109_clk_out, sw_109_data_out, sw_109_scan_out, sw_109_latch_out;
    scan_wrapper_341528610027340372 #(.NUM_IOS(8)) scan_wrapper_341528610027340372_109 (
        .clk_in          (sw_108_clk_out),
        .data_in         (sw_108_data_out),
        .scan_select_in  (sw_108_scan_out),
        .latch_enable_in (sw_108_latch_out),
        .clk_out         (sw_109_clk_out),
        .data_out        (sw_109_data_out),
        .scan_select_out (sw_109_scan_out),
        .latch_enable_out(sw_109_latch_out)
    );

    // [110] https://github.com/goran-mahovlic/tinytapeout-verilog-piano
    wire sw_110_clk_out, sw_110_data_out, sw_110_scan_out, sw_110_latch_out;
    scan_wrapper_341424636358034002 #(.NUM_IOS(8)) scan_wrapper_341424636358034002_110 (
        .clk_in          (sw_109_clk_out),
        .data_in         (sw_109_data_out),
        .scan_select_in  (sw_109_scan_out),
        .latch_enable_in (sw_109_latch_out),
        .clk_out         (sw_110_clk_out),
        .data_out        (sw_110_data_out),
        .scan_select_out (sw_110_scan_out),
        .latch_enable_out(sw_110_latch_out)
    );

    // [111] https://github.com/andars/universal-turing-machine-aw7s8
    wire sw_111_clk_out, sw_111_data_out, sw_111_scan_out, sw_111_latch_out;
    scan_wrapper_341717091617866324 #(.NUM_IOS(8)) scan_wrapper_341717091617866324_111 (
        .clk_in          (sw_110_clk_out),
        .data_in         (sw_110_data_out),
        .scan_select_in  (sw_110_scan_out),
        .latch_enable_in (sw_110_latch_out),
        .clk_out         (sw_111_clk_out),
        .data_out        (sw_111_data_out),
        .scan_select_out (sw_111_scan_out),
        .latch_enable_out(sw_111_latch_out)
    );

    // [112] https://github.com/marcusmueller/hamming74-tapeout
    wire sw_112_clk_out, sw_112_data_out, sw_112_scan_out, sw_112_latch_out;
    scan_wrapper_hamming74 #(.NUM_IOS(8)) scan_wrapper_hamming74_112 (
        .clk_in          (sw_111_clk_out),
        .data_in         (sw_111_data_out),
        .scan_select_in  (sw_111_scan_out),
        .latch_enable_in (sw_111_latch_out),
        .clk_out         (sw_112_clk_out),
        .data_out        (sw_112_data_out),
        .scan_select_out (sw_112_scan_out),
        .latch_enable_out(sw_112_latch_out)
    );

    // [113] https://github.com/13arn/tinytapeout_counter_steamdeck
    wire sw_113_clk_out, sw_113_data_out, sw_113_scan_out, sw_113_latch_out;
    scan_wrapper_341541108650607187 #(.NUM_IOS(8)) scan_wrapper_341541108650607187_113 (
        .clk_in          (sw_112_clk_out),
        .data_in         (sw_112_data_out),
        .scan_select_in  (sw_112_scan_out),
        .latch_enable_in (sw_112_latch_out),
        .clk_out         (sw_113_clk_out),
        .data_out        (sw_113_data_out),
        .scan_select_out (sw_113_scan_out),
        .latch_enable_out(sw_113_latch_out)
    );

    // [114] https://github.com/johshoff/tinytapeout-verilog
    wire sw_114_clk_out, sw_114_data_out, sw_114_scan_out, sw_114_latch_out;
    scan_wrapper_341360223723717202 #(.NUM_IOS(8)) scan_wrapper_341360223723717202_114 (
        .clk_in          (sw_113_clk_out),
        .data_in         (sw_113_data_out),
        .scan_select_in  (sw_113_scan_out),
        .latch_enable_in (sw_113_latch_out),
        .clk_out         (sw_114_clk_out),
        .data_out        (sw_114_data_out),
        .scan_select_out (sw_114_scan_out),
        .latch_enable_out(sw_114_latch_out)
    );

    // [115] https://github.com/cy384/seven-segment-with-adder
    wire sw_115_clk_out, sw_115_data_out, sw_115_scan_out, sw_115_latch_out;
    scan_wrapper_341546888233747026 #(.NUM_IOS(8)) scan_wrapper_341546888233747026_115 (
        .clk_in          (sw_114_clk_out),
        .data_in         (sw_114_data_out),
        .scan_select_in  (sw_114_scan_out),
        .latch_enable_in (sw_114_latch_out),
        .clk_out         (sw_115_clk_out),
        .data_out        (sw_115_data_out),
        .scan_select_out (sw_115_scan_out),
        .latch_enable_out(sw_115_latch_out)
    );

    // [116] https://github.com/georgerennie/tinytapeout-wokwi-cd4518
    wire sw_116_clk_out, sw_116_data_out, sw_116_scan_out, sw_116_latch_out;
    scan_wrapper_340979268609638995 #(.NUM_IOS(8)) scan_wrapper_340979268609638995_116 (
        .clk_in          (sw_115_clk_out),
        .data_in         (sw_115_data_out),
        .scan_select_in  (sw_115_scan_out),
        .latch_enable_in (sw_115_latch_out),
        .clk_out         (sw_116_clk_out),
        .data_out        (sw_116_data_out),
        .scan_select_out (sw_116_scan_out),
        .latch_enable_out(sw_116_latch_out)
    );

    // [117] https://github.com/ElectricPotato/tinytapeout-picture-printer-b
    wire sw_117_clk_out, sw_117_data_out, sw_117_scan_out, sw_117_latch_out;
    scan_wrapper_341542971476279892 #(.NUM_IOS(8)) scan_wrapper_341542971476279892_117 (
        .clk_in          (sw_116_clk_out),
        .data_in         (sw_116_data_out),
        .scan_select_in  (sw_116_scan_out),
        .latch_enable_in (sw_116_latch_out),
        .clk_out         (sw_117_clk_out),
        .data_out        (sw_117_data_out),
        .scan_select_out (sw_117_scan_out),
        .latch_enable_out(sw_117_latch_out)
    );

    // [118] https://github.com/theFestest/tinytapeout-simple-invert8
    wire sw_118_clk_out, sw_118_data_out, sw_118_scan_out, sw_118_latch_out;
    scan_wrapper_341556236196512338 #(.NUM_IOS(8)) scan_wrapper_341556236196512338_118 (
        .clk_in          (sw_117_clk_out),
        .data_in         (sw_117_data_out),
        .scan_select_in  (sw_117_scan_out),
        .latch_enable_in (sw_117_latch_out),
        .clk_out         (sw_118_clk_out),
        .data_out        (sw_118_data_out),
        .scan_select_out (sw_118_scan_out),
        .latch_enable_out(sw_118_latch_out)
    );

    // [119] https://github.com/ArsenioDev/CustomSiliconTest
    wire sw_119_clk_out, sw_119_data_out, sw_119_scan_out, sw_119_latch_out;
    scan_wrapper_341558189536313940 #(.NUM_IOS(8)) scan_wrapper_341558189536313940_119 (
        .clk_in          (sw_118_clk_out),
        .data_in         (sw_118_data_out),
        .scan_select_in  (sw_118_scan_out),
        .latch_enable_in (sw_118_latch_out),
        .clk_out         (sw_119_clk_out),
        .data_out        (sw_119_data_out),
        .scan_select_out (sw_119_scan_out),
        .latch_enable_out(sw_119_latch_out)
    );

    // [120] https://github.com/mgargano/tinytapeout_alu_with_4bit_7segmetdisplay_decoder
    wire sw_120_clk_out, sw_120_data_out, sw_120_scan_out, sw_120_latch_out;
    scan_wrapper_341538994733974098 #(.NUM_IOS(8)) scan_wrapper_341538994733974098_120 (
        .clk_in          (sw_119_clk_out),
        .data_in         (sw_119_data_out),
        .scan_select_in  (sw_119_scan_out),
        .latch_enable_in (sw_119_latch_out),
        .clk_out         (sw_120_clk_out),
        .data_out        (sw_120_data_out),
        .scan_select_out (sw_120_scan_out),
        .latch_enable_out(sw_120_latch_out)
    );

    // [121] https://github.com/theFestest/tinytapeout-4x4-ram
    wire sw_121_clk_out, sw_121_data_out, sw_121_scan_out, sw_121_latch_out;
    scan_wrapper_341557831870186068 #(.NUM_IOS(8)) scan_wrapper_341557831870186068_121 (
        .clk_in          (sw_120_clk_out),
        .data_in         (sw_120_data_out),
        .scan_select_in  (sw_120_scan_out),
        .latch_enable_in (sw_120_latch_out),
        .clk_out         (sw_121_clk_out),
        .data_out        (sw_121_data_out),
        .scan_select_out (sw_121_scan_out),
        .latch_enable_out(sw_121_latch_out)
    );

    // [122] https://github.com/michael-christen/wokwi-verilog-asic-experiment
    wire sw_122_clk_out, sw_122_data_out, sw_122_scan_out, sw_122_latch_out;
    scan_wrapper_341569483755749970 #(.NUM_IOS(8)) scan_wrapper_341569483755749970_122 (
        .clk_in          (sw_121_clk_out),
        .data_in         (sw_121_data_out),
        .scan_select_in  (sw_121_scan_out),
        .latch_enable_in (sw_121_latch_out),
        .clk_out         (sw_122_clk_out),
        .data_out        (sw_122_data_out),
        .scan_select_out (sw_122_scan_out),
        .latch_enable_out(sw_122_latch_out)
    );

    // [123] https://github.com/craigcc-frii/tinytapeout_craig
    wire sw_123_clk_out, sw_123_data_out, sw_123_scan_out, sw_123_latch_out;
    scan_wrapper_341573751072096850 #(.NUM_IOS(8)) scan_wrapper_341573751072096850_123 (
        .clk_in          (sw_122_clk_out),
        .data_in         (sw_122_data_out),
        .scan_select_in  (sw_122_scan_out),
        .latch_enable_in (sw_122_latch_out),
        .clk_out         (sw_123_clk_out),
        .data_out        (sw_123_data_out),
        .scan_select_out (sw_123_scan_out),
        .latch_enable_out(sw_123_latch_out)
    );

    // [124] https://github.com/youngpines/r2rdac_tinytapeout_demo
    wire sw_124_clk_out, sw_124_data_out, sw_124_scan_out, sw_124_latch_out;
    scan_wrapper_341571228858843732 #(.NUM_IOS(8)) scan_wrapper_341571228858843732_124 (
        .clk_in          (sw_123_clk_out),
        .data_in         (sw_123_data_out),
        .scan_select_in  (sw_123_scan_out),
        .latch_enable_in (sw_123_latch_out),
        .clk_out         (sw_124_clk_out),
        .data_out        (sw_124_data_out),
        .scan_select_out (sw_124_scan_out),
        .latch_enable_out(sw_124_latch_out)
    );

    // [125] https://github.com/toybuilder/learn-tinytapeout
    wire sw_125_clk_out, sw_125_data_out, sw_125_scan_out, sw_125_latch_out;
    scan_wrapper_341490465660469844 #(.NUM_IOS(8)) scan_wrapper_341490465660469844_125 (
        .clk_in          (sw_124_clk_out),
        .data_in         (sw_124_data_out),
        .scan_select_in  (sw_124_scan_out),
        .latch_enable_in (sw_124_latch_out),
        .clk_out         (sw_125_clk_out),
        .data_out        (sw_125_data_out),
        .scan_select_out (sw_125_scan_out),
        .latch_enable_out(sw_125_latch_out)
    );

    // [126] https://github.com/eggsactly/tinytapeout_demo
    wire sw_126_clk_out, sw_126_data_out, sw_126_scan_out, sw_126_latch_out;
    scan_wrapper_341581732833657427 #(.NUM_IOS(8)) scan_wrapper_341581732833657427_126 (
        .clk_in          (sw_125_clk_out),
        .data_in         (sw_125_data_out),
        .scan_select_in  (sw_125_scan_out),
        .latch_enable_in (sw_125_latch_out),
        .clk_out         (sw_126_clk_out),
        .data_out        (sw_126_data_out),
        .scan_select_out (sw_126_scan_out),
        .latch_enable_out(sw_126_latch_out)
    );

    // [127] https://github.com/gsegura96/tinytapeout-chisel
    wire sw_127_clk_out, sw_127_data_out, sw_127_scan_out, sw_127_latch_out;
    scan_wrapper_341457494561784402 #(.NUM_IOS(8)) scan_wrapper_341457494561784402_127 (
        .clk_in          (sw_126_clk_out),
        .data_in         (sw_126_data_out),
        .scan_select_in  (sw_126_scan_out),
        .latch_enable_in (sw_126_latch_out),
        .clk_out         (sw_127_clk_out),
        .data_out        (sw_127_data_out),
        .scan_select_out (sw_127_scan_out),
        .latch_enable_out(sw_127_latch_out)
    );

    // [128] https://github.com/abf149/fbna_like_verilog_abf149
    wire sw_128_clk_out, sw_128_data_out, sw_128_scan_out, sw_128_latch_out;
    scan_wrapper_341590933015364178 #(.NUM_IOS(8)) scan_wrapper_341590933015364178_128 (
        .clk_in          (sw_127_clk_out),
        .data_in         (sw_127_data_out),
        .scan_select_in  (sw_127_scan_out),
        .latch_enable_in (sw_127_latch_out),
        .clk_out         (sw_128_clk_out),
        .data_out        (sw_128_data_out),
        .scan_select_out (sw_128_scan_out),
        .latch_enable_out(sw_128_latch_out)
    );

    // [129] https://github.com/MC-SecPat/tinytapeout_chi2shares
    wire sw_129_clk_out, sw_129_data_out, sw_129_scan_out, sw_129_latch_out;
    scan_wrapper_341589685194195540 #(.NUM_IOS(8)) scan_wrapper_341589685194195540_129 (
        .clk_in          (sw_128_clk_out),
        .data_in         (sw_128_data_out),
        .scan_select_in  (sw_128_scan_out),
        .latch_enable_in (sw_128_latch_out),
        .clk_out         (sw_129_clk_out),
        .data_out        (sw_129_data_out),
        .scan_select_out (sw_129_scan_out),
        .latch_enable_out(sw_129_latch_out)
    );

    // [130] https://github.com/MC-SecPat/tinytapeout_chi3shares
    wire sw_130_clk_out, sw_130_data_out, sw_130_scan_out, sw_130_latch_out;
    scan_wrapper_341608574336631379 #(.NUM_IOS(8)) scan_wrapper_341608574336631379_130 (
        .clk_in          (sw_129_clk_out),
        .data_in         (sw_129_data_out),
        .scan_select_in  (sw_129_scan_out),
        .latch_enable_in (sw_129_latch_out),
        .clk_out         (sw_130_clk_out),
        .data_out        (sw_130_data_out),
        .scan_select_out (sw_130_scan_out),
        .latch_enable_out(sw_130_latch_out)
    );

    // [131] https://github.com/Adil8442/tiny_tapeout_test
    wire sw_131_clk_out, sw_131_data_out, sw_131_scan_out, sw_131_latch_out;
    scan_wrapper_341608297106768466 #(.NUM_IOS(8)) scan_wrapper_341608297106768466_131 (
        .clk_in          (sw_130_clk_out),
        .data_in         (sw_130_data_out),
        .scan_select_in  (sw_130_scan_out),
        .latch_enable_in (sw_130_latch_out),
        .clk_out         (sw_131_clk_out),
        .data_out        (sw_131_data_out),
        .scan_select_out (sw_131_scan_out),
        .latch_enable_out(sw_131_latch_out)
    );

    // [132] https://github.com/mattvenn/tinytapeout-341802448429515346
    wire sw_132_clk_out, sw_132_data_out, sw_132_scan_out, sw_132_latch_out;
    scan_wrapper_341802448429515346 #(.NUM_IOS(8)) scan_wrapper_341802448429515346_132 (
        .clk_in          (sw_131_clk_out),
        .data_in         (sw_131_data_out),
        .scan_select_in  (sw_131_scan_out),
        .latch_enable_in (sw_131_latch_out),
        .clk_out         (sw_132_clk_out),
        .data_out        (sw_132_data_out),
        .scan_select_out (sw_132_scan_out),
        .latch_enable_out(sw_132_latch_out)
    );

    // [133] https://github.com/r4d10n/tinytapeout-HELLo-3orLd-7seg
    wire sw_133_clk_out, sw_133_data_out, sw_133_scan_out, sw_133_latch_out;
    scan_wrapper_341609034095264340 #(.NUM_IOS(8)) scan_wrapper_341609034095264340_133 (
        .clk_in          (sw_132_clk_out),
        .data_in         (sw_132_data_out),
        .scan_select_in  (sw_132_scan_out),
        .latch_enable_in (sw_132_latch_out),
        .clk_out         (sw_133_clk_out),
        .data_out        (sw_133_data_out),
        .scan_select_out (sw_133_scan_out),
        .latch_enable_out(sw_133_latch_out)
    );

    // [134] https://github.com/proppy/tinytapeout-xls-graydec
    wire sw_134_clk_out, sw_134_data_out, sw_134_scan_out, sw_134_latch_out;
    scan_wrapper_341617722294010450 #(.NUM_IOS(8)) scan_wrapper_341617722294010450_134 (
        .clk_in          (sw_133_clk_out),
        .data_in         (sw_133_data_out),
        .scan_select_in  (sw_133_scan_out),
        .latch_enable_in (sw_133_latch_out),
        .clk_out         (sw_134_clk_out),
        .data_out        (sw_134_data_out),
        .scan_select_out (sw_134_scan_out),
        .latch_enable_out(sw_134_latch_out)
    );

    // [135] https://github.com/prabaldutta/tinytapeout_adi
    wire sw_135_clk_out, sw_135_data_out, sw_135_scan_out, sw_135_latch_out;
    scan_wrapper_341613097060926036 #(.NUM_IOS(8)) scan_wrapper_341613097060926036_135 (
        .clk_in          (sw_134_clk_out),
        .data_in         (sw_134_data_out),
        .scan_select_in  (sw_134_scan_out),
        .latch_enable_in (sw_134_latch_out),
        .clk_out         (sw_135_clk_out),
        .data_out        (sw_135_data_out),
        .scan_select_out (sw_135_scan_out),
        .latch_enable_out(sw_135_latch_out)
    );

    // [136] https://github.com/maehw/wokwi-verilog-gds-wolf-goat-cabbage
    wire sw_136_clk_out, sw_136_data_out, sw_136_scan_out, sw_136_latch_out;
    scan_wrapper_341614346808328788 #(.NUM_IOS(8)) scan_wrapper_341614346808328788_136 (
        .clk_in          (sw_135_clk_out),
        .data_in         (sw_135_data_out),
        .scan_select_in  (sw_135_scan_out),
        .latch_enable_in (sw_135_latch_out),
        .clk_out         (sw_136_clk_out),
        .data_out        (sw_136_data_out),
        .scan_select_out (sw_136_scan_out),
        .latch_enable_out(sw_136_latch_out)
    );

    // [137] https://github.com/ThorKn/tinytapeout_pattern_player
    wire sw_137_clk_out, sw_137_data_out, sw_137_scan_out, sw_137_latch_out;
    scan_wrapper_341620484740219475 #(.NUM_IOS(8)) scan_wrapper_341620484740219475_137 (
        .clk_in          (sw_136_clk_out),
        .data_in         (sw_136_data_out),
        .scan_select_in  (sw_136_scan_out),
        .latch_enable_in (sw_136_latch_out),
        .clk_out         (sw_137_clk_out),
        .data_out        (sw_137_data_out),
        .scan_select_out (sw_137_scan_out),
        .latch_enable_out(sw_137_latch_out)
    );

    // [138] https://github.com/rigobertoruiz98/cts_fsm
    wire sw_138_clk_out, sw_138_data_out, sw_138_scan_out, sw_138_latch_out;
    scan_wrapper_341624400621077076 #(.NUM_IOS(8)) scan_wrapper_341624400621077076_138 (
        .clk_in          (sw_137_clk_out),
        .data_in         (sw_137_data_out),
        .scan_select_in  (sw_137_scan_out),
        .latch_enable_in (sw_137_latch_out),
        .clk_out         (sw_138_clk_out),
        .data_out        (sw_138_data_out),
        .scan_select_out (sw_138_scan_out),
        .latch_enable_out(sw_138_latch_out)
    );

    // [139] https://github.com/rajarshiroy/tinytapout0_rajarshi
    wire sw_139_clk_out, sw_139_data_out, sw_139_scan_out, sw_139_latch_out;
    scan_wrapper_341614536664547922 #(.NUM_IOS(8)) scan_wrapper_341614536664547922_139 (
        .clk_in          (sw_138_clk_out),
        .data_in         (sw_138_data_out),
        .scan_select_in  (sw_138_scan_out),
        .latch_enable_in (sw_138_latch_out),
        .clk_out         (sw_139_clk_out),
        .data_out        (sw_139_data_out),
        .scan_select_out (sw_139_scan_out),
        .latch_enable_out(sw_139_latch_out)
    );

    // [140] https://github.com/BarsMonster/MicroASIC
    wire sw_140_clk_out, sw_140_data_out, sw_140_scan_out, sw_140_latch_out;
    scan_wrapper_341567111632519764 #(.NUM_IOS(8)) scan_wrapper_341567111632519764_140 (
        .clk_in          (sw_139_clk_out),
        .data_in         (sw_139_data_out),
        .scan_select_in  (sw_139_scan_out),
        .latch_enable_in (sw_139_latch_out),
        .clk_out         (sw_140_clk_out),
        .data_out        (sw_140_data_out),
        .scan_select_out (sw_140_scan_out),
        .latch_enable_out(sw_140_latch_out)
    );

    // [141] https://github.com/cpldcpu/TinyTapeout_TrainLED
    wire sw_141_clk_out, sw_141_data_out, sw_141_scan_out, sw_141_latch_out;
    scan_wrapper_341631485498884690 #(.NUM_IOS(8)) scan_wrapper_341631485498884690_141 (
        .clk_in          (sw_140_clk_out),
        .data_in         (sw_140_data_out),
        .scan_select_in  (sw_140_scan_out),
        .latch_enable_in (sw_140_latch_out),
        .clk_out         (sw_141_clk_out),
        .data_out        (sw_141_data_out),
        .scan_select_out (sw_141_scan_out),
        .latch_enable_out(sw_141_latch_out)
    );

    // [142] https://github.com/malkam03/tinytapeout-game-of-life
    wire sw_142_clk_out, sw_142_data_out, sw_142_scan_out, sw_142_latch_out;
    scan_wrapper_341632596577354323 #(.NUM_IOS(8)) scan_wrapper_341632596577354323_142 (
        .clk_in          (sw_141_clk_out),
        .data_in         (sw_141_data_out),
        .scan_select_in  (sw_141_scan_out),
        .latch_enable_in (sw_141_latch_out),
        .clk_out         (sw_142_clk_out),
        .data_out        (sw_142_data_out),
        .scan_select_out (sw_142_scan_out),
        .latch_enable_out(sw_142_latch_out)
    );

    // [143] https://github.com/BarsMonster/MicroAsicV
    wire sw_143_clk_out, sw_143_data_out, sw_143_scan_out, sw_143_latch_out;
    scan_wrapper_341628725785264722 #(.NUM_IOS(8)) scan_wrapper_341628725785264722_143 (
        .clk_in          (sw_142_clk_out),
        .data_in         (sw_142_data_out),
        .scan_select_in  (sw_142_scan_out),
        .latch_enable_in (sw_142_latch_out),
        .clk_out         (sw_143_clk_out),
        .data_out        (sw_143_data_out),
        .scan_select_out (sw_143_scan_out),
        .latch_enable_out(sw_143_latch_out)
    );

    // [144] https://github.com/maehw/wokwi-verilog-gds-lowspeed-tiny-uart
    wire sw_144_clk_out, sw_144_data_out, sw_144_scan_out, sw_144_latch_out;
    scan_wrapper_341631511790879314 #(.NUM_IOS(8)) scan_wrapper_341631511790879314_144 (
        .clk_in          (sw_143_clk_out),
        .data_in         (sw_143_data_out),
        .scan_select_in  (sw_143_scan_out),
        .latch_enable_in (sw_143_latch_out),
        .clk_out         (sw_144_clk_out),
        .data_out        (sw_144_data_out),
        .scan_select_out (sw_144_scan_out),
        .latch_enable_out(sw_144_latch_out)
    );

    // [145] https://github.com/smunaut/tinytapeout-smolram
    wire sw_145_clk_out, sw_145_data_out, sw_145_scan_out, sw_145_latch_out;
    scan_wrapper_341426151397261906 #(.NUM_IOS(8)) scan_wrapper_341426151397261906_145 (
        .clk_in          (sw_144_clk_out),
        .data_in         (sw_144_data_out),
        .scan_select_in  (sw_144_scan_out),
        .latch_enable_in (sw_144_latch_out),
        .clk_out         (sw_145_clk_out),
        .data_out        (sw_145_data_out),
        .scan_select_out (sw_145_scan_out),
        .latch_enable_out(sw_145_latch_out)
    );

    // [146] https://github.com/sirejdua/6bit-cellular-automata-tinytapeout
    wire sw_146_clk_out, sw_146_data_out, sw_146_scan_out, sw_146_latch_out;
    scan_wrapper_341629415144292948 #(.NUM_IOS(8)) scan_wrapper_341629415144292948_146 (
        .clk_in          (sw_145_clk_out),
        .data_in         (sw_145_data_out),
        .scan_select_in  (sw_145_scan_out),
        .latch_enable_in (sw_145_latch_out),
        .clk_out         (sw_146_clk_out),
        .data_out        (sw_146_data_out),
        .scan_select_out (sw_146_scan_out),
        .latch_enable_out(sw_146_latch_out)
    );

    // [147] https://github.com/DuaneSand/TinyTapeout-Hello
    wire sw_147_clk_out, sw_147_data_out, sw_147_scan_out, sw_147_latch_out;
    scan_wrapper_341637831098106450 #(.NUM_IOS(8)) scan_wrapper_341637831098106450_147 (
        .clk_in          (sw_146_clk_out),
        .data_in         (sw_146_data_out),
        .scan_select_in  (sw_146_scan_out),
        .latch_enable_in (sw_146_latch_out),
        .clk_out         (sw_147_clk_out),
        .data_out        (sw_147_data_out),
        .scan_select_out (sw_147_scan_out),
        .latch_enable_out(sw_147_latch_out)
    );

    // [148] https://github.com/tzachari/tinytapeout-lab11
    wire sw_148_clk_out, sw_148_data_out, sw_148_scan_out, sw_148_latch_out;
    scan_wrapper_341631644820570706 #(.NUM_IOS(8)) scan_wrapper_341631644820570706_148 (
        .clk_in          (sw_147_clk_out),
        .data_in         (sw_147_data_out),
        .scan_select_in  (sw_147_scan_out),
        .latch_enable_in (sw_147_latch_out),
        .clk_out         (sw_148_clk_out),
        .data_out        (sw_148_data_out),
        .scan_select_out (sw_148_scan_out),
        .latch_enable_out(sw_148_latch_out)
    );

    // [149] https://github.com/mattvenn/tinytapeout-marc
    wire sw_149_clk_out, sw_149_data_out, sw_149_scan_out, sw_149_latch_out;
    scan_wrapper_340596276030603858 #(.NUM_IOS(8)) scan_wrapper_340596276030603858_149 (
        .clk_in          (sw_148_clk_out),
        .data_in         (sw_148_data_out),
        .scan_select_in  (sw_148_scan_out),
        .latch_enable_in (sw_148_latch_out),
        .clk_out         (sw_149_clk_out),
        .data_out        (sw_149_data_out),
        .scan_select_out (sw_149_scan_out),
        .latch_enable_out(sw_149_latch_out)
    );

    // [150] https://github.com/mattvenn/tinytapeout-laura
    wire sw_150_clk_out, sw_150_data_out, sw_150_scan_out, sw_150_latch_out;
    scan_wrapper_341678527574180436 #(.NUM_IOS(8)) scan_wrapper_341678527574180436_150 (
        .clk_in          (sw_149_clk_out),
        .data_in         (sw_149_data_out),
        .scan_select_in  (sw_149_scan_out),
        .latch_enable_in (sw_149_latch_out),
        .clk_out         (sw_150_clk_out),
        .data_out        (sw_150_data_out),
        .scan_select_out (sw_150_scan_out),
        .latch_enable_out(sw_150_latch_out)
    );

    // [151] https://github.com/mattvenn/wokwi_filler
    wire sw_151_clk_out, sw_151_data_out, sw_151_scan_out, sw_151_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_151 (
        .clk_in          (sw_150_clk_out),
        .data_in         (sw_150_data_out),
        .scan_select_in  (sw_150_scan_out),
        .latch_enable_in (sw_150_latch_out),
        .clk_out         (sw_151_clk_out),
        .data_out        (sw_151_data_out),
        .scan_select_out (sw_151_scan_out),
        .latch_enable_out(sw_151_latch_out)
    );

    // [152] https://github.com/mattvenn/wokwi_filler
    wire sw_152_clk_out, sw_152_data_out, sw_152_scan_out, sw_152_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_152 (
        .clk_in          (sw_151_clk_out),
        .data_in         (sw_151_data_out),
        .scan_select_in  (sw_151_scan_out),
        .latch_enable_in (sw_151_latch_out),
        .clk_out         (sw_152_clk_out),
        .data_out        (sw_152_data_out),
        .scan_select_out (sw_152_scan_out),
        .latch_enable_out(sw_152_latch_out)
    );

    // [153] https://github.com/mattvenn/wokwi_filler
    wire sw_153_clk_out, sw_153_data_out, sw_153_scan_out, sw_153_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_153 (
        .clk_in          (sw_152_clk_out),
        .data_in         (sw_152_data_out),
        .scan_select_in  (sw_152_scan_out),
        .latch_enable_in (sw_152_latch_out),
        .clk_out         (sw_153_clk_out),
        .data_out        (sw_153_data_out),
        .scan_select_out (sw_153_scan_out),
        .latch_enable_out(sw_153_latch_out)
    );

    // [154] https://github.com/mattvenn/wokwi_filler
    wire sw_154_clk_out, sw_154_data_out, sw_154_scan_out, sw_154_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_154 (
        .clk_in          (sw_153_clk_out),
        .data_in         (sw_153_data_out),
        .scan_select_in  (sw_153_scan_out),
        .latch_enable_in (sw_153_latch_out),
        .clk_out         (sw_154_clk_out),
        .data_out        (sw_154_data_out),
        .scan_select_out (sw_154_scan_out),
        .latch_enable_out(sw_154_latch_out)
    );

    // [155] https://github.com/mattvenn/wokwi_filler
    wire sw_155_clk_out, sw_155_data_out, sw_155_scan_out, sw_155_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_155 (
        .clk_in          (sw_154_clk_out),
        .data_in         (sw_154_data_out),
        .scan_select_in  (sw_154_scan_out),
        .latch_enable_in (sw_154_latch_out),
        .clk_out         (sw_155_clk_out),
        .data_out        (sw_155_data_out),
        .scan_select_out (sw_155_scan_out),
        .latch_enable_out(sw_155_latch_out)
    );

    // [156] https://github.com/mattvenn/wokwi_filler
    wire sw_156_clk_out, sw_156_data_out, sw_156_scan_out, sw_156_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_156 (
        .clk_in          (sw_155_clk_out),
        .data_in         (sw_155_data_out),
        .scan_select_in  (sw_155_scan_out),
        .latch_enable_in (sw_155_latch_out),
        .clk_out         (sw_156_clk_out),
        .data_out        (sw_156_data_out),
        .scan_select_out (sw_156_scan_out),
        .latch_enable_out(sw_156_latch_out)
    );

    // [157] https://github.com/mattvenn/wokwi_filler
    wire sw_157_clk_out, sw_157_data_out, sw_157_scan_out, sw_157_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_157 (
        .clk_in          (sw_156_clk_out),
        .data_in         (sw_156_data_out),
        .scan_select_in  (sw_156_scan_out),
        .latch_enable_in (sw_156_latch_out),
        .clk_out         (sw_157_clk_out),
        .data_out        (sw_157_data_out),
        .scan_select_out (sw_157_scan_out),
        .latch_enable_out(sw_157_latch_out)
    );

    // [158] https://github.com/mattvenn/wokwi_filler
    wire sw_158_clk_out, sw_158_data_out, sw_158_scan_out, sw_158_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_158 (
        .clk_in          (sw_157_clk_out),
        .data_in         (sw_157_data_out),
        .scan_select_in  (sw_157_scan_out),
        .latch_enable_in (sw_157_latch_out),
        .clk_out         (sw_158_clk_out),
        .data_out        (sw_158_data_out),
        .scan_select_out (sw_158_scan_out),
        .latch_enable_out(sw_158_latch_out)
    );

    // [159] https://github.com/mattvenn/wokwi_filler
    wire sw_159_clk_out, sw_159_data_out, sw_159_scan_out, sw_159_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_159 (
        .clk_in          (sw_158_clk_out),
        .data_in         (sw_158_data_out),
        .scan_select_in  (sw_158_scan_out),
        .latch_enable_in (sw_158_latch_out),
        .clk_out         (sw_159_clk_out),
        .data_out        (sw_159_data_out),
        .scan_select_out (sw_159_scan_out),
        .latch_enable_out(sw_159_latch_out)
    );

    // [160] https://github.com/mattvenn/wokwi_filler
    wire sw_160_clk_out, sw_160_data_out, sw_160_scan_out, sw_160_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_160 (
        .clk_in          (sw_159_clk_out),
        .data_in         (sw_159_data_out),
        .scan_select_in  (sw_159_scan_out),
        .latch_enable_in (sw_159_latch_out),
        .clk_out         (sw_160_clk_out),
        .data_out        (sw_160_data_out),
        .scan_select_out (sw_160_scan_out),
        .latch_enable_out(sw_160_latch_out)
    );

    // [161] https://github.com/mattvenn/wokwi_filler
    wire sw_161_clk_out, sw_161_data_out, sw_161_scan_out, sw_161_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_161 (
        .clk_in          (sw_160_clk_out),
        .data_in         (sw_160_data_out),
        .scan_select_in  (sw_160_scan_out),
        .latch_enable_in (sw_160_latch_out),
        .clk_out         (sw_161_clk_out),
        .data_out        (sw_161_data_out),
        .scan_select_out (sw_161_scan_out),
        .latch_enable_out(sw_161_latch_out)
    );

    // [162] https://github.com/mattvenn/wokwi_filler
    wire sw_162_clk_out, sw_162_data_out, sw_162_scan_out, sw_162_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_162 (
        .clk_in          (sw_161_clk_out),
        .data_in         (sw_161_data_out),
        .scan_select_in  (sw_161_scan_out),
        .latch_enable_in (sw_161_latch_out),
        .clk_out         (sw_162_clk_out),
        .data_out        (sw_162_data_out),
        .scan_select_out (sw_162_scan_out),
        .latch_enable_out(sw_162_latch_out)
    );

    // [163] https://github.com/mattvenn/wokwi_filler
    wire sw_163_clk_out, sw_163_data_out, sw_163_scan_out, sw_163_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_163 (
        .clk_in          (sw_162_clk_out),
        .data_in         (sw_162_data_out),
        .scan_select_in  (sw_162_scan_out),
        .latch_enable_in (sw_162_latch_out),
        .clk_out         (sw_163_clk_out),
        .data_out        (sw_163_data_out),
        .scan_select_out (sw_163_scan_out),
        .latch_enable_out(sw_163_latch_out)
    );

    // [164] https://github.com/mattvenn/wokwi_filler
    wire sw_164_clk_out, sw_164_data_out, sw_164_scan_out, sw_164_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_164 (
        .clk_in          (sw_163_clk_out),
        .data_in         (sw_163_data_out),
        .scan_select_in  (sw_163_scan_out),
        .latch_enable_in (sw_163_latch_out),
        .clk_out         (sw_164_clk_out),
        .data_out        (sw_164_data_out),
        .scan_select_out (sw_164_scan_out),
        .latch_enable_out(sw_164_latch_out)
    );

    // [165] https://github.com/mattvenn/wokwi_filler
    wire sw_165_clk_out, sw_165_data_out, sw_165_scan_out, sw_165_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_165 (
        .clk_in          (sw_164_clk_out),
        .data_in         (sw_164_data_out),
        .scan_select_in  (sw_164_scan_out),
        .latch_enable_in (sw_164_latch_out),
        .clk_out         (sw_165_clk_out),
        .data_out        (sw_165_data_out),
        .scan_select_out (sw_165_scan_out),
        .latch_enable_out(sw_165_latch_out)
    );

    // [166] https://github.com/mattvenn/wokwi_filler
    wire sw_166_clk_out, sw_166_data_out, sw_166_scan_out, sw_166_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_166 (
        .clk_in          (sw_165_clk_out),
        .data_in         (sw_165_data_out),
        .scan_select_in  (sw_165_scan_out),
        .latch_enable_in (sw_165_latch_out),
        .clk_out         (sw_166_clk_out),
        .data_out        (sw_166_data_out),
        .scan_select_out (sw_166_scan_out),
        .latch_enable_out(sw_166_latch_out)
    );

    // [167] https://github.com/mattvenn/wokwi_filler
    wire sw_167_clk_out, sw_167_data_out, sw_167_scan_out, sw_167_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_167 (
        .clk_in          (sw_166_clk_out),
        .data_in         (sw_166_data_out),
        .scan_select_in  (sw_166_scan_out),
        .latch_enable_in (sw_166_latch_out),
        .clk_out         (sw_167_clk_out),
        .data_out        (sw_167_data_out),
        .scan_select_out (sw_167_scan_out),
        .latch_enable_out(sw_167_latch_out)
    );

    // [168] https://github.com/mattvenn/wokwi_filler
    wire sw_168_clk_out, sw_168_data_out, sw_168_scan_out, sw_168_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_168 (
        .clk_in          (sw_167_clk_out),
        .data_in         (sw_167_data_out),
        .scan_select_in  (sw_167_scan_out),
        .latch_enable_in (sw_167_latch_out),
        .clk_out         (sw_168_clk_out),
        .data_out        (sw_168_data_out),
        .scan_select_out (sw_168_scan_out),
        .latch_enable_out(sw_168_latch_out)
    );

    // [169] https://github.com/mattvenn/wokwi_filler
    wire sw_169_clk_out, sw_169_data_out, sw_169_scan_out, sw_169_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_169 (
        .clk_in          (sw_168_clk_out),
        .data_in         (sw_168_data_out),
        .scan_select_in  (sw_168_scan_out),
        .latch_enable_in (sw_168_latch_out),
        .clk_out         (sw_169_clk_out),
        .data_out        (sw_169_data_out),
        .scan_select_out (sw_169_scan_out),
        .latch_enable_out(sw_169_latch_out)
    );

    // [170] https://github.com/mattvenn/wokwi_filler
    wire sw_170_clk_out, sw_170_data_out, sw_170_scan_out, sw_170_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_170 (
        .clk_in          (sw_169_clk_out),
        .data_in         (sw_169_data_out),
        .scan_select_in  (sw_169_scan_out),
        .latch_enable_in (sw_169_latch_out),
        .clk_out         (sw_170_clk_out),
        .data_out        (sw_170_data_out),
        .scan_select_out (sw_170_scan_out),
        .latch_enable_out(sw_170_latch_out)
    );

    // [171] https://github.com/mattvenn/wokwi_filler
    wire sw_171_clk_out, sw_171_data_out, sw_171_scan_out, sw_171_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_171 (
        .clk_in          (sw_170_clk_out),
        .data_in         (sw_170_data_out),
        .scan_select_in  (sw_170_scan_out),
        .latch_enable_in (sw_170_latch_out),
        .clk_out         (sw_171_clk_out),
        .data_out        (sw_171_data_out),
        .scan_select_out (sw_171_scan_out),
        .latch_enable_out(sw_171_latch_out)
    );

    // [172] https://github.com/mattvenn/wokwi_filler
    wire sw_172_clk_out, sw_172_data_out, sw_172_scan_out, sw_172_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_172 (
        .clk_in          (sw_171_clk_out),
        .data_in         (sw_171_data_out),
        .scan_select_in  (sw_171_scan_out),
        .latch_enable_in (sw_171_latch_out),
        .clk_out         (sw_172_clk_out),
        .data_out        (sw_172_data_out),
        .scan_select_out (sw_172_scan_out),
        .latch_enable_out(sw_172_latch_out)
    );

    // [173] https://github.com/mattvenn/wokwi_filler
    wire sw_173_clk_out, sw_173_data_out, sw_173_scan_out, sw_173_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_173 (
        .clk_in          (sw_172_clk_out),
        .data_in         (sw_172_data_out),
        .scan_select_in  (sw_172_scan_out),
        .latch_enable_in (sw_172_latch_out),
        .clk_out         (sw_173_clk_out),
        .data_out        (sw_173_data_out),
        .scan_select_out (sw_173_scan_out),
        .latch_enable_out(sw_173_latch_out)
    );

    // [174] https://github.com/mattvenn/wokwi_filler
    wire sw_174_clk_out, sw_174_data_out, sw_174_scan_out, sw_174_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_174 (
        .clk_in          (sw_173_clk_out),
        .data_in         (sw_173_data_out),
        .scan_select_in  (sw_173_scan_out),
        .latch_enable_in (sw_173_latch_out),
        .clk_out         (sw_174_clk_out),
        .data_out        (sw_174_data_out),
        .scan_select_out (sw_174_scan_out),
        .latch_enable_out(sw_174_latch_out)
    );

    // [175] https://github.com/mattvenn/wokwi_filler
    wire sw_175_clk_out, sw_175_data_out, sw_175_scan_out, sw_175_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_175 (
        .clk_in          (sw_174_clk_out),
        .data_in         (sw_174_data_out),
        .scan_select_in  (sw_174_scan_out),
        .latch_enable_in (sw_174_latch_out),
        .clk_out         (sw_175_clk_out),
        .data_out        (sw_175_data_out),
        .scan_select_out (sw_175_scan_out),
        .latch_enable_out(sw_175_latch_out)
    );

    // [176] https://github.com/mattvenn/wokwi_filler
    wire sw_176_clk_out, sw_176_data_out, sw_176_scan_out, sw_176_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_176 (
        .clk_in          (sw_175_clk_out),
        .data_in         (sw_175_data_out),
        .scan_select_in  (sw_175_scan_out),
        .latch_enable_in (sw_175_latch_out),
        .clk_out         (sw_176_clk_out),
        .data_out        (sw_176_data_out),
        .scan_select_out (sw_176_scan_out),
        .latch_enable_out(sw_176_latch_out)
    );

    // [177] https://github.com/mattvenn/wokwi_filler
    wire sw_177_clk_out, sw_177_data_out, sw_177_scan_out, sw_177_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_177 (
        .clk_in          (sw_176_clk_out),
        .data_in         (sw_176_data_out),
        .scan_select_in  (sw_176_scan_out),
        .latch_enable_in (sw_176_latch_out),
        .clk_out         (sw_177_clk_out),
        .data_out        (sw_177_data_out),
        .scan_select_out (sw_177_scan_out),
        .latch_enable_out(sw_177_latch_out)
    );

    // [178] https://github.com/mattvenn/wokwi_filler
    wire sw_178_clk_out, sw_178_data_out, sw_178_scan_out, sw_178_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_178 (
        .clk_in          (sw_177_clk_out),
        .data_in         (sw_177_data_out),
        .scan_select_in  (sw_177_scan_out),
        .latch_enable_in (sw_177_latch_out),
        .clk_out         (sw_178_clk_out),
        .data_out        (sw_178_data_out),
        .scan_select_out (sw_178_scan_out),
        .latch_enable_out(sw_178_latch_out)
    );

    // [179] https://github.com/mattvenn/wokwi_filler
    wire sw_179_clk_out, sw_179_data_out, sw_179_scan_out, sw_179_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_179 (
        .clk_in          (sw_178_clk_out),
        .data_in         (sw_178_data_out),
        .scan_select_in  (sw_178_scan_out),
        .latch_enable_in (sw_178_latch_out),
        .clk_out         (sw_179_clk_out),
        .data_out        (sw_179_data_out),
        .scan_select_out (sw_179_scan_out),
        .latch_enable_out(sw_179_latch_out)
    );

    // [180] https://github.com/mattvenn/wokwi_filler
    wire sw_180_clk_out, sw_180_data_out, sw_180_scan_out, sw_180_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_180 (
        .clk_in          (sw_179_clk_out),
        .data_in         (sw_179_data_out),
        .scan_select_in  (sw_179_scan_out),
        .latch_enable_in (sw_179_latch_out),
        .clk_out         (sw_180_clk_out),
        .data_out        (sw_180_data_out),
        .scan_select_out (sw_180_scan_out),
        .latch_enable_out(sw_180_latch_out)
    );

    // [181] https://github.com/mattvenn/wokwi_filler
    wire sw_181_clk_out, sw_181_data_out, sw_181_scan_out, sw_181_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_181 (
        .clk_in          (sw_180_clk_out),
        .data_in         (sw_180_data_out),
        .scan_select_in  (sw_180_scan_out),
        .latch_enable_in (sw_180_latch_out),
        .clk_out         (sw_181_clk_out),
        .data_out        (sw_181_data_out),
        .scan_select_out (sw_181_scan_out),
        .latch_enable_out(sw_181_latch_out)
    );

    // [182] https://github.com/mattvenn/wokwi_filler
    wire sw_182_clk_out, sw_182_data_out, sw_182_scan_out, sw_182_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_182 (
        .clk_in          (sw_181_clk_out),
        .data_in         (sw_181_data_out),
        .scan_select_in  (sw_181_scan_out),
        .latch_enable_in (sw_181_latch_out),
        .clk_out         (sw_182_clk_out),
        .data_out        (sw_182_data_out),
        .scan_select_out (sw_182_scan_out),
        .latch_enable_out(sw_182_latch_out)
    );

    // [183] https://github.com/mattvenn/wokwi_filler
    wire sw_183_clk_out, sw_183_data_out, sw_183_scan_out, sw_183_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_183 (
        .clk_in          (sw_182_clk_out),
        .data_in         (sw_182_data_out),
        .scan_select_in  (sw_182_scan_out),
        .latch_enable_in (sw_182_latch_out),
        .clk_out         (sw_183_clk_out),
        .data_out        (sw_183_data_out),
        .scan_select_out (sw_183_scan_out),
        .latch_enable_out(sw_183_latch_out)
    );

    // [184] https://github.com/mattvenn/wokwi_filler
    wire sw_184_clk_out, sw_184_data_out, sw_184_scan_out, sw_184_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_184 (
        .clk_in          (sw_183_clk_out),
        .data_in         (sw_183_data_out),
        .scan_select_in  (sw_183_scan_out),
        .latch_enable_in (sw_183_latch_out),
        .clk_out         (sw_184_clk_out),
        .data_out        (sw_184_data_out),
        .scan_select_out (sw_184_scan_out),
        .latch_enable_out(sw_184_latch_out)
    );

    // [185] https://github.com/mattvenn/wokwi_filler
    wire sw_185_clk_out, sw_185_data_out, sw_185_scan_out, sw_185_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_185 (
        .clk_in          (sw_184_clk_out),
        .data_in         (sw_184_data_out),
        .scan_select_in  (sw_184_scan_out),
        .latch_enable_in (sw_184_latch_out),
        .clk_out         (sw_185_clk_out),
        .data_out        (sw_185_data_out),
        .scan_select_out (sw_185_scan_out),
        .latch_enable_out(sw_185_latch_out)
    );

    // [186] https://github.com/mattvenn/wokwi_filler
    wire sw_186_clk_out, sw_186_data_out, sw_186_scan_out, sw_186_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_186 (
        .clk_in          (sw_185_clk_out),
        .data_in         (sw_185_data_out),
        .scan_select_in  (sw_185_scan_out),
        .latch_enable_in (sw_185_latch_out),
        .clk_out         (sw_186_clk_out),
        .data_out        (sw_186_data_out),
        .scan_select_out (sw_186_scan_out),
        .latch_enable_out(sw_186_latch_out)
    );

    // [187] https://github.com/mattvenn/wokwi_filler
    wire sw_187_clk_out, sw_187_data_out, sw_187_scan_out, sw_187_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_187 (
        .clk_in          (sw_186_clk_out),
        .data_in         (sw_186_data_out),
        .scan_select_in  (sw_186_scan_out),
        .latch_enable_in (sw_186_latch_out),
        .clk_out         (sw_187_clk_out),
        .data_out        (sw_187_data_out),
        .scan_select_out (sw_187_scan_out),
        .latch_enable_out(sw_187_latch_out)
    );

    // [188] https://github.com/mattvenn/wokwi_filler
    wire sw_188_clk_out, sw_188_data_out, sw_188_scan_out, sw_188_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_188 (
        .clk_in          (sw_187_clk_out),
        .data_in         (sw_187_data_out),
        .scan_select_in  (sw_187_scan_out),
        .latch_enable_in (sw_187_latch_out),
        .clk_out         (sw_188_clk_out),
        .data_out        (sw_188_data_out),
        .scan_select_out (sw_188_scan_out),
        .latch_enable_out(sw_188_latch_out)
    );

    // [189] https://github.com/mattvenn/wokwi_filler
    wire sw_189_clk_out, sw_189_data_out, sw_189_scan_out, sw_189_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_189 (
        .clk_in          (sw_188_clk_out),
        .data_in         (sw_188_data_out),
        .scan_select_in  (sw_188_scan_out),
        .latch_enable_in (sw_188_latch_out),
        .clk_out         (sw_189_clk_out),
        .data_out        (sw_189_data_out),
        .scan_select_out (sw_189_scan_out),
        .latch_enable_out(sw_189_latch_out)
    );

    // [190] https://github.com/mattvenn/wokwi_filler
    wire sw_190_clk_out, sw_190_data_out, sw_190_scan_out, sw_190_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_190 (
        .clk_in          (sw_189_clk_out),
        .data_in         (sw_189_data_out),
        .scan_select_in  (sw_189_scan_out),
        .latch_enable_in (sw_189_latch_out),
        .clk_out         (sw_190_clk_out),
        .data_out        (sw_190_data_out),
        .scan_select_out (sw_190_scan_out),
        .latch_enable_out(sw_190_latch_out)
    );

    // [191] https://github.com/mattvenn/wokwi_filler
    wire sw_191_clk_out, sw_191_data_out, sw_191_scan_out, sw_191_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_191 (
        .clk_in          (sw_190_clk_out),
        .data_in         (sw_190_data_out),
        .scan_select_in  (sw_190_scan_out),
        .latch_enable_in (sw_190_latch_out),
        .clk_out         (sw_191_clk_out),
        .data_out        (sw_191_data_out),
        .scan_select_out (sw_191_scan_out),
        .latch_enable_out(sw_191_latch_out)
    );

    // [192] https://github.com/mattvenn/wokwi_filler
    wire sw_192_clk_out, sw_192_data_out, sw_192_scan_out, sw_192_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_192 (
        .clk_in          (sw_191_clk_out),
        .data_in         (sw_191_data_out),
        .scan_select_in  (sw_191_scan_out),
        .latch_enable_in (sw_191_latch_out),
        .clk_out         (sw_192_clk_out),
        .data_out        (sw_192_data_out),
        .scan_select_out (sw_192_scan_out),
        .latch_enable_out(sw_192_latch_out)
    );

    // [193] https://github.com/mattvenn/wokwi_filler
    wire sw_193_clk_out, sw_193_data_out, sw_193_scan_out, sw_193_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_193 (
        .clk_in          (sw_192_clk_out),
        .data_in         (sw_192_data_out),
        .scan_select_in  (sw_192_scan_out),
        .latch_enable_in (sw_192_latch_out),
        .clk_out         (sw_193_clk_out),
        .data_out        (sw_193_data_out),
        .scan_select_out (sw_193_scan_out),
        .latch_enable_out(sw_193_latch_out)
    );

    // [194] https://github.com/mattvenn/wokwi_filler
    wire sw_194_clk_out, sw_194_data_out, sw_194_scan_out, sw_194_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_194 (
        .clk_in          (sw_193_clk_out),
        .data_in         (sw_193_data_out),
        .scan_select_in  (sw_193_scan_out),
        .latch_enable_in (sw_193_latch_out),
        .clk_out         (sw_194_clk_out),
        .data_out        (sw_194_data_out),
        .scan_select_out (sw_194_scan_out),
        .latch_enable_out(sw_194_latch_out)
    );

    // [195] https://github.com/mattvenn/wokwi_filler
    wire sw_195_clk_out, sw_195_data_out, sw_195_scan_out, sw_195_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_195 (
        .clk_in          (sw_194_clk_out),
        .data_in         (sw_194_data_out),
        .scan_select_in  (sw_194_scan_out),
        .latch_enable_in (sw_194_latch_out),
        .clk_out         (sw_195_clk_out),
        .data_out        (sw_195_data_out),
        .scan_select_out (sw_195_scan_out),
        .latch_enable_out(sw_195_latch_out)
    );

    // [196] https://github.com/mattvenn/wokwi_filler
    wire sw_196_clk_out, sw_196_data_out, sw_196_scan_out, sw_196_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_196 (
        .clk_in          (sw_195_clk_out),
        .data_in         (sw_195_data_out),
        .scan_select_in  (sw_195_scan_out),
        .latch_enable_in (sw_195_latch_out),
        .clk_out         (sw_196_clk_out),
        .data_out        (sw_196_data_out),
        .scan_select_out (sw_196_scan_out),
        .latch_enable_out(sw_196_latch_out)
    );

    // [197] https://github.com/mattvenn/wokwi_filler
    wire sw_197_clk_out, sw_197_data_out, sw_197_scan_out, sw_197_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_197 (
        .clk_in          (sw_196_clk_out),
        .data_in         (sw_196_data_out),
        .scan_select_in  (sw_196_scan_out),
        .latch_enable_in (sw_196_latch_out),
        .clk_out         (sw_197_clk_out),
        .data_out        (sw_197_data_out),
        .scan_select_out (sw_197_scan_out),
        .latch_enable_out(sw_197_latch_out)
    );

    // [198] https://github.com/mattvenn/wokwi_filler
    wire sw_198_clk_out, sw_198_data_out, sw_198_scan_out, sw_198_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_198 (
        .clk_in          (sw_197_clk_out),
        .data_in         (sw_197_data_out),
        .scan_select_in  (sw_197_scan_out),
        .latch_enable_in (sw_197_latch_out),
        .clk_out         (sw_198_clk_out),
        .data_out        (sw_198_data_out),
        .scan_select_out (sw_198_scan_out),
        .latch_enable_out(sw_198_latch_out)
    );

    // [199] https://github.com/mattvenn/wokwi_filler
    wire sw_199_clk_out, sw_199_data_out, sw_199_scan_out, sw_199_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_199 (
        .clk_in          (sw_198_clk_out),
        .data_in         (sw_198_data_out),
        .scan_select_in  (sw_198_scan_out),
        .latch_enable_in (sw_198_latch_out),
        .clk_out         (sw_199_clk_out),
        .data_out        (sw_199_data_out),
        .scan_select_out (sw_199_scan_out),
        .latch_enable_out(sw_199_latch_out)
    );

    // [200] https://github.com/mattvenn/wokwi_filler
    wire sw_200_clk_out, sw_200_data_out, sw_200_scan_out, sw_200_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_200 (
        .clk_in          (sw_199_clk_out),
        .data_in         (sw_199_data_out),
        .scan_select_in  (sw_199_scan_out),
        .latch_enable_in (sw_199_latch_out),
        .clk_out         (sw_200_clk_out),
        .data_out        (sw_200_data_out),
        .scan_select_out (sw_200_scan_out),
        .latch_enable_out(sw_200_latch_out)
    );

    // [201] https://github.com/mattvenn/wokwi_filler
    wire sw_201_clk_out, sw_201_data_out, sw_201_scan_out, sw_201_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_201 (
        .clk_in          (sw_200_clk_out),
        .data_in         (sw_200_data_out),
        .scan_select_in  (sw_200_scan_out),
        .latch_enable_in (sw_200_latch_out),
        .clk_out         (sw_201_clk_out),
        .data_out        (sw_201_data_out),
        .scan_select_out (sw_201_scan_out),
        .latch_enable_out(sw_201_latch_out)
    );

    // [202] https://github.com/mattvenn/wokwi_filler
    wire sw_202_clk_out, sw_202_data_out, sw_202_scan_out, sw_202_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_202 (
        .clk_in          (sw_201_clk_out),
        .data_in         (sw_201_data_out),
        .scan_select_in  (sw_201_scan_out),
        .latch_enable_in (sw_201_latch_out),
        .clk_out         (sw_202_clk_out),
        .data_out        (sw_202_data_out),
        .scan_select_out (sw_202_scan_out),
        .latch_enable_out(sw_202_latch_out)
    );

    // [203] https://github.com/mattvenn/wokwi_filler
    wire sw_203_clk_out, sw_203_data_out, sw_203_scan_out, sw_203_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_203 (
        .clk_in          (sw_202_clk_out),
        .data_in         (sw_202_data_out),
        .scan_select_in  (sw_202_scan_out),
        .latch_enable_in (sw_202_latch_out),
        .clk_out         (sw_203_clk_out),
        .data_out        (sw_203_data_out),
        .scan_select_out (sw_203_scan_out),
        .latch_enable_out(sw_203_latch_out)
    );

    // [204] https://github.com/mattvenn/wokwi_filler
    wire sw_204_clk_out, sw_204_data_out, sw_204_scan_out, sw_204_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_204 (
        .clk_in          (sw_203_clk_out),
        .data_in         (sw_203_data_out),
        .scan_select_in  (sw_203_scan_out),
        .latch_enable_in (sw_203_latch_out),
        .clk_out         (sw_204_clk_out),
        .data_out        (sw_204_data_out),
        .scan_select_out (sw_204_scan_out),
        .latch_enable_out(sw_204_latch_out)
    );

    // [205] https://github.com/mattvenn/wokwi_filler
    wire sw_205_clk_out, sw_205_data_out, sw_205_scan_out, sw_205_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_205 (
        .clk_in          (sw_204_clk_out),
        .data_in         (sw_204_data_out),
        .scan_select_in  (sw_204_scan_out),
        .latch_enable_in (sw_204_latch_out),
        .clk_out         (sw_205_clk_out),
        .data_out        (sw_205_data_out),
        .scan_select_out (sw_205_scan_out),
        .latch_enable_out(sw_205_latch_out)
    );

    // [206] https://github.com/mattvenn/wokwi_filler
    wire sw_206_clk_out, sw_206_data_out, sw_206_scan_out, sw_206_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_206 (
        .clk_in          (sw_205_clk_out),
        .data_in         (sw_205_data_out),
        .scan_select_in  (sw_205_scan_out),
        .latch_enable_in (sw_205_latch_out),
        .clk_out         (sw_206_clk_out),
        .data_out        (sw_206_data_out),
        .scan_select_out (sw_206_scan_out),
        .latch_enable_out(sw_206_latch_out)
    );

    // [207] https://github.com/mattvenn/wokwi_filler
    wire sw_207_clk_out, sw_207_data_out, sw_207_scan_out, sw_207_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_207 (
        .clk_in          (sw_206_clk_out),
        .data_in         (sw_206_data_out),
        .scan_select_in  (sw_206_scan_out),
        .latch_enable_in (sw_206_latch_out),
        .clk_out         (sw_207_clk_out),
        .data_out        (sw_207_data_out),
        .scan_select_out (sw_207_scan_out),
        .latch_enable_out(sw_207_latch_out)
    );

    // [208] https://github.com/mattvenn/wokwi_filler
    wire sw_208_clk_out, sw_208_data_out, sw_208_scan_out, sw_208_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_208 (
        .clk_in          (sw_207_clk_out),
        .data_in         (sw_207_data_out),
        .scan_select_in  (sw_207_scan_out),
        .latch_enable_in (sw_207_latch_out),
        .clk_out         (sw_208_clk_out),
        .data_out        (sw_208_data_out),
        .scan_select_out (sw_208_scan_out),
        .latch_enable_out(sw_208_latch_out)
    );

    // [209] https://github.com/mattvenn/wokwi_filler
    wire sw_209_clk_out, sw_209_data_out, sw_209_scan_out, sw_209_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_209 (
        .clk_in          (sw_208_clk_out),
        .data_in         (sw_208_data_out),
        .scan_select_in  (sw_208_scan_out),
        .latch_enable_in (sw_208_latch_out),
        .clk_out         (sw_209_clk_out),
        .data_out        (sw_209_data_out),
        .scan_select_out (sw_209_scan_out),
        .latch_enable_out(sw_209_latch_out)
    );

    // [210] https://github.com/mattvenn/wokwi_filler
    wire sw_210_clk_out, sw_210_data_out, sw_210_scan_out, sw_210_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_210 (
        .clk_in          (sw_209_clk_out),
        .data_in         (sw_209_data_out),
        .scan_select_in  (sw_209_scan_out),
        .latch_enable_in (sw_209_latch_out),
        .clk_out         (sw_210_clk_out),
        .data_out        (sw_210_data_out),
        .scan_select_out (sw_210_scan_out),
        .latch_enable_out(sw_210_latch_out)
    );

    // [211] https://github.com/mattvenn/wokwi_filler
    wire sw_211_clk_out, sw_211_data_out, sw_211_scan_out, sw_211_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_211 (
        .clk_in          (sw_210_clk_out),
        .data_in         (sw_210_data_out),
        .scan_select_in  (sw_210_scan_out),
        .latch_enable_in (sw_210_latch_out),
        .clk_out         (sw_211_clk_out),
        .data_out        (sw_211_data_out),
        .scan_select_out (sw_211_scan_out),
        .latch_enable_out(sw_211_latch_out)
    );

    // [212] https://github.com/mattvenn/wokwi_filler
    wire sw_212_clk_out, sw_212_data_out, sw_212_scan_out, sw_212_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_212 (
        .clk_in          (sw_211_clk_out),
        .data_in         (sw_211_data_out),
        .scan_select_in  (sw_211_scan_out),
        .latch_enable_in (sw_211_latch_out),
        .clk_out         (sw_212_clk_out),
        .data_out        (sw_212_data_out),
        .scan_select_out (sw_212_scan_out),
        .latch_enable_out(sw_212_latch_out)
    );

    // [213] https://github.com/mattvenn/wokwi_filler
    wire sw_213_clk_out, sw_213_data_out, sw_213_scan_out, sw_213_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_213 (
        .clk_in          (sw_212_clk_out),
        .data_in         (sw_212_data_out),
        .scan_select_in  (sw_212_scan_out),
        .latch_enable_in (sw_212_latch_out),
        .clk_out         (sw_213_clk_out),
        .data_out        (sw_213_data_out),
        .scan_select_out (sw_213_scan_out),
        .latch_enable_out(sw_213_latch_out)
    );

    // [214] https://github.com/mattvenn/wokwi_filler
    wire sw_214_clk_out, sw_214_data_out, sw_214_scan_out, sw_214_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_214 (
        .clk_in          (sw_213_clk_out),
        .data_in         (sw_213_data_out),
        .scan_select_in  (sw_213_scan_out),
        .latch_enable_in (sw_213_latch_out),
        .clk_out         (sw_214_clk_out),
        .data_out        (sw_214_data_out),
        .scan_select_out (sw_214_scan_out),
        .latch_enable_out(sw_214_latch_out)
    );

    // [215] https://github.com/mattvenn/wokwi_filler
    wire sw_215_clk_out, sw_215_data_out, sw_215_scan_out, sw_215_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_215 (
        .clk_in          (sw_214_clk_out),
        .data_in         (sw_214_data_out),
        .scan_select_in  (sw_214_scan_out),
        .latch_enable_in (sw_214_latch_out),
        .clk_out         (sw_215_clk_out),
        .data_out        (sw_215_data_out),
        .scan_select_out (sw_215_scan_out),
        .latch_enable_out(sw_215_latch_out)
    );

    // [216] https://github.com/mattvenn/wokwi_filler
    wire sw_216_clk_out, sw_216_data_out, sw_216_scan_out, sw_216_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_216 (
        .clk_in          (sw_215_clk_out),
        .data_in         (sw_215_data_out),
        .scan_select_in  (sw_215_scan_out),
        .latch_enable_in (sw_215_latch_out),
        .clk_out         (sw_216_clk_out),
        .data_out        (sw_216_data_out),
        .scan_select_out (sw_216_scan_out),
        .latch_enable_out(sw_216_latch_out)
    );

    // [217] https://github.com/mattvenn/wokwi_filler
    wire sw_217_clk_out, sw_217_data_out, sw_217_scan_out, sw_217_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_217 (
        .clk_in          (sw_216_clk_out),
        .data_in         (sw_216_data_out),
        .scan_select_in  (sw_216_scan_out),
        .latch_enable_in (sw_216_latch_out),
        .clk_out         (sw_217_clk_out),
        .data_out        (sw_217_data_out),
        .scan_select_out (sw_217_scan_out),
        .latch_enable_out(sw_217_latch_out)
    );

    // [218] https://github.com/mattvenn/wokwi_filler
    wire sw_218_clk_out, sw_218_data_out, sw_218_scan_out, sw_218_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_218 (
        .clk_in          (sw_217_clk_out),
        .data_in         (sw_217_data_out),
        .scan_select_in  (sw_217_scan_out),
        .latch_enable_in (sw_217_latch_out),
        .clk_out         (sw_218_clk_out),
        .data_out        (sw_218_data_out),
        .scan_select_out (sw_218_scan_out),
        .latch_enable_out(sw_218_latch_out)
    );

    // [219] https://github.com/mattvenn/wokwi_filler
    wire sw_219_clk_out, sw_219_data_out, sw_219_scan_out, sw_219_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_219 (
        .clk_in          (sw_218_clk_out),
        .data_in         (sw_218_data_out),
        .scan_select_in  (sw_218_scan_out),
        .latch_enable_in (sw_218_latch_out),
        .clk_out         (sw_219_clk_out),
        .data_out        (sw_219_data_out),
        .scan_select_out (sw_219_scan_out),
        .latch_enable_out(sw_219_latch_out)
    );

    // [220] https://github.com/mattvenn/wokwi_filler
    wire sw_220_clk_out, sw_220_data_out, sw_220_scan_out, sw_220_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_220 (
        .clk_in          (sw_219_clk_out),
        .data_in         (sw_219_data_out),
        .scan_select_in  (sw_219_scan_out),
        .latch_enable_in (sw_219_latch_out),
        .clk_out         (sw_220_clk_out),
        .data_out        (sw_220_data_out),
        .scan_select_out (sw_220_scan_out),
        .latch_enable_out(sw_220_latch_out)
    );

    // [221] https://github.com/mattvenn/wokwi_filler
    wire sw_221_clk_out, sw_221_data_out, sw_221_scan_out, sw_221_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_221 (
        .clk_in          (sw_220_clk_out),
        .data_in         (sw_220_data_out),
        .scan_select_in  (sw_220_scan_out),
        .latch_enable_in (sw_220_latch_out),
        .clk_out         (sw_221_clk_out),
        .data_out        (sw_221_data_out),
        .scan_select_out (sw_221_scan_out),
        .latch_enable_out(sw_221_latch_out)
    );

    // [222] https://github.com/mattvenn/wokwi_filler
    wire sw_222_clk_out, sw_222_data_out, sw_222_scan_out, sw_222_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_222 (
        .clk_in          (sw_221_clk_out),
        .data_in         (sw_221_data_out),
        .scan_select_in  (sw_221_scan_out),
        .latch_enable_in (sw_221_latch_out),
        .clk_out         (sw_222_clk_out),
        .data_out        (sw_222_data_out),
        .scan_select_out (sw_222_scan_out),
        .latch_enable_out(sw_222_latch_out)
    );

    // [223] https://github.com/mattvenn/wokwi_filler
    wire sw_223_clk_out, sw_223_data_out, sw_223_scan_out, sw_223_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_223 (
        .clk_in          (sw_222_clk_out),
        .data_in         (sw_222_data_out),
        .scan_select_in  (sw_222_scan_out),
        .latch_enable_in (sw_222_latch_out),
        .clk_out         (sw_223_clk_out),
        .data_out        (sw_223_data_out),
        .scan_select_out (sw_223_scan_out),
        .latch_enable_out(sw_223_latch_out)
    );

    // [224] https://github.com/mattvenn/wokwi_filler
    wire sw_224_clk_out, sw_224_data_out, sw_224_scan_out, sw_224_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_224 (
        .clk_in          (sw_223_clk_out),
        .data_in         (sw_223_data_out),
        .scan_select_in  (sw_223_scan_out),
        .latch_enable_in (sw_223_latch_out),
        .clk_out         (sw_224_clk_out),
        .data_out        (sw_224_data_out),
        .scan_select_out (sw_224_scan_out),
        .latch_enable_out(sw_224_latch_out)
    );

    // [225] https://github.com/mattvenn/wokwi_filler
    wire sw_225_clk_out, sw_225_data_out, sw_225_scan_out, sw_225_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_225 (
        .clk_in          (sw_224_clk_out),
        .data_in         (sw_224_data_out),
        .scan_select_in  (sw_224_scan_out),
        .latch_enable_in (sw_224_latch_out),
        .clk_out         (sw_225_clk_out),
        .data_out        (sw_225_data_out),
        .scan_select_out (sw_225_scan_out),
        .latch_enable_out(sw_225_latch_out)
    );

    // [226] https://github.com/mattvenn/wokwi_filler
    wire sw_226_clk_out, sw_226_data_out, sw_226_scan_out, sw_226_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_226 (
        .clk_in          (sw_225_clk_out),
        .data_in         (sw_225_data_out),
        .scan_select_in  (sw_225_scan_out),
        .latch_enable_in (sw_225_latch_out),
        .clk_out         (sw_226_clk_out),
        .data_out        (sw_226_data_out),
        .scan_select_out (sw_226_scan_out),
        .latch_enable_out(sw_226_latch_out)
    );

    // [227] https://github.com/mattvenn/wokwi_filler
    wire sw_227_clk_out, sw_227_data_out, sw_227_scan_out, sw_227_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_227 (
        .clk_in          (sw_226_clk_out),
        .data_in         (sw_226_data_out),
        .scan_select_in  (sw_226_scan_out),
        .latch_enable_in (sw_226_latch_out),
        .clk_out         (sw_227_clk_out),
        .data_out        (sw_227_data_out),
        .scan_select_out (sw_227_scan_out),
        .latch_enable_out(sw_227_latch_out)
    );

    // [228] https://github.com/mattvenn/wokwi_filler
    wire sw_228_clk_out, sw_228_data_out, sw_228_scan_out, sw_228_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_228 (
        .clk_in          (sw_227_clk_out),
        .data_in         (sw_227_data_out),
        .scan_select_in  (sw_227_scan_out),
        .latch_enable_in (sw_227_latch_out),
        .clk_out         (sw_228_clk_out),
        .data_out        (sw_228_data_out),
        .scan_select_out (sw_228_scan_out),
        .latch_enable_out(sw_228_latch_out)
    );

    // [229] https://github.com/mattvenn/wokwi_filler
    wire sw_229_clk_out, sw_229_data_out, sw_229_scan_out, sw_229_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_229 (
        .clk_in          (sw_228_clk_out),
        .data_in         (sw_228_data_out),
        .scan_select_in  (sw_228_scan_out),
        .latch_enable_in (sw_228_latch_out),
        .clk_out         (sw_229_clk_out),
        .data_out        (sw_229_data_out),
        .scan_select_out (sw_229_scan_out),
        .latch_enable_out(sw_229_latch_out)
    );

    // [230] https://github.com/mattvenn/wokwi_filler
    wire sw_230_clk_out, sw_230_data_out, sw_230_scan_out, sw_230_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_230 (
        .clk_in          (sw_229_clk_out),
        .data_in         (sw_229_data_out),
        .scan_select_in  (sw_229_scan_out),
        .latch_enable_in (sw_229_latch_out),
        .clk_out         (sw_230_clk_out),
        .data_out        (sw_230_data_out),
        .scan_select_out (sw_230_scan_out),
        .latch_enable_out(sw_230_latch_out)
    );

    // [231] https://github.com/mattvenn/wokwi_filler
    wire sw_231_clk_out, sw_231_data_out, sw_231_scan_out, sw_231_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_231 (
        .clk_in          (sw_230_clk_out),
        .data_in         (sw_230_data_out),
        .scan_select_in  (sw_230_scan_out),
        .latch_enable_in (sw_230_latch_out),
        .clk_out         (sw_231_clk_out),
        .data_out        (sw_231_data_out),
        .scan_select_out (sw_231_scan_out),
        .latch_enable_out(sw_231_latch_out)
    );

    // [232] https://github.com/mattvenn/wokwi_filler
    wire sw_232_clk_out, sw_232_data_out, sw_232_scan_out, sw_232_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_232 (
        .clk_in          (sw_231_clk_out),
        .data_in         (sw_231_data_out),
        .scan_select_in  (sw_231_scan_out),
        .latch_enable_in (sw_231_latch_out),
        .clk_out         (sw_232_clk_out),
        .data_out        (sw_232_data_out),
        .scan_select_out (sw_232_scan_out),
        .latch_enable_out(sw_232_latch_out)
    );

    // [233] https://github.com/mattvenn/wokwi_filler
    wire sw_233_clk_out, sw_233_data_out, sw_233_scan_out, sw_233_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_233 (
        .clk_in          (sw_232_clk_out),
        .data_in         (sw_232_data_out),
        .scan_select_in  (sw_232_scan_out),
        .latch_enable_in (sw_232_latch_out),
        .clk_out         (sw_233_clk_out),
        .data_out        (sw_233_data_out),
        .scan_select_out (sw_233_scan_out),
        .latch_enable_out(sw_233_latch_out)
    );

    // [234] https://github.com/mattvenn/wokwi_filler
    wire sw_234_clk_out, sw_234_data_out, sw_234_scan_out, sw_234_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_234 (
        .clk_in          (sw_233_clk_out),
        .data_in         (sw_233_data_out),
        .scan_select_in  (sw_233_scan_out),
        .latch_enable_in (sw_233_latch_out),
        .clk_out         (sw_234_clk_out),
        .data_out        (sw_234_data_out),
        .scan_select_out (sw_234_scan_out),
        .latch_enable_out(sw_234_latch_out)
    );

    // [235] https://github.com/mattvenn/wokwi_filler
    wire sw_235_clk_out, sw_235_data_out, sw_235_scan_out, sw_235_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_235 (
        .clk_in          (sw_234_clk_out),
        .data_in         (sw_234_data_out),
        .scan_select_in  (sw_234_scan_out),
        .latch_enable_in (sw_234_latch_out),
        .clk_out         (sw_235_clk_out),
        .data_out        (sw_235_data_out),
        .scan_select_out (sw_235_scan_out),
        .latch_enable_out(sw_235_latch_out)
    );

    // [236] https://github.com/mattvenn/wokwi_filler
    wire sw_236_clk_out, sw_236_data_out, sw_236_scan_out, sw_236_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_236 (
        .clk_in          (sw_235_clk_out),
        .data_in         (sw_235_data_out),
        .scan_select_in  (sw_235_scan_out),
        .latch_enable_in (sw_235_latch_out),
        .clk_out         (sw_236_clk_out),
        .data_out        (sw_236_data_out),
        .scan_select_out (sw_236_scan_out),
        .latch_enable_out(sw_236_latch_out)
    );

    // [237] https://github.com/mattvenn/wokwi_filler
    wire sw_237_clk_out, sw_237_data_out, sw_237_scan_out, sw_237_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_237 (
        .clk_in          (sw_236_clk_out),
        .data_in         (sw_236_data_out),
        .scan_select_in  (sw_236_scan_out),
        .latch_enable_in (sw_236_latch_out),
        .clk_out         (sw_237_clk_out),
        .data_out        (sw_237_data_out),
        .scan_select_out (sw_237_scan_out),
        .latch_enable_out(sw_237_latch_out)
    );

    // [238] https://github.com/mattvenn/wokwi_filler
    wire sw_238_clk_out, sw_238_data_out, sw_238_scan_out, sw_238_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_238 (
        .clk_in          (sw_237_clk_out),
        .data_in         (sw_237_data_out),
        .scan_select_in  (sw_237_scan_out),
        .latch_enable_in (sw_237_latch_out),
        .clk_out         (sw_238_clk_out),
        .data_out        (sw_238_data_out),
        .scan_select_out (sw_238_scan_out),
        .latch_enable_out(sw_238_latch_out)
    );

    // [239] https://github.com/mattvenn/wokwi_filler
    wire sw_239_clk_out, sw_239_data_out, sw_239_scan_out, sw_239_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_239 (
        .clk_in          (sw_238_clk_out),
        .data_in         (sw_238_data_out),
        .scan_select_in  (sw_238_scan_out),
        .latch_enable_in (sw_238_latch_out),
        .clk_out         (sw_239_clk_out),
        .data_out        (sw_239_data_out),
        .scan_select_out (sw_239_scan_out),
        .latch_enable_out(sw_239_latch_out)
    );

    // [240] https://github.com/mattvenn/wokwi_filler
    wire sw_240_clk_out, sw_240_data_out, sw_240_scan_out, sw_240_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_240 (
        .clk_in          (sw_239_clk_out),
        .data_in         (sw_239_data_out),
        .scan_select_in  (sw_239_scan_out),
        .latch_enable_in (sw_239_latch_out),
        .clk_out         (sw_240_clk_out),
        .data_out        (sw_240_data_out),
        .scan_select_out (sw_240_scan_out),
        .latch_enable_out(sw_240_latch_out)
    );

    // [241] https://github.com/mattvenn/wokwi_filler
    wire sw_241_clk_out, sw_241_data_out, sw_241_scan_out, sw_241_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_241 (
        .clk_in          (sw_240_clk_out),
        .data_in         (sw_240_data_out),
        .scan_select_in  (sw_240_scan_out),
        .latch_enable_in (sw_240_latch_out),
        .clk_out         (sw_241_clk_out),
        .data_out        (sw_241_data_out),
        .scan_select_out (sw_241_scan_out),
        .latch_enable_out(sw_241_latch_out)
    );

    // [242] https://github.com/mattvenn/wokwi_filler
    wire sw_242_clk_out, sw_242_data_out, sw_242_scan_out, sw_242_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_242 (
        .clk_in          (sw_241_clk_out),
        .data_in         (sw_241_data_out),
        .scan_select_in  (sw_241_scan_out),
        .latch_enable_in (sw_241_latch_out),
        .clk_out         (sw_242_clk_out),
        .data_out        (sw_242_data_out),
        .scan_select_out (sw_242_scan_out),
        .latch_enable_out(sw_242_latch_out)
    );

    // [243] https://github.com/mattvenn/wokwi_filler
    wire sw_243_clk_out, sw_243_data_out, sw_243_scan_out, sw_243_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_243 (
        .clk_in          (sw_242_clk_out),
        .data_in         (sw_242_data_out),
        .scan_select_in  (sw_242_scan_out),
        .latch_enable_in (sw_242_latch_out),
        .clk_out         (sw_243_clk_out),
        .data_out        (sw_243_data_out),
        .scan_select_out (sw_243_scan_out),
        .latch_enable_out(sw_243_latch_out)
    );

    // [244] https://github.com/mattvenn/wokwi_filler
    wire sw_244_clk_out, sw_244_data_out, sw_244_scan_out, sw_244_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_244 (
        .clk_in          (sw_243_clk_out),
        .data_in         (sw_243_data_out),
        .scan_select_in  (sw_243_scan_out),
        .latch_enable_in (sw_243_latch_out),
        .clk_out         (sw_244_clk_out),
        .data_out        (sw_244_data_out),
        .scan_select_out (sw_244_scan_out),
        .latch_enable_out(sw_244_latch_out)
    );

    // [245] https://github.com/mattvenn/wokwi_filler
    wire sw_245_clk_out, sw_245_data_out, sw_245_scan_out, sw_245_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_245 (
        .clk_in          (sw_244_clk_out),
        .data_in         (sw_244_data_out),
        .scan_select_in  (sw_244_scan_out),
        .latch_enable_in (sw_244_latch_out),
        .clk_out         (sw_245_clk_out),
        .data_out        (sw_245_data_out),
        .scan_select_out (sw_245_scan_out),
        .latch_enable_out(sw_245_latch_out)
    );

    // [246] https://github.com/mattvenn/wokwi_filler
    wire sw_246_clk_out, sw_246_data_out, sw_246_scan_out, sw_246_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_246 (
        .clk_in          (sw_245_clk_out),
        .data_in         (sw_245_data_out),
        .scan_select_in  (sw_245_scan_out),
        .latch_enable_in (sw_245_latch_out),
        .clk_out         (sw_246_clk_out),
        .data_out        (sw_246_data_out),
        .scan_select_out (sw_246_scan_out),
        .latch_enable_out(sw_246_latch_out)
    );

    // [247] https://github.com/mattvenn/wokwi_filler
    wire sw_247_clk_out, sw_247_data_out, sw_247_scan_out, sw_247_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_247 (
        .clk_in          (sw_246_clk_out),
        .data_in         (sw_246_data_out),
        .scan_select_in  (sw_246_scan_out),
        .latch_enable_in (sw_246_latch_out),
        .clk_out         (sw_247_clk_out),
        .data_out        (sw_247_data_out),
        .scan_select_out (sw_247_scan_out),
        .latch_enable_out(sw_247_latch_out)
    );

    // [248] https://github.com/mattvenn/wokwi_filler
    wire sw_248_clk_out, sw_248_data_out, sw_248_scan_out, sw_248_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_248 (
        .clk_in          (sw_247_clk_out),
        .data_in         (sw_247_data_out),
        .scan_select_in  (sw_247_scan_out),
        .latch_enable_in (sw_247_latch_out),
        .clk_out         (sw_248_clk_out),
        .data_out        (sw_248_data_out),
        .scan_select_out (sw_248_scan_out),
        .latch_enable_out(sw_248_latch_out)
    );

    // [249] https://github.com/mattvenn/wokwi_filler
    wire sw_249_clk_out, sw_249_data_out, sw_249_scan_out, sw_249_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_249 (
        .clk_in          (sw_248_clk_out),
        .data_in         (sw_248_data_out),
        .scan_select_in  (sw_248_scan_out),
        .latch_enable_in (sw_248_latch_out),
        .clk_out         (sw_249_clk_out),
        .data_out        (sw_249_data_out),
        .scan_select_out (sw_249_scan_out),
        .latch_enable_out(sw_249_latch_out)
    );

    // [250] https://github.com/mattvenn/wokwi_filler
    wire sw_250_clk_out, sw_250_data_out, sw_250_scan_out, sw_250_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_250 (
        .clk_in          (sw_249_clk_out),
        .data_in         (sw_249_data_out),
        .scan_select_in  (sw_249_scan_out),
        .latch_enable_in (sw_249_latch_out),
        .clk_out         (sw_250_clk_out),
        .data_out        (sw_250_data_out),
        .scan_select_out (sw_250_scan_out),
        .latch_enable_out(sw_250_latch_out)
    );

    // [251] https://github.com/mattvenn/wokwi_filler
    wire sw_251_clk_out, sw_251_data_out, sw_251_scan_out, sw_251_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_251 (
        .clk_in          (sw_250_clk_out),
        .data_in         (sw_250_data_out),
        .scan_select_in  (sw_250_scan_out),
        .latch_enable_in (sw_250_latch_out),
        .clk_out         (sw_251_clk_out),
        .data_out        (sw_251_data_out),
        .scan_select_out (sw_251_scan_out),
        .latch_enable_out(sw_251_latch_out)
    );

    // [252] https://github.com/mattvenn/wokwi_filler
    wire sw_252_clk_out, sw_252_data_out, sw_252_scan_out, sw_252_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_252 (
        .clk_in          (sw_251_clk_out),
        .data_in         (sw_251_data_out),
        .scan_select_in  (sw_251_scan_out),
        .latch_enable_in (sw_251_latch_out),
        .clk_out         (sw_252_clk_out),
        .data_out        (sw_252_data_out),
        .scan_select_out (sw_252_scan_out),
        .latch_enable_out(sw_252_latch_out)
    );

    // [253] https://github.com/mattvenn/wokwi_filler
    wire sw_253_clk_out, sw_253_data_out, sw_253_scan_out, sw_253_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_253 (
        .clk_in          (sw_252_clk_out),
        .data_in         (sw_252_data_out),
        .scan_select_in  (sw_252_scan_out),
        .latch_enable_in (sw_252_latch_out),
        .clk_out         (sw_253_clk_out),
        .data_out        (sw_253_data_out),
        .scan_select_out (sw_253_scan_out),
        .latch_enable_out(sw_253_latch_out)
    );

    // [254] https://github.com/mattvenn/wokwi_filler
    wire sw_254_clk_out, sw_254_data_out, sw_254_scan_out, sw_254_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_254 (
        .clk_in          (sw_253_clk_out),
        .data_in         (sw_253_data_out),
        .scan_select_in  (sw_253_scan_out),
        .latch_enable_in (sw_253_latch_out),
        .clk_out         (sw_254_clk_out),
        .data_out        (sw_254_data_out),
        .scan_select_out (sw_254_scan_out),
        .latch_enable_out(sw_254_latch_out)
    );

    // [255] https://github.com/mattvenn/wokwi_filler
    wire sw_255_clk_out, sw_255_data_out, sw_255_scan_out, sw_255_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_255 (
        .clk_in          (sw_254_clk_out),
        .data_in         (sw_254_data_out),
        .scan_select_in  (sw_254_scan_out),
        .latch_enable_in (sw_254_latch_out),
        .clk_out         (sw_255_clk_out),
        .data_out        (sw_255_data_out),
        .scan_select_out (sw_255_scan_out),
        .latch_enable_out(sw_255_latch_out)
    );

    // [256] https://github.com/mattvenn/wokwi_filler
    wire sw_256_clk_out, sw_256_data_out, sw_256_scan_out, sw_256_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_256 (
        .clk_in          (sw_255_clk_out),
        .data_in         (sw_255_data_out),
        .scan_select_in  (sw_255_scan_out),
        .latch_enable_in (sw_255_latch_out),
        .clk_out         (sw_256_clk_out),
        .data_out        (sw_256_data_out),
        .scan_select_out (sw_256_scan_out),
        .latch_enable_out(sw_256_latch_out)
    );

    // [257] https://github.com/mattvenn/wokwi_filler
    wire sw_257_clk_out, sw_257_data_out, sw_257_scan_out, sw_257_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_257 (
        .clk_in          (sw_256_clk_out),
        .data_in         (sw_256_data_out),
        .scan_select_in  (sw_256_scan_out),
        .latch_enable_in (sw_256_latch_out),
        .clk_out         (sw_257_clk_out),
        .data_out        (sw_257_data_out),
        .scan_select_out (sw_257_scan_out),
        .latch_enable_out(sw_257_latch_out)
    );

    // [258] https://github.com/mattvenn/wokwi_filler
    wire sw_258_clk_out, sw_258_data_out, sw_258_scan_out, sw_258_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_258 (
        .clk_in          (sw_257_clk_out),
        .data_in         (sw_257_data_out),
        .scan_select_in  (sw_257_scan_out),
        .latch_enable_in (sw_257_latch_out),
        .clk_out         (sw_258_clk_out),
        .data_out        (sw_258_data_out),
        .scan_select_out (sw_258_scan_out),
        .latch_enable_out(sw_258_latch_out)
    );

    // [259] https://github.com/mattvenn/wokwi_filler
    wire sw_259_clk_out, sw_259_data_out, sw_259_scan_out, sw_259_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_259 (
        .clk_in          (sw_258_clk_out),
        .data_in         (sw_258_data_out),
        .scan_select_in  (sw_258_scan_out),
        .latch_enable_in (sw_258_latch_out),
        .clk_out         (sw_259_clk_out),
        .data_out        (sw_259_data_out),
        .scan_select_out (sw_259_scan_out),
        .latch_enable_out(sw_259_latch_out)
    );

    // [260] https://github.com/mattvenn/wokwi_filler
    wire sw_260_clk_out, sw_260_data_out, sw_260_scan_out, sw_260_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_260 (
        .clk_in          (sw_259_clk_out),
        .data_in         (sw_259_data_out),
        .scan_select_in  (sw_259_scan_out),
        .latch_enable_in (sw_259_latch_out),
        .clk_out         (sw_260_clk_out),
        .data_out        (sw_260_data_out),
        .scan_select_out (sw_260_scan_out),
        .latch_enable_out(sw_260_latch_out)
    );

    // [261] https://github.com/mattvenn/wokwi_filler
    wire sw_261_clk_out, sw_261_data_out, sw_261_scan_out, sw_261_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_261 (
        .clk_in          (sw_260_clk_out),
        .data_in         (sw_260_data_out),
        .scan_select_in  (sw_260_scan_out),
        .latch_enable_in (sw_260_latch_out),
        .clk_out         (sw_261_clk_out),
        .data_out        (sw_261_data_out),
        .scan_select_out (sw_261_scan_out),
        .latch_enable_out(sw_261_latch_out)
    );

    // [262] https://github.com/mattvenn/wokwi_filler
    wire sw_262_clk_out, sw_262_data_out, sw_262_scan_out, sw_262_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_262 (
        .clk_in          (sw_261_clk_out),
        .data_in         (sw_261_data_out),
        .scan_select_in  (sw_261_scan_out),
        .latch_enable_in (sw_261_latch_out),
        .clk_out         (sw_262_clk_out),
        .data_out        (sw_262_data_out),
        .scan_select_out (sw_262_scan_out),
        .latch_enable_out(sw_262_latch_out)
    );

    // [263] https://github.com/mattvenn/wokwi_filler
    wire sw_263_clk_out, sw_263_data_out, sw_263_scan_out, sw_263_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_263 (
        .clk_in          (sw_262_clk_out),
        .data_in         (sw_262_data_out),
        .scan_select_in  (sw_262_scan_out),
        .latch_enable_in (sw_262_latch_out),
        .clk_out         (sw_263_clk_out),
        .data_out        (sw_263_data_out),
        .scan_select_out (sw_263_scan_out),
        .latch_enable_out(sw_263_latch_out)
    );

    // [264] https://github.com/mattvenn/wokwi_filler
    wire sw_264_clk_out, sw_264_data_out, sw_264_scan_out, sw_264_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_264 (
        .clk_in          (sw_263_clk_out),
        .data_in         (sw_263_data_out),
        .scan_select_in  (sw_263_scan_out),
        .latch_enable_in (sw_263_latch_out),
        .clk_out         (sw_264_clk_out),
        .data_out        (sw_264_data_out),
        .scan_select_out (sw_264_scan_out),
        .latch_enable_out(sw_264_latch_out)
    );

    // [265] https://github.com/mattvenn/wokwi_filler
    wire sw_265_clk_out, sw_265_data_out, sw_265_scan_out, sw_265_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_265 (
        .clk_in          (sw_264_clk_out),
        .data_in         (sw_264_data_out),
        .scan_select_in  (sw_264_scan_out),
        .latch_enable_in (sw_264_latch_out),
        .clk_out         (sw_265_clk_out),
        .data_out        (sw_265_data_out),
        .scan_select_out (sw_265_scan_out),
        .latch_enable_out(sw_265_latch_out)
    );

    // [266] https://github.com/mattvenn/wokwi_filler
    wire sw_266_clk_out, sw_266_data_out, sw_266_scan_out, sw_266_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_266 (
        .clk_in          (sw_265_clk_out),
        .data_in         (sw_265_data_out),
        .scan_select_in  (sw_265_scan_out),
        .latch_enable_in (sw_265_latch_out),
        .clk_out         (sw_266_clk_out),
        .data_out        (sw_266_data_out),
        .scan_select_out (sw_266_scan_out),
        .latch_enable_out(sw_266_latch_out)
    );

    // [267] https://github.com/mattvenn/wokwi_filler
    wire sw_267_clk_out, sw_267_data_out, sw_267_scan_out, sw_267_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_267 (
        .clk_in          (sw_266_clk_out),
        .data_in         (sw_266_data_out),
        .scan_select_in  (sw_266_scan_out),
        .latch_enable_in (sw_266_latch_out),
        .clk_out         (sw_267_clk_out),
        .data_out        (sw_267_data_out),
        .scan_select_out (sw_267_scan_out),
        .latch_enable_out(sw_267_latch_out)
    );

    // [268] https://github.com/mattvenn/wokwi_filler
    wire sw_268_clk_out, sw_268_data_out, sw_268_scan_out, sw_268_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_268 (
        .clk_in          (sw_267_clk_out),
        .data_in         (sw_267_data_out),
        .scan_select_in  (sw_267_scan_out),
        .latch_enable_in (sw_267_latch_out),
        .clk_out         (sw_268_clk_out),
        .data_out        (sw_268_data_out),
        .scan_select_out (sw_268_scan_out),
        .latch_enable_out(sw_268_latch_out)
    );

    // [269] https://github.com/mattvenn/wokwi_filler
    wire sw_269_clk_out, sw_269_data_out, sw_269_scan_out, sw_269_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_269 (
        .clk_in          (sw_268_clk_out),
        .data_in         (sw_268_data_out),
        .scan_select_in  (sw_268_scan_out),
        .latch_enable_in (sw_268_latch_out),
        .clk_out         (sw_269_clk_out),
        .data_out        (sw_269_data_out),
        .scan_select_out (sw_269_scan_out),
        .latch_enable_out(sw_269_latch_out)
    );

    // [270] https://github.com/mattvenn/wokwi_filler
    wire sw_270_clk_out, sw_270_data_out, sw_270_scan_out, sw_270_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_270 (
        .clk_in          (sw_269_clk_out),
        .data_in         (sw_269_data_out),
        .scan_select_in  (sw_269_scan_out),
        .latch_enable_in (sw_269_latch_out),
        .clk_out         (sw_270_clk_out),
        .data_out        (sw_270_data_out),
        .scan_select_out (sw_270_scan_out),
        .latch_enable_out(sw_270_latch_out)
    );

    // [271] https://github.com/mattvenn/wokwi_filler
    wire sw_271_clk_out, sw_271_data_out, sw_271_scan_out, sw_271_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_271 (
        .clk_in          (sw_270_clk_out),
        .data_in         (sw_270_data_out),
        .scan_select_in  (sw_270_scan_out),
        .latch_enable_in (sw_270_latch_out),
        .clk_out         (sw_271_clk_out),
        .data_out        (sw_271_data_out),
        .scan_select_out (sw_271_scan_out),
        .latch_enable_out(sw_271_latch_out)
    );

    // [272] https://github.com/mattvenn/wokwi_filler
    wire sw_272_clk_out, sw_272_data_out, sw_272_scan_out, sw_272_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_272 (
        .clk_in          (sw_271_clk_out),
        .data_in         (sw_271_data_out),
        .scan_select_in  (sw_271_scan_out),
        .latch_enable_in (sw_271_latch_out),
        .clk_out         (sw_272_clk_out),
        .data_out        (sw_272_data_out),
        .scan_select_out (sw_272_scan_out),
        .latch_enable_out(sw_272_latch_out)
    );

    // [273] https://github.com/mattvenn/wokwi_filler
    wire sw_273_clk_out, sw_273_data_out, sw_273_scan_out, sw_273_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_273 (
        .clk_in          (sw_272_clk_out),
        .data_in         (sw_272_data_out),
        .scan_select_in  (sw_272_scan_out),
        .latch_enable_in (sw_272_latch_out),
        .clk_out         (sw_273_clk_out),
        .data_out        (sw_273_data_out),
        .scan_select_out (sw_273_scan_out),
        .latch_enable_out(sw_273_latch_out)
    );

    // [274] https://github.com/mattvenn/wokwi_filler
    wire sw_274_clk_out, sw_274_data_out, sw_274_scan_out, sw_274_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_274 (
        .clk_in          (sw_273_clk_out),
        .data_in         (sw_273_data_out),
        .scan_select_in  (sw_273_scan_out),
        .latch_enable_in (sw_273_latch_out),
        .clk_out         (sw_274_clk_out),
        .data_out        (sw_274_data_out),
        .scan_select_out (sw_274_scan_out),
        .latch_enable_out(sw_274_latch_out)
    );

    // [275] https://github.com/mattvenn/wokwi_filler
    wire sw_275_clk_out, sw_275_data_out, sw_275_scan_out, sw_275_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_275 (
        .clk_in          (sw_274_clk_out),
        .data_in         (sw_274_data_out),
        .scan_select_in  (sw_274_scan_out),
        .latch_enable_in (sw_274_latch_out),
        .clk_out         (sw_275_clk_out),
        .data_out        (sw_275_data_out),
        .scan_select_out (sw_275_scan_out),
        .latch_enable_out(sw_275_latch_out)
    );

    // [276] https://github.com/mattvenn/wokwi_filler
    wire sw_276_clk_out, sw_276_data_out, sw_276_scan_out, sw_276_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_276 (
        .clk_in          (sw_275_clk_out),
        .data_in         (sw_275_data_out),
        .scan_select_in  (sw_275_scan_out),
        .latch_enable_in (sw_275_latch_out),
        .clk_out         (sw_276_clk_out),
        .data_out        (sw_276_data_out),
        .scan_select_out (sw_276_scan_out),
        .latch_enable_out(sw_276_latch_out)
    );

    // [277] https://github.com/mattvenn/wokwi_filler
    wire sw_277_clk_out, sw_277_data_out, sw_277_scan_out, sw_277_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_277 (
        .clk_in          (sw_276_clk_out),
        .data_in         (sw_276_data_out),
        .scan_select_in  (sw_276_scan_out),
        .latch_enable_in (sw_276_latch_out),
        .clk_out         (sw_277_clk_out),
        .data_out        (sw_277_data_out),
        .scan_select_out (sw_277_scan_out),
        .latch_enable_out(sw_277_latch_out)
    );

    // [278] https://github.com/mattvenn/wokwi_filler
    wire sw_278_clk_out, sw_278_data_out, sw_278_scan_out, sw_278_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_278 (
        .clk_in          (sw_277_clk_out),
        .data_in         (sw_277_data_out),
        .scan_select_in  (sw_277_scan_out),
        .latch_enable_in (sw_277_latch_out),
        .clk_out         (sw_278_clk_out),
        .data_out        (sw_278_data_out),
        .scan_select_out (sw_278_scan_out),
        .latch_enable_out(sw_278_latch_out)
    );

    // [279] https://github.com/mattvenn/wokwi_filler
    wire sw_279_clk_out, sw_279_data_out, sw_279_scan_out, sw_279_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_279 (
        .clk_in          (sw_278_clk_out),
        .data_in         (sw_278_data_out),
        .scan_select_in  (sw_278_scan_out),
        .latch_enable_in (sw_278_latch_out),
        .clk_out         (sw_279_clk_out),
        .data_out        (sw_279_data_out),
        .scan_select_out (sw_279_scan_out),
        .latch_enable_out(sw_279_latch_out)
    );

    // [280] https://github.com/mattvenn/wokwi_filler
    wire sw_280_clk_out, sw_280_data_out, sw_280_scan_out, sw_280_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_280 (
        .clk_in          (sw_279_clk_out),
        .data_in         (sw_279_data_out),
        .scan_select_in  (sw_279_scan_out),
        .latch_enable_in (sw_279_latch_out),
        .clk_out         (sw_280_clk_out),
        .data_out        (sw_280_data_out),
        .scan_select_out (sw_280_scan_out),
        .latch_enable_out(sw_280_latch_out)
    );

    // [281] https://github.com/mattvenn/wokwi_filler
    wire sw_281_clk_out, sw_281_data_out, sw_281_scan_out, sw_281_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_281 (
        .clk_in          (sw_280_clk_out),
        .data_in         (sw_280_data_out),
        .scan_select_in  (sw_280_scan_out),
        .latch_enable_in (sw_280_latch_out),
        .clk_out         (sw_281_clk_out),
        .data_out        (sw_281_data_out),
        .scan_select_out (sw_281_scan_out),
        .latch_enable_out(sw_281_latch_out)
    );

    // [282] https://github.com/mattvenn/wokwi_filler
    wire sw_282_clk_out, sw_282_data_out, sw_282_scan_out, sw_282_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_282 (
        .clk_in          (sw_281_clk_out),
        .data_in         (sw_281_data_out),
        .scan_select_in  (sw_281_scan_out),
        .latch_enable_in (sw_281_latch_out),
        .clk_out         (sw_282_clk_out),
        .data_out        (sw_282_data_out),
        .scan_select_out (sw_282_scan_out),
        .latch_enable_out(sw_282_latch_out)
    );

    // [283] https://github.com/mattvenn/wokwi_filler
    wire sw_283_clk_out, sw_283_data_out, sw_283_scan_out, sw_283_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_283 (
        .clk_in          (sw_282_clk_out),
        .data_in         (sw_282_data_out),
        .scan_select_in  (sw_282_scan_out),
        .latch_enable_in (sw_282_latch_out),
        .clk_out         (sw_283_clk_out),
        .data_out        (sw_283_data_out),
        .scan_select_out (sw_283_scan_out),
        .latch_enable_out(sw_283_latch_out)
    );

    // [284] https://github.com/mattvenn/wokwi_filler
    wire sw_284_clk_out, sw_284_data_out, sw_284_scan_out, sw_284_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_284 (
        .clk_in          (sw_283_clk_out),
        .data_in         (sw_283_data_out),
        .scan_select_in  (sw_283_scan_out),
        .latch_enable_in (sw_283_latch_out),
        .clk_out         (sw_284_clk_out),
        .data_out        (sw_284_data_out),
        .scan_select_out (sw_284_scan_out),
        .latch_enable_out(sw_284_latch_out)
    );

    // [285] https://github.com/mattvenn/wokwi_filler
    wire sw_285_clk_out, sw_285_data_out, sw_285_scan_out, sw_285_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_285 (
        .clk_in          (sw_284_clk_out),
        .data_in         (sw_284_data_out),
        .scan_select_in  (sw_284_scan_out),
        .latch_enable_in (sw_284_latch_out),
        .clk_out         (sw_285_clk_out),
        .data_out        (sw_285_data_out),
        .scan_select_out (sw_285_scan_out),
        .latch_enable_out(sw_285_latch_out)
    );

    // [286] https://github.com/mattvenn/wokwi_filler
    wire sw_286_clk_out, sw_286_data_out, sw_286_scan_out, sw_286_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_286 (
        .clk_in          (sw_285_clk_out),
        .data_in         (sw_285_data_out),
        .scan_select_in  (sw_285_scan_out),
        .latch_enable_in (sw_285_latch_out),
        .clk_out         (sw_286_clk_out),
        .data_out        (sw_286_data_out),
        .scan_select_out (sw_286_scan_out),
        .latch_enable_out(sw_286_latch_out)
    );

    // [287] https://github.com/mattvenn/wokwi_filler
    wire sw_287_clk_out, sw_287_data_out, sw_287_scan_out, sw_287_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_287 (
        .clk_in          (sw_286_clk_out),
        .data_in         (sw_286_data_out),
        .scan_select_in  (sw_286_scan_out),
        .latch_enable_in (sw_286_latch_out),
        .clk_out         (sw_287_clk_out),
        .data_out        (sw_287_data_out),
        .scan_select_out (sw_287_scan_out),
        .latch_enable_out(sw_287_latch_out)
    );

    // [288] https://github.com/mattvenn/wokwi_filler
    wire sw_288_clk_out, sw_288_data_out, sw_288_scan_out, sw_288_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_288 (
        .clk_in          (sw_287_clk_out),
        .data_in         (sw_287_data_out),
        .scan_select_in  (sw_287_scan_out),
        .latch_enable_in (sw_287_latch_out),
        .clk_out         (sw_288_clk_out),
        .data_out        (sw_288_data_out),
        .scan_select_out (sw_288_scan_out),
        .latch_enable_out(sw_288_latch_out)
    );

    // [289] https://github.com/mattvenn/wokwi_filler
    wire sw_289_clk_out, sw_289_data_out, sw_289_scan_out, sw_289_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_289 (
        .clk_in          (sw_288_clk_out),
        .data_in         (sw_288_data_out),
        .scan_select_in  (sw_288_scan_out),
        .latch_enable_in (sw_288_latch_out),
        .clk_out         (sw_289_clk_out),
        .data_out        (sw_289_data_out),
        .scan_select_out (sw_289_scan_out),
        .latch_enable_out(sw_289_latch_out)
    );

    // [290] https://github.com/mattvenn/wokwi_filler
    wire sw_290_clk_out, sw_290_data_out, sw_290_scan_out, sw_290_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_290 (
        .clk_in          (sw_289_clk_out),
        .data_in         (sw_289_data_out),
        .scan_select_in  (sw_289_scan_out),
        .latch_enable_in (sw_289_latch_out),
        .clk_out         (sw_290_clk_out),
        .data_out        (sw_290_data_out),
        .scan_select_out (sw_290_scan_out),
        .latch_enable_out(sw_290_latch_out)
    );

    // [291] https://github.com/mattvenn/wokwi_filler
    wire sw_291_clk_out, sw_291_data_out, sw_291_scan_out, sw_291_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_291 (
        .clk_in          (sw_290_clk_out),
        .data_in         (sw_290_data_out),
        .scan_select_in  (sw_290_scan_out),
        .latch_enable_in (sw_290_latch_out),
        .clk_out         (sw_291_clk_out),
        .data_out        (sw_291_data_out),
        .scan_select_out (sw_291_scan_out),
        .latch_enable_out(sw_291_latch_out)
    );

    // [292] https://github.com/mattvenn/wokwi_filler
    wire sw_292_clk_out, sw_292_data_out, sw_292_scan_out, sw_292_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_292 (
        .clk_in          (sw_291_clk_out),
        .data_in         (sw_291_data_out),
        .scan_select_in  (sw_291_scan_out),
        .latch_enable_in (sw_291_latch_out),
        .clk_out         (sw_292_clk_out),
        .data_out        (sw_292_data_out),
        .scan_select_out (sw_292_scan_out),
        .latch_enable_out(sw_292_latch_out)
    );

    // [293] https://github.com/mattvenn/wokwi_filler
    wire sw_293_clk_out, sw_293_data_out, sw_293_scan_out, sw_293_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_293 (
        .clk_in          (sw_292_clk_out),
        .data_in         (sw_292_data_out),
        .scan_select_in  (sw_292_scan_out),
        .latch_enable_in (sw_292_latch_out),
        .clk_out         (sw_293_clk_out),
        .data_out        (sw_293_data_out),
        .scan_select_out (sw_293_scan_out),
        .latch_enable_out(sw_293_latch_out)
    );

    // [294] https://github.com/mattvenn/wokwi_filler
    wire sw_294_clk_out, sw_294_data_out, sw_294_scan_out, sw_294_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_294 (
        .clk_in          (sw_293_clk_out),
        .data_in         (sw_293_data_out),
        .scan_select_in  (sw_293_scan_out),
        .latch_enable_in (sw_293_latch_out),
        .clk_out         (sw_294_clk_out),
        .data_out        (sw_294_data_out),
        .scan_select_out (sw_294_scan_out),
        .latch_enable_out(sw_294_latch_out)
    );

    // [295] https://github.com/mattvenn/wokwi_filler
    wire sw_295_clk_out, sw_295_data_out, sw_295_scan_out, sw_295_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_295 (
        .clk_in          (sw_294_clk_out),
        .data_in         (sw_294_data_out),
        .scan_select_in  (sw_294_scan_out),
        .latch_enable_in (sw_294_latch_out),
        .clk_out         (sw_295_clk_out),
        .data_out        (sw_295_data_out),
        .scan_select_out (sw_295_scan_out),
        .latch_enable_out(sw_295_latch_out)
    );

    // [296] https://github.com/mattvenn/wokwi_filler
    wire sw_296_clk_out, sw_296_data_out, sw_296_scan_out, sw_296_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_296 (
        .clk_in          (sw_295_clk_out),
        .data_in         (sw_295_data_out),
        .scan_select_in  (sw_295_scan_out),
        .latch_enable_in (sw_295_latch_out),
        .clk_out         (sw_296_clk_out),
        .data_out        (sw_296_data_out),
        .scan_select_out (sw_296_scan_out),
        .latch_enable_out(sw_296_latch_out)
    );

    // [297] https://github.com/mattvenn/wokwi_filler
    wire sw_297_clk_out, sw_297_data_out, sw_297_scan_out, sw_297_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_297 (
        .clk_in          (sw_296_clk_out),
        .data_in         (sw_296_data_out),
        .scan_select_in  (sw_296_scan_out),
        .latch_enable_in (sw_296_latch_out),
        .clk_out         (sw_297_clk_out),
        .data_out        (sw_297_data_out),
        .scan_select_out (sw_297_scan_out),
        .latch_enable_out(sw_297_latch_out)
    );

    // [298] https://github.com/mattvenn/wokwi_filler
    wire sw_298_clk_out, sw_298_data_out, sw_298_scan_out, sw_298_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_298 (
        .clk_in          (sw_297_clk_out),
        .data_in         (sw_297_data_out),
        .scan_select_in  (sw_297_scan_out),
        .latch_enable_in (sw_297_latch_out),
        .clk_out         (sw_298_clk_out),
        .data_out        (sw_298_data_out),
        .scan_select_out (sw_298_scan_out),
        .latch_enable_out(sw_298_latch_out)
    );

    // [299] https://github.com/mattvenn/wokwi_filler
    wire sw_299_clk_out, sw_299_data_out, sw_299_scan_out, sw_299_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_299 (
        .clk_in          (sw_298_clk_out),
        .data_in         (sw_298_data_out),
        .scan_select_in  (sw_298_scan_out),
        .latch_enable_in (sw_298_latch_out),
        .clk_out         (sw_299_clk_out),
        .data_out        (sw_299_data_out),
        .scan_select_out (sw_299_scan_out),
        .latch_enable_out(sw_299_latch_out)
    );

    // [300] https://github.com/mattvenn/wokwi_filler
    wire sw_300_clk_out, sw_300_data_out, sw_300_scan_out, sw_300_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_300 (
        .clk_in          (sw_299_clk_out),
        .data_in         (sw_299_data_out),
        .scan_select_in  (sw_299_scan_out),
        .latch_enable_in (sw_299_latch_out),
        .clk_out         (sw_300_clk_out),
        .data_out        (sw_300_data_out),
        .scan_select_out (sw_300_scan_out),
        .latch_enable_out(sw_300_latch_out)
    );

    // [301] https://github.com/mattvenn/wokwi_filler
    wire sw_301_clk_out, sw_301_data_out, sw_301_scan_out, sw_301_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_301 (
        .clk_in          (sw_300_clk_out),
        .data_in         (sw_300_data_out),
        .scan_select_in  (sw_300_scan_out),
        .latch_enable_in (sw_300_latch_out),
        .clk_out         (sw_301_clk_out),
        .data_out        (sw_301_data_out),
        .scan_select_out (sw_301_scan_out),
        .latch_enable_out(sw_301_latch_out)
    );

    // [302] https://github.com/mattvenn/wokwi_filler
    wire sw_302_clk_out, sw_302_data_out, sw_302_scan_out, sw_302_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_302 (
        .clk_in          (sw_301_clk_out),
        .data_in         (sw_301_data_out),
        .scan_select_in  (sw_301_scan_out),
        .latch_enable_in (sw_301_latch_out),
        .clk_out         (sw_302_clk_out),
        .data_out        (sw_302_data_out),
        .scan_select_out (sw_302_scan_out),
        .latch_enable_out(sw_302_latch_out)
    );

    // [303] https://github.com/mattvenn/wokwi_filler
    wire sw_303_clk_out, sw_303_data_out, sw_303_scan_out, sw_303_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_303 (
        .clk_in          (sw_302_clk_out),
        .data_in         (sw_302_data_out),
        .scan_select_in  (sw_302_scan_out),
        .latch_enable_in (sw_302_latch_out),
        .clk_out         (sw_303_clk_out),
        .data_out        (sw_303_data_out),
        .scan_select_out (sw_303_scan_out),
        .latch_enable_out(sw_303_latch_out)
    );

    // [304] https://github.com/mattvenn/wokwi_filler
    wire sw_304_clk_out, sw_304_data_out, sw_304_scan_out, sw_304_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_304 (
        .clk_in          (sw_303_clk_out),
        .data_in         (sw_303_data_out),
        .scan_select_in  (sw_303_scan_out),
        .latch_enable_in (sw_303_latch_out),
        .clk_out         (sw_304_clk_out),
        .data_out        (sw_304_data_out),
        .scan_select_out (sw_304_scan_out),
        .latch_enable_out(sw_304_latch_out)
    );

    // [305] https://github.com/mattvenn/wokwi_filler
    wire sw_305_clk_out, sw_305_data_out, sw_305_scan_out, sw_305_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_305 (
        .clk_in          (sw_304_clk_out),
        .data_in         (sw_304_data_out),
        .scan_select_in  (sw_304_scan_out),
        .latch_enable_in (sw_304_latch_out),
        .clk_out         (sw_305_clk_out),
        .data_out        (sw_305_data_out),
        .scan_select_out (sw_305_scan_out),
        .latch_enable_out(sw_305_latch_out)
    );

    // [306] https://github.com/mattvenn/wokwi_filler
    wire sw_306_clk_out, sw_306_data_out, sw_306_scan_out, sw_306_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_306 (
        .clk_in          (sw_305_clk_out),
        .data_in         (sw_305_data_out),
        .scan_select_in  (sw_305_scan_out),
        .latch_enable_in (sw_305_latch_out),
        .clk_out         (sw_306_clk_out),
        .data_out        (sw_306_data_out),
        .scan_select_out (sw_306_scan_out),
        .latch_enable_out(sw_306_latch_out)
    );

    // [307] https://github.com/mattvenn/wokwi_filler
    wire sw_307_clk_out, sw_307_data_out, sw_307_scan_out, sw_307_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_307 (
        .clk_in          (sw_306_clk_out),
        .data_in         (sw_306_data_out),
        .scan_select_in  (sw_306_scan_out),
        .latch_enable_in (sw_306_latch_out),
        .clk_out         (sw_307_clk_out),
        .data_out        (sw_307_data_out),
        .scan_select_out (sw_307_scan_out),
        .latch_enable_out(sw_307_latch_out)
    );

    // [308] https://github.com/mattvenn/wokwi_filler
    wire sw_308_clk_out, sw_308_data_out, sw_308_scan_out, sw_308_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_308 (
        .clk_in          (sw_307_clk_out),
        .data_in         (sw_307_data_out),
        .scan_select_in  (sw_307_scan_out),
        .latch_enable_in (sw_307_latch_out),
        .clk_out         (sw_308_clk_out),
        .data_out        (sw_308_data_out),
        .scan_select_out (sw_308_scan_out),
        .latch_enable_out(sw_308_latch_out)
    );

    // [309] https://github.com/mattvenn/wokwi_filler
    wire sw_309_clk_out, sw_309_data_out, sw_309_scan_out, sw_309_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_309 (
        .clk_in          (sw_308_clk_out),
        .data_in         (sw_308_data_out),
        .scan_select_in  (sw_308_scan_out),
        .latch_enable_in (sw_308_latch_out),
        .clk_out         (sw_309_clk_out),
        .data_out        (sw_309_data_out),
        .scan_select_out (sw_309_scan_out),
        .latch_enable_out(sw_309_latch_out)
    );

    // [310] https://github.com/mattvenn/wokwi_filler
    wire sw_310_clk_out, sw_310_data_out, sw_310_scan_out, sw_310_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_310 (
        .clk_in          (sw_309_clk_out),
        .data_in         (sw_309_data_out),
        .scan_select_in  (sw_309_scan_out),
        .latch_enable_in (sw_309_latch_out),
        .clk_out         (sw_310_clk_out),
        .data_out        (sw_310_data_out),
        .scan_select_out (sw_310_scan_out),
        .latch_enable_out(sw_310_latch_out)
    );

    // [311] https://github.com/mattvenn/wokwi_filler
    wire sw_311_clk_out, sw_311_data_out, sw_311_scan_out, sw_311_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_311 (
        .clk_in          (sw_310_clk_out),
        .data_in         (sw_310_data_out),
        .scan_select_in  (sw_310_scan_out),
        .latch_enable_in (sw_310_latch_out),
        .clk_out         (sw_311_clk_out),
        .data_out        (sw_311_data_out),
        .scan_select_out (sw_311_scan_out),
        .latch_enable_out(sw_311_latch_out)
    );

    // [312] https://github.com/mattvenn/wokwi_filler
    wire sw_312_clk_out, sw_312_data_out, sw_312_scan_out, sw_312_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_312 (
        .clk_in          (sw_311_clk_out),
        .data_in         (sw_311_data_out),
        .scan_select_in  (sw_311_scan_out),
        .latch_enable_in (sw_311_latch_out),
        .clk_out         (sw_312_clk_out),
        .data_out        (sw_312_data_out),
        .scan_select_out (sw_312_scan_out),
        .latch_enable_out(sw_312_latch_out)
    );

    // [313] https://github.com/mattvenn/wokwi_filler
    wire sw_313_clk_out, sw_313_data_out, sw_313_scan_out, sw_313_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_313 (
        .clk_in          (sw_312_clk_out),
        .data_in         (sw_312_data_out),
        .scan_select_in  (sw_312_scan_out),
        .latch_enable_in (sw_312_latch_out),
        .clk_out         (sw_313_clk_out),
        .data_out        (sw_313_data_out),
        .scan_select_out (sw_313_scan_out),
        .latch_enable_out(sw_313_latch_out)
    );

    // [314] https://github.com/mattvenn/wokwi_filler
    wire sw_314_clk_out, sw_314_data_out, sw_314_scan_out, sw_314_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_314 (
        .clk_in          (sw_313_clk_out),
        .data_in         (sw_313_data_out),
        .scan_select_in  (sw_313_scan_out),
        .latch_enable_in (sw_313_latch_out),
        .clk_out         (sw_314_clk_out),
        .data_out        (sw_314_data_out),
        .scan_select_out (sw_314_scan_out),
        .latch_enable_out(sw_314_latch_out)
    );

    // [315] https://github.com/mattvenn/wokwi_filler
    wire sw_315_clk_out, sw_315_data_out, sw_315_scan_out, sw_315_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_315 (
        .clk_in          (sw_314_clk_out),
        .data_in         (sw_314_data_out),
        .scan_select_in  (sw_314_scan_out),
        .latch_enable_in (sw_314_latch_out),
        .clk_out         (sw_315_clk_out),
        .data_out        (sw_315_data_out),
        .scan_select_out (sw_315_scan_out),
        .latch_enable_out(sw_315_latch_out)
    );

    // [316] https://github.com/mattvenn/wokwi_filler
    wire sw_316_clk_out, sw_316_data_out, sw_316_scan_out, sw_316_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_316 (
        .clk_in          (sw_315_clk_out),
        .data_in         (sw_315_data_out),
        .scan_select_in  (sw_315_scan_out),
        .latch_enable_in (sw_315_latch_out),
        .clk_out         (sw_316_clk_out),
        .data_out        (sw_316_data_out),
        .scan_select_out (sw_316_scan_out),
        .latch_enable_out(sw_316_latch_out)
    );

    // [317] https://github.com/mattvenn/wokwi_filler
    wire sw_317_clk_out, sw_317_data_out, sw_317_scan_out, sw_317_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_317 (
        .clk_in          (sw_316_clk_out),
        .data_in         (sw_316_data_out),
        .scan_select_in  (sw_316_scan_out),
        .latch_enable_in (sw_316_latch_out),
        .clk_out         (sw_317_clk_out),
        .data_out        (sw_317_data_out),
        .scan_select_out (sw_317_scan_out),
        .latch_enable_out(sw_317_latch_out)
    );

    // [318] https://github.com/mattvenn/wokwi_filler
    wire sw_318_clk_out, sw_318_data_out, sw_318_scan_out, sw_318_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_318 (
        .clk_in          (sw_317_clk_out),
        .data_in         (sw_317_data_out),
        .scan_select_in  (sw_317_scan_out),
        .latch_enable_in (sw_317_latch_out),
        .clk_out         (sw_318_clk_out),
        .data_out        (sw_318_data_out),
        .scan_select_out (sw_318_scan_out),
        .latch_enable_out(sw_318_latch_out)
    );

    // [319] https://github.com/mattvenn/wokwi_filler
    wire sw_319_clk_out, sw_319_data_out, sw_319_scan_out, sw_319_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_319 (
        .clk_in          (sw_318_clk_out),
        .data_in         (sw_318_data_out),
        .scan_select_in  (sw_318_scan_out),
        .latch_enable_in (sw_318_latch_out),
        .clk_out         (sw_319_clk_out),
        .data_out        (sw_319_data_out),
        .scan_select_out (sw_319_scan_out),
        .latch_enable_out(sw_319_latch_out)
    );

    // [320] https://github.com/mattvenn/wokwi_filler
    wire sw_320_clk_out, sw_320_data_out, sw_320_scan_out, sw_320_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_320 (
        .clk_in          (sw_319_clk_out),
        .data_in         (sw_319_data_out),
        .scan_select_in  (sw_319_scan_out),
        .latch_enable_in (sw_319_latch_out),
        .clk_out         (sw_320_clk_out),
        .data_out        (sw_320_data_out),
        .scan_select_out (sw_320_scan_out),
        .latch_enable_out(sw_320_latch_out)
    );

    // [321] https://github.com/mattvenn/wokwi_filler
    wire sw_321_clk_out, sw_321_data_out, sw_321_scan_out, sw_321_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_321 (
        .clk_in          (sw_320_clk_out),
        .data_in         (sw_320_data_out),
        .scan_select_in  (sw_320_scan_out),
        .latch_enable_in (sw_320_latch_out),
        .clk_out         (sw_321_clk_out),
        .data_out        (sw_321_data_out),
        .scan_select_out (sw_321_scan_out),
        .latch_enable_out(sw_321_latch_out)
    );

    // [322] https://github.com/mattvenn/wokwi_filler
    wire sw_322_clk_out, sw_322_data_out, sw_322_scan_out, sw_322_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_322 (
        .clk_in          (sw_321_clk_out),
        .data_in         (sw_321_data_out),
        .scan_select_in  (sw_321_scan_out),
        .latch_enable_in (sw_321_latch_out),
        .clk_out         (sw_322_clk_out),
        .data_out        (sw_322_data_out),
        .scan_select_out (sw_322_scan_out),
        .latch_enable_out(sw_322_latch_out)
    );

    // [323] https://github.com/mattvenn/wokwi_filler
    wire sw_323_clk_out, sw_323_data_out, sw_323_scan_out, sw_323_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_323 (
        .clk_in          (sw_322_clk_out),
        .data_in         (sw_322_data_out),
        .scan_select_in  (sw_322_scan_out),
        .latch_enable_in (sw_322_latch_out),
        .clk_out         (sw_323_clk_out),
        .data_out        (sw_323_data_out),
        .scan_select_out (sw_323_scan_out),
        .latch_enable_out(sw_323_latch_out)
    );

    // [324] https://github.com/mattvenn/wokwi_filler
    wire sw_324_clk_out, sw_324_data_out, sw_324_scan_out, sw_324_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_324 (
        .clk_in          (sw_323_clk_out),
        .data_in         (sw_323_data_out),
        .scan_select_in  (sw_323_scan_out),
        .latch_enable_in (sw_323_latch_out),
        .clk_out         (sw_324_clk_out),
        .data_out        (sw_324_data_out),
        .scan_select_out (sw_324_scan_out),
        .latch_enable_out(sw_324_latch_out)
    );

    // [325] https://github.com/mattvenn/wokwi_filler
    wire sw_325_clk_out, sw_325_data_out, sw_325_scan_out, sw_325_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_325 (
        .clk_in          (sw_324_clk_out),
        .data_in         (sw_324_data_out),
        .scan_select_in  (sw_324_scan_out),
        .latch_enable_in (sw_324_latch_out),
        .clk_out         (sw_325_clk_out),
        .data_out        (sw_325_data_out),
        .scan_select_out (sw_325_scan_out),
        .latch_enable_out(sw_325_latch_out)
    );

    // [326] https://github.com/mattvenn/wokwi_filler
    wire sw_326_clk_out, sw_326_data_out, sw_326_scan_out, sw_326_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_326 (
        .clk_in          (sw_325_clk_out),
        .data_in         (sw_325_data_out),
        .scan_select_in  (sw_325_scan_out),
        .latch_enable_in (sw_325_latch_out),
        .clk_out         (sw_326_clk_out),
        .data_out        (sw_326_data_out),
        .scan_select_out (sw_326_scan_out),
        .latch_enable_out(sw_326_latch_out)
    );

    // [327] https://github.com/mattvenn/wokwi_filler
    wire sw_327_clk_out, sw_327_data_out, sw_327_scan_out, sw_327_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_327 (
        .clk_in          (sw_326_clk_out),
        .data_in         (sw_326_data_out),
        .scan_select_in  (sw_326_scan_out),
        .latch_enable_in (sw_326_latch_out),
        .clk_out         (sw_327_clk_out),
        .data_out        (sw_327_data_out),
        .scan_select_out (sw_327_scan_out),
        .latch_enable_out(sw_327_latch_out)
    );

    // [328] https://github.com/mattvenn/wokwi_filler
    wire sw_328_clk_out, sw_328_data_out, sw_328_scan_out, sw_328_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_328 (
        .clk_in          (sw_327_clk_out),
        .data_in         (sw_327_data_out),
        .scan_select_in  (sw_327_scan_out),
        .latch_enable_in (sw_327_latch_out),
        .clk_out         (sw_328_clk_out),
        .data_out        (sw_328_data_out),
        .scan_select_out (sw_328_scan_out),
        .latch_enable_out(sw_328_latch_out)
    );

    // [329] https://github.com/mattvenn/wokwi_filler
    wire sw_329_clk_out, sw_329_data_out, sw_329_scan_out, sw_329_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_329 (
        .clk_in          (sw_328_clk_out),
        .data_in         (sw_328_data_out),
        .scan_select_in  (sw_328_scan_out),
        .latch_enable_in (sw_328_latch_out),
        .clk_out         (sw_329_clk_out),
        .data_out        (sw_329_data_out),
        .scan_select_out (sw_329_scan_out),
        .latch_enable_out(sw_329_latch_out)
    );

    // [330] https://github.com/mattvenn/wokwi_filler
    wire sw_330_clk_out, sw_330_data_out, sw_330_scan_out, sw_330_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_330 (
        .clk_in          (sw_329_clk_out),
        .data_in         (sw_329_data_out),
        .scan_select_in  (sw_329_scan_out),
        .latch_enable_in (sw_329_latch_out),
        .clk_out         (sw_330_clk_out),
        .data_out        (sw_330_data_out),
        .scan_select_out (sw_330_scan_out),
        .latch_enable_out(sw_330_latch_out)
    );

    // [331] https://github.com/mattvenn/wokwi_filler
    wire sw_331_clk_out, sw_331_data_out, sw_331_scan_out, sw_331_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_331 (
        .clk_in          (sw_330_clk_out),
        .data_in         (sw_330_data_out),
        .scan_select_in  (sw_330_scan_out),
        .latch_enable_in (sw_330_latch_out),
        .clk_out         (sw_331_clk_out),
        .data_out        (sw_331_data_out),
        .scan_select_out (sw_331_scan_out),
        .latch_enable_out(sw_331_latch_out)
    );

    // [332] https://github.com/mattvenn/wokwi_filler
    wire sw_332_clk_out, sw_332_data_out, sw_332_scan_out, sw_332_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_332 (
        .clk_in          (sw_331_clk_out),
        .data_in         (sw_331_data_out),
        .scan_select_in  (sw_331_scan_out),
        .latch_enable_in (sw_331_latch_out),
        .clk_out         (sw_332_clk_out),
        .data_out        (sw_332_data_out),
        .scan_select_out (sw_332_scan_out),
        .latch_enable_out(sw_332_latch_out)
    );

    // [333] https://github.com/mattvenn/wokwi_filler
    wire sw_333_clk_out, sw_333_data_out, sw_333_scan_out, sw_333_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_333 (
        .clk_in          (sw_332_clk_out),
        .data_in         (sw_332_data_out),
        .scan_select_in  (sw_332_scan_out),
        .latch_enable_in (sw_332_latch_out),
        .clk_out         (sw_333_clk_out),
        .data_out        (sw_333_data_out),
        .scan_select_out (sw_333_scan_out),
        .latch_enable_out(sw_333_latch_out)
    );

    // [334] https://github.com/mattvenn/wokwi_filler
    wire sw_334_clk_out, sw_334_data_out, sw_334_scan_out, sw_334_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_334 (
        .clk_in          (sw_333_clk_out),
        .data_in         (sw_333_data_out),
        .scan_select_in  (sw_333_scan_out),
        .latch_enable_in (sw_333_latch_out),
        .clk_out         (sw_334_clk_out),
        .data_out        (sw_334_data_out),
        .scan_select_out (sw_334_scan_out),
        .latch_enable_out(sw_334_latch_out)
    );

    // [335] https://github.com/mattvenn/wokwi_filler
    wire sw_335_clk_out, sw_335_data_out, sw_335_scan_out, sw_335_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_335 (
        .clk_in          (sw_334_clk_out),
        .data_in         (sw_334_data_out),
        .scan_select_in  (sw_334_scan_out),
        .latch_enable_in (sw_334_latch_out),
        .clk_out         (sw_335_clk_out),
        .data_out        (sw_335_data_out),
        .scan_select_out (sw_335_scan_out),
        .latch_enable_out(sw_335_latch_out)
    );

    // [336] https://github.com/mattvenn/wokwi_filler
    wire sw_336_clk_out, sw_336_data_out, sw_336_scan_out, sw_336_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_336 (
        .clk_in          (sw_335_clk_out),
        .data_in         (sw_335_data_out),
        .scan_select_in  (sw_335_scan_out),
        .latch_enable_in (sw_335_latch_out),
        .clk_out         (sw_336_clk_out),
        .data_out        (sw_336_data_out),
        .scan_select_out (sw_336_scan_out),
        .latch_enable_out(sw_336_latch_out)
    );

    // [337] https://github.com/mattvenn/wokwi_filler
    wire sw_337_clk_out, sw_337_data_out, sw_337_scan_out, sw_337_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_337 (
        .clk_in          (sw_336_clk_out),
        .data_in         (sw_336_data_out),
        .scan_select_in  (sw_336_scan_out),
        .latch_enable_in (sw_336_latch_out),
        .clk_out         (sw_337_clk_out),
        .data_out        (sw_337_data_out),
        .scan_select_out (sw_337_scan_out),
        .latch_enable_out(sw_337_latch_out)
    );

    // [338] https://github.com/mattvenn/wokwi_filler
    wire sw_338_clk_out, sw_338_data_out, sw_338_scan_out, sw_338_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_338 (
        .clk_in          (sw_337_clk_out),
        .data_in         (sw_337_data_out),
        .scan_select_in  (sw_337_scan_out),
        .latch_enable_in (sw_337_latch_out),
        .clk_out         (sw_338_clk_out),
        .data_out        (sw_338_data_out),
        .scan_select_out (sw_338_scan_out),
        .latch_enable_out(sw_338_latch_out)
    );

    // [339] https://github.com/mattvenn/wokwi_filler
    wire sw_339_clk_out, sw_339_data_out, sw_339_scan_out, sw_339_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_339 (
        .clk_in          (sw_338_clk_out),
        .data_in         (sw_338_data_out),
        .scan_select_in  (sw_338_scan_out),
        .latch_enable_in (sw_338_latch_out),
        .clk_out         (sw_339_clk_out),
        .data_out        (sw_339_data_out),
        .scan_select_out (sw_339_scan_out),
        .latch_enable_out(sw_339_latch_out)
    );

    // [340] https://github.com/mattvenn/wokwi_filler
    wire sw_340_clk_out, sw_340_data_out, sw_340_scan_out, sw_340_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_340 (
        .clk_in          (sw_339_clk_out),
        .data_in         (sw_339_data_out),
        .scan_select_in  (sw_339_scan_out),
        .latch_enable_in (sw_339_latch_out),
        .clk_out         (sw_340_clk_out),
        .data_out        (sw_340_data_out),
        .scan_select_out (sw_340_scan_out),
        .latch_enable_out(sw_340_latch_out)
    );

    // [341] https://github.com/mattvenn/wokwi_filler
    wire sw_341_clk_out, sw_341_data_out, sw_341_scan_out, sw_341_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_341 (
        .clk_in          (sw_340_clk_out),
        .data_in         (sw_340_data_out),
        .scan_select_in  (sw_340_scan_out),
        .latch_enable_in (sw_340_latch_out),
        .clk_out         (sw_341_clk_out),
        .data_out        (sw_341_data_out),
        .scan_select_out (sw_341_scan_out),
        .latch_enable_out(sw_341_latch_out)
    );

    // [342] https://github.com/mattvenn/wokwi_filler
    wire sw_342_clk_out, sw_342_data_out, sw_342_scan_out, sw_342_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_342 (
        .clk_in          (sw_341_clk_out),
        .data_in         (sw_341_data_out),
        .scan_select_in  (sw_341_scan_out),
        .latch_enable_in (sw_341_latch_out),
        .clk_out         (sw_342_clk_out),
        .data_out        (sw_342_data_out),
        .scan_select_out (sw_342_scan_out),
        .latch_enable_out(sw_342_latch_out)
    );

    // [343] https://github.com/mattvenn/wokwi_filler
    wire sw_343_clk_out, sw_343_data_out, sw_343_scan_out, sw_343_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_343 (
        .clk_in          (sw_342_clk_out),
        .data_in         (sw_342_data_out),
        .scan_select_in  (sw_342_scan_out),
        .latch_enable_in (sw_342_latch_out),
        .clk_out         (sw_343_clk_out),
        .data_out        (sw_343_data_out),
        .scan_select_out (sw_343_scan_out),
        .latch_enable_out(sw_343_latch_out)
    );

    // [344] https://github.com/mattvenn/wokwi_filler
    wire sw_344_clk_out, sw_344_data_out, sw_344_scan_out, sw_344_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_344 (
        .clk_in          (sw_343_clk_out),
        .data_in         (sw_343_data_out),
        .scan_select_in  (sw_343_scan_out),
        .latch_enable_in (sw_343_latch_out),
        .clk_out         (sw_344_clk_out),
        .data_out        (sw_344_data_out),
        .scan_select_out (sw_344_scan_out),
        .latch_enable_out(sw_344_latch_out)
    );

    // [345] https://github.com/mattvenn/wokwi_filler
    wire sw_345_clk_out, sw_345_data_out, sw_345_scan_out, sw_345_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_345 (
        .clk_in          (sw_344_clk_out),
        .data_in         (sw_344_data_out),
        .scan_select_in  (sw_344_scan_out),
        .latch_enable_in (sw_344_latch_out),
        .clk_out         (sw_345_clk_out),
        .data_out        (sw_345_data_out),
        .scan_select_out (sw_345_scan_out),
        .latch_enable_out(sw_345_latch_out)
    );

    // [346] https://github.com/mattvenn/wokwi_filler
    wire sw_346_clk_out, sw_346_data_out, sw_346_scan_out, sw_346_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_346 (
        .clk_in          (sw_345_clk_out),
        .data_in         (sw_345_data_out),
        .scan_select_in  (sw_345_scan_out),
        .latch_enable_in (sw_345_latch_out),
        .clk_out         (sw_346_clk_out),
        .data_out        (sw_346_data_out),
        .scan_select_out (sw_346_scan_out),
        .latch_enable_out(sw_346_latch_out)
    );

    // [347] https://github.com/mattvenn/wokwi_filler
    wire sw_347_clk_out, sw_347_data_out, sw_347_scan_out, sw_347_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_347 (
        .clk_in          (sw_346_clk_out),
        .data_in         (sw_346_data_out),
        .scan_select_in  (sw_346_scan_out),
        .latch_enable_in (sw_346_latch_out),
        .clk_out         (sw_347_clk_out),
        .data_out        (sw_347_data_out),
        .scan_select_out (sw_347_scan_out),
        .latch_enable_out(sw_347_latch_out)
    );

    // [348] https://github.com/mattvenn/wokwi_filler
    wire sw_348_clk_out, sw_348_data_out, sw_348_scan_out, sw_348_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_348 (
        .clk_in          (sw_347_clk_out),
        .data_in         (sw_347_data_out),
        .scan_select_in  (sw_347_scan_out),
        .latch_enable_in (sw_347_latch_out),
        .clk_out         (sw_348_clk_out),
        .data_out        (sw_348_data_out),
        .scan_select_out (sw_348_scan_out),
        .latch_enable_out(sw_348_latch_out)
    );

    // [349] https://github.com/mattvenn/wokwi_filler
    wire sw_349_clk_out, sw_349_data_out, sw_349_scan_out, sw_349_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_349 (
        .clk_in          (sw_348_clk_out),
        .data_in         (sw_348_data_out),
        .scan_select_in  (sw_348_scan_out),
        .latch_enable_in (sw_348_latch_out),
        .clk_out         (sw_349_clk_out),
        .data_out        (sw_349_data_out),
        .scan_select_out (sw_349_scan_out),
        .latch_enable_out(sw_349_latch_out)
    );

    // [350] https://github.com/mattvenn/wokwi_filler
    wire sw_350_clk_out, sw_350_data_out, sw_350_scan_out, sw_350_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_350 (
        .clk_in          (sw_349_clk_out),
        .data_in         (sw_349_data_out),
        .scan_select_in  (sw_349_scan_out),
        .latch_enable_in (sw_349_latch_out),
        .clk_out         (sw_350_clk_out),
        .data_out        (sw_350_data_out),
        .scan_select_out (sw_350_scan_out),
        .latch_enable_out(sw_350_latch_out)
    );

    // [351] https://github.com/mattvenn/wokwi_filler
    wire sw_351_clk_out, sw_351_data_out, sw_351_scan_out, sw_351_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_351 (
        .clk_in          (sw_350_clk_out),
        .data_in         (sw_350_data_out),
        .scan_select_in  (sw_350_scan_out),
        .latch_enable_in (sw_350_latch_out),
        .clk_out         (sw_351_clk_out),
        .data_out        (sw_351_data_out),
        .scan_select_out (sw_351_scan_out),
        .latch_enable_out(sw_351_latch_out)
    );

    // [352] https://github.com/mattvenn/wokwi_filler
    wire sw_352_clk_out, sw_352_data_out, sw_352_scan_out, sw_352_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_352 (
        .clk_in          (sw_351_clk_out),
        .data_in         (sw_351_data_out),
        .scan_select_in  (sw_351_scan_out),
        .latch_enable_in (sw_351_latch_out),
        .clk_out         (sw_352_clk_out),
        .data_out        (sw_352_data_out),
        .scan_select_out (sw_352_scan_out),
        .latch_enable_out(sw_352_latch_out)
    );

    // [353] https://github.com/mattvenn/wokwi_filler
    wire sw_353_clk_out, sw_353_data_out, sw_353_scan_out, sw_353_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_353 (
        .clk_in          (sw_352_clk_out),
        .data_in         (sw_352_data_out),
        .scan_select_in  (sw_352_scan_out),
        .latch_enable_in (sw_352_latch_out),
        .clk_out         (sw_353_clk_out),
        .data_out        (sw_353_data_out),
        .scan_select_out (sw_353_scan_out),
        .latch_enable_out(sw_353_latch_out)
    );

    // [354] https://github.com/mattvenn/wokwi_filler
    wire sw_354_clk_out, sw_354_data_out, sw_354_scan_out, sw_354_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_354 (
        .clk_in          (sw_353_clk_out),
        .data_in         (sw_353_data_out),
        .scan_select_in  (sw_353_scan_out),
        .latch_enable_in (sw_353_latch_out),
        .clk_out         (sw_354_clk_out),
        .data_out        (sw_354_data_out),
        .scan_select_out (sw_354_scan_out),
        .latch_enable_out(sw_354_latch_out)
    );

    // [355] https://github.com/mattvenn/wokwi_filler
    wire sw_355_clk_out, sw_355_data_out, sw_355_scan_out, sw_355_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_355 (
        .clk_in          (sw_354_clk_out),
        .data_in         (sw_354_data_out),
        .scan_select_in  (sw_354_scan_out),
        .latch_enable_in (sw_354_latch_out),
        .clk_out         (sw_355_clk_out),
        .data_out        (sw_355_data_out),
        .scan_select_out (sw_355_scan_out),
        .latch_enable_out(sw_355_latch_out)
    );

    // [356] https://github.com/mattvenn/wokwi_filler
    wire sw_356_clk_out, sw_356_data_out, sw_356_scan_out, sw_356_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_356 (
        .clk_in          (sw_355_clk_out),
        .data_in         (sw_355_data_out),
        .scan_select_in  (sw_355_scan_out),
        .latch_enable_in (sw_355_latch_out),
        .clk_out         (sw_356_clk_out),
        .data_out        (sw_356_data_out),
        .scan_select_out (sw_356_scan_out),
        .latch_enable_out(sw_356_latch_out)
    );

    // [357] https://github.com/mattvenn/wokwi_filler
    wire sw_357_clk_out, sw_357_data_out, sw_357_scan_out, sw_357_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_357 (
        .clk_in          (sw_356_clk_out),
        .data_in         (sw_356_data_out),
        .scan_select_in  (sw_356_scan_out),
        .latch_enable_in (sw_356_latch_out),
        .clk_out         (sw_357_clk_out),
        .data_out        (sw_357_data_out),
        .scan_select_out (sw_357_scan_out),
        .latch_enable_out(sw_357_latch_out)
    );

    // [358] https://github.com/mattvenn/wokwi_filler
    wire sw_358_clk_out, sw_358_data_out, sw_358_scan_out, sw_358_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_358 (
        .clk_in          (sw_357_clk_out),
        .data_in         (sw_357_data_out),
        .scan_select_in  (sw_357_scan_out),
        .latch_enable_in (sw_357_latch_out),
        .clk_out         (sw_358_clk_out),
        .data_out        (sw_358_data_out),
        .scan_select_out (sw_358_scan_out),
        .latch_enable_out(sw_358_latch_out)
    );

    // [359] https://github.com/mattvenn/wokwi_filler
    wire sw_359_clk_out, sw_359_data_out, sw_359_scan_out, sw_359_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_359 (
        .clk_in          (sw_358_clk_out),
        .data_in         (sw_358_data_out),
        .scan_select_in  (sw_358_scan_out),
        .latch_enable_in (sw_358_latch_out),
        .clk_out         (sw_359_clk_out),
        .data_out        (sw_359_data_out),
        .scan_select_out (sw_359_scan_out),
        .latch_enable_out(sw_359_latch_out)
    );

    // [360] https://github.com/mattvenn/wokwi_filler
    wire sw_360_clk_out, sw_360_data_out, sw_360_scan_out, sw_360_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_360 (
        .clk_in          (sw_359_clk_out),
        .data_in         (sw_359_data_out),
        .scan_select_in  (sw_359_scan_out),
        .latch_enable_in (sw_359_latch_out),
        .clk_out         (sw_360_clk_out),
        .data_out        (sw_360_data_out),
        .scan_select_out (sw_360_scan_out),
        .latch_enable_out(sw_360_latch_out)
    );

    // [361] https://github.com/mattvenn/wokwi_filler
    wire sw_361_clk_out, sw_361_data_out, sw_361_scan_out, sw_361_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_361 (
        .clk_in          (sw_360_clk_out),
        .data_in         (sw_360_data_out),
        .scan_select_in  (sw_360_scan_out),
        .latch_enable_in (sw_360_latch_out),
        .clk_out         (sw_361_clk_out),
        .data_out        (sw_361_data_out),
        .scan_select_out (sw_361_scan_out),
        .latch_enable_out(sw_361_latch_out)
    );

    // [362] https://github.com/mattvenn/wokwi_filler
    wire sw_362_clk_out, sw_362_data_out, sw_362_scan_out, sw_362_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_362 (
        .clk_in          (sw_361_clk_out),
        .data_in         (sw_361_data_out),
        .scan_select_in  (sw_361_scan_out),
        .latch_enable_in (sw_361_latch_out),
        .clk_out         (sw_362_clk_out),
        .data_out        (sw_362_data_out),
        .scan_select_out (sw_362_scan_out),
        .latch_enable_out(sw_362_latch_out)
    );

    // [363] https://github.com/mattvenn/wokwi_filler
    wire sw_363_clk_out, sw_363_data_out, sw_363_scan_out, sw_363_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_363 (
        .clk_in          (sw_362_clk_out),
        .data_in         (sw_362_data_out),
        .scan_select_in  (sw_362_scan_out),
        .latch_enable_in (sw_362_latch_out),
        .clk_out         (sw_363_clk_out),
        .data_out        (sw_363_data_out),
        .scan_select_out (sw_363_scan_out),
        .latch_enable_out(sw_363_latch_out)
    );

    // [364] https://github.com/mattvenn/wokwi_filler
    wire sw_364_clk_out, sw_364_data_out, sw_364_scan_out, sw_364_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_364 (
        .clk_in          (sw_363_clk_out),
        .data_in         (sw_363_data_out),
        .scan_select_in  (sw_363_scan_out),
        .latch_enable_in (sw_363_latch_out),
        .clk_out         (sw_364_clk_out),
        .data_out        (sw_364_data_out),
        .scan_select_out (sw_364_scan_out),
        .latch_enable_out(sw_364_latch_out)
    );

    // [365] https://github.com/mattvenn/wokwi_filler
    wire sw_365_clk_out, sw_365_data_out, sw_365_scan_out, sw_365_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_365 (
        .clk_in          (sw_364_clk_out),
        .data_in         (sw_364_data_out),
        .scan_select_in  (sw_364_scan_out),
        .latch_enable_in (sw_364_latch_out),
        .clk_out         (sw_365_clk_out),
        .data_out        (sw_365_data_out),
        .scan_select_out (sw_365_scan_out),
        .latch_enable_out(sw_365_latch_out)
    );

    // [366] https://github.com/mattvenn/wokwi_filler
    wire sw_366_clk_out, sw_366_data_out, sw_366_scan_out, sw_366_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_366 (
        .clk_in          (sw_365_clk_out),
        .data_in         (sw_365_data_out),
        .scan_select_in  (sw_365_scan_out),
        .latch_enable_in (sw_365_latch_out),
        .clk_out         (sw_366_clk_out),
        .data_out        (sw_366_data_out),
        .scan_select_out (sw_366_scan_out),
        .latch_enable_out(sw_366_latch_out)
    );

    // [367] https://github.com/mattvenn/wokwi_filler
    wire sw_367_clk_out, sw_367_data_out, sw_367_scan_out, sw_367_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_367 (
        .clk_in          (sw_366_clk_out),
        .data_in         (sw_366_data_out),
        .scan_select_in  (sw_366_scan_out),
        .latch_enable_in (sw_366_latch_out),
        .clk_out         (sw_367_clk_out),
        .data_out        (sw_367_data_out),
        .scan_select_out (sw_367_scan_out),
        .latch_enable_out(sw_367_latch_out)
    );

    // [368] https://github.com/mattvenn/wokwi_filler
    wire sw_368_clk_out, sw_368_data_out, sw_368_scan_out, sw_368_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_368 (
        .clk_in          (sw_367_clk_out),
        .data_in         (sw_367_data_out),
        .scan_select_in  (sw_367_scan_out),
        .latch_enable_in (sw_367_latch_out),
        .clk_out         (sw_368_clk_out),
        .data_out        (sw_368_data_out),
        .scan_select_out (sw_368_scan_out),
        .latch_enable_out(sw_368_latch_out)
    );

    // [369] https://github.com/mattvenn/wokwi_filler
    wire sw_369_clk_out, sw_369_data_out, sw_369_scan_out, sw_369_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_369 (
        .clk_in          (sw_368_clk_out),
        .data_in         (sw_368_data_out),
        .scan_select_in  (sw_368_scan_out),
        .latch_enable_in (sw_368_latch_out),
        .clk_out         (sw_369_clk_out),
        .data_out        (sw_369_data_out),
        .scan_select_out (sw_369_scan_out),
        .latch_enable_out(sw_369_latch_out)
    );

    // [370] https://github.com/mattvenn/wokwi_filler
    wire sw_370_clk_out, sw_370_data_out, sw_370_scan_out, sw_370_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_370 (
        .clk_in          (sw_369_clk_out),
        .data_in         (sw_369_data_out),
        .scan_select_in  (sw_369_scan_out),
        .latch_enable_in (sw_369_latch_out),
        .clk_out         (sw_370_clk_out),
        .data_out        (sw_370_data_out),
        .scan_select_out (sw_370_scan_out),
        .latch_enable_out(sw_370_latch_out)
    );

    // [371] https://github.com/mattvenn/wokwi_filler
    wire sw_371_clk_out, sw_371_data_out, sw_371_scan_out, sw_371_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_371 (
        .clk_in          (sw_370_clk_out),
        .data_in         (sw_370_data_out),
        .scan_select_in  (sw_370_scan_out),
        .latch_enable_in (sw_370_latch_out),
        .clk_out         (sw_371_clk_out),
        .data_out        (sw_371_data_out),
        .scan_select_out (sw_371_scan_out),
        .latch_enable_out(sw_371_latch_out)
    );

    // [372] https://github.com/mattvenn/wokwi_filler
    wire sw_372_clk_out, sw_372_data_out, sw_372_scan_out, sw_372_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_372 (
        .clk_in          (sw_371_clk_out),
        .data_in         (sw_371_data_out),
        .scan_select_in  (sw_371_scan_out),
        .latch_enable_in (sw_371_latch_out),
        .clk_out         (sw_372_clk_out),
        .data_out        (sw_372_data_out),
        .scan_select_out (sw_372_scan_out),
        .latch_enable_out(sw_372_latch_out)
    );

    // [373] https://github.com/mattvenn/wokwi_filler
    wire sw_373_clk_out, sw_373_data_out, sw_373_scan_out, sw_373_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_373 (
        .clk_in          (sw_372_clk_out),
        .data_in         (sw_372_data_out),
        .scan_select_in  (sw_372_scan_out),
        .latch_enable_in (sw_372_latch_out),
        .clk_out         (sw_373_clk_out),
        .data_out        (sw_373_data_out),
        .scan_select_out (sw_373_scan_out),
        .latch_enable_out(sw_373_latch_out)
    );

    // [374] https://github.com/mattvenn/wokwi_filler
    wire sw_374_clk_out, sw_374_data_out, sw_374_scan_out, sw_374_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_374 (
        .clk_in          (sw_373_clk_out),
        .data_in         (sw_373_data_out),
        .scan_select_in  (sw_373_scan_out),
        .latch_enable_in (sw_373_latch_out),
        .clk_out         (sw_374_clk_out),
        .data_out        (sw_374_data_out),
        .scan_select_out (sw_374_scan_out),
        .latch_enable_out(sw_374_latch_out)
    );

    // [375] https://github.com/mattvenn/wokwi_filler
    wire sw_375_clk_out, sw_375_data_out, sw_375_scan_out, sw_375_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_375 (
        .clk_in          (sw_374_clk_out),
        .data_in         (sw_374_data_out),
        .scan_select_in  (sw_374_scan_out),
        .latch_enable_in (sw_374_latch_out),
        .clk_out         (sw_375_clk_out),
        .data_out        (sw_375_data_out),
        .scan_select_out (sw_375_scan_out),
        .latch_enable_out(sw_375_latch_out)
    );

    // [376] https://github.com/mattvenn/wokwi_filler
    wire sw_376_clk_out, sw_376_data_out, sw_376_scan_out, sw_376_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_376 (
        .clk_in          (sw_375_clk_out),
        .data_in         (sw_375_data_out),
        .scan_select_in  (sw_375_scan_out),
        .latch_enable_in (sw_375_latch_out),
        .clk_out         (sw_376_clk_out),
        .data_out        (sw_376_data_out),
        .scan_select_out (sw_376_scan_out),
        .latch_enable_out(sw_376_latch_out)
    );

    // [377] https://github.com/mattvenn/wokwi_filler
    wire sw_377_clk_out, sw_377_data_out, sw_377_scan_out, sw_377_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_377 (
        .clk_in          (sw_376_clk_out),
        .data_in         (sw_376_data_out),
        .scan_select_in  (sw_376_scan_out),
        .latch_enable_in (sw_376_latch_out),
        .clk_out         (sw_377_clk_out),
        .data_out        (sw_377_data_out),
        .scan_select_out (sw_377_scan_out),
        .latch_enable_out(sw_377_latch_out)
    );

    // [378] https://github.com/mattvenn/wokwi_filler
    wire sw_378_clk_out, sw_378_data_out, sw_378_scan_out, sw_378_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_378 (
        .clk_in          (sw_377_clk_out),
        .data_in         (sw_377_data_out),
        .scan_select_in  (sw_377_scan_out),
        .latch_enable_in (sw_377_latch_out),
        .clk_out         (sw_378_clk_out),
        .data_out        (sw_378_data_out),
        .scan_select_out (sw_378_scan_out),
        .latch_enable_out(sw_378_latch_out)
    );

    // [379] https://github.com/mattvenn/wokwi_filler
    wire sw_379_clk_out, sw_379_data_out, sw_379_scan_out, sw_379_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_379 (
        .clk_in          (sw_378_clk_out),
        .data_in         (sw_378_data_out),
        .scan_select_in  (sw_378_scan_out),
        .latch_enable_in (sw_378_latch_out),
        .clk_out         (sw_379_clk_out),
        .data_out        (sw_379_data_out),
        .scan_select_out (sw_379_scan_out),
        .latch_enable_out(sw_379_latch_out)
    );

    // [380] https://github.com/mattvenn/wokwi_filler
    wire sw_380_clk_out, sw_380_data_out, sw_380_scan_out, sw_380_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_380 (
        .clk_in          (sw_379_clk_out),
        .data_in         (sw_379_data_out),
        .scan_select_in  (sw_379_scan_out),
        .latch_enable_in (sw_379_latch_out),
        .clk_out         (sw_380_clk_out),
        .data_out        (sw_380_data_out),
        .scan_select_out (sw_380_scan_out),
        .latch_enable_out(sw_380_latch_out)
    );

    // [381] https://github.com/mattvenn/wokwi_filler
    wire sw_381_clk_out, sw_381_data_out, sw_381_scan_out, sw_381_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_381 (
        .clk_in          (sw_380_clk_out),
        .data_in         (sw_380_data_out),
        .scan_select_in  (sw_380_scan_out),
        .latch_enable_in (sw_380_latch_out),
        .clk_out         (sw_381_clk_out),
        .data_out        (sw_381_data_out),
        .scan_select_out (sw_381_scan_out),
        .latch_enable_out(sw_381_latch_out)
    );

    // [382] https://github.com/mattvenn/wokwi_filler
    wire sw_382_clk_out, sw_382_data_out, sw_382_scan_out, sw_382_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_382 (
        .clk_in          (sw_381_clk_out),
        .data_in         (sw_381_data_out),
        .scan_select_in  (sw_381_scan_out),
        .latch_enable_in (sw_381_latch_out),
        .clk_out         (sw_382_clk_out),
        .data_out        (sw_382_data_out),
        .scan_select_out (sw_382_scan_out),
        .latch_enable_out(sw_382_latch_out)
    );

    // [383] https://github.com/mattvenn/wokwi_filler
    wire sw_383_clk_out, sw_383_data_out, sw_383_scan_out, sw_383_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_383 (
        .clk_in          (sw_382_clk_out),
        .data_in         (sw_382_data_out),
        .scan_select_in  (sw_382_scan_out),
        .latch_enable_in (sw_382_latch_out),
        .clk_out         (sw_383_clk_out),
        .data_out        (sw_383_data_out),
        .scan_select_out (sw_383_scan_out),
        .latch_enable_out(sw_383_latch_out)
    );

    // [384] https://github.com/mattvenn/wokwi_filler
    wire sw_384_clk_out, sw_384_data_out, sw_384_scan_out, sw_384_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_384 (
        .clk_in          (sw_383_clk_out),
        .data_in         (sw_383_data_out),
        .scan_select_in  (sw_383_scan_out),
        .latch_enable_in (sw_383_latch_out),
        .clk_out         (sw_384_clk_out),
        .data_out        (sw_384_data_out),
        .scan_select_out (sw_384_scan_out),
        .latch_enable_out(sw_384_latch_out)
    );

    // [385] https://github.com/mattvenn/wokwi_filler
    wire sw_385_clk_out, sw_385_data_out, sw_385_scan_out, sw_385_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_385 (
        .clk_in          (sw_384_clk_out),
        .data_in         (sw_384_data_out),
        .scan_select_in  (sw_384_scan_out),
        .latch_enable_in (sw_384_latch_out),
        .clk_out         (sw_385_clk_out),
        .data_out        (sw_385_data_out),
        .scan_select_out (sw_385_scan_out),
        .latch_enable_out(sw_385_latch_out)
    );

    // [386] https://github.com/mattvenn/wokwi_filler
    wire sw_386_clk_out, sw_386_data_out, sw_386_scan_out, sw_386_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_386 (
        .clk_in          (sw_385_clk_out),
        .data_in         (sw_385_data_out),
        .scan_select_in  (sw_385_scan_out),
        .latch_enable_in (sw_385_latch_out),
        .clk_out         (sw_386_clk_out),
        .data_out        (sw_386_data_out),
        .scan_select_out (sw_386_scan_out),
        .latch_enable_out(sw_386_latch_out)
    );

    // [387] https://github.com/mattvenn/wokwi_filler
    wire sw_387_clk_out, sw_387_data_out, sw_387_scan_out, sw_387_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_387 (
        .clk_in          (sw_386_clk_out),
        .data_in         (sw_386_data_out),
        .scan_select_in  (sw_386_scan_out),
        .latch_enable_in (sw_386_latch_out),
        .clk_out         (sw_387_clk_out),
        .data_out        (sw_387_data_out),
        .scan_select_out (sw_387_scan_out),
        .latch_enable_out(sw_387_latch_out)
    );

    // [388] https://github.com/mattvenn/wokwi_filler
    wire sw_388_clk_out, sw_388_data_out, sw_388_scan_out, sw_388_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_388 (
        .clk_in          (sw_387_clk_out),
        .data_in         (sw_387_data_out),
        .scan_select_in  (sw_387_scan_out),
        .latch_enable_in (sw_387_latch_out),
        .clk_out         (sw_388_clk_out),
        .data_out        (sw_388_data_out),
        .scan_select_out (sw_388_scan_out),
        .latch_enable_out(sw_388_latch_out)
    );

    // [389] https://github.com/mattvenn/wokwi_filler
    wire sw_389_clk_out, sw_389_data_out, sw_389_scan_out, sw_389_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_389 (
        .clk_in          (sw_388_clk_out),
        .data_in         (sw_388_data_out),
        .scan_select_in  (sw_388_scan_out),
        .latch_enable_in (sw_388_latch_out),
        .clk_out         (sw_389_clk_out),
        .data_out        (sw_389_data_out),
        .scan_select_out (sw_389_scan_out),
        .latch_enable_out(sw_389_latch_out)
    );

    // [390] https://github.com/mattvenn/wokwi_filler
    wire sw_390_clk_out, sw_390_data_out, sw_390_scan_out, sw_390_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_390 (
        .clk_in          (sw_389_clk_out),
        .data_in         (sw_389_data_out),
        .scan_select_in  (sw_389_scan_out),
        .latch_enable_in (sw_389_latch_out),
        .clk_out         (sw_390_clk_out),
        .data_out        (sw_390_data_out),
        .scan_select_out (sw_390_scan_out),
        .latch_enable_out(sw_390_latch_out)
    );

    // [391] https://github.com/mattvenn/wokwi_filler
    wire sw_391_clk_out, sw_391_data_out, sw_391_scan_out, sw_391_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_391 (
        .clk_in          (sw_390_clk_out),
        .data_in         (sw_390_data_out),
        .scan_select_in  (sw_390_scan_out),
        .latch_enable_in (sw_390_latch_out),
        .clk_out         (sw_391_clk_out),
        .data_out        (sw_391_data_out),
        .scan_select_out (sw_391_scan_out),
        .latch_enable_out(sw_391_latch_out)
    );

    // [392] https://github.com/mattvenn/wokwi_filler
    wire sw_392_clk_out, sw_392_data_out, sw_392_scan_out, sw_392_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_392 (
        .clk_in          (sw_391_clk_out),
        .data_in         (sw_391_data_out),
        .scan_select_in  (sw_391_scan_out),
        .latch_enable_in (sw_391_latch_out),
        .clk_out         (sw_392_clk_out),
        .data_out        (sw_392_data_out),
        .scan_select_out (sw_392_scan_out),
        .latch_enable_out(sw_392_latch_out)
    );

    // [393] https://github.com/mattvenn/wokwi_filler
    wire sw_393_clk_out, sw_393_data_out, sw_393_scan_out, sw_393_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_393 (
        .clk_in          (sw_392_clk_out),
        .data_in         (sw_392_data_out),
        .scan_select_in  (sw_392_scan_out),
        .latch_enable_in (sw_392_latch_out),
        .clk_out         (sw_393_clk_out),
        .data_out        (sw_393_data_out),
        .scan_select_out (sw_393_scan_out),
        .latch_enable_out(sw_393_latch_out)
    );

    // [394] https://github.com/mattvenn/wokwi_filler
    wire sw_394_clk_out, sw_394_data_out, sw_394_scan_out, sw_394_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_394 (
        .clk_in          (sw_393_clk_out),
        .data_in         (sw_393_data_out),
        .scan_select_in  (sw_393_scan_out),
        .latch_enable_in (sw_393_latch_out),
        .clk_out         (sw_394_clk_out),
        .data_out        (sw_394_data_out),
        .scan_select_out (sw_394_scan_out),
        .latch_enable_out(sw_394_latch_out)
    );

    // [395] https://github.com/mattvenn/wokwi_filler
    wire sw_395_clk_out, sw_395_data_out, sw_395_scan_out, sw_395_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_395 (
        .clk_in          (sw_394_clk_out),
        .data_in         (sw_394_data_out),
        .scan_select_in  (sw_394_scan_out),
        .latch_enable_in (sw_394_latch_out),
        .clk_out         (sw_395_clk_out),
        .data_out        (sw_395_data_out),
        .scan_select_out (sw_395_scan_out),
        .latch_enable_out(sw_395_latch_out)
    );

    // [396] https://github.com/mattvenn/wokwi_filler
    wire sw_396_clk_out, sw_396_data_out, sw_396_scan_out, sw_396_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_396 (
        .clk_in          (sw_395_clk_out),
        .data_in         (sw_395_data_out),
        .scan_select_in  (sw_395_scan_out),
        .latch_enable_in (sw_395_latch_out),
        .clk_out         (sw_396_clk_out),
        .data_out        (sw_396_data_out),
        .scan_select_out (sw_396_scan_out),
        .latch_enable_out(sw_396_latch_out)
    );

    // [397] https://github.com/mattvenn/wokwi_filler
    wire sw_397_clk_out, sw_397_data_out, sw_397_scan_out, sw_397_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_397 (
        .clk_in          (sw_396_clk_out),
        .data_in         (sw_396_data_out),
        .scan_select_in  (sw_396_scan_out),
        .latch_enable_in (sw_396_latch_out),
        .clk_out         (sw_397_clk_out),
        .data_out        (sw_397_data_out),
        .scan_select_out (sw_397_scan_out),
        .latch_enable_out(sw_397_latch_out)
    );

    // [398] https://github.com/mattvenn/wokwi_filler
    wire sw_398_clk_out, sw_398_data_out, sw_398_scan_out, sw_398_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_398 (
        .clk_in          (sw_397_clk_out),
        .data_in         (sw_397_data_out),
        .scan_select_in  (sw_397_scan_out),
        .latch_enable_in (sw_397_latch_out),
        .clk_out         (sw_398_clk_out),
        .data_out        (sw_398_data_out),
        .scan_select_out (sw_398_scan_out),
        .latch_enable_out(sw_398_latch_out)
    );

    // [399] https://github.com/mattvenn/wokwi_filler
    wire sw_399_clk_out, sw_399_data_out, sw_399_scan_out, sw_399_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_399 (
        .clk_in          (sw_398_clk_out),
        .data_in         (sw_398_data_out),
        .scan_select_in  (sw_398_scan_out),
        .latch_enable_in (sw_398_latch_out),
        .clk_out         (sw_399_clk_out),
        .data_out        (sw_399_data_out),
        .scan_select_out (sw_399_scan_out),
        .latch_enable_out(sw_399_latch_out)
    );

    // [400] https://github.com/mattvenn/wokwi_filler
    wire sw_400_clk_out, sw_400_data_out, sw_400_scan_out, sw_400_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_400 (
        .clk_in          (sw_399_clk_out),
        .data_in         (sw_399_data_out),
        .scan_select_in  (sw_399_scan_out),
        .latch_enable_in (sw_399_latch_out),
        .clk_out         (sw_400_clk_out),
        .data_out        (sw_400_data_out),
        .scan_select_out (sw_400_scan_out),
        .latch_enable_out(sw_400_latch_out)
    );

    // [401] https://github.com/mattvenn/wokwi_filler
    wire sw_401_clk_out, sw_401_data_out, sw_401_scan_out, sw_401_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_401 (
        .clk_in          (sw_400_clk_out),
        .data_in         (sw_400_data_out),
        .scan_select_in  (sw_400_scan_out),
        .latch_enable_in (sw_400_latch_out),
        .clk_out         (sw_401_clk_out),
        .data_out        (sw_401_data_out),
        .scan_select_out (sw_401_scan_out),
        .latch_enable_out(sw_401_latch_out)
    );

    // [402] https://github.com/mattvenn/wokwi_filler
    wire sw_402_clk_out, sw_402_data_out, sw_402_scan_out, sw_402_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_402 (
        .clk_in          (sw_401_clk_out),
        .data_in         (sw_401_data_out),
        .scan_select_in  (sw_401_scan_out),
        .latch_enable_in (sw_401_latch_out),
        .clk_out         (sw_402_clk_out),
        .data_out        (sw_402_data_out),
        .scan_select_out (sw_402_scan_out),
        .latch_enable_out(sw_402_latch_out)
    );

    // [403] https://github.com/mattvenn/wokwi_filler
    wire sw_403_clk_out, sw_403_data_out, sw_403_scan_out, sw_403_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_403 (
        .clk_in          (sw_402_clk_out),
        .data_in         (sw_402_data_out),
        .scan_select_in  (sw_402_scan_out),
        .latch_enable_in (sw_402_latch_out),
        .clk_out         (sw_403_clk_out),
        .data_out        (sw_403_data_out),
        .scan_select_out (sw_403_scan_out),
        .latch_enable_out(sw_403_latch_out)
    );

    // [404] https://github.com/mattvenn/wokwi_filler
    wire sw_404_clk_out, sw_404_data_out, sw_404_scan_out, sw_404_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_404 (
        .clk_in          (sw_403_clk_out),
        .data_in         (sw_403_data_out),
        .scan_select_in  (sw_403_scan_out),
        .latch_enable_in (sw_403_latch_out),
        .clk_out         (sw_404_clk_out),
        .data_out        (sw_404_data_out),
        .scan_select_out (sw_404_scan_out),
        .latch_enable_out(sw_404_latch_out)
    );

    // [405] https://github.com/mattvenn/wokwi_filler
    wire sw_405_clk_out, sw_405_data_out, sw_405_scan_out, sw_405_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_405 (
        .clk_in          (sw_404_clk_out),
        .data_in         (sw_404_data_out),
        .scan_select_in  (sw_404_scan_out),
        .latch_enable_in (sw_404_latch_out),
        .clk_out         (sw_405_clk_out),
        .data_out        (sw_405_data_out),
        .scan_select_out (sw_405_scan_out),
        .latch_enable_out(sw_405_latch_out)
    );

    // [406] https://github.com/mattvenn/wokwi_filler
    wire sw_406_clk_out, sw_406_data_out, sw_406_scan_out, sw_406_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_406 (
        .clk_in          (sw_405_clk_out),
        .data_in         (sw_405_data_out),
        .scan_select_in  (sw_405_scan_out),
        .latch_enable_in (sw_405_latch_out),
        .clk_out         (sw_406_clk_out),
        .data_out        (sw_406_data_out),
        .scan_select_out (sw_406_scan_out),
        .latch_enable_out(sw_406_latch_out)
    );

    // [407] https://github.com/mattvenn/wokwi_filler
    wire sw_407_clk_out, sw_407_data_out, sw_407_scan_out, sw_407_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_407 (
        .clk_in          (sw_406_clk_out),
        .data_in         (sw_406_data_out),
        .scan_select_in  (sw_406_scan_out),
        .latch_enable_in (sw_406_latch_out),
        .clk_out         (sw_407_clk_out),
        .data_out        (sw_407_data_out),
        .scan_select_out (sw_407_scan_out),
        .latch_enable_out(sw_407_latch_out)
    );

    // [408] https://github.com/mattvenn/wokwi_filler
    wire sw_408_clk_out, sw_408_data_out, sw_408_scan_out, sw_408_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_408 (
        .clk_in          (sw_407_clk_out),
        .data_in         (sw_407_data_out),
        .scan_select_in  (sw_407_scan_out),
        .latch_enable_in (sw_407_latch_out),
        .clk_out         (sw_408_clk_out),
        .data_out        (sw_408_data_out),
        .scan_select_out (sw_408_scan_out),
        .latch_enable_out(sw_408_latch_out)
    );

    // [409] https://github.com/mattvenn/wokwi_filler
    wire sw_409_clk_out, sw_409_data_out, sw_409_scan_out, sw_409_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_409 (
        .clk_in          (sw_408_clk_out),
        .data_in         (sw_408_data_out),
        .scan_select_in  (sw_408_scan_out),
        .latch_enable_in (sw_408_latch_out),
        .clk_out         (sw_409_clk_out),
        .data_out        (sw_409_data_out),
        .scan_select_out (sw_409_scan_out),
        .latch_enable_out(sw_409_latch_out)
    );

    // [410] https://github.com/mattvenn/wokwi_filler
    wire sw_410_clk_out, sw_410_data_out, sw_410_scan_out, sw_410_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_410 (
        .clk_in          (sw_409_clk_out),
        .data_in         (sw_409_data_out),
        .scan_select_in  (sw_409_scan_out),
        .latch_enable_in (sw_409_latch_out),
        .clk_out         (sw_410_clk_out),
        .data_out        (sw_410_data_out),
        .scan_select_out (sw_410_scan_out),
        .latch_enable_out(sw_410_latch_out)
    );

    // [411] https://github.com/mattvenn/wokwi_filler
    wire sw_411_clk_out, sw_411_data_out, sw_411_scan_out, sw_411_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_411 (
        .clk_in          (sw_410_clk_out),
        .data_in         (sw_410_data_out),
        .scan_select_in  (sw_410_scan_out),
        .latch_enable_in (sw_410_latch_out),
        .clk_out         (sw_411_clk_out),
        .data_out        (sw_411_data_out),
        .scan_select_out (sw_411_scan_out),
        .latch_enable_out(sw_411_latch_out)
    );

    // [412] https://github.com/mattvenn/wokwi_filler
    wire sw_412_clk_out, sw_412_data_out, sw_412_scan_out, sw_412_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_412 (
        .clk_in          (sw_411_clk_out),
        .data_in         (sw_411_data_out),
        .scan_select_in  (sw_411_scan_out),
        .latch_enable_in (sw_411_latch_out),
        .clk_out         (sw_412_clk_out),
        .data_out        (sw_412_data_out),
        .scan_select_out (sw_412_scan_out),
        .latch_enable_out(sw_412_latch_out)
    );

    // [413] https://github.com/mattvenn/wokwi_filler
    wire sw_413_clk_out, sw_413_data_out, sw_413_scan_out, sw_413_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_413 (
        .clk_in          (sw_412_clk_out),
        .data_in         (sw_412_data_out),
        .scan_select_in  (sw_412_scan_out),
        .latch_enable_in (sw_412_latch_out),
        .clk_out         (sw_413_clk_out),
        .data_out        (sw_413_data_out),
        .scan_select_out (sw_413_scan_out),
        .latch_enable_out(sw_413_latch_out)
    );

    // [414] https://github.com/mattvenn/wokwi_filler
    wire sw_414_clk_out, sw_414_data_out, sw_414_scan_out, sw_414_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_414 (
        .clk_in          (sw_413_clk_out),
        .data_in         (sw_413_data_out),
        .scan_select_in  (sw_413_scan_out),
        .latch_enable_in (sw_413_latch_out),
        .clk_out         (sw_414_clk_out),
        .data_out        (sw_414_data_out),
        .scan_select_out (sw_414_scan_out),
        .latch_enable_out(sw_414_latch_out)
    );

    // [415] https://github.com/mattvenn/wokwi_filler
    wire sw_415_clk_out, sw_415_data_out, sw_415_scan_out, sw_415_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_415 (
        .clk_in          (sw_414_clk_out),
        .data_in         (sw_414_data_out),
        .scan_select_in  (sw_414_scan_out),
        .latch_enable_in (sw_414_latch_out),
        .clk_out         (sw_415_clk_out),
        .data_out        (sw_415_data_out),
        .scan_select_out (sw_415_scan_out),
        .latch_enable_out(sw_415_latch_out)
    );

    // [416] https://github.com/mattvenn/wokwi_filler
    wire sw_416_clk_out, sw_416_data_out, sw_416_scan_out, sw_416_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_416 (
        .clk_in          (sw_415_clk_out),
        .data_in         (sw_415_data_out),
        .scan_select_in  (sw_415_scan_out),
        .latch_enable_in (sw_415_latch_out),
        .clk_out         (sw_416_clk_out),
        .data_out        (sw_416_data_out),
        .scan_select_out (sw_416_scan_out),
        .latch_enable_out(sw_416_latch_out)
    );

    // [417] https://github.com/mattvenn/wokwi_filler
    wire sw_417_clk_out, sw_417_data_out, sw_417_scan_out, sw_417_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_417 (
        .clk_in          (sw_416_clk_out),
        .data_in         (sw_416_data_out),
        .scan_select_in  (sw_416_scan_out),
        .latch_enable_in (sw_416_latch_out),
        .clk_out         (sw_417_clk_out),
        .data_out        (sw_417_data_out),
        .scan_select_out (sw_417_scan_out),
        .latch_enable_out(sw_417_latch_out)
    );

    // [418] https://github.com/mattvenn/wokwi_filler
    wire sw_418_clk_out, sw_418_data_out, sw_418_scan_out, sw_418_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_418 (
        .clk_in          (sw_417_clk_out),
        .data_in         (sw_417_data_out),
        .scan_select_in  (sw_417_scan_out),
        .latch_enable_in (sw_417_latch_out),
        .clk_out         (sw_418_clk_out),
        .data_out        (sw_418_data_out),
        .scan_select_out (sw_418_scan_out),
        .latch_enable_out(sw_418_latch_out)
    );

    // [419] https://github.com/mattvenn/wokwi_filler
    wire sw_419_clk_out, sw_419_data_out, sw_419_scan_out, sw_419_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_419 (
        .clk_in          (sw_418_clk_out),
        .data_in         (sw_418_data_out),
        .scan_select_in  (sw_418_scan_out),
        .latch_enable_in (sw_418_latch_out),
        .clk_out         (sw_419_clk_out),
        .data_out        (sw_419_data_out),
        .scan_select_out (sw_419_scan_out),
        .latch_enable_out(sw_419_latch_out)
    );

    // [420] https://github.com/mattvenn/wokwi_filler
    wire sw_420_clk_out, sw_420_data_out, sw_420_scan_out, sw_420_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_420 (
        .clk_in          (sw_419_clk_out),
        .data_in         (sw_419_data_out),
        .scan_select_in  (sw_419_scan_out),
        .latch_enable_in (sw_419_latch_out),
        .clk_out         (sw_420_clk_out),
        .data_out        (sw_420_data_out),
        .scan_select_out (sw_420_scan_out),
        .latch_enable_out(sw_420_latch_out)
    );

    // [421] https://github.com/mattvenn/wokwi_filler
    wire sw_421_clk_out, sw_421_data_out, sw_421_scan_out, sw_421_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_421 (
        .clk_in          (sw_420_clk_out),
        .data_in         (sw_420_data_out),
        .scan_select_in  (sw_420_scan_out),
        .latch_enable_in (sw_420_latch_out),
        .clk_out         (sw_421_clk_out),
        .data_out        (sw_421_data_out),
        .scan_select_out (sw_421_scan_out),
        .latch_enable_out(sw_421_latch_out)
    );

    // [422] https://github.com/mattvenn/wokwi_filler
    wire sw_422_clk_out, sw_422_data_out, sw_422_scan_out, sw_422_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_422 (
        .clk_in          (sw_421_clk_out),
        .data_in         (sw_421_data_out),
        .scan_select_in  (sw_421_scan_out),
        .latch_enable_in (sw_421_latch_out),
        .clk_out         (sw_422_clk_out),
        .data_out        (sw_422_data_out),
        .scan_select_out (sw_422_scan_out),
        .latch_enable_out(sw_422_latch_out)
    );

    // [423] https://github.com/mattvenn/wokwi_filler
    wire sw_423_clk_out, sw_423_data_out, sw_423_scan_out, sw_423_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_423 (
        .clk_in          (sw_422_clk_out),
        .data_in         (sw_422_data_out),
        .scan_select_in  (sw_422_scan_out),
        .latch_enable_in (sw_422_latch_out),
        .clk_out         (sw_423_clk_out),
        .data_out        (sw_423_data_out),
        .scan_select_out (sw_423_scan_out),
        .latch_enable_out(sw_423_latch_out)
    );

    // [424] https://github.com/mattvenn/wokwi_filler
    wire sw_424_clk_out, sw_424_data_out, sw_424_scan_out, sw_424_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_424 (
        .clk_in          (sw_423_clk_out),
        .data_in         (sw_423_data_out),
        .scan_select_in  (sw_423_scan_out),
        .latch_enable_in (sw_423_latch_out),
        .clk_out         (sw_424_clk_out),
        .data_out        (sw_424_data_out),
        .scan_select_out (sw_424_scan_out),
        .latch_enable_out(sw_424_latch_out)
    );

    // [425] https://github.com/mattvenn/wokwi_filler
    wire sw_425_clk_out, sw_425_data_out, sw_425_scan_out, sw_425_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_425 (
        .clk_in          (sw_424_clk_out),
        .data_in         (sw_424_data_out),
        .scan_select_in  (sw_424_scan_out),
        .latch_enable_in (sw_424_latch_out),
        .clk_out         (sw_425_clk_out),
        .data_out        (sw_425_data_out),
        .scan_select_out (sw_425_scan_out),
        .latch_enable_out(sw_425_latch_out)
    );

    // [426] https://github.com/mattvenn/wokwi_filler
    wire sw_426_clk_out, sw_426_data_out, sw_426_scan_out, sw_426_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_426 (
        .clk_in          (sw_425_clk_out),
        .data_in         (sw_425_data_out),
        .scan_select_in  (sw_425_scan_out),
        .latch_enable_in (sw_425_latch_out),
        .clk_out         (sw_426_clk_out),
        .data_out        (sw_426_data_out),
        .scan_select_out (sw_426_scan_out),
        .latch_enable_out(sw_426_latch_out)
    );

    // [427] https://github.com/mattvenn/wokwi_filler
    wire sw_427_clk_out, sw_427_data_out, sw_427_scan_out, sw_427_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_427 (
        .clk_in          (sw_426_clk_out),
        .data_in         (sw_426_data_out),
        .scan_select_in  (sw_426_scan_out),
        .latch_enable_in (sw_426_latch_out),
        .clk_out         (sw_427_clk_out),
        .data_out        (sw_427_data_out),
        .scan_select_out (sw_427_scan_out),
        .latch_enable_out(sw_427_latch_out)
    );

    // [428] https://github.com/mattvenn/wokwi_filler
    wire sw_428_clk_out, sw_428_data_out, sw_428_scan_out, sw_428_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_428 (
        .clk_in          (sw_427_clk_out),
        .data_in         (sw_427_data_out),
        .scan_select_in  (sw_427_scan_out),
        .latch_enable_in (sw_427_latch_out),
        .clk_out         (sw_428_clk_out),
        .data_out        (sw_428_data_out),
        .scan_select_out (sw_428_scan_out),
        .latch_enable_out(sw_428_latch_out)
    );

    // [429] https://github.com/mattvenn/wokwi_filler
    wire sw_429_clk_out, sw_429_data_out, sw_429_scan_out, sw_429_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_429 (
        .clk_in          (sw_428_clk_out),
        .data_in         (sw_428_data_out),
        .scan_select_in  (sw_428_scan_out),
        .latch_enable_in (sw_428_latch_out),
        .clk_out         (sw_429_clk_out),
        .data_out        (sw_429_data_out),
        .scan_select_out (sw_429_scan_out),
        .latch_enable_out(sw_429_latch_out)
    );

    // [430] https://github.com/mattvenn/wokwi_filler
    wire sw_430_clk_out, sw_430_data_out, sw_430_scan_out, sw_430_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_430 (
        .clk_in          (sw_429_clk_out),
        .data_in         (sw_429_data_out),
        .scan_select_in  (sw_429_scan_out),
        .latch_enable_in (sw_429_latch_out),
        .clk_out         (sw_430_clk_out),
        .data_out        (sw_430_data_out),
        .scan_select_out (sw_430_scan_out),
        .latch_enable_out(sw_430_latch_out)
    );

    // [431] https://github.com/mattvenn/wokwi_filler
    wire sw_431_clk_out, sw_431_data_out, sw_431_scan_out, sw_431_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_431 (
        .clk_in          (sw_430_clk_out),
        .data_in         (sw_430_data_out),
        .scan_select_in  (sw_430_scan_out),
        .latch_enable_in (sw_430_latch_out),
        .clk_out         (sw_431_clk_out),
        .data_out        (sw_431_data_out),
        .scan_select_out (sw_431_scan_out),
        .latch_enable_out(sw_431_latch_out)
    );

    // [432] https://github.com/mattvenn/wokwi_filler
    wire sw_432_clk_out, sw_432_data_out, sw_432_scan_out, sw_432_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_432 (
        .clk_in          (sw_431_clk_out),
        .data_in         (sw_431_data_out),
        .scan_select_in  (sw_431_scan_out),
        .latch_enable_in (sw_431_latch_out),
        .clk_out         (sw_432_clk_out),
        .data_out        (sw_432_data_out),
        .scan_select_out (sw_432_scan_out),
        .latch_enable_out(sw_432_latch_out)
    );

    // [433] https://github.com/mattvenn/wokwi_filler
    wire sw_433_clk_out, sw_433_data_out, sw_433_scan_out, sw_433_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_433 (
        .clk_in          (sw_432_clk_out),
        .data_in         (sw_432_data_out),
        .scan_select_in  (sw_432_scan_out),
        .latch_enable_in (sw_432_latch_out),
        .clk_out         (sw_433_clk_out),
        .data_out        (sw_433_data_out),
        .scan_select_out (sw_433_scan_out),
        .latch_enable_out(sw_433_latch_out)
    );

    // [434] https://github.com/mattvenn/wokwi_filler
    wire sw_434_clk_out, sw_434_data_out, sw_434_scan_out, sw_434_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_434 (
        .clk_in          (sw_433_clk_out),
        .data_in         (sw_433_data_out),
        .scan_select_in  (sw_433_scan_out),
        .latch_enable_in (sw_433_latch_out),
        .clk_out         (sw_434_clk_out),
        .data_out        (sw_434_data_out),
        .scan_select_out (sw_434_scan_out),
        .latch_enable_out(sw_434_latch_out)
    );

    // [435] https://github.com/mattvenn/wokwi_filler
    wire sw_435_clk_out, sw_435_data_out, sw_435_scan_out, sw_435_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_435 (
        .clk_in          (sw_434_clk_out),
        .data_in         (sw_434_data_out),
        .scan_select_in  (sw_434_scan_out),
        .latch_enable_in (sw_434_latch_out),
        .clk_out         (sw_435_clk_out),
        .data_out        (sw_435_data_out),
        .scan_select_out (sw_435_scan_out),
        .latch_enable_out(sw_435_latch_out)
    );

    // [436] https://github.com/mattvenn/wokwi_filler
    wire sw_436_clk_out, sw_436_data_out, sw_436_scan_out, sw_436_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_436 (
        .clk_in          (sw_435_clk_out),
        .data_in         (sw_435_data_out),
        .scan_select_in  (sw_435_scan_out),
        .latch_enable_in (sw_435_latch_out),
        .clk_out         (sw_436_clk_out),
        .data_out        (sw_436_data_out),
        .scan_select_out (sw_436_scan_out),
        .latch_enable_out(sw_436_latch_out)
    );

    // [437] https://github.com/mattvenn/wokwi_filler
    wire sw_437_clk_out, sw_437_data_out, sw_437_scan_out, sw_437_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_437 (
        .clk_in          (sw_436_clk_out),
        .data_in         (sw_436_data_out),
        .scan_select_in  (sw_436_scan_out),
        .latch_enable_in (sw_436_latch_out),
        .clk_out         (sw_437_clk_out),
        .data_out        (sw_437_data_out),
        .scan_select_out (sw_437_scan_out),
        .latch_enable_out(sw_437_latch_out)
    );

    // [438] https://github.com/mattvenn/wokwi_filler
    wire sw_438_clk_out, sw_438_data_out, sw_438_scan_out, sw_438_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_438 (
        .clk_in          (sw_437_clk_out),
        .data_in         (sw_437_data_out),
        .scan_select_in  (sw_437_scan_out),
        .latch_enable_in (sw_437_latch_out),
        .clk_out         (sw_438_clk_out),
        .data_out        (sw_438_data_out),
        .scan_select_out (sw_438_scan_out),
        .latch_enable_out(sw_438_latch_out)
    );

    // [439] https://github.com/mattvenn/wokwi_filler
    wire sw_439_clk_out, sw_439_data_out, sw_439_scan_out, sw_439_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_439 (
        .clk_in          (sw_438_clk_out),
        .data_in         (sw_438_data_out),
        .scan_select_in  (sw_438_scan_out),
        .latch_enable_in (sw_438_latch_out),
        .clk_out         (sw_439_clk_out),
        .data_out        (sw_439_data_out),
        .scan_select_out (sw_439_scan_out),
        .latch_enable_out(sw_439_latch_out)
    );

    // [440] https://github.com/mattvenn/wokwi_filler
    wire sw_440_clk_out, sw_440_data_out, sw_440_scan_out, sw_440_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_440 (
        .clk_in          (sw_439_clk_out),
        .data_in         (sw_439_data_out),
        .scan_select_in  (sw_439_scan_out),
        .latch_enable_in (sw_439_latch_out),
        .clk_out         (sw_440_clk_out),
        .data_out        (sw_440_data_out),
        .scan_select_out (sw_440_scan_out),
        .latch_enable_out(sw_440_latch_out)
    );

    // [441] https://github.com/mattvenn/wokwi_filler
    wire sw_441_clk_out, sw_441_data_out, sw_441_scan_out, sw_441_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_441 (
        .clk_in          (sw_440_clk_out),
        .data_in         (sw_440_data_out),
        .scan_select_in  (sw_440_scan_out),
        .latch_enable_in (sw_440_latch_out),
        .clk_out         (sw_441_clk_out),
        .data_out        (sw_441_data_out),
        .scan_select_out (sw_441_scan_out),
        .latch_enable_out(sw_441_latch_out)
    );

    // [442] https://github.com/mattvenn/wokwi_filler
    wire sw_442_clk_out, sw_442_data_out, sw_442_scan_out, sw_442_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_442 (
        .clk_in          (sw_441_clk_out),
        .data_in         (sw_441_data_out),
        .scan_select_in  (sw_441_scan_out),
        .latch_enable_in (sw_441_latch_out),
        .clk_out         (sw_442_clk_out),
        .data_out        (sw_442_data_out),
        .scan_select_out (sw_442_scan_out),
        .latch_enable_out(sw_442_latch_out)
    );

    // [443] https://github.com/mattvenn/wokwi_filler
    wire sw_443_clk_out, sw_443_data_out, sw_443_scan_out, sw_443_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_443 (
        .clk_in          (sw_442_clk_out),
        .data_in         (sw_442_data_out),
        .scan_select_in  (sw_442_scan_out),
        .latch_enable_in (sw_442_latch_out),
        .clk_out         (sw_443_clk_out),
        .data_out        (sw_443_data_out),
        .scan_select_out (sw_443_scan_out),
        .latch_enable_out(sw_443_latch_out)
    );

    // [444] https://github.com/mattvenn/wokwi_filler
    wire sw_444_clk_out, sw_444_data_out, sw_444_scan_out, sw_444_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_444 (
        .clk_in          (sw_443_clk_out),
        .data_in         (sw_443_data_out),
        .scan_select_in  (sw_443_scan_out),
        .latch_enable_in (sw_443_latch_out),
        .clk_out         (sw_444_clk_out),
        .data_out        (sw_444_data_out),
        .scan_select_out (sw_444_scan_out),
        .latch_enable_out(sw_444_latch_out)
    );

    // [445] https://github.com/mattvenn/wokwi_filler
    wire sw_445_clk_out, sw_445_data_out, sw_445_scan_out, sw_445_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_445 (
        .clk_in          (sw_444_clk_out),
        .data_in         (sw_444_data_out),
        .scan_select_in  (sw_444_scan_out),
        .latch_enable_in (sw_444_latch_out),
        .clk_out         (sw_445_clk_out),
        .data_out        (sw_445_data_out),
        .scan_select_out (sw_445_scan_out),
        .latch_enable_out(sw_445_latch_out)
    );

    // [446] https://github.com/mattvenn/wokwi_filler
    wire sw_446_clk_out, sw_446_data_out, sw_446_scan_out, sw_446_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_446 (
        .clk_in          (sw_445_clk_out),
        .data_in         (sw_445_data_out),
        .scan_select_in  (sw_445_scan_out),
        .latch_enable_in (sw_445_latch_out),
        .clk_out         (sw_446_clk_out),
        .data_out        (sw_446_data_out),
        .scan_select_out (sw_446_scan_out),
        .latch_enable_out(sw_446_latch_out)
    );

    // [447] https://github.com/mattvenn/wokwi_filler
    wire sw_447_clk_out, sw_447_data_out, sw_447_scan_out, sw_447_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_447 (
        .clk_in          (sw_446_clk_out),
        .data_in         (sw_446_data_out),
        .scan_select_in  (sw_446_scan_out),
        .latch_enable_in (sw_446_latch_out),
        .clk_out         (sw_447_clk_out),
        .data_out        (sw_447_data_out),
        .scan_select_out (sw_447_scan_out),
        .latch_enable_out(sw_447_latch_out)
    );

    // [448] https://github.com/mattvenn/wokwi_filler
    wire sw_448_clk_out, sw_448_data_out, sw_448_scan_out, sw_448_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_448 (
        .clk_in          (sw_447_clk_out),
        .data_in         (sw_447_data_out),
        .scan_select_in  (sw_447_scan_out),
        .latch_enable_in (sw_447_latch_out),
        .clk_out         (sw_448_clk_out),
        .data_out        (sw_448_data_out),
        .scan_select_out (sw_448_scan_out),
        .latch_enable_out(sw_448_latch_out)
    );

    // [449] https://github.com/mattvenn/wokwi_filler
    wire sw_449_clk_out, sw_449_data_out, sw_449_scan_out, sw_449_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_449 (
        .clk_in          (sw_448_clk_out),
        .data_in         (sw_448_data_out),
        .scan_select_in  (sw_448_scan_out),
        .latch_enable_in (sw_448_latch_out),
        .clk_out         (sw_449_clk_out),
        .data_out        (sw_449_data_out),
        .scan_select_out (sw_449_scan_out),
        .latch_enable_out(sw_449_latch_out)
    );

    // [450] https://github.com/mattvenn/wokwi_filler
    wire sw_450_clk_out, sw_450_data_out, sw_450_scan_out, sw_450_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_450 (
        .clk_in          (sw_449_clk_out),
        .data_in         (sw_449_data_out),
        .scan_select_in  (sw_449_scan_out),
        .latch_enable_in (sw_449_latch_out),
        .clk_out         (sw_450_clk_out),
        .data_out        (sw_450_data_out),
        .scan_select_out (sw_450_scan_out),
        .latch_enable_out(sw_450_latch_out)
    );

    // [451] https://github.com/mattvenn/wokwi_filler
    wire sw_451_clk_out, sw_451_data_out, sw_451_scan_out, sw_451_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_451 (
        .clk_in          (sw_450_clk_out),
        .data_in         (sw_450_data_out),
        .scan_select_in  (sw_450_scan_out),
        .latch_enable_in (sw_450_latch_out),
        .clk_out         (sw_451_clk_out),
        .data_out        (sw_451_data_out),
        .scan_select_out (sw_451_scan_out),
        .latch_enable_out(sw_451_latch_out)
    );

    // [452] https://github.com/mattvenn/wokwi_filler
    wire sw_452_clk_out, sw_452_data_out, sw_452_scan_out, sw_452_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_452 (
        .clk_in          (sw_451_clk_out),
        .data_in         (sw_451_data_out),
        .scan_select_in  (sw_451_scan_out),
        .latch_enable_in (sw_451_latch_out),
        .clk_out         (sw_452_clk_out),
        .data_out        (sw_452_data_out),
        .scan_select_out (sw_452_scan_out),
        .latch_enable_out(sw_452_latch_out)
    );

    // [453] https://github.com/mattvenn/wokwi_filler
    wire sw_453_clk_out, sw_453_data_out, sw_453_scan_out, sw_453_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_453 (
        .clk_in          (sw_452_clk_out),
        .data_in         (sw_452_data_out),
        .scan_select_in  (sw_452_scan_out),
        .latch_enable_in (sw_452_latch_out),
        .clk_out         (sw_453_clk_out),
        .data_out        (sw_453_data_out),
        .scan_select_out (sw_453_scan_out),
        .latch_enable_out(sw_453_latch_out)
    );

    // [454] https://github.com/mattvenn/wokwi_filler
    wire sw_454_clk_out, sw_454_data_out, sw_454_scan_out, sw_454_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_454 (
        .clk_in          (sw_453_clk_out),
        .data_in         (sw_453_data_out),
        .scan_select_in  (sw_453_scan_out),
        .latch_enable_in (sw_453_latch_out),
        .clk_out         (sw_454_clk_out),
        .data_out        (sw_454_data_out),
        .scan_select_out (sw_454_scan_out),
        .latch_enable_out(sw_454_latch_out)
    );

    // [455] https://github.com/mattvenn/wokwi_filler
    wire sw_455_clk_out, sw_455_data_out, sw_455_scan_out, sw_455_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_455 (
        .clk_in          (sw_454_clk_out),
        .data_in         (sw_454_data_out),
        .scan_select_in  (sw_454_scan_out),
        .latch_enable_in (sw_454_latch_out),
        .clk_out         (sw_455_clk_out),
        .data_out        (sw_455_data_out),
        .scan_select_out (sw_455_scan_out),
        .latch_enable_out(sw_455_latch_out)
    );

    // [456] https://github.com/mattvenn/wokwi_filler
    wire sw_456_clk_out, sw_456_data_out, sw_456_scan_out, sw_456_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_456 (
        .clk_in          (sw_455_clk_out),
        .data_in         (sw_455_data_out),
        .scan_select_in  (sw_455_scan_out),
        .latch_enable_in (sw_455_latch_out),
        .clk_out         (sw_456_clk_out),
        .data_out        (sw_456_data_out),
        .scan_select_out (sw_456_scan_out),
        .latch_enable_out(sw_456_latch_out)
    );

    // [457] https://github.com/mattvenn/wokwi_filler
    wire sw_457_clk_out, sw_457_data_out, sw_457_scan_out, sw_457_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_457 (
        .clk_in          (sw_456_clk_out),
        .data_in         (sw_456_data_out),
        .scan_select_in  (sw_456_scan_out),
        .latch_enable_in (sw_456_latch_out),
        .clk_out         (sw_457_clk_out),
        .data_out        (sw_457_data_out),
        .scan_select_out (sw_457_scan_out),
        .latch_enable_out(sw_457_latch_out)
    );

    // [458] https://github.com/mattvenn/wokwi_filler
    wire sw_458_clk_out, sw_458_data_out, sw_458_scan_out, sw_458_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_458 (
        .clk_in          (sw_457_clk_out),
        .data_in         (sw_457_data_out),
        .scan_select_in  (sw_457_scan_out),
        .latch_enable_in (sw_457_latch_out),
        .clk_out         (sw_458_clk_out),
        .data_out        (sw_458_data_out),
        .scan_select_out (sw_458_scan_out),
        .latch_enable_out(sw_458_latch_out)
    );

    // [459] https://github.com/mattvenn/wokwi_filler
    wire sw_459_clk_out, sw_459_data_out, sw_459_scan_out, sw_459_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_459 (
        .clk_in          (sw_458_clk_out),
        .data_in         (sw_458_data_out),
        .scan_select_in  (sw_458_scan_out),
        .latch_enable_in (sw_458_latch_out),
        .clk_out         (sw_459_clk_out),
        .data_out        (sw_459_data_out),
        .scan_select_out (sw_459_scan_out),
        .latch_enable_out(sw_459_latch_out)
    );

    // [460] https://github.com/mattvenn/wokwi_filler
    wire sw_460_clk_out, sw_460_data_out, sw_460_scan_out, sw_460_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_460 (
        .clk_in          (sw_459_clk_out),
        .data_in         (sw_459_data_out),
        .scan_select_in  (sw_459_scan_out),
        .latch_enable_in (sw_459_latch_out),
        .clk_out         (sw_460_clk_out),
        .data_out        (sw_460_data_out),
        .scan_select_out (sw_460_scan_out),
        .latch_enable_out(sw_460_latch_out)
    );

    // [461] https://github.com/mattvenn/wokwi_filler
    wire sw_461_clk_out, sw_461_data_out, sw_461_scan_out, sw_461_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_461 (
        .clk_in          (sw_460_clk_out),
        .data_in         (sw_460_data_out),
        .scan_select_in  (sw_460_scan_out),
        .latch_enable_in (sw_460_latch_out),
        .clk_out         (sw_461_clk_out),
        .data_out        (sw_461_data_out),
        .scan_select_out (sw_461_scan_out),
        .latch_enable_out(sw_461_latch_out)
    );

    // [462] https://github.com/mattvenn/wokwi_filler
    wire sw_462_clk_out, sw_462_data_out, sw_462_scan_out, sw_462_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_462 (
        .clk_in          (sw_461_clk_out),
        .data_in         (sw_461_data_out),
        .scan_select_in  (sw_461_scan_out),
        .latch_enable_in (sw_461_latch_out),
        .clk_out         (sw_462_clk_out),
        .data_out        (sw_462_data_out),
        .scan_select_out (sw_462_scan_out),
        .latch_enable_out(sw_462_latch_out)
    );

    // [463] https://github.com/mattvenn/wokwi_filler
    wire sw_463_clk_out, sw_463_data_out, sw_463_scan_out, sw_463_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_463 (
        .clk_in          (sw_462_clk_out),
        .data_in         (sw_462_data_out),
        .scan_select_in  (sw_462_scan_out),
        .latch_enable_in (sw_462_latch_out),
        .clk_out         (sw_463_clk_out),
        .data_out        (sw_463_data_out),
        .scan_select_out (sw_463_scan_out),
        .latch_enable_out(sw_463_latch_out)
    );

    // [464] https://github.com/mattvenn/wokwi_filler
    wire sw_464_clk_out, sw_464_data_out, sw_464_scan_out, sw_464_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_464 (
        .clk_in          (sw_463_clk_out),
        .data_in         (sw_463_data_out),
        .scan_select_in  (sw_463_scan_out),
        .latch_enable_in (sw_463_latch_out),
        .clk_out         (sw_464_clk_out),
        .data_out        (sw_464_data_out),
        .scan_select_out (sw_464_scan_out),
        .latch_enable_out(sw_464_latch_out)
    );

    // [465] https://github.com/mattvenn/wokwi_filler
    wire sw_465_clk_out, sw_465_data_out, sw_465_scan_out, sw_465_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_465 (
        .clk_in          (sw_464_clk_out),
        .data_in         (sw_464_data_out),
        .scan_select_in  (sw_464_scan_out),
        .latch_enable_in (sw_464_latch_out),
        .clk_out         (sw_465_clk_out),
        .data_out        (sw_465_data_out),
        .scan_select_out (sw_465_scan_out),
        .latch_enable_out(sw_465_latch_out)
    );

    // [466] https://github.com/mattvenn/wokwi_filler
    wire sw_466_clk_out, sw_466_data_out, sw_466_scan_out, sw_466_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_466 (
        .clk_in          (sw_465_clk_out),
        .data_in         (sw_465_data_out),
        .scan_select_in  (sw_465_scan_out),
        .latch_enable_in (sw_465_latch_out),
        .clk_out         (sw_466_clk_out),
        .data_out        (sw_466_data_out),
        .scan_select_out (sw_466_scan_out),
        .latch_enable_out(sw_466_latch_out)
    );

    // [467] https://github.com/mattvenn/wokwi_filler
    wire sw_467_clk_out, sw_467_data_out, sw_467_scan_out, sw_467_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_467 (
        .clk_in          (sw_466_clk_out),
        .data_in         (sw_466_data_out),
        .scan_select_in  (sw_466_scan_out),
        .latch_enable_in (sw_466_latch_out),
        .clk_out         (sw_467_clk_out),
        .data_out        (sw_467_data_out),
        .scan_select_out (sw_467_scan_out),
        .latch_enable_out(sw_467_latch_out)
    );

    // [468] https://github.com/mattvenn/wokwi_filler
    wire sw_468_clk_out, sw_468_data_out, sw_468_scan_out, sw_468_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_468 (
        .clk_in          (sw_467_clk_out),
        .data_in         (sw_467_data_out),
        .scan_select_in  (sw_467_scan_out),
        .latch_enable_in (sw_467_latch_out),
        .clk_out         (sw_468_clk_out),
        .data_out        (sw_468_data_out),
        .scan_select_out (sw_468_scan_out),
        .latch_enable_out(sw_468_latch_out)
    );

    // [469] https://github.com/mattvenn/wokwi_filler
    wire sw_469_clk_out, sw_469_data_out, sw_469_scan_out, sw_469_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_469 (
        .clk_in          (sw_468_clk_out),
        .data_in         (sw_468_data_out),
        .scan_select_in  (sw_468_scan_out),
        .latch_enable_in (sw_468_latch_out),
        .clk_out         (sw_469_clk_out),
        .data_out        (sw_469_data_out),
        .scan_select_out (sw_469_scan_out),
        .latch_enable_out(sw_469_latch_out)
    );

    // [470] https://github.com/mattvenn/wokwi_filler
    wire sw_470_clk_out, sw_470_data_out, sw_470_scan_out, sw_470_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_470 (
        .clk_in          (sw_469_clk_out),
        .data_in         (sw_469_data_out),
        .scan_select_in  (sw_469_scan_out),
        .latch_enable_in (sw_469_latch_out),
        .clk_out         (sw_470_clk_out),
        .data_out        (sw_470_data_out),
        .scan_select_out (sw_470_scan_out),
        .latch_enable_out(sw_470_latch_out)
    );

    // [471] https://github.com/mattvenn/wokwi_filler
    wire sw_471_clk_out, sw_471_data_out, sw_471_scan_out, sw_471_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_471 (
        .clk_in          (sw_470_clk_out),
        .data_in         (sw_470_data_out),
        .scan_select_in  (sw_470_scan_out),
        .latch_enable_in (sw_470_latch_out),
        .clk_out         (sw_471_clk_out),
        .data_out        (sw_471_data_out),
        .scan_select_out (sw_471_scan_out),
        .latch_enable_out(sw_471_latch_out)
    );

    // [472] https://github.com/mattvenn/wokwi_filler
    wire sw_472_clk_out, sw_472_data_out, sw_472_scan_out, sw_472_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_472 (
        .clk_in          (sw_471_clk_out),
        .data_in         (sw_471_data_out),
        .scan_select_in  (sw_471_scan_out),
        .latch_enable_in (sw_471_latch_out),
        .clk_out         (sw_472_clk_out),
        .data_out        (sw_472_data_out),
        .scan_select_out (sw_472_scan_out),
        .latch_enable_out(sw_472_latch_out)
    );

    // [473] https://github.com/mattvenn/wokwi_filler
    wire sw_473_clk_out, sw_473_data_out, sw_473_scan_out, sw_473_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_473 (
        .clk_in          (sw_472_clk_out),
        .data_in         (sw_472_data_out),
        .scan_select_in  (sw_472_scan_out),
        .latch_enable_in (sw_472_latch_out),
        .clk_out         (sw_473_clk_out),
        .data_out        (sw_473_data_out),
        .scan_select_out (sw_473_scan_out),
        .latch_enable_out(sw_473_latch_out)
    );

    // [474] https://github.com/mattvenn/wokwi_filler
    wire sw_474_clk_out, sw_474_data_out, sw_474_scan_out, sw_474_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_474 (
        .clk_in          (sw_473_clk_out),
        .data_in         (sw_473_data_out),
        .scan_select_in  (sw_473_scan_out),
        .latch_enable_in (sw_473_latch_out),
        .clk_out         (sw_474_clk_out),
        .data_out        (sw_474_data_out),
        .scan_select_out (sw_474_scan_out),
        .latch_enable_out(sw_474_latch_out)
    );

    // [475] https://github.com/mattvenn/wokwi_filler
    wire sw_475_clk_out, sw_475_data_out, sw_475_scan_out, sw_475_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_475 (
        .clk_in          (sw_474_clk_out),
        .data_in         (sw_474_data_out),
        .scan_select_in  (sw_474_scan_out),
        .latch_enable_in (sw_474_latch_out),
        .clk_out         (sw_475_clk_out),
        .data_out        (sw_475_data_out),
        .scan_select_out (sw_475_scan_out),
        .latch_enable_out(sw_475_latch_out)
    );

    // [476] https://github.com/mattvenn/wokwi_filler
    wire sw_476_clk_out, sw_476_data_out, sw_476_scan_out, sw_476_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_476 (
        .clk_in          (sw_475_clk_out),
        .data_in         (sw_475_data_out),
        .scan_select_in  (sw_475_scan_out),
        .latch_enable_in (sw_475_latch_out),
        .clk_out         (sw_476_clk_out),
        .data_out        (sw_476_data_out),
        .scan_select_out (sw_476_scan_out),
        .latch_enable_out(sw_476_latch_out)
    );

    // [477] https://github.com/mattvenn/wokwi_filler
    wire sw_477_clk_out, sw_477_data_out, sw_477_scan_out, sw_477_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_477 (
        .clk_in          (sw_476_clk_out),
        .data_in         (sw_476_data_out),
        .scan_select_in  (sw_476_scan_out),
        .latch_enable_in (sw_476_latch_out),
        .clk_out         (sw_477_clk_out),
        .data_out        (sw_477_data_out),
        .scan_select_out (sw_477_scan_out),
        .latch_enable_out(sw_477_latch_out)
    );

    // [478] https://github.com/mattvenn/wokwi_filler
    wire sw_478_clk_out, sw_478_data_out, sw_478_scan_out, sw_478_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_478 (
        .clk_in          (sw_477_clk_out),
        .data_in         (sw_477_data_out),
        .scan_select_in  (sw_477_scan_out),
        .latch_enable_in (sw_477_latch_out),
        .clk_out         (sw_478_clk_out),
        .data_out        (sw_478_data_out),
        .scan_select_out (sw_478_scan_out),
        .latch_enable_out(sw_478_latch_out)
    );

    // [479] https://github.com/mattvenn/wokwi_filler
    wire sw_479_clk_out, sw_479_data_out, sw_479_scan_out, sw_479_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_479 (
        .clk_in          (sw_478_clk_out),
        .data_in         (sw_478_data_out),
        .scan_select_in  (sw_478_scan_out),
        .latch_enable_in (sw_478_latch_out),
        .clk_out         (sw_479_clk_out),
        .data_out        (sw_479_data_out),
        .scan_select_out (sw_479_scan_out),
        .latch_enable_out(sw_479_latch_out)
    );

    // [480] https://github.com/mattvenn/wokwi_filler
    wire sw_480_clk_out, sw_480_data_out, sw_480_scan_out, sw_480_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_480 (
        .clk_in          (sw_479_clk_out),
        .data_in         (sw_479_data_out),
        .scan_select_in  (sw_479_scan_out),
        .latch_enable_in (sw_479_latch_out),
        .clk_out         (sw_480_clk_out),
        .data_out        (sw_480_data_out),
        .scan_select_out (sw_480_scan_out),
        .latch_enable_out(sw_480_latch_out)
    );

    // [481] https://github.com/mattvenn/wokwi_filler
    wire sw_481_clk_out, sw_481_data_out, sw_481_scan_out, sw_481_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_481 (
        .clk_in          (sw_480_clk_out),
        .data_in         (sw_480_data_out),
        .scan_select_in  (sw_480_scan_out),
        .latch_enable_in (sw_480_latch_out),
        .clk_out         (sw_481_clk_out),
        .data_out        (sw_481_data_out),
        .scan_select_out (sw_481_scan_out),
        .latch_enable_out(sw_481_latch_out)
    );

    // [482] https://github.com/mattvenn/wokwi_filler
    wire sw_482_clk_out, sw_482_data_out, sw_482_scan_out, sw_482_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_482 (
        .clk_in          (sw_481_clk_out),
        .data_in         (sw_481_data_out),
        .scan_select_in  (sw_481_scan_out),
        .latch_enable_in (sw_481_latch_out),
        .clk_out         (sw_482_clk_out),
        .data_out        (sw_482_data_out),
        .scan_select_out (sw_482_scan_out),
        .latch_enable_out(sw_482_latch_out)
    );

    // [483] https://github.com/mattvenn/wokwi_filler
    wire sw_483_clk_out, sw_483_data_out, sw_483_scan_out, sw_483_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_483 (
        .clk_in          (sw_482_clk_out),
        .data_in         (sw_482_data_out),
        .scan_select_in  (sw_482_scan_out),
        .latch_enable_in (sw_482_latch_out),
        .clk_out         (sw_483_clk_out),
        .data_out        (sw_483_data_out),
        .scan_select_out (sw_483_scan_out),
        .latch_enable_out(sw_483_latch_out)
    );

    // [484] https://github.com/mattvenn/wokwi_filler
    wire sw_484_clk_out, sw_484_data_out, sw_484_scan_out, sw_484_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_484 (
        .clk_in          (sw_483_clk_out),
        .data_in         (sw_483_data_out),
        .scan_select_in  (sw_483_scan_out),
        .latch_enable_in (sw_483_latch_out),
        .clk_out         (sw_484_clk_out),
        .data_out        (sw_484_data_out),
        .scan_select_out (sw_484_scan_out),
        .latch_enable_out(sw_484_latch_out)
    );

    // [485] https://github.com/mattvenn/wokwi_filler
    wire sw_485_clk_out, sw_485_data_out, sw_485_scan_out, sw_485_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_485 (
        .clk_in          (sw_484_clk_out),
        .data_in         (sw_484_data_out),
        .scan_select_in  (sw_484_scan_out),
        .latch_enable_in (sw_484_latch_out),
        .clk_out         (sw_485_clk_out),
        .data_out        (sw_485_data_out),
        .scan_select_out (sw_485_scan_out),
        .latch_enable_out(sw_485_latch_out)
    );

    // [486] https://github.com/mattvenn/wokwi_filler
    wire sw_486_clk_out, sw_486_data_out, sw_486_scan_out, sw_486_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_486 (
        .clk_in          (sw_485_clk_out),
        .data_in         (sw_485_data_out),
        .scan_select_in  (sw_485_scan_out),
        .latch_enable_in (sw_485_latch_out),
        .clk_out         (sw_486_clk_out),
        .data_out        (sw_486_data_out),
        .scan_select_out (sw_486_scan_out),
        .latch_enable_out(sw_486_latch_out)
    );

    // [487] https://github.com/mattvenn/wokwi_filler
    wire sw_487_clk_out, sw_487_data_out, sw_487_scan_out, sw_487_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_487 (
        .clk_in          (sw_486_clk_out),
        .data_in         (sw_486_data_out),
        .scan_select_in  (sw_486_scan_out),
        .latch_enable_in (sw_486_latch_out),
        .clk_out         (sw_487_clk_out),
        .data_out        (sw_487_data_out),
        .scan_select_out (sw_487_scan_out),
        .latch_enable_out(sw_487_latch_out)
    );

    // [488] https://github.com/mattvenn/wokwi_filler
    wire sw_488_clk_out, sw_488_data_out, sw_488_scan_out, sw_488_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_488 (
        .clk_in          (sw_487_clk_out),
        .data_in         (sw_487_data_out),
        .scan_select_in  (sw_487_scan_out),
        .latch_enable_in (sw_487_latch_out),
        .clk_out         (sw_488_clk_out),
        .data_out        (sw_488_data_out),
        .scan_select_out (sw_488_scan_out),
        .latch_enable_out(sw_488_latch_out)
    );

    // [489] https://github.com/mattvenn/wokwi_filler
    wire sw_489_clk_out, sw_489_data_out, sw_489_scan_out, sw_489_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_489 (
        .clk_in          (sw_488_clk_out),
        .data_in         (sw_488_data_out),
        .scan_select_in  (sw_488_scan_out),
        .latch_enable_in (sw_488_latch_out),
        .clk_out         (sw_489_clk_out),
        .data_out        (sw_489_data_out),
        .scan_select_out (sw_489_scan_out),
        .latch_enable_out(sw_489_latch_out)
    );

    // [490] https://github.com/mattvenn/wokwi_filler
    wire sw_490_clk_out, sw_490_data_out, sw_490_scan_out, sw_490_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_490 (
        .clk_in          (sw_489_clk_out),
        .data_in         (sw_489_data_out),
        .scan_select_in  (sw_489_scan_out),
        .latch_enable_in (sw_489_latch_out),
        .clk_out         (sw_490_clk_out),
        .data_out        (sw_490_data_out),
        .scan_select_out (sw_490_scan_out),
        .latch_enable_out(sw_490_latch_out)
    );

    // [491] https://github.com/mattvenn/wokwi_filler
    wire sw_491_clk_out, sw_491_data_out, sw_491_scan_out, sw_491_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_491 (
        .clk_in          (sw_490_clk_out),
        .data_in         (sw_490_data_out),
        .scan_select_in  (sw_490_scan_out),
        .latch_enable_in (sw_490_latch_out),
        .clk_out         (sw_491_clk_out),
        .data_out        (sw_491_data_out),
        .scan_select_out (sw_491_scan_out),
        .latch_enable_out(sw_491_latch_out)
    );

    // [492] https://github.com/mattvenn/wokwi_filler
    wire sw_492_clk_out, sw_492_data_out, sw_492_scan_out, sw_492_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_492 (
        .clk_in          (sw_491_clk_out),
        .data_in         (sw_491_data_out),
        .scan_select_in  (sw_491_scan_out),
        .latch_enable_in (sw_491_latch_out),
        .clk_out         (sw_492_clk_out),
        .data_out        (sw_492_data_out),
        .scan_select_out (sw_492_scan_out),
        .latch_enable_out(sw_492_latch_out)
    );

    // [493] https://github.com/mattvenn/wokwi_filler
    wire sw_493_clk_out, sw_493_data_out, sw_493_scan_out, sw_493_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_493 (
        .clk_in          (sw_492_clk_out),
        .data_in         (sw_492_data_out),
        .scan_select_in  (sw_492_scan_out),
        .latch_enable_in (sw_492_latch_out),
        .clk_out         (sw_493_clk_out),
        .data_out        (sw_493_data_out),
        .scan_select_out (sw_493_scan_out),
        .latch_enable_out(sw_493_latch_out)
    );

    // [494] https://github.com/mattvenn/wokwi_filler
    wire sw_494_clk_out, sw_494_data_out, sw_494_scan_out, sw_494_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_494 (
        .clk_in          (sw_493_clk_out),
        .data_in         (sw_493_data_out),
        .scan_select_in  (sw_493_scan_out),
        .latch_enable_in (sw_493_latch_out),
        .clk_out         (sw_494_clk_out),
        .data_out        (sw_494_data_out),
        .scan_select_out (sw_494_scan_out),
        .latch_enable_out(sw_494_latch_out)
    );

    // [495] https://github.com/mattvenn/wokwi_filler
    wire sw_495_clk_out, sw_495_data_out, sw_495_scan_out, sw_495_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_495 (
        .clk_in          (sw_494_clk_out),
        .data_in         (sw_494_data_out),
        .scan_select_in  (sw_494_scan_out),
        .latch_enable_in (sw_494_latch_out),
        .clk_out         (sw_495_clk_out),
        .data_out        (sw_495_data_out),
        .scan_select_out (sw_495_scan_out),
        .latch_enable_out(sw_495_latch_out)
    );

    // [496] https://github.com/mattvenn/wokwi_filler
    wire sw_496_clk_out, sw_496_data_out, sw_496_scan_out, sw_496_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_496 (
        .clk_in          (sw_495_clk_out),
        .data_in         (sw_495_data_out),
        .scan_select_in  (sw_495_scan_out),
        .latch_enable_in (sw_495_latch_out),
        .clk_out         (sw_496_clk_out),
        .data_out        (sw_496_data_out),
        .scan_select_out (sw_496_scan_out),
        .latch_enable_out(sw_496_latch_out)
    );

    // [497] https://github.com/mattvenn/wokwi_filler
    wire sw_497_clk_out, sw_497_data_out, sw_497_scan_out, sw_497_latch_out;
    scan_wrapper_339501025136214612 #(.NUM_IOS(8)) scan_wrapper_339501025136214612_497 (
        .clk_in          (sw_496_clk_out),
        .data_in         (sw_496_data_out),
        .scan_select_in  (sw_496_scan_out),
        .latch_enable_in (sw_496_latch_out),
        .clk_out         (sw_497_clk_out),
        .data_out        (sw_497_data_out),
        .scan_select_out (sw_497_scan_out),
        .latch_enable_out(sw_497_latch_out)
    );

    // Connect final signals back to the scan controller
    assign sc_clk_in  = sw_497_clk_out;
    assign sc_data_in = sw_497_data_out;

    // end of module instantiation

endmodule	// user_project_wrapper
`default_nettype wire
