    // end of module instantiation

endmodule	// user_project_wrapper
`default_nettype wire
