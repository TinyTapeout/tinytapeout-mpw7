VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO scan_wrapper_341631511790879314
  CLASS BLOCK ;
  FOREIGN scan_wrapper_341631511790879314 ;
  ORIGIN 0.000 0.000 ;
  SIZE 105.000 BY 105.000 ;
  PIN clk_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 101.000 103.410 105.000 ;
    END
  END clk_in
  PIN clk_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END clk_out
  PIN data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.000 51.040 105.000 51.640 ;
    END
  END data_in
  PIN data_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END data_out
  PIN latch_enable_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END latch_enable_in
  PIN latch_enable_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 101.000 0.370 105.000 ;
    END
  END latch_enable_out
  PIN scan_select_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 101.000 51.890 105.000 ;
    END
  END scan_select_in
  PIN scan_select_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END scan_select_out
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 16.465 10.640 18.065 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.955 10.640 41.555 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.445 10.640 65.045 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 86.935 10.640 88.535 92.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 28.210 10.640 29.810 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.700 10.640 53.300 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.190 10.640 76.790 92.720 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 99.360 92.565 ;
      LAYER met1 ;
        RECT 0.070 10.640 103.430 92.720 ;
      LAYER met2 ;
        RECT 0.650 100.720 51.330 101.730 ;
        RECT 52.170 100.720 102.850 101.730 ;
        RECT 0.100 4.280 103.400 100.720 ;
        RECT 0.650 4.000 51.330 4.280 ;
        RECT 52.170 4.000 102.850 4.280 ;
      LAYER met3 ;
        RECT 4.000 52.040 101.000 92.645 ;
        RECT 4.400 50.640 100.600 52.040 ;
        RECT 4.000 10.715 101.000 50.640 ;
  END
END scan_wrapper_341631511790879314
END LIBRARY

