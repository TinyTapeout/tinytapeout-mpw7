magic
tech sky130B
magscale 1 2
timestamp 1662135081
<< metal1 >>
rect 36538 700612 36544 700664
rect 36596 700652 36602 700664
rect 105446 700652 105452 700664
rect 36596 700624 105452 700652
rect 36596 700612 36602 700624
rect 105446 700612 105452 700624
rect 105504 700612 105510 700664
rect 71038 700544 71044 700596
rect 71096 700584 71102 700596
rect 267642 700584 267648 700596
rect 71096 700556 267648 700584
rect 71096 700544 71102 700556
rect 267642 700544 267648 700556
rect 267700 700544 267706 700596
rect 13446 700476 13452 700528
rect 13504 700516 13510 700528
rect 300118 700516 300124 700528
rect 13504 700488 300124 700516
rect 13504 700476 13510 700488
rect 300118 700476 300124 700488
rect 300176 700476 300182 700528
rect 322198 700476 322204 700528
rect 322256 700516 322262 700528
rect 332502 700516 332508 700528
rect 322256 700488 332508 700516
rect 322256 700476 322262 700488
rect 332502 700476 332508 700488
rect 332560 700476 332566 700528
rect 65518 700408 65524 700460
rect 65576 700448 65582 700460
rect 137830 700448 137836 700460
rect 65576 700420 137836 700448
rect 65576 700408 65582 700420
rect 137830 700408 137836 700420
rect 137888 700408 137894 700460
rect 153838 700408 153844 700460
rect 153896 700448 153902 700460
rect 170306 700448 170312 700460
rect 153896 700420 170312 700448
rect 153896 700408 153902 700420
rect 170306 700408 170312 700420
rect 170364 700408 170370 700460
rect 204898 700408 204904 700460
rect 204956 700448 204962 700460
rect 494790 700448 494796 700460
rect 204956 700420 494796 700448
rect 204956 700408 204962 700420
rect 494790 700408 494796 700420
rect 494848 700408 494854 700460
rect 64138 700340 64144 700392
rect 64196 700380 64202 700392
rect 364978 700380 364984 700392
rect 64196 700352 364984 700380
rect 64196 700340 64202 700352
rect 364978 700340 364984 700352
rect 365036 700340 365042 700392
rect 378778 700340 378784 700392
rect 378836 700380 378842 700392
rect 397454 700380 397460 700392
rect 378836 700352 397460 700380
rect 378836 700340 378842 700352
rect 397454 700340 397460 700352
rect 397512 700340 397518 700392
rect 518158 700340 518164 700392
rect 518216 700380 518222 700392
rect 527174 700380 527180 700392
rect 518216 700352 527180 700380
rect 518216 700340 518222 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 64230 700272 64236 700324
rect 64288 700312 64294 700324
rect 202782 700312 202788 700324
rect 64288 700284 202788 700312
rect 64288 700272 64294 700284
rect 202782 700272 202788 700284
rect 202840 700272 202846 700324
rect 233878 700272 233884 700324
rect 233936 700312 233942 700324
rect 559650 700312 559656 700324
rect 233936 700284 559656 700312
rect 233936 700272 233942 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 40494 699932 40500 699984
rect 40552 699972 40558 699984
rect 42058 699972 42064 699984
rect 40552 699944 42064 699972
rect 40552 699932 40558 699944
rect 42058 699932 42064 699944
rect 42116 699932 42122 699984
rect 65610 699660 65616 699712
rect 65668 699700 65674 699712
rect 72970 699700 72976 699712
rect 65668 699672 72976 699700
rect 65668 699660 65674 699672
rect 72970 699660 72976 699672
rect 73028 699660 73034 699712
rect 65702 696940 65708 696992
rect 65760 696980 65766 696992
rect 580166 696980 580172 696992
rect 65760 696952 580172 696980
rect 65760 696940 65766 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 212350 686060 212356 686112
rect 212408 686100 212414 686112
rect 232682 686100 232688 686112
rect 212408 686072 232688 686100
rect 212408 686060 212414 686072
rect 232682 686060 232688 686072
rect 232740 686060 232746 686112
rect 296346 686060 296352 686112
rect 296404 686100 296410 686112
rect 316770 686100 316776 686112
rect 296404 686072 316776 686100
rect 296404 686060 296410 686072
rect 316770 686060 316776 686072
rect 316828 686060 316834 686112
rect 408034 686060 408040 686112
rect 408092 686100 408098 686112
rect 428642 686100 428648 686112
rect 408092 686072 428648 686100
rect 408092 686060 408098 686072
rect 428642 686060 428648 686072
rect 428700 686060 428706 686112
rect 492030 686060 492036 686112
rect 492088 686100 492094 686112
rect 512730 686100 512736 686112
rect 492088 686072 512736 686100
rect 492088 686060 492094 686072
rect 512730 686060 512736 686072
rect 512788 686060 512794 686112
rect 148318 685992 148324 686044
rect 148376 686032 148382 686044
rect 165706 686032 165712 686044
rect 148376 686004 165712 686032
rect 148376 685992 148382 686004
rect 165706 685992 165712 686004
rect 165764 685992 165770 686044
rect 175458 685992 175464 686044
rect 175516 686032 175522 686044
rect 193674 686032 193680 686044
rect 175516 686004 193680 686032
rect 175516 685992 175522 686004
rect 193674 685992 193680 686004
rect 193732 685992 193738 686044
rect 203518 685992 203524 686044
rect 203576 686032 203582 686044
rect 221366 686032 221372 686044
rect 203576 686004 221372 686032
rect 203576 685992 203582 686004
rect 221366 685992 221372 686004
rect 221424 685992 221430 686044
rect 260098 685992 260104 686044
rect 260156 686032 260162 686044
rect 277670 686032 277676 686044
rect 260156 686004 277676 686032
rect 260156 685992 260162 686004
rect 277670 685992 277676 686004
rect 277728 685992 277734 686044
rect 287514 685992 287520 686044
rect 287572 686032 287578 686044
rect 305362 686032 305368 686044
rect 287572 686004 305368 686032
rect 287572 685992 287578 686004
rect 305362 685992 305368 686004
rect 305420 685992 305426 686044
rect 345658 685992 345664 686044
rect 345716 686032 345722 686044
rect 361666 686032 361672 686044
rect 345716 686004 361672 686032
rect 345716 685992 345722 686004
rect 361666 685992 361672 686004
rect 361724 685992 361730 686044
rect 371510 685992 371516 686044
rect 371568 686032 371574 686044
rect 389358 686032 389364 686044
rect 371568 686004 389364 686032
rect 371568 685992 371574 686004
rect 389358 685992 389364 686004
rect 389416 685992 389422 686044
rect 399478 685992 399484 686044
rect 399536 686032 399542 686044
rect 417694 686032 417700 686044
rect 399536 686004 417700 686032
rect 399536 685992 399542 686004
rect 417694 685992 417700 686004
rect 417752 685992 417758 686044
rect 456058 685992 456064 686044
rect 456116 686032 456122 686044
rect 473354 686032 473360 686044
rect 456116 686004 473360 686032
rect 456116 685992 456122 686004
rect 473354 685992 473360 686004
rect 473412 685992 473418 686044
rect 483474 685992 483480 686044
rect 483532 686032 483538 686044
rect 501690 686032 501696 686044
rect 483532 686004 501696 686032
rect 483532 685992 483538 686004
rect 501690 685992 501696 686004
rect 501748 685992 501754 686044
rect 36722 685924 36728 685976
rect 36780 685964 36786 685976
rect 53650 685964 53656 685976
rect 36780 685936 53656 685964
rect 36780 685924 36786 685936
rect 53650 685924 53656 685936
rect 53708 685924 53714 685976
rect 64322 685924 64328 685976
rect 64380 685964 64386 685976
rect 81434 685964 81440 685976
rect 64380 685936 81440 685964
rect 64380 685924 64386 685936
rect 81434 685924 81440 685936
rect 81492 685924 81498 685976
rect 91462 685924 91468 685976
rect 91520 685964 91526 685976
rect 109678 685964 109684 685976
rect 91520 685936 109684 685964
rect 91520 685924 91526 685936
rect 109678 685924 109684 685936
rect 109736 685924 109742 685976
rect 119430 685924 119436 685976
rect 119488 685964 119494 685976
rect 137646 685964 137652 685976
rect 119488 685936 137652 685964
rect 119488 685924 119494 685936
rect 137646 685924 137652 685936
rect 137704 685924 137710 685976
rect 156322 685924 156328 685976
rect 156380 685964 156386 685976
rect 178678 685964 178684 685976
rect 156380 685936 178684 685964
rect 156380 685924 156386 685936
rect 178678 685924 178684 685936
rect 178736 685924 178742 685976
rect 232590 685924 232596 685976
rect 232648 685964 232654 685976
rect 249702 685964 249708 685976
rect 232648 685936 249708 685964
rect 232648 685924 232654 685936
rect 249702 685924 249708 685936
rect 249760 685924 249766 685976
rect 268010 685924 268016 685976
rect 268068 685964 268074 685976
rect 287698 685964 287704 685976
rect 268068 685936 287704 685964
rect 268068 685924 268074 685936
rect 287698 685924 287704 685936
rect 287756 685924 287762 685976
rect 315482 685924 315488 685976
rect 315540 685964 315546 685976
rect 333698 685964 333704 685976
rect 315540 685936 333704 685964
rect 315540 685924 315546 685936
rect 333698 685924 333704 685936
rect 333756 685924 333762 685976
rect 352006 685924 352012 685976
rect 352064 685964 352070 685976
rect 374638 685964 374644 685976
rect 352064 685936 374644 685964
rect 352064 685924 352070 685936
rect 374638 685924 374644 685936
rect 374696 685924 374702 685976
rect 428550 685924 428556 685976
rect 428608 685964 428614 685976
rect 445662 685964 445668 685976
rect 428608 685936 445668 685964
rect 428608 685924 428614 685936
rect 445662 685924 445668 685936
rect 445720 685924 445726 685976
rect 464338 685924 464344 685976
rect 464396 685964 464402 685976
rect 483658 685964 483664 685976
rect 464396 685936 483664 685964
rect 464396 685924 464402 685936
rect 483658 685924 483664 685936
rect 483716 685924 483722 685976
rect 511442 685924 511448 685976
rect 511500 685964 511506 685976
rect 529658 685964 529664 685976
rect 511500 685936 529664 685964
rect 511500 685924 511506 685936
rect 529658 685924 529664 685936
rect 529716 685924 529722 685976
rect 541618 685924 541624 685976
rect 541676 685964 541682 685976
rect 557534 685964 557540 685976
rect 541676 685936 557540 685964
rect 541676 685924 541682 685936
rect 557534 685924 557540 685936
rect 557592 685924 557598 685976
rect 16114 685856 16120 685908
rect 16172 685896 16178 685908
rect 25682 685896 25688 685908
rect 16172 685868 25688 685896
rect 16172 685856 16178 685868
rect 25682 685856 25688 685868
rect 25740 685856 25746 685908
rect 36630 685856 36636 685908
rect 36688 685896 36694 685908
rect 63310 685896 63316 685908
rect 36688 685868 63316 685896
rect 36688 685856 36694 685868
rect 63310 685856 63316 685868
rect 63368 685856 63374 685908
rect 66898 685856 66904 685908
rect 66956 685896 66962 685908
rect 91094 685896 91100 685908
rect 66956 685868 91100 685896
rect 66956 685856 66962 685868
rect 91094 685856 91100 685868
rect 91152 685856 91158 685908
rect 93118 685856 93124 685908
rect 93176 685896 93182 685908
rect 119338 685896 119344 685908
rect 93176 685868 119344 685896
rect 93176 685856 93182 685868
rect 119338 685856 119344 685868
rect 119396 685856 119402 685908
rect 122098 685856 122104 685908
rect 122156 685896 122162 685908
rect 147306 685896 147312 685908
rect 122156 685868 147312 685896
rect 122156 685856 122162 685868
rect 147306 685856 147312 685868
rect 147364 685856 147370 685908
rect 148410 685856 148416 685908
rect 148468 685896 148474 685908
rect 175366 685896 175372 685908
rect 148468 685868 175372 685896
rect 148468 685856 148474 685868
rect 175366 685856 175372 685868
rect 175424 685856 175430 685908
rect 177298 685856 177304 685908
rect 177356 685896 177362 685908
rect 203334 685896 203340 685908
rect 177356 685868 203340 685896
rect 177356 685856 177362 685868
rect 203334 685856 203340 685868
rect 203392 685856 203398 685908
rect 204990 685856 204996 685908
rect 205048 685896 205054 685908
rect 231026 685896 231032 685908
rect 205048 685868 231032 685896
rect 205048 685856 205054 685868
rect 231026 685856 231032 685868
rect 231084 685856 231090 685908
rect 232498 685856 232504 685908
rect 232556 685896 232562 685908
rect 259362 685896 259368 685908
rect 232556 685868 259368 685896
rect 232556 685856 232562 685868
rect 259362 685856 259368 685868
rect 259420 685856 259426 685908
rect 260190 685856 260196 685908
rect 260248 685896 260254 685908
rect 287330 685896 287336 685908
rect 260248 685868 287336 685896
rect 260248 685856 260254 685868
rect 287330 685856 287336 685868
rect 287388 685856 287394 685908
rect 289078 685856 289084 685908
rect 289136 685896 289142 685908
rect 315022 685896 315028 685908
rect 289136 685868 315028 685896
rect 289136 685856 289142 685868
rect 315022 685856 315028 685868
rect 315080 685856 315086 685908
rect 316678 685856 316684 685908
rect 316736 685896 316742 685908
rect 343358 685896 343364 685908
rect 316736 685868 343364 685896
rect 316736 685856 316742 685868
rect 343358 685856 343364 685868
rect 343416 685856 343422 685908
rect 344278 685856 344284 685908
rect 344336 685896 344342 685908
rect 371326 685896 371332 685908
rect 344336 685868 371332 685896
rect 344336 685856 344342 685868
rect 371326 685856 371332 685868
rect 371384 685856 371390 685908
rect 373258 685856 373264 685908
rect 373316 685896 373322 685908
rect 399018 685896 399024 685908
rect 373316 685868 399024 685896
rect 373316 685856 373322 685868
rect 399018 685856 399024 685868
rect 399076 685856 399082 685908
rect 400858 685856 400864 685908
rect 400916 685896 400922 685908
rect 427354 685896 427360 685908
rect 400916 685868 427360 685896
rect 400916 685856 400922 685868
rect 427354 685856 427360 685868
rect 427412 685856 427418 685908
rect 428458 685856 428464 685908
rect 428516 685896 428522 685908
rect 455322 685896 455328 685908
rect 428516 685868 455328 685896
rect 428516 685856 428522 685868
rect 455322 685856 455328 685868
rect 455380 685856 455386 685908
rect 456150 685856 456156 685908
rect 456208 685896 456214 685908
rect 483014 685896 483020 685908
rect 456208 685868 483020 685896
rect 456208 685856 456214 685868
rect 483014 685856 483020 685868
rect 483072 685856 483078 685908
rect 485038 685856 485044 685908
rect 485096 685896 485102 685908
rect 511350 685896 511356 685908
rect 485096 685868 511356 685896
rect 485096 685856 485102 685868
rect 511350 685856 511356 685868
rect 511408 685856 511414 685908
rect 512638 685856 512644 685908
rect 512696 685896 512702 685908
rect 539318 685896 539324 685908
rect 512696 685868 539324 685896
rect 512696 685856 512702 685868
rect 539318 685856 539324 685868
rect 539376 685856 539382 685908
rect 540238 685856 540244 685908
rect 540296 685896 540302 685908
rect 567194 685896 567200 685908
rect 540296 685868 567200 685896
rect 540296 685856 540302 685868
rect 567194 685856 567200 685868
rect 567252 685856 567258 685908
rect 15838 683272 15844 683324
rect 15896 683312 15902 683324
rect 16114 683312 16120 683324
rect 15896 683284 16120 683312
rect 15896 683272 15902 683284
rect 16114 683272 16120 683284
rect 16172 683272 16178 683324
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 43438 683244 43444 683256
rect 3476 683216 43444 683244
rect 3476 683204 3482 683216
rect 43438 683204 43444 683216
rect 43496 683204 43502 683256
rect 182082 683204 182088 683256
rect 182140 683244 182146 683256
rect 233234 683244 233240 683256
rect 182140 683216 233240 683244
rect 182140 683204 182146 683216
rect 233234 683204 233240 683216
rect 233292 683204 233298 683256
rect 350442 683204 350448 683256
rect 350500 683244 350506 683256
rect 401594 683244 401600 683256
rect 350500 683216 401600 683244
rect 350500 683204 350506 683216
rect 401594 683204 401600 683216
rect 401652 683204 401658 683256
rect 42702 683136 42708 683188
rect 42760 683176 42766 683188
rect 93854 683176 93860 683188
rect 42760 683148 93860 683176
rect 42760 683136 42766 683148
rect 93854 683136 93860 683148
rect 93912 683136 93918 683188
rect 97902 683136 97908 683188
rect 97960 683176 97966 683188
rect 149054 683176 149060 683188
rect 97960 683148 149060 683176
rect 97960 683136 97966 683148
rect 149054 683136 149060 683148
rect 149112 683136 149118 683188
rect 154482 683136 154488 683188
rect 154540 683176 154546 683188
rect 205634 683176 205640 683188
rect 154540 683148 205640 683176
rect 154540 683136 154546 683148
rect 205634 683136 205640 683148
rect 205692 683136 205698 683188
rect 238662 683136 238668 683188
rect 238720 683176 238726 683188
rect 289814 683176 289820 683188
rect 238720 683148 289820 683176
rect 238720 683136 238726 683148
rect 289814 683136 289820 683148
rect 289872 683136 289878 683188
rect 293862 683136 293868 683188
rect 293920 683176 293926 683188
rect 345014 683176 345020 683188
rect 293920 683148 345020 683176
rect 293920 683136 293926 683148
rect 345014 683136 345020 683148
rect 345072 683136 345078 683188
rect 378042 683136 378048 683188
rect 378100 683176 378106 683188
rect 429286 683176 429292 683188
rect 378100 683148 429292 683176
rect 378100 683136 378106 683148
rect 429286 683136 429292 683148
rect 429344 683136 429350 683188
rect 434622 683136 434628 683188
rect 434680 683176 434686 683188
rect 485774 683176 485780 683188
rect 434680 683148 485780 683176
rect 434680 683136 434686 683148
rect 485774 683136 485780 683148
rect 485832 683136 485838 683188
rect 489822 683136 489828 683188
rect 489880 683176 489886 683188
rect 542354 683176 542360 683188
rect 489880 683148 542360 683176
rect 489880 683136 489886 683148
rect 542354 683136 542360 683148
rect 542412 683136 542418 683188
rect 542998 673752 543004 673804
rect 543056 673792 543062 673804
rect 545114 673792 545120 673804
rect 543056 673764 545120 673792
rect 543056 673752 543062 673764
rect 545114 673752 545120 673764
rect 545172 673752 545178 673804
rect 63586 668720 63592 668772
rect 63644 668760 63650 668772
rect 64322 668760 64328 668772
rect 63644 668732 64328 668760
rect 63644 668720 63650 668732
rect 64322 668720 64328 668732
rect 64380 668720 64386 668772
rect 428642 665796 428648 665848
rect 428700 665836 428706 665848
rect 435726 665836 435732 665848
rect 428700 665808 435732 665836
rect 428700 665796 428706 665808
rect 435726 665796 435732 665808
rect 435784 665796 435790 665848
rect 287698 665456 287704 665508
rect 287756 665496 287762 665508
rect 295702 665496 295708 665508
rect 287756 665468 295708 665496
rect 287756 665456 287762 665468
rect 295702 665456 295708 665468
rect 295760 665456 295766 665508
rect 316770 665456 316776 665508
rect 316828 665496 316834 665508
rect 323670 665496 323676 665508
rect 316828 665468 323676 665496
rect 316828 665456 316834 665468
rect 323670 665456 323676 665468
rect 323728 665456 323734 665508
rect 232682 665252 232688 665304
rect 232740 665292 232746 665304
rect 239766 665292 239772 665304
rect 232740 665264 239772 665292
rect 232740 665252 232746 665264
rect 239766 665252 239772 665264
rect 239824 665252 239830 665304
rect 483658 665252 483664 665304
rect 483716 665292 483722 665304
rect 491662 665292 491668 665304
rect 483716 665264 491668 665292
rect 483716 665252 483722 665264
rect 491662 665252 491668 665264
rect 491720 665252 491726 665304
rect 512730 665252 512736 665304
rect 512788 665292 512794 665304
rect 519630 665292 519636 665304
rect 512788 665264 519636 665292
rect 512788 665252 512794 665264
rect 519630 665252 519636 665264
rect 519688 665252 519694 665304
rect 13630 665116 13636 665168
rect 13688 665156 13694 665168
rect 66254 665156 66260 665168
rect 13688 665128 66260 665156
rect 13688 665116 13694 665128
rect 66254 665116 66260 665128
rect 66312 665116 66318 665168
rect 70302 665116 70308 665168
rect 70360 665156 70366 665168
rect 121454 665156 121460 665168
rect 70360 665128 121460 665156
rect 70360 665116 70366 665128
rect 121454 665116 121460 665128
rect 121512 665116 121518 665168
rect 126882 665116 126888 665168
rect 126940 665156 126946 665168
rect 178034 665156 178040 665168
rect 126940 665128 178040 665156
rect 126940 665116 126946 665128
rect 178034 665116 178040 665128
rect 178092 665116 178098 665168
rect 209682 665116 209688 665168
rect 209740 665156 209746 665168
rect 262214 665156 262220 665168
rect 209740 665128 262220 665156
rect 209740 665116 209746 665128
rect 262214 665116 262220 665128
rect 262272 665116 262278 665168
rect 266262 665116 266268 665168
rect 266320 665156 266326 665168
rect 317414 665156 317420 665168
rect 266320 665128 317420 665156
rect 266320 665116 266326 665128
rect 317414 665116 317420 665128
rect 317472 665116 317478 665168
rect 322842 665116 322848 665168
rect 322900 665156 322906 665168
rect 373994 665156 374000 665168
rect 322900 665128 374000 665156
rect 322900 665116 322906 665128
rect 373994 665116 374000 665128
rect 374052 665116 374058 665168
rect 405642 665116 405648 665168
rect 405700 665156 405706 665168
rect 458174 665156 458180 665168
rect 405700 665128 458180 665156
rect 405700 665116 405706 665128
rect 458174 665116 458180 665128
rect 458232 665116 458238 665168
rect 462222 665116 462228 665168
rect 462280 665156 462286 665168
rect 513374 665156 513380 665168
rect 462280 665128 513380 665156
rect 462280 665116 462286 665128
rect 513374 665116 513380 665128
rect 513432 665116 513438 665168
rect 518802 665116 518808 665168
rect 518860 665156 518866 665168
rect 569954 665156 569960 665168
rect 518860 665128 569960 665156
rect 518860 665116 518866 665128
rect 569954 665116 569960 665128
rect 570012 665116 570018 665168
rect 343542 665048 343548 665100
rect 343600 665088 343606 665100
rect 345658 665088 345664 665100
rect 343600 665060 345664 665088
rect 343600 665048 343606 665060
rect 345658 665048 345664 665060
rect 345716 665048 345722 665100
rect 427722 665048 427728 665100
rect 427780 665088 427786 665100
rect 428550 665088 428556 665100
rect 427780 665060 428556 665088
rect 427780 665048 427786 665060
rect 428550 665048 428556 665060
rect 428608 665048 428614 665100
rect 35250 664708 35256 664760
rect 35308 664748 35314 664760
rect 36722 664748 36728 664760
rect 35308 664720 36728 664748
rect 35308 664708 35314 664720
rect 36722 664708 36728 664720
rect 36780 664708 36786 664760
rect 15838 664096 15844 664148
rect 15896 664136 15902 664148
rect 16574 664136 16580 664148
rect 15896 664108 16580 664136
rect 15896 664096 15902 664108
rect 16574 664096 16580 664108
rect 16632 664096 16638 664148
rect 231578 663688 231584 663740
rect 231636 663728 231642 663740
rect 232590 663728 232596 663740
rect 231636 663700 232596 663728
rect 231636 663688 231642 663700
rect 232590 663688 232596 663700
rect 232648 663688 232654 663740
rect 539318 663688 539324 663740
rect 539376 663728 539382 663740
rect 541618 663728 541624 663740
rect 539376 663700 541624 663728
rect 539376 663688 539382 663700
rect 541618 663688 541624 663700
rect 541676 663688 541682 663740
rect 71866 662328 71872 662380
rect 71924 662368 71930 662380
rect 100018 662368 100024 662380
rect 71924 662340 100024 662368
rect 71924 662328 71930 662340
rect 100018 662328 100024 662340
rect 100076 662328 100082 662380
rect 127710 662368 127716 662380
rect 103486 662340 127716 662368
rect 25682 662260 25688 662312
rect 25740 662300 25746 662312
rect 36630 662300 36636 662312
rect 25740 662272 36636 662300
rect 25740 662260 25746 662272
rect 36630 662260 36636 662272
rect 36688 662260 36694 662312
rect 42886 662260 42892 662312
rect 42944 662300 42950 662312
rect 42944 662272 45554 662300
rect 42944 662260 42950 662272
rect 15286 662192 15292 662244
rect 15344 662232 15350 662244
rect 43622 662232 43628 662244
rect 15344 662204 43628 662232
rect 15344 662192 15350 662204
rect 43622 662192 43628 662204
rect 43680 662192 43686 662244
rect 45526 662232 45554 662272
rect 53742 662260 53748 662312
rect 53800 662300 53806 662312
rect 66898 662300 66904 662312
rect 53800 662272 66904 662300
rect 53800 662260 53806 662272
rect 66898 662260 66904 662272
rect 66956 662260 66962 662312
rect 81986 662260 81992 662312
rect 82044 662300 82050 662312
rect 93118 662300 93124 662312
rect 82044 662272 93124 662300
rect 82044 662260 82050 662272
rect 93118 662260 93124 662272
rect 93176 662260 93182 662312
rect 99466 662260 99472 662312
rect 99524 662300 99530 662312
rect 103486 662300 103514 662340
rect 127710 662328 127716 662340
rect 127768 662328 127774 662380
rect 165982 662328 165988 662380
rect 166040 662368 166046 662380
rect 177298 662368 177304 662380
rect 166040 662340 177304 662368
rect 166040 662328 166046 662340
rect 177298 662328 177304 662340
rect 177356 662328 177362 662380
rect 178678 662328 178684 662380
rect 178736 662368 178742 662380
rect 184014 662368 184020 662380
rect 178736 662340 184020 662368
rect 178736 662328 178742 662340
rect 184014 662328 184020 662340
rect 184072 662328 184078 662380
rect 211706 662368 211712 662380
rect 190426 662340 211712 662368
rect 99524 662272 103514 662300
rect 99524 662260 99530 662272
rect 109678 662260 109684 662312
rect 109736 662300 109742 662312
rect 122098 662300 122104 662312
rect 109736 662272 122104 662300
rect 109736 662260 109742 662272
rect 122098 662260 122104 662272
rect 122156 662260 122162 662312
rect 137922 662260 137928 662312
rect 137980 662300 137986 662312
rect 148410 662300 148416 662312
rect 137980 662272 148416 662300
rect 137980 662260 137986 662272
rect 148410 662260 148416 662272
rect 148468 662260 148474 662312
rect 183646 662260 183652 662312
rect 183704 662300 183710 662312
rect 190426 662300 190454 662340
rect 211706 662328 211712 662340
rect 211764 662328 211770 662380
rect 277670 662328 277676 662380
rect 277728 662368 277734 662380
rect 289078 662368 289084 662380
rect 277728 662340 289084 662368
rect 277728 662328 277734 662340
rect 289078 662328 289084 662340
rect 289136 662328 289142 662380
rect 306006 662328 306012 662380
rect 306064 662368 306070 662380
rect 316678 662368 316684 662380
rect 306064 662340 316684 662368
rect 306064 662328 306070 662340
rect 316678 662328 316684 662340
rect 316736 662328 316742 662380
rect 361666 662328 361672 662380
rect 361724 662368 361730 662380
rect 373258 662368 373264 662380
rect 361724 662340 373264 662368
rect 361724 662328 361730 662340
rect 373258 662328 373264 662340
rect 373316 662328 373322 662380
rect 379606 662328 379612 662380
rect 379664 662368 379670 662380
rect 408034 662368 408040 662380
rect 379664 662340 408040 662368
rect 379664 662328 379670 662340
rect 408034 662328 408040 662340
rect 408092 662328 408098 662380
rect 473998 662328 474004 662380
rect 474056 662368 474062 662380
rect 485038 662368 485044 662380
rect 474056 662340 485044 662368
rect 474056 662328 474062 662340
rect 485038 662328 485044 662340
rect 485096 662328 485102 662380
rect 501690 662328 501696 662380
rect 501748 662368 501754 662380
rect 512638 662368 512644 662380
rect 501748 662340 512644 662368
rect 501748 662328 501754 662340
rect 512638 662328 512644 662340
rect 512696 662328 512702 662380
rect 183704 662272 190454 662300
rect 183704 662260 183710 662272
rect 193674 662260 193680 662312
rect 193732 662300 193738 662312
rect 204990 662300 204996 662312
rect 193732 662272 204996 662300
rect 193732 662260 193738 662272
rect 204990 662260 204996 662272
rect 205048 662260 205054 662312
rect 222010 662260 222016 662312
rect 222068 662300 222074 662312
rect 232498 662300 232504 662312
rect 222068 662272 232504 662300
rect 222068 662260 222074 662272
rect 232498 662260 232504 662272
rect 232556 662260 232562 662312
rect 249610 662260 249616 662312
rect 249668 662300 249674 662312
rect 260190 662300 260196 662312
rect 249668 662272 260196 662300
rect 249668 662260 249674 662272
rect 260190 662260 260196 662272
rect 260248 662260 260254 662312
rect 333882 662260 333888 662312
rect 333940 662300 333946 662312
rect 344278 662300 344284 662312
rect 333940 662272 344284 662300
rect 333940 662260 333946 662272
rect 344278 662260 344284 662272
rect 344336 662260 344342 662312
rect 374638 662260 374644 662312
rect 374696 662300 374702 662312
rect 379698 662300 379704 662312
rect 374696 662272 379704 662300
rect 374696 662260 374702 662272
rect 379698 662260 379704 662272
rect 379756 662260 379762 662312
rect 390002 662260 390008 662312
rect 390060 662300 390066 662312
rect 400858 662300 400864 662312
rect 390060 662272 400864 662300
rect 390060 662260 390066 662272
rect 400858 662260 400864 662272
rect 400916 662260 400922 662312
rect 417694 662260 417700 662312
rect 417752 662300 417758 662312
rect 428458 662300 428464 662312
rect 417752 662272 428464 662300
rect 417752 662260 417758 662272
rect 428458 662260 428464 662272
rect 428516 662260 428522 662312
rect 445662 662260 445668 662312
rect 445720 662300 445726 662312
rect 456150 662300 456156 662312
rect 445720 662272 456156 662300
rect 445720 662260 445726 662272
rect 456150 662260 456156 662272
rect 456208 662260 456214 662312
rect 529658 662260 529664 662312
rect 529716 662300 529722 662312
rect 540238 662300 540244 662312
rect 529716 662272 540244 662300
rect 529716 662260 529722 662272
rect 540238 662260 540244 662272
rect 540296 662260 540302 662312
rect 71958 662232 71964 662244
rect 45526 662204 71964 662232
rect 71958 662192 71964 662204
rect 72016 662192 72022 662244
rect 127066 662192 127072 662244
rect 127124 662232 127130 662244
rect 155954 662232 155960 662244
rect 127124 662204 155960 662232
rect 127124 662192 127130 662204
rect 155954 662192 155960 662204
rect 156012 662192 156018 662244
rect 238846 662192 238852 662244
rect 238904 662232 238910 662244
rect 268010 662232 268016 662244
rect 238904 662204 268016 662232
rect 238904 662192 238910 662204
rect 268010 662192 268016 662204
rect 268068 662192 268074 662244
rect 323026 662192 323032 662244
rect 323084 662232 323090 662244
rect 352006 662232 352012 662244
rect 323084 662204 352012 662232
rect 323084 662192 323090 662204
rect 352006 662192 352012 662204
rect 352064 662192 352070 662244
rect 434806 662192 434812 662244
rect 434864 662232 434870 662244
rect 463786 662232 463792 662244
rect 434864 662204 463792 662232
rect 434864 662192 434870 662204
rect 463786 662192 463792 662204
rect 463844 662192 463850 662244
rect 518986 662192 518992 662244
rect 519044 662232 519050 662244
rect 547874 662232 547880 662244
rect 519044 662204 547880 662232
rect 519044 662192 519050 662204
rect 547874 662192 547880 662204
rect 547932 662192 547938 662244
rect 13630 661648 13636 661700
rect 13688 661688 13694 661700
rect 557534 661688 557540 661700
rect 13688 661660 557540 661688
rect 13688 661648 13694 661660
rect 557534 661648 557540 661660
rect 557592 661648 557598 661700
rect 267826 658452 267832 658504
rect 267884 658492 267890 658504
rect 267884 658464 277394 658492
rect 267884 658452 267890 658464
rect 71130 658384 71136 658436
rect 71188 658424 71194 658436
rect 82262 658424 82268 658436
rect 71188 658396 82268 658424
rect 71188 658384 71194 658396
rect 82262 658384 82268 658396
rect 82320 658384 82326 658436
rect 99466 658384 99472 658436
rect 99524 658424 99530 658436
rect 100386 658424 100392 658436
rect 99524 658396 100392 658424
rect 99524 658384 99530 658396
rect 100386 658384 100392 658396
rect 100444 658384 100450 658436
rect 183646 658384 183652 658436
rect 183704 658424 183710 658436
rect 222286 658424 222292 658436
rect 183704 658396 222292 658424
rect 183704 658384 183710 658396
rect 222286 658384 222292 658396
rect 222344 658384 222350 658436
rect 266998 658384 267004 658436
rect 267056 658424 267062 658436
rect 267056 658396 271276 658424
rect 267056 658384 267062 658396
rect 26234 658316 26240 658368
rect 26292 658356 26298 658368
rect 35434 658356 35440 658368
rect 26292 658328 35440 658356
rect 26292 658316 26298 658328
rect 35434 658316 35440 658328
rect 35492 658316 35498 658368
rect 36630 658316 36636 658368
rect 36688 658356 36694 658368
rect 53926 658356 53932 658368
rect 36688 658328 53932 658356
rect 36688 658316 36694 658328
rect 53926 658316 53932 658328
rect 53984 658316 53990 658368
rect 71866 658316 71872 658368
rect 71924 658356 71930 658368
rect 109954 658356 109960 658368
rect 71924 658328 109960 658356
rect 71924 658316 71930 658328
rect 109954 658316 109960 658328
rect 110012 658316 110018 658368
rect 124858 658316 124864 658368
rect 124916 658356 124922 658368
rect 128630 658356 128636 658368
rect 124916 658328 128636 658356
rect 124916 658316 124922 658328
rect 128630 658316 128636 658328
rect 128688 658316 128694 658368
rect 151078 658316 151084 658368
rect 151136 658356 151142 658368
rect 156598 658356 156604 658368
rect 151136 658328 156604 658356
rect 151136 658316 151142 658328
rect 156598 658316 156604 658328
rect 156656 658316 156662 658368
rect 182818 658316 182824 658368
rect 182876 658356 182882 658368
rect 193950 658356 193956 658368
rect 182876 658328 193956 658356
rect 182876 658316 182882 658328
rect 193950 658316 193956 658328
rect 194008 658316 194014 658368
rect 232498 658316 232504 658368
rect 232556 658356 232562 658368
rect 232556 658328 248414 658356
rect 232556 658316 232562 658328
rect 66898 658248 66904 658300
rect 66956 658288 66962 658300
rect 72602 658288 72608 658300
rect 66956 658260 72608 658288
rect 66956 658248 66962 658260
rect 72602 658248 72608 658260
rect 72660 658248 72666 658300
rect 93118 658248 93124 658300
rect 93176 658288 93182 658300
rect 100294 658288 100300 658300
rect 93176 658260 100300 658288
rect 93176 658248 93182 658260
rect 100294 658248 100300 658260
rect 100352 658248 100358 658300
rect 100386 658248 100392 658300
rect 100444 658288 100450 658300
rect 138290 658288 138296 658300
rect 100444 658260 138296 658288
rect 100444 658248 100450 658260
rect 138290 658248 138296 658260
rect 138348 658248 138354 658300
rect 149698 658248 149704 658300
rect 149756 658288 149762 658300
rect 166258 658288 166264 658300
rect 149756 658260 166264 658288
rect 149756 658248 149762 658260
rect 166258 658248 166264 658260
rect 166316 658248 166322 658300
rect 177298 658248 177304 658300
rect 177356 658288 177362 658300
rect 184290 658288 184296 658300
rect 177356 658260 184296 658288
rect 177356 658248 177362 658260
rect 184290 658248 184296 658260
rect 184348 658248 184354 658300
rect 233970 658248 233976 658300
rect 234028 658288 234034 658300
rect 240594 658288 240600 658300
rect 234028 658260 240600 658288
rect 234028 658248 234034 658260
rect 240594 658248 240600 658260
rect 240652 658248 240658 658300
rect 248386 658288 248414 658328
rect 250254 658288 250260 658300
rect 248386 658260 250260 658288
rect 250254 658248 250260 658260
rect 250312 658248 250318 658300
rect 261478 658248 261484 658300
rect 261536 658288 261542 658300
rect 268286 658288 268292 658300
rect 261536 658260 268292 658288
rect 261536 658248 261542 658260
rect 268286 658248 268292 658260
rect 268344 658248 268350 658300
rect 271248 658288 271276 658396
rect 277366 658356 277394 658464
rect 295426 658384 295432 658436
rect 295484 658424 295490 658436
rect 334250 658424 334256 658436
rect 295484 658396 334256 658424
rect 295484 658384 295490 658396
rect 334250 658384 334256 658396
rect 334308 658384 334314 658436
rect 352006 658384 352012 658436
rect 352064 658424 352070 658436
rect 352064 658396 364334 658424
rect 352064 658384 352070 658396
rect 306282 658356 306288 658368
rect 277366 658328 306288 658356
rect 306282 658316 306288 658328
rect 306340 658316 306346 658368
rect 347038 658316 347044 658368
rect 347096 658356 347102 658368
rect 361942 658356 361948 658368
rect 347096 658328 361948 658356
rect 347096 658316 347102 658328
rect 361942 658316 361948 658328
rect 362000 658316 362006 658368
rect 364306 658356 364334 658396
rect 379606 658384 379612 658436
rect 379664 658424 379670 658436
rect 418246 658424 418252 658436
rect 379664 658396 418252 658424
rect 379664 658384 379670 658396
rect 418246 658384 418252 658396
rect 418304 658384 418310 658436
rect 463786 658384 463792 658436
rect 463844 658424 463850 658436
rect 463844 658396 470594 658424
rect 463844 658384 463850 658396
rect 390278 658356 390284 658368
rect 364306 658328 390284 658356
rect 390278 658316 390284 658328
rect 390336 658316 390342 658368
rect 400858 658316 400864 658368
rect 400916 658356 400922 658368
rect 408586 658356 408592 658368
rect 400916 658328 408592 658356
rect 400916 658316 400922 658328
rect 408586 658316 408592 658328
rect 408644 658316 408650 658368
rect 429838 658316 429844 658368
rect 429896 658356 429902 658368
rect 436278 658356 436284 658368
rect 429896 658328 436284 658356
rect 429896 658316 429902 658328
rect 436278 658316 436284 658328
rect 436336 658316 436342 658368
rect 457438 658316 457444 658368
rect 457496 658356 457502 658368
rect 464614 658356 464620 658368
rect 457496 658328 464620 658356
rect 457496 658316 457502 658328
rect 464614 658316 464620 658328
rect 464672 658316 464678 658368
rect 470566 658356 470594 658396
rect 491386 658384 491392 658436
rect 491444 658424 491450 658436
rect 529934 658424 529940 658436
rect 491444 658396 529940 658424
rect 491444 658384 491450 658396
rect 529934 658384 529940 658396
rect 529992 658384 529998 658436
rect 502242 658356 502248 658368
rect 470566 658328 502248 658356
rect 502242 658316 502248 658328
rect 502300 658316 502306 658368
rect 512638 658316 512644 658368
rect 512696 658356 512702 658368
rect 520274 658356 520280 658368
rect 512696 658328 520280 658356
rect 512696 658316 512702 658328
rect 520274 658316 520280 658328
rect 520332 658316 520338 658368
rect 541618 658316 541624 658368
rect 541676 658356 541682 658368
rect 541676 658328 557534 658356
rect 541676 658316 541682 658328
rect 277946 658288 277952 658300
rect 271248 658260 277952 658288
rect 277946 658248 277952 658260
rect 278004 658248 278010 658300
rect 289078 658248 289084 658300
rect 289136 658288 289142 658300
rect 296622 658288 296628 658300
rect 289136 658260 296628 658288
rect 289136 658248 289142 658260
rect 296622 658248 296628 658260
rect 296680 658248 296686 658300
rect 318058 658248 318064 658300
rect 318116 658288 318122 658300
rect 324590 658288 324596 658300
rect 318116 658260 324596 658288
rect 318116 658248 318122 658260
rect 324590 658248 324596 658260
rect 324648 658248 324654 658300
rect 348418 658248 348424 658300
rect 348476 658288 348482 658300
rect 352282 658288 352288 658300
rect 348476 658260 352288 658288
rect 348476 658248 348482 658260
rect 352282 658248 352288 658260
rect 352340 658248 352346 658300
rect 373258 658248 373264 658300
rect 373316 658288 373322 658300
rect 380618 658288 380624 658300
rect 373316 658260 380624 658288
rect 373316 658248 373322 658260
rect 380618 658248 380624 658260
rect 380676 658248 380682 658300
rect 428458 658248 428464 658300
rect 428516 658288 428522 658300
rect 445938 658288 445944 658300
rect 428516 658260 445944 658288
rect 428516 658248 428522 658260
rect 445938 658248 445944 658260
rect 445996 658248 446002 658300
rect 462958 658248 462964 658300
rect 463016 658288 463022 658300
rect 474274 658288 474280 658300
rect 463016 658260 474280 658288
rect 463016 658248 463022 658260
rect 474274 658248 474280 658260
rect 474332 658248 474338 658300
rect 485038 658248 485044 658300
rect 485096 658288 485102 658300
rect 492582 658288 492588 658300
rect 485096 658260 492588 658288
rect 485096 658248 485102 658260
rect 492582 658248 492588 658260
rect 492640 658248 492646 658300
rect 544378 658248 544384 658300
rect 544436 658288 544442 658300
rect 548610 658288 548616 658300
rect 544436 658260 548616 658288
rect 544436 658248 544442 658260
rect 548610 658248 548616 658260
rect 548668 658248 548674 658300
rect 557506 658288 557534 658328
rect 558270 658288 558276 658300
rect 557506 658260 558276 658288
rect 558270 658248 558276 658260
rect 558328 658248 558334 658300
rect 2774 657500 2780 657552
rect 2832 657540 2838 657552
rect 6178 657540 6184 657552
rect 2832 657512 6184 657540
rect 2832 657500 2838 657512
rect 6178 657500 6184 657512
rect 6236 657500 6242 657552
rect 120166 656208 120172 656260
rect 120224 656248 120230 656260
rect 122098 656248 122104 656260
rect 120224 656220 122104 656248
rect 120224 656208 120230 656220
rect 122098 656208 122104 656220
rect 122156 656208 122162 656260
rect 210418 656208 210424 656260
rect 210476 656248 210482 656260
rect 212350 656248 212356 656260
rect 210476 656220 212356 656248
rect 210476 656208 210482 656220
rect 212350 656208 212356 656220
rect 212408 656208 212414 656260
rect 512086 656208 512092 656260
rect 512144 656248 512150 656260
rect 514018 656248 514024 656260
rect 512144 656220 514024 656248
rect 512144 656208 512150 656220
rect 514018 656208 514024 656220
rect 514076 656208 514082 656260
rect 184382 655664 184388 655716
rect 184440 655704 184446 655716
rect 233234 655704 233240 655716
rect 184440 655676 233240 655704
rect 184440 655664 184446 655676
rect 233234 655664 233240 655676
rect 233292 655664 233298 655716
rect 350442 655664 350448 655716
rect 350500 655704 350506 655716
rect 401594 655704 401600 655716
rect 350500 655676 401600 655704
rect 350500 655664 350506 655676
rect 401594 655664 401600 655676
rect 401652 655664 401658 655716
rect 464430 655664 464436 655716
rect 464488 655704 464494 655716
rect 513374 655704 513380 655716
rect 464488 655676 513380 655704
rect 464488 655664 464494 655676
rect 513374 655664 513380 655676
rect 513432 655664 513438 655716
rect 42702 655596 42708 655648
rect 42760 655636 42766 655648
rect 93854 655636 93860 655648
rect 42760 655608 93860 655636
rect 42760 655596 42766 655608
rect 93854 655596 93860 655608
rect 93912 655596 93918 655648
rect 97902 655596 97908 655648
rect 97960 655636 97966 655648
rect 149054 655636 149060 655648
rect 97960 655608 149060 655636
rect 97960 655596 97966 655608
rect 149054 655596 149060 655608
rect 149112 655596 149118 655648
rect 156414 655596 156420 655648
rect 156472 655636 156478 655648
rect 205634 655636 205640 655648
rect 156472 655608 205640 655636
rect 156472 655596 156478 655608
rect 205634 655596 205640 655608
rect 205692 655596 205698 655648
rect 238662 655596 238668 655648
rect 238720 655636 238726 655648
rect 289814 655636 289820 655648
rect 238720 655608 289820 655636
rect 238720 655596 238726 655608
rect 289814 655596 289820 655608
rect 289872 655596 289878 655648
rect 293862 655596 293868 655648
rect 293920 655636 293926 655648
rect 345014 655636 345020 655648
rect 293920 655608 345020 655636
rect 293920 655596 293926 655608
rect 345014 655596 345020 655608
rect 345072 655596 345078 655648
rect 378042 655596 378048 655648
rect 378100 655636 378106 655648
rect 429286 655636 429292 655648
rect 378100 655608 429292 655636
rect 378100 655596 378106 655608
rect 429286 655596 429292 655608
rect 429344 655596 429350 655648
rect 436462 655596 436468 655648
rect 436520 655636 436526 655648
rect 485774 655636 485780 655648
rect 436520 655608 485780 655636
rect 436520 655596 436526 655608
rect 485774 655596 485780 655608
rect 485832 655596 485838 655648
rect 518802 655596 518808 655648
rect 518860 655636 518866 655648
rect 569954 655636 569960 655648
rect 518860 655608 569960 655636
rect 518860 655596 518866 655608
rect 569954 655596 569960 655608
rect 570012 655596 570018 655648
rect 13722 655528 13728 655580
rect 13780 655568 13786 655580
rect 66254 655568 66260 655580
rect 13780 655540 66260 655568
rect 13780 655528 13786 655540
rect 66254 655528 66260 655540
rect 66312 655528 66318 655580
rect 70302 655528 70308 655580
rect 70360 655568 70366 655580
rect 121454 655568 121460 655580
rect 70360 655540 121460 655568
rect 70360 655528 70366 655540
rect 121454 655528 121460 655540
rect 121512 655528 121518 655580
rect 126882 655528 126888 655580
rect 126940 655568 126946 655580
rect 178034 655568 178040 655580
rect 126940 655540 178040 655568
rect 126940 655528 126946 655540
rect 178034 655528 178040 655540
rect 178092 655528 178098 655580
rect 209682 655528 209688 655580
rect 209740 655568 209746 655580
rect 262214 655568 262220 655580
rect 209740 655540 262220 655568
rect 209740 655528 209746 655540
rect 262214 655528 262220 655540
rect 262272 655528 262278 655580
rect 266262 655528 266268 655580
rect 266320 655568 266326 655580
rect 317414 655568 317420 655580
rect 266320 655540 317420 655568
rect 266320 655528 266326 655540
rect 317414 655528 317420 655540
rect 317472 655528 317478 655580
rect 322842 655528 322848 655580
rect 322900 655568 322906 655580
rect 373994 655568 374000 655580
rect 322900 655540 374000 655568
rect 322900 655528 322906 655540
rect 373994 655528 374000 655540
rect 374052 655528 374058 655580
rect 408402 655528 408408 655580
rect 408460 655568 408466 655580
rect 458174 655568 458180 655580
rect 408460 655540 458180 655568
rect 408460 655528 408466 655540
rect 458174 655528 458180 655540
rect 458232 655528 458238 655580
rect 489822 655528 489828 655580
rect 489880 655568 489886 655580
rect 542354 655568 542360 655580
rect 489880 655540 542360 655568
rect 489880 655528 489886 655540
rect 542354 655528 542360 655540
rect 542412 655528 542418 655580
rect 400306 655188 400312 655240
rect 400364 655228 400370 655240
rect 400950 655228 400956 655240
rect 400364 655200 400956 655228
rect 400364 655188 400370 655200
rect 400950 655188 400956 655200
rect 401008 655188 401014 655240
rect 204254 654304 204260 654356
rect 204312 654344 204318 654356
rect 204990 654344 204996 654356
rect 204312 654316 204996 654344
rect 204312 654304 204318 654316
rect 204990 654304 204996 654316
rect 205048 654304 205054 654356
rect 434622 654032 434628 654084
rect 434680 654072 434686 654084
rect 436462 654072 436468 654084
rect 434680 654044 436468 654072
rect 434680 654032 434686 654044
rect 436462 654032 436468 654044
rect 436520 654032 436526 654084
rect 15194 634720 15200 634772
rect 15252 634760 15258 634772
rect 35894 634760 35900 634772
rect 15252 634732 35900 634760
rect 15252 634720 15258 634732
rect 35894 634720 35900 634732
rect 35952 634720 35958 634772
rect 36078 634720 36084 634772
rect 36136 634760 36142 634772
rect 63586 634760 63592 634772
rect 36136 634732 63592 634760
rect 36136 634720 36142 634732
rect 63586 634720 63592 634732
rect 63644 634720 63650 634772
rect 64046 634720 64052 634772
rect 64104 634760 64110 634772
rect 91922 634760 91928 634772
rect 64104 634732 91928 634760
rect 64104 634720 64110 634732
rect 91922 634720 91928 634732
rect 91980 634720 91986 634772
rect 92106 634720 92112 634772
rect 92164 634760 92170 634772
rect 119614 634760 119620 634772
rect 92164 634732 119620 634760
rect 92164 634720 92170 634732
rect 119614 634720 119620 634732
rect 119672 634720 119678 634772
rect 122098 634720 122104 634772
rect 122156 634760 122162 634772
rect 147950 634760 147956 634772
rect 122156 634732 147956 634760
rect 122156 634720 122162 634732
rect 147950 634720 147956 634732
rect 148008 634720 148014 634772
rect 148042 634720 148048 634772
rect 148100 634760 148106 634772
rect 175918 634760 175924 634772
rect 148100 634732 175924 634760
rect 148100 634720 148106 634732
rect 175918 634720 175924 634732
rect 175976 634720 175982 634772
rect 176102 634720 176108 634772
rect 176160 634760 176166 634772
rect 203610 634760 203616 634772
rect 176160 634732 203616 634760
rect 176160 634720 176166 634732
rect 203610 634720 203616 634732
rect 203668 634720 203674 634772
rect 204990 634720 204996 634772
rect 205048 634760 205054 634772
rect 231946 634760 231952 634772
rect 205048 634732 231952 634760
rect 205048 634720 205054 634732
rect 231946 634720 231952 634732
rect 232004 634720 232010 634772
rect 232038 634720 232044 634772
rect 232096 634760 232102 634772
rect 259914 634760 259920 634772
rect 232096 634732 259920 634760
rect 232096 634720 232102 634732
rect 259914 634720 259920 634732
rect 259972 634720 259978 634772
rect 260098 634720 260104 634772
rect 260156 634760 260162 634772
rect 287606 634760 287612 634772
rect 260156 634732 287612 634760
rect 260156 634720 260162 634732
rect 287606 634720 287612 634732
rect 287664 634720 287670 634772
rect 288066 634720 288072 634772
rect 288124 634760 288130 634772
rect 315942 634760 315948 634772
rect 288124 634732 315948 634760
rect 288124 634720 288130 634732
rect 315942 634720 315948 634732
rect 316000 634720 316006 634772
rect 316678 634720 316684 634772
rect 316736 634760 316742 634772
rect 343910 634760 343916 634772
rect 316736 634732 343916 634760
rect 316736 634720 316742 634732
rect 343910 634720 343916 634732
rect 343968 634720 343974 634772
rect 344094 634720 344100 634772
rect 344152 634760 344158 634772
rect 371602 634760 371608 634772
rect 344152 634732 371608 634760
rect 344152 634720 344158 634732
rect 371602 634720 371608 634732
rect 371660 634720 371666 634772
rect 372062 634720 372068 634772
rect 372120 634760 372126 634772
rect 399938 634760 399944 634772
rect 372120 634732 399944 634760
rect 372120 634720 372126 634732
rect 399938 634720 399944 634732
rect 399996 634720 400002 634772
rect 400950 634720 400956 634772
rect 401008 634760 401014 634772
rect 427906 634760 427912 634772
rect 401008 634732 427912 634760
rect 401008 634720 401014 634732
rect 427906 634720 427912 634732
rect 427964 634720 427970 634772
rect 428090 634720 428096 634772
rect 428148 634760 428154 634772
rect 455598 634760 455604 634772
rect 428148 634732 455604 634760
rect 428148 634720 428154 634732
rect 455598 634720 455604 634732
rect 455656 634720 455662 634772
rect 456058 634720 456064 634772
rect 456116 634760 456122 634772
rect 483934 634760 483940 634772
rect 456116 634732 483940 634760
rect 456116 634720 456122 634732
rect 483934 634720 483940 634732
rect 483992 634720 483998 634772
rect 484026 634720 484032 634772
rect 484084 634760 484090 634772
rect 511902 634760 511908 634772
rect 484084 634732 511908 634760
rect 484084 634720 484090 634732
rect 511902 634720 511908 634732
rect 511960 634720 511966 634772
rect 514018 634720 514024 634772
rect 514076 634760 514082 634772
rect 539594 634760 539600 634772
rect 514076 634732 539600 634760
rect 514076 634720 514082 634732
rect 539594 634720 539600 634732
rect 539652 634720 539658 634772
rect 540054 634720 540060 634772
rect 540112 634760 540118 634772
rect 567930 634760 567936 634772
rect 540112 634732 567936 634760
rect 540112 634720 540118 634732
rect 567930 634720 567936 634732
rect 567988 634720 567994 634772
rect 16574 634652 16580 634704
rect 16632 634692 16638 634704
rect 36630 634692 36636 634704
rect 16632 634664 36636 634692
rect 16632 634652 16638 634664
rect 36630 634652 36636 634664
rect 36688 634652 36694 634704
rect 44910 634652 44916 634704
rect 44968 634692 44974 634704
rect 71130 634692 71136 634704
rect 44968 634664 71136 634692
rect 44968 634652 44974 634664
rect 71130 634652 71136 634664
rect 71188 634652 71194 634704
rect 82262 634652 82268 634704
rect 82320 634692 82326 634704
rect 93118 634692 93124 634704
rect 82320 634664 93124 634692
rect 82320 634652 82326 634664
rect 93118 634652 93124 634664
rect 93176 634652 93182 634704
rect 110322 634652 110328 634704
rect 110380 634692 110386 634704
rect 124858 634692 124864 634704
rect 110380 634664 124864 634692
rect 110380 634652 110386 634664
rect 124858 634652 124864 634664
rect 124916 634652 124922 634704
rect 128630 634652 128636 634704
rect 128688 634692 128694 634704
rect 149698 634692 149704 634704
rect 128688 634664 149704 634692
rect 128688 634652 128694 634664
rect 149698 634652 149704 634664
rect 149756 634652 149762 634704
rect 156598 634652 156604 634704
rect 156656 634692 156662 634704
rect 182818 634692 182824 634704
rect 156656 634664 182824 634692
rect 156656 634652 156662 634664
rect 182818 634652 182824 634664
rect 182876 634652 182882 634704
rect 194502 634652 194508 634704
rect 194560 634692 194566 634704
rect 210418 634692 210424 634704
rect 194560 634664 210424 634692
rect 194560 634652 194566 634664
rect 210418 634652 210424 634664
rect 210476 634652 210482 634704
rect 212626 634652 212632 634704
rect 212684 634692 212690 634704
rect 232498 634692 232504 634704
rect 212684 634664 232504 634692
rect 212684 634652 212690 634664
rect 232498 634652 232504 634664
rect 232556 634652 232562 634704
rect 240594 634652 240600 634704
rect 240652 634692 240658 634704
rect 266998 634692 267004 634704
rect 240652 634664 267004 634692
rect 240652 634652 240658 634664
rect 266998 634652 267004 634664
rect 267056 634652 267062 634704
rect 278590 634652 278596 634704
rect 278648 634692 278654 634704
rect 289078 634692 289084 634704
rect 278648 634664 289084 634692
rect 278648 634652 278654 634664
rect 289078 634652 289084 634664
rect 289136 634652 289142 634704
rect 306282 634652 306288 634704
rect 306340 634692 306346 634704
rect 318058 634692 318064 634704
rect 306340 634664 318064 634692
rect 306340 634652 306346 634664
rect 318058 634652 318064 634664
rect 318116 634652 318122 634704
rect 324590 634652 324596 634704
rect 324648 634692 324654 634704
rect 347038 634692 347044 634704
rect 324648 634664 347044 634692
rect 324648 634652 324654 634664
rect 347038 634652 347044 634664
rect 347096 634652 347102 634704
rect 362586 634652 362592 634704
rect 362644 634692 362650 634704
rect 373258 634692 373264 634704
rect 362644 634664 373264 634692
rect 362644 634652 362650 634664
rect 373258 634652 373264 634664
rect 373316 634652 373322 634704
rect 390278 634652 390284 634704
rect 390336 634692 390342 634704
rect 400858 634692 400864 634704
rect 390336 634664 400864 634692
rect 390336 634652 390342 634664
rect 400858 634652 400864 634664
rect 400916 634652 400922 634704
rect 408586 634652 408592 634704
rect 408644 634692 408650 634704
rect 428458 634692 428464 634704
rect 408644 634664 428464 634692
rect 408644 634652 408650 634664
rect 428458 634652 428464 634664
rect 428516 634652 428522 634704
rect 436922 634652 436928 634704
rect 436980 634692 436986 634704
rect 462958 634692 462964 634704
rect 436980 634664 462964 634692
rect 436980 634652 436986 634664
rect 462958 634652 462964 634664
rect 463016 634652 463022 634704
rect 474274 634652 474280 634704
rect 474332 634692 474338 634704
rect 485038 634692 485044 634704
rect 474332 634664 485044 634692
rect 474332 634652 474338 634664
rect 485038 634652 485044 634664
rect 485096 634652 485102 634704
rect 502242 634652 502248 634704
rect 502300 634692 502306 634704
rect 512638 634692 512644 634704
rect 502300 634664 512644 634692
rect 502300 634652 502306 634664
rect 512638 634652 512644 634664
rect 512696 634652 512702 634704
rect 520918 634652 520924 634704
rect 520976 634692 520982 634704
rect 541618 634692 541624 634704
rect 520976 634664 541624 634692
rect 520976 634652 520982 634664
rect 541618 634652 541624 634664
rect 541676 634652 541682 634704
rect 26234 634584 26240 634636
rect 26292 634624 26298 634636
rect 43530 634624 43536 634636
rect 26292 634596 43536 634624
rect 26292 634584 26298 634596
rect 43530 634584 43536 634596
rect 43588 634584 43594 634636
rect 54570 634584 54576 634636
rect 54628 634624 54634 634636
rect 66898 634624 66904 634636
rect 54628 634596 66904 634624
rect 54628 634584 54634 634596
rect 66898 634584 66904 634596
rect 66956 634584 66962 634636
rect 138290 634584 138296 634636
rect 138348 634624 138354 634636
rect 151078 634624 151084 634636
rect 138348 634596 151084 634624
rect 138348 634584 138354 634596
rect 151078 634584 151084 634596
rect 151136 634584 151142 634636
rect 166258 634584 166264 634636
rect 166316 634624 166322 634636
rect 177298 634624 177304 634636
rect 166316 634596 177304 634624
rect 166316 634584 166322 634596
rect 177298 634584 177304 634596
rect 177356 634584 177362 634636
rect 222286 634584 222292 634636
rect 222344 634624 222350 634636
rect 233970 634624 233976 634636
rect 222344 634596 233976 634624
rect 222344 634584 222350 634596
rect 233970 634584 233976 634596
rect 234028 634584 234034 634636
rect 250254 634584 250260 634636
rect 250312 634624 250318 634636
rect 261478 634624 261484 634636
rect 250312 634596 261484 634624
rect 250312 634584 250318 634596
rect 261478 634584 261484 634596
rect 261536 634584 261542 634636
rect 334250 634584 334256 634636
rect 334308 634624 334314 634636
rect 348418 634624 348424 634636
rect 334308 634596 348424 634624
rect 334308 634584 334314 634596
rect 348418 634584 348424 634596
rect 348476 634584 348482 634636
rect 418246 634584 418252 634636
rect 418304 634624 418310 634636
rect 429838 634624 429844 634636
rect 418304 634596 429844 634624
rect 418304 634584 418310 634596
rect 429838 634584 429844 634596
rect 429896 634584 429902 634636
rect 446582 634584 446588 634636
rect 446640 634624 446646 634636
rect 457438 634624 457444 634636
rect 446640 634596 457444 634624
rect 446640 634584 446646 634596
rect 457438 634584 457444 634596
rect 457496 634584 457502 634636
rect 530578 634584 530584 634636
rect 530636 634624 530642 634636
rect 544378 634624 544384 634636
rect 530636 634596 544384 634624
rect 530636 634584 530642 634596
rect 544378 634584 544384 634596
rect 544436 634584 544442 634636
rect 558270 634040 558276 634092
rect 558328 634080 558334 634092
rect 567470 634080 567476 634092
rect 558328 634052 567476 634080
rect 558328 634040 558334 634052
rect 567470 634040 567476 634052
rect 567528 634040 567534 634092
rect 548334 632680 548340 632732
rect 548392 632720 548398 632732
rect 568022 632720 568028 632732
rect 548392 632692 568028 632720
rect 548392 632680 548398 632692
rect 568022 632680 568028 632692
rect 568080 632680 568086 632732
rect 212350 632272 212356 632324
rect 212408 632312 212414 632324
rect 232682 632312 232688 632324
rect 212408 632284 232688 632312
rect 212408 632272 212414 632284
rect 232682 632272 232688 632284
rect 232740 632272 232746 632324
rect 296346 632272 296352 632324
rect 296404 632312 296410 632324
rect 316770 632312 316776 632324
rect 296404 632284 316776 632312
rect 296404 632272 296410 632284
rect 316770 632272 316776 632284
rect 316828 632272 316834 632324
rect 408034 632272 408040 632324
rect 408092 632312 408098 632324
rect 428642 632312 428648 632324
rect 408092 632284 428648 632312
rect 408092 632272 408098 632284
rect 428642 632272 428648 632284
rect 428700 632272 428706 632324
rect 492030 632272 492036 632324
rect 492088 632312 492094 632324
rect 512730 632312 512736 632324
rect 492088 632284 512736 632312
rect 492088 632272 492094 632284
rect 512730 632272 512736 632284
rect 512788 632272 512794 632324
rect 148318 632204 148324 632256
rect 148376 632244 148382 632256
rect 165706 632244 165712 632256
rect 148376 632216 165712 632244
rect 148376 632204 148382 632216
rect 165706 632204 165712 632216
rect 165764 632204 165770 632256
rect 175458 632204 175464 632256
rect 175516 632244 175522 632256
rect 193674 632244 193680 632256
rect 175516 632216 193680 632244
rect 175516 632204 175522 632216
rect 193674 632204 193680 632216
rect 193732 632204 193738 632256
rect 203518 632204 203524 632256
rect 203576 632244 203582 632256
rect 221366 632244 221372 632256
rect 203576 632216 221372 632244
rect 203576 632204 203582 632216
rect 221366 632204 221372 632216
rect 221424 632204 221430 632256
rect 260098 632204 260104 632256
rect 260156 632244 260162 632256
rect 277670 632244 277676 632256
rect 260156 632216 277676 632244
rect 260156 632204 260162 632216
rect 277670 632204 277676 632216
rect 277728 632204 277734 632256
rect 287514 632204 287520 632256
rect 287572 632244 287578 632256
rect 305362 632244 305368 632256
rect 287572 632216 305368 632244
rect 287572 632204 287578 632216
rect 305362 632204 305368 632216
rect 305420 632204 305426 632256
rect 345658 632204 345664 632256
rect 345716 632244 345722 632256
rect 361666 632244 361672 632256
rect 345716 632216 361672 632244
rect 345716 632204 345722 632216
rect 361666 632204 361672 632216
rect 361724 632204 361730 632256
rect 371510 632204 371516 632256
rect 371568 632244 371574 632256
rect 389358 632244 389364 632256
rect 371568 632216 389364 632244
rect 371568 632204 371574 632216
rect 389358 632204 389364 632216
rect 389416 632204 389422 632256
rect 399478 632204 399484 632256
rect 399536 632244 399542 632256
rect 417694 632244 417700 632256
rect 399536 632216 417700 632244
rect 399536 632204 399542 632216
rect 417694 632204 417700 632216
rect 417752 632204 417758 632256
rect 456150 632204 456156 632256
rect 456208 632244 456214 632256
rect 473354 632244 473360 632256
rect 456208 632216 473360 632244
rect 456208 632204 456214 632216
rect 473354 632204 473360 632216
rect 473412 632204 473418 632256
rect 483474 632204 483480 632256
rect 483532 632244 483538 632256
rect 501690 632244 501696 632256
rect 483532 632216 501696 632244
rect 483532 632204 483538 632216
rect 501690 632204 501696 632216
rect 501748 632204 501754 632256
rect 36722 632136 36728 632188
rect 36780 632176 36786 632188
rect 53650 632176 53656 632188
rect 36780 632148 53656 632176
rect 36780 632136 36786 632148
rect 53650 632136 53656 632148
rect 53708 632136 53714 632188
rect 64322 632136 64328 632188
rect 64380 632176 64386 632188
rect 81434 632176 81440 632188
rect 64380 632148 81440 632176
rect 64380 632136 64386 632148
rect 81434 632136 81440 632148
rect 81492 632136 81498 632188
rect 91462 632136 91468 632188
rect 91520 632176 91526 632188
rect 109678 632176 109684 632188
rect 91520 632148 109684 632176
rect 91520 632136 91526 632148
rect 109678 632136 109684 632148
rect 109736 632136 109742 632188
rect 119430 632136 119436 632188
rect 119488 632176 119494 632188
rect 137646 632176 137652 632188
rect 119488 632148 137652 632176
rect 119488 632136 119494 632148
rect 137646 632136 137652 632148
rect 137704 632136 137710 632188
rect 156322 632136 156328 632188
rect 156380 632176 156386 632188
rect 178678 632176 178684 632188
rect 156380 632148 178684 632176
rect 156380 632136 156386 632148
rect 178678 632136 178684 632148
rect 178736 632136 178742 632188
rect 232498 632136 232504 632188
rect 232556 632176 232562 632188
rect 249702 632176 249708 632188
rect 232556 632148 249708 632176
rect 232556 632136 232562 632148
rect 249702 632136 249708 632148
rect 249760 632136 249766 632188
rect 268010 632136 268016 632188
rect 268068 632176 268074 632188
rect 287698 632176 287704 632188
rect 268068 632148 287704 632176
rect 268068 632136 268074 632148
rect 287698 632136 287704 632148
rect 287756 632136 287762 632188
rect 315482 632136 315488 632188
rect 315540 632176 315546 632188
rect 333698 632176 333704 632188
rect 315540 632148 333704 632176
rect 315540 632136 315546 632148
rect 333698 632136 333704 632148
rect 333756 632136 333762 632188
rect 352006 632136 352012 632188
rect 352064 632176 352070 632188
rect 374638 632176 374644 632188
rect 352064 632148 374644 632176
rect 352064 632136 352070 632148
rect 374638 632136 374644 632148
rect 374696 632136 374702 632188
rect 428458 632136 428464 632188
rect 428516 632176 428522 632188
rect 445662 632176 445668 632188
rect 428516 632148 445668 632176
rect 428516 632136 428522 632148
rect 445662 632136 445668 632148
rect 445720 632136 445726 632188
rect 464338 632136 464344 632188
rect 464396 632176 464402 632188
rect 483658 632176 483664 632188
rect 464396 632148 483664 632176
rect 464396 632136 464402 632148
rect 483658 632136 483664 632148
rect 483716 632136 483722 632188
rect 511442 632136 511448 632188
rect 511500 632176 511506 632188
rect 529658 632176 529664 632188
rect 511500 632148 529664 632176
rect 511500 632136 511506 632148
rect 529658 632136 529664 632148
rect 529716 632136 529722 632188
rect 541618 632136 541624 632188
rect 541676 632176 541682 632188
rect 557534 632176 557540 632188
rect 541676 632148 557540 632176
rect 541676 632136 541682 632148
rect 557534 632136 557540 632148
rect 557592 632136 557598 632188
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 14458 632108 14464 632120
rect 3476 632080 14464 632108
rect 3476 632068 3482 632080
rect 14458 632068 14464 632080
rect 14516 632068 14522 632120
rect 16114 632068 16120 632120
rect 16172 632108 16178 632120
rect 25682 632108 25688 632120
rect 16172 632080 25688 632108
rect 16172 632068 16178 632080
rect 25682 632068 25688 632080
rect 25740 632068 25746 632120
rect 36630 632068 36636 632120
rect 36688 632108 36694 632120
rect 63310 632108 63316 632120
rect 36688 632080 63316 632108
rect 36688 632068 36694 632080
rect 63310 632068 63316 632080
rect 63368 632068 63374 632120
rect 66898 632068 66904 632120
rect 66956 632108 66962 632120
rect 91094 632108 91100 632120
rect 66956 632080 91100 632108
rect 66956 632068 66962 632080
rect 91094 632068 91100 632080
rect 91152 632068 91158 632120
rect 93118 632068 93124 632120
rect 93176 632108 93182 632120
rect 119338 632108 119344 632120
rect 93176 632080 119344 632108
rect 93176 632068 93182 632080
rect 119338 632068 119344 632080
rect 119396 632068 119402 632120
rect 124858 632068 124864 632120
rect 124916 632108 124922 632120
rect 147306 632108 147312 632120
rect 124916 632080 147312 632108
rect 124916 632068 124922 632080
rect 147306 632068 147312 632080
rect 147364 632068 147370 632120
rect 148410 632068 148416 632120
rect 148468 632108 148474 632120
rect 175366 632108 175372 632120
rect 148468 632080 175372 632108
rect 148468 632068 148474 632080
rect 175366 632068 175372 632080
rect 175424 632068 175430 632120
rect 177298 632068 177304 632120
rect 177356 632108 177362 632120
rect 203334 632108 203340 632120
rect 177356 632080 203340 632108
rect 177356 632068 177362 632080
rect 203334 632068 203340 632080
rect 203392 632068 203398 632120
rect 204990 632068 204996 632120
rect 205048 632108 205054 632120
rect 231026 632108 231032 632120
rect 205048 632080 231032 632108
rect 205048 632068 205054 632080
rect 231026 632068 231032 632080
rect 231084 632068 231090 632120
rect 232590 632068 232596 632120
rect 232648 632108 232654 632120
rect 259362 632108 259368 632120
rect 232648 632080 259368 632108
rect 232648 632068 232654 632080
rect 259362 632068 259368 632080
rect 259420 632068 259426 632120
rect 260190 632068 260196 632120
rect 260248 632108 260254 632120
rect 287330 632108 287336 632120
rect 260248 632080 287336 632108
rect 260248 632068 260254 632080
rect 287330 632068 287336 632080
rect 287388 632068 287394 632120
rect 289078 632068 289084 632120
rect 289136 632108 289142 632120
rect 315022 632108 315028 632120
rect 289136 632080 315028 632108
rect 289136 632068 289142 632080
rect 315022 632068 315028 632080
rect 315080 632068 315086 632120
rect 316678 632068 316684 632120
rect 316736 632108 316742 632120
rect 343358 632108 343364 632120
rect 316736 632080 343364 632108
rect 316736 632068 316742 632080
rect 343358 632068 343364 632080
rect 343416 632068 343422 632120
rect 344278 632068 344284 632120
rect 344336 632108 344342 632120
rect 371326 632108 371332 632120
rect 344336 632080 371332 632108
rect 344336 632068 344342 632080
rect 371326 632068 371332 632080
rect 371384 632068 371390 632120
rect 373258 632068 373264 632120
rect 373316 632108 373322 632120
rect 399018 632108 399024 632120
rect 373316 632080 399024 632108
rect 373316 632068 373322 632080
rect 399018 632068 399024 632080
rect 399076 632068 399082 632120
rect 400858 632068 400864 632120
rect 400916 632108 400922 632120
rect 427354 632108 427360 632120
rect 400916 632080 427360 632108
rect 400916 632068 400922 632080
rect 427354 632068 427360 632080
rect 427412 632068 427418 632120
rect 428550 632068 428556 632120
rect 428608 632108 428614 632120
rect 455322 632108 455328 632120
rect 428608 632080 455328 632108
rect 428608 632068 428614 632080
rect 455322 632068 455328 632080
rect 455380 632068 455386 632120
rect 456058 632068 456064 632120
rect 456116 632108 456122 632120
rect 483014 632108 483020 632120
rect 456116 632080 483020 632108
rect 456116 632068 456122 632080
rect 483014 632068 483020 632080
rect 483072 632068 483078 632120
rect 485038 632068 485044 632120
rect 485096 632108 485102 632120
rect 511350 632108 511356 632120
rect 485096 632080 511356 632108
rect 485096 632068 485102 632080
rect 511350 632068 511356 632080
rect 511408 632068 511414 632120
rect 512638 632068 512644 632120
rect 512696 632108 512702 632120
rect 539318 632108 539324 632120
rect 512696 632080 539324 632108
rect 512696 632068 512702 632080
rect 539318 632068 539324 632080
rect 539376 632068 539382 632120
rect 540238 632068 540244 632120
rect 540296 632108 540302 632120
rect 567194 632108 567200 632120
rect 540296 632080 567200 632108
rect 540296 632068 540302 632080
rect 567194 632068 567200 632080
rect 567252 632068 567258 632120
rect 15838 629280 15844 629332
rect 15896 629320 15902 629332
rect 16114 629320 16120 629332
rect 15896 629292 16120 629320
rect 15896 629280 15902 629292
rect 16114 629280 16120 629292
rect 16172 629280 16178 629332
rect 42886 627240 42892 627292
rect 42944 627280 42950 627292
rect 43622 627280 43628 627292
rect 42944 627252 43628 627280
rect 42944 627240 42950 627252
rect 43622 627240 43628 627252
rect 43680 627240 43686 627292
rect 63586 612756 63592 612808
rect 63644 612796 63650 612808
rect 64322 612796 64328 612808
rect 63644 612768 64328 612796
rect 63644 612756 63650 612768
rect 64322 612756 64328 612768
rect 64380 612756 64386 612808
rect 455690 612756 455696 612808
rect 455748 612796 455754 612808
rect 456150 612796 456156 612808
rect 455748 612768 456156 612796
rect 455748 612756 455754 612768
rect 456150 612756 456156 612768
rect 456208 612756 456214 612808
rect 428642 612008 428648 612060
rect 428700 612048 428706 612060
rect 435726 612048 435732 612060
rect 428700 612020 435732 612048
rect 428700 612008 428706 612020
rect 435726 612008 435732 612020
rect 435784 612008 435790 612060
rect 232682 611940 232688 611992
rect 232740 611980 232746 611992
rect 239766 611980 239772 611992
rect 232740 611952 239772 611980
rect 232740 611940 232746 611952
rect 239766 611940 239772 611952
rect 239824 611940 239830 611992
rect 287698 611872 287704 611924
rect 287756 611912 287762 611924
rect 295702 611912 295708 611924
rect 287756 611884 295708 611912
rect 287756 611872 287762 611884
rect 295702 611872 295708 611884
rect 295760 611872 295766 611924
rect 316770 611872 316776 611924
rect 316828 611912 316834 611924
rect 323670 611912 323676 611924
rect 316828 611884 323676 611912
rect 316828 611872 316834 611884
rect 323670 611872 323676 611884
rect 323728 611872 323734 611924
rect 483658 611736 483664 611788
rect 483716 611776 483722 611788
rect 491662 611776 491668 611788
rect 483716 611748 491668 611776
rect 483716 611736 483722 611748
rect 491662 611736 491668 611748
rect 491720 611736 491726 611788
rect 512730 611736 512736 611788
rect 512788 611776 512794 611788
rect 519630 611776 519636 611788
rect 512788 611748 519636 611776
rect 512788 611736 512794 611748
rect 519630 611736 519636 611748
rect 519688 611736 519694 611788
rect 13538 611260 13544 611312
rect 13596 611300 13602 611312
rect 66254 611300 66260 611312
rect 13596 611272 66260 611300
rect 13596 611260 13602 611272
rect 66254 611260 66260 611272
rect 66312 611260 66318 611312
rect 70302 611260 70308 611312
rect 70360 611300 70366 611312
rect 121454 611300 121460 611312
rect 70360 611272 121460 611300
rect 70360 611260 70366 611272
rect 121454 611260 121460 611272
rect 121512 611260 121518 611312
rect 126882 611260 126888 611312
rect 126940 611300 126946 611312
rect 178034 611300 178040 611312
rect 126940 611272 178040 611300
rect 126940 611260 126946 611272
rect 178034 611260 178040 611272
rect 178092 611260 178098 611312
rect 209682 611260 209688 611312
rect 209740 611300 209746 611312
rect 262214 611300 262220 611312
rect 209740 611272 262220 611300
rect 209740 611260 209746 611272
rect 262214 611260 262220 611272
rect 262272 611260 262278 611312
rect 266262 611260 266268 611312
rect 266320 611300 266326 611312
rect 317414 611300 317420 611312
rect 266320 611272 317420 611300
rect 266320 611260 266326 611272
rect 317414 611260 317420 611272
rect 317472 611260 317478 611312
rect 322842 611260 322848 611312
rect 322900 611300 322906 611312
rect 373994 611300 374000 611312
rect 322900 611272 374000 611300
rect 322900 611260 322906 611272
rect 373994 611260 374000 611272
rect 374052 611260 374058 611312
rect 405642 611260 405648 611312
rect 405700 611300 405706 611312
rect 458174 611300 458180 611312
rect 405700 611272 458180 611300
rect 405700 611260 405706 611272
rect 458174 611260 458180 611272
rect 458232 611260 458238 611312
rect 489822 611260 489828 611312
rect 489880 611300 489886 611312
rect 489880 611272 539364 611300
rect 489880 611260 489886 611272
rect 42702 611192 42708 611244
rect 42760 611232 42766 611244
rect 93854 611232 93860 611244
rect 42760 611204 93860 611232
rect 42760 611192 42766 611204
rect 93854 611192 93860 611204
rect 93912 611192 93918 611244
rect 97902 611192 97908 611244
rect 97960 611232 97966 611244
rect 149054 611232 149060 611244
rect 97960 611204 149060 611232
rect 97960 611192 97966 611204
rect 149054 611192 149060 611204
rect 149112 611192 149118 611244
rect 154482 611192 154488 611244
rect 154540 611232 154546 611244
rect 205634 611232 205640 611244
rect 154540 611204 205640 611232
rect 154540 611192 154546 611204
rect 205634 611192 205640 611204
rect 205692 611192 205698 611244
rect 238662 611192 238668 611244
rect 238720 611232 238726 611244
rect 289814 611232 289820 611244
rect 238720 611204 289820 611232
rect 238720 611192 238726 611204
rect 289814 611192 289820 611204
rect 289872 611192 289878 611244
rect 293862 611192 293868 611244
rect 293920 611232 293926 611244
rect 345014 611232 345020 611244
rect 293920 611204 345020 611232
rect 293920 611192 293926 611204
rect 345014 611192 345020 611204
rect 345072 611192 345078 611244
rect 378042 611192 378048 611244
rect 378100 611232 378106 611244
rect 429286 611232 429292 611244
rect 378100 611204 429292 611232
rect 378100 611192 378106 611204
rect 429286 611192 429292 611204
rect 429344 611192 429350 611244
rect 434622 611192 434628 611244
rect 434680 611232 434686 611244
rect 485774 611232 485780 611244
rect 434680 611204 485780 611232
rect 434680 611192 434686 611204
rect 485774 611192 485780 611204
rect 485832 611192 485838 611244
rect 518802 611192 518808 611244
rect 518860 611232 518866 611244
rect 518860 611204 528554 611232
rect 518860 611192 518866 611204
rect 182082 611124 182088 611176
rect 182140 611164 182146 611176
rect 233234 611164 233240 611176
rect 182140 611136 233240 611164
rect 182140 611124 182146 611136
rect 233234 611124 233240 611136
rect 233292 611124 233298 611176
rect 350442 611124 350448 611176
rect 350500 611164 350506 611176
rect 401594 611164 401600 611176
rect 350500 611136 401600 611164
rect 350500 611124 350506 611136
rect 401594 611124 401600 611136
rect 401652 611124 401658 611176
rect 462222 611124 462228 611176
rect 462280 611164 462286 611176
rect 513374 611164 513380 611176
rect 462280 611136 513380 611164
rect 462280 611124 462286 611136
rect 513374 611124 513380 611136
rect 513432 611124 513438 611176
rect 528526 611096 528554 611204
rect 539336 611164 539364 611272
rect 539502 611260 539508 611312
rect 539560 611300 539566 611312
rect 541618 611300 541624 611312
rect 539560 611272 541624 611300
rect 539560 611260 539566 611272
rect 541618 611260 541624 611272
rect 541676 611260 541682 611312
rect 569954 611232 569960 611244
rect 547846 611204 569960 611232
rect 542354 611164 542360 611176
rect 539336 611136 542360 611164
rect 542354 611124 542360 611136
rect 542412 611124 542418 611176
rect 547846 611096 547874 611204
rect 569954 611192 569960 611204
rect 570012 611192 570018 611244
rect 528526 611068 547874 611096
rect 15838 610648 15844 610700
rect 15896 610688 15902 610700
rect 16574 610688 16580 610700
rect 15896 610660 16580 610688
rect 15896 610648 15902 610660
rect 16574 610648 16580 610660
rect 16632 610648 16638 610700
rect 35250 610648 35256 610700
rect 35308 610688 35314 610700
rect 36722 610688 36728 610700
rect 35308 610660 36728 610688
rect 35308 610648 35314 610660
rect 36722 610648 36728 610660
rect 36780 610648 36786 610700
rect 547874 610648 547880 610700
rect 547932 610688 547938 610700
rect 548150 610688 548156 610700
rect 547932 610660 548156 610688
rect 547932 610648 547938 610660
rect 548150 610648 548156 610660
rect 548208 610648 548214 610700
rect 71866 608540 71872 608592
rect 71924 608580 71930 608592
rect 100018 608580 100024 608592
rect 71924 608552 100024 608580
rect 71924 608540 71930 608552
rect 100018 608540 100024 608552
rect 100076 608540 100082 608592
rect 127986 608580 127992 608592
rect 103486 608552 127992 608580
rect 25682 608472 25688 608524
rect 25740 608512 25746 608524
rect 36630 608512 36636 608524
rect 25740 608484 36636 608512
rect 25740 608472 25746 608484
rect 36630 608472 36636 608484
rect 36688 608472 36694 608524
rect 42886 608472 42892 608524
rect 42944 608512 42950 608524
rect 42944 608484 45554 608512
rect 42944 608472 42950 608484
rect 15286 608404 15292 608456
rect 15344 608444 15350 608456
rect 43990 608444 43996 608456
rect 15344 608416 43996 608444
rect 15344 608404 15350 608416
rect 43990 608404 43996 608416
rect 44048 608404 44054 608456
rect 45526 608444 45554 608484
rect 53650 608472 53656 608524
rect 53708 608512 53714 608524
rect 66898 608512 66904 608524
rect 53708 608484 66904 608512
rect 53708 608472 53714 608484
rect 66898 608472 66904 608484
rect 66956 608472 66962 608524
rect 81986 608472 81992 608524
rect 82044 608512 82050 608524
rect 93118 608512 93124 608524
rect 82044 608484 93124 608512
rect 82044 608472 82050 608484
rect 93118 608472 93124 608484
rect 93176 608472 93182 608524
rect 99466 608472 99472 608524
rect 99524 608512 99530 608524
rect 103486 608512 103514 608552
rect 127986 608540 127992 608552
rect 128044 608540 128050 608592
rect 165982 608540 165988 608592
rect 166040 608580 166046 608592
rect 177298 608580 177304 608592
rect 166040 608552 177304 608580
rect 166040 608540 166046 608552
rect 177298 608540 177304 608552
rect 177356 608540 177362 608592
rect 178678 608540 178684 608592
rect 178736 608580 178742 608592
rect 184014 608580 184020 608592
rect 178736 608552 184020 608580
rect 178736 608540 178742 608552
rect 184014 608540 184020 608552
rect 184072 608540 184078 608592
rect 211706 608580 211712 608592
rect 190426 608552 211712 608580
rect 99524 608484 103514 608512
rect 99524 608472 99530 608484
rect 109678 608472 109684 608524
rect 109736 608512 109742 608524
rect 124858 608512 124864 608524
rect 109736 608484 124864 608512
rect 109736 608472 109742 608484
rect 124858 608472 124864 608484
rect 124916 608472 124922 608524
rect 137646 608472 137652 608524
rect 137704 608512 137710 608524
rect 148410 608512 148416 608524
rect 137704 608484 148416 608512
rect 137704 608472 137710 608484
rect 148410 608472 148416 608484
rect 148468 608472 148474 608524
rect 183646 608472 183652 608524
rect 183704 608512 183710 608524
rect 190426 608512 190454 608552
rect 211706 608540 211712 608552
rect 211764 608540 211770 608592
rect 277670 608540 277676 608592
rect 277728 608580 277734 608592
rect 289078 608580 289084 608592
rect 277728 608552 289084 608580
rect 277728 608540 277734 608552
rect 289078 608540 289084 608552
rect 289136 608540 289142 608592
rect 306006 608540 306012 608592
rect 306064 608580 306070 608592
rect 316678 608580 316684 608592
rect 306064 608552 316684 608580
rect 306064 608540 306070 608552
rect 316678 608540 316684 608552
rect 316736 608540 316742 608592
rect 343358 608540 343364 608592
rect 343416 608580 343422 608592
rect 345658 608580 345664 608592
rect 343416 608552 345664 608580
rect 343416 608540 343422 608552
rect 345658 608540 345664 608552
rect 345716 608540 345722 608592
rect 361666 608540 361672 608592
rect 361724 608580 361730 608592
rect 373258 608580 373264 608592
rect 361724 608552 373264 608580
rect 361724 608540 361730 608552
rect 373258 608540 373264 608552
rect 373316 608540 373322 608592
rect 379606 608540 379612 608592
rect 379664 608580 379670 608592
rect 408034 608580 408040 608592
rect 379664 608552 408040 608580
rect 379664 608540 379670 608552
rect 408034 608540 408040 608552
rect 408092 608540 408098 608592
rect 473998 608540 474004 608592
rect 474056 608580 474062 608592
rect 485038 608580 485044 608592
rect 474056 608552 485044 608580
rect 474056 608540 474062 608552
rect 485038 608540 485044 608552
rect 485096 608540 485102 608592
rect 501690 608540 501696 608592
rect 501748 608580 501754 608592
rect 512638 608580 512644 608592
rect 501748 608552 512644 608580
rect 501748 608540 501754 608552
rect 512638 608540 512644 608552
rect 512696 608540 512702 608592
rect 548150 608540 548156 608592
rect 548208 608580 548214 608592
rect 557534 608580 557540 608592
rect 548208 608552 557540 608580
rect 548208 608540 548214 608552
rect 557534 608540 557540 608552
rect 557592 608540 557598 608592
rect 183704 608484 190454 608512
rect 183704 608472 183710 608484
rect 193674 608472 193680 608524
rect 193732 608512 193738 608524
rect 204990 608512 204996 608524
rect 193732 608484 204996 608512
rect 193732 608472 193738 608484
rect 204990 608472 204996 608484
rect 205048 608472 205054 608524
rect 222010 608472 222016 608524
rect 222068 608512 222074 608524
rect 232590 608512 232596 608524
rect 222068 608484 232596 608512
rect 222068 608472 222074 608484
rect 232590 608472 232596 608484
rect 232648 608472 232654 608524
rect 249702 608472 249708 608524
rect 249760 608512 249766 608524
rect 260190 608512 260196 608524
rect 249760 608484 260196 608512
rect 249760 608472 249766 608484
rect 260190 608472 260196 608484
rect 260248 608472 260254 608524
rect 333698 608472 333704 608524
rect 333756 608512 333762 608524
rect 344278 608512 344284 608524
rect 333756 608484 344284 608512
rect 333756 608472 333762 608484
rect 344278 608472 344284 608484
rect 344336 608472 344342 608524
rect 374638 608472 374644 608524
rect 374696 608512 374702 608524
rect 379698 608512 379704 608524
rect 374696 608484 379704 608512
rect 374696 608472 374702 608484
rect 379698 608472 379704 608484
rect 379756 608472 379762 608524
rect 390002 608472 390008 608524
rect 390060 608512 390066 608524
rect 400858 608512 400864 608524
rect 390060 608484 400864 608512
rect 390060 608472 390066 608484
rect 400858 608472 400864 608484
rect 400916 608472 400922 608524
rect 417694 608472 417700 608524
rect 417752 608512 417758 608524
rect 428550 608512 428556 608524
rect 417752 608484 428556 608512
rect 417752 608472 417758 608484
rect 428550 608472 428556 608484
rect 428608 608472 428614 608524
rect 445662 608472 445668 608524
rect 445720 608512 445726 608524
rect 456058 608512 456064 608524
rect 445720 608484 456064 608512
rect 445720 608472 445726 608484
rect 456058 608472 456064 608484
rect 456116 608472 456122 608524
rect 529658 608472 529664 608524
rect 529716 608512 529722 608524
rect 540238 608512 540244 608524
rect 529716 608484 540244 608512
rect 529716 608472 529722 608484
rect 540238 608472 540244 608484
rect 540296 608472 540302 608524
rect 72050 608444 72056 608456
rect 45526 608416 72056 608444
rect 72050 608404 72056 608416
rect 72108 608404 72114 608456
rect 127066 608404 127072 608456
rect 127124 608444 127130 608456
rect 156046 608444 156052 608456
rect 127124 608416 156052 608444
rect 127124 608404 127130 608416
rect 156046 608404 156052 608416
rect 156104 608404 156110 608456
rect 238846 608404 238852 608456
rect 238904 608444 238910 608456
rect 268010 608444 268016 608456
rect 238904 608416 268016 608444
rect 238904 608404 238910 608416
rect 268010 608404 268016 608416
rect 268068 608404 268074 608456
rect 323026 608404 323032 608456
rect 323084 608444 323090 608456
rect 352006 608444 352012 608456
rect 323084 608416 352012 608444
rect 323084 608404 323090 608416
rect 352006 608404 352012 608416
rect 352064 608404 352070 608456
rect 434806 608404 434812 608456
rect 434864 608444 434870 608456
rect 463694 608444 463700 608456
rect 434864 608416 463700 608444
rect 434864 608404 434870 608416
rect 463694 608404 463700 608416
rect 463752 608404 463758 608456
rect 518986 608404 518992 608456
rect 519044 608444 519050 608456
rect 547874 608444 547880 608456
rect 519044 608416 547880 608444
rect 519044 608404 519050 608416
rect 547874 608404 547880 608416
rect 547932 608404 547938 608456
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 11698 605860 11704 605872
rect 3292 605832 11704 605860
rect 3292 605820 3298 605832
rect 11698 605820 11704 605832
rect 11756 605820 11762 605872
rect 71130 604596 71136 604648
rect 71188 604636 71194 604648
rect 82262 604636 82268 604648
rect 71188 604608 82268 604636
rect 71188 604596 71194 604608
rect 82262 604596 82268 604608
rect 82320 604596 82326 604648
rect 99466 604596 99472 604648
rect 99524 604636 99530 604648
rect 100386 604636 100392 604648
rect 99524 604608 100392 604636
rect 99524 604596 99530 604608
rect 100386 604596 100392 604608
rect 100444 604596 100450 604648
rect 183646 604596 183652 604648
rect 183704 604636 183710 604648
rect 222286 604636 222292 604648
rect 183704 604608 222292 604636
rect 183704 604596 183710 604608
rect 222286 604596 222292 604608
rect 222344 604596 222350 604648
rect 266998 604596 267004 604648
rect 267056 604636 267062 604648
rect 277946 604636 277952 604648
rect 267056 604608 277952 604636
rect 267056 604596 267062 604608
rect 277946 604596 277952 604608
rect 278004 604596 278010 604648
rect 295426 604596 295432 604648
rect 295484 604636 295490 604648
rect 334250 604636 334256 604648
rect 295484 604608 334256 604636
rect 295484 604596 295490 604608
rect 334250 604596 334256 604608
rect 334308 604596 334314 604648
rect 352006 604596 352012 604648
rect 352064 604636 352070 604648
rect 352064 604608 364334 604636
rect 352064 604596 352070 604608
rect 36630 604528 36636 604580
rect 36688 604568 36694 604580
rect 53926 604568 53932 604580
rect 36688 604540 53932 604568
rect 36688 604528 36694 604540
rect 53926 604528 53932 604540
rect 53984 604528 53990 604580
rect 71866 604528 71872 604580
rect 71924 604568 71930 604580
rect 109954 604568 109960 604580
rect 71924 604540 109960 604568
rect 71924 604528 71930 604540
rect 109954 604528 109960 604540
rect 110012 604528 110018 604580
rect 151078 604528 151084 604580
rect 151136 604568 151142 604580
rect 156598 604568 156604 604580
rect 151136 604540 156604 604568
rect 151136 604528 151142 604540
rect 156598 604528 156604 604540
rect 156656 604528 156662 604580
rect 182818 604528 182824 604580
rect 182876 604568 182882 604580
rect 193950 604568 193956 604580
rect 182876 604540 193956 604568
rect 182876 604528 182882 604540
rect 193950 604528 193956 604540
rect 194008 604528 194014 604580
rect 232498 604528 232504 604580
rect 232556 604568 232562 604580
rect 232556 604540 248414 604568
rect 232556 604528 232562 604540
rect 26234 604460 26240 604512
rect 26292 604500 26298 604512
rect 35434 604500 35440 604512
rect 26292 604472 35440 604500
rect 26292 604460 26298 604472
rect 35434 604460 35440 604472
rect 35492 604460 35498 604512
rect 66898 604460 66904 604512
rect 66956 604500 66962 604512
rect 72602 604500 72608 604512
rect 66956 604472 72608 604500
rect 66956 604460 66962 604472
rect 72602 604460 72608 604472
rect 72660 604460 72666 604512
rect 93118 604460 93124 604512
rect 93176 604500 93182 604512
rect 100294 604500 100300 604512
rect 93176 604472 100300 604500
rect 93176 604460 93182 604472
rect 100294 604460 100300 604472
rect 100352 604460 100358 604512
rect 100386 604460 100392 604512
rect 100444 604500 100450 604512
rect 138290 604500 138296 604512
rect 100444 604472 138296 604500
rect 100444 604460 100450 604472
rect 138290 604460 138296 604472
rect 138348 604460 138354 604512
rect 149698 604460 149704 604512
rect 149756 604500 149762 604512
rect 166258 604500 166264 604512
rect 149756 604472 166264 604500
rect 149756 604460 149762 604472
rect 166258 604460 166264 604472
rect 166316 604460 166322 604512
rect 177298 604460 177304 604512
rect 177356 604500 177362 604512
rect 184290 604500 184296 604512
rect 177356 604472 184296 604500
rect 177356 604460 177362 604472
rect 184290 604460 184296 604472
rect 184348 604460 184354 604512
rect 233970 604460 233976 604512
rect 234028 604500 234034 604512
rect 240594 604500 240600 604512
rect 234028 604472 240600 604500
rect 234028 604460 234034 604472
rect 240594 604460 240600 604472
rect 240652 604460 240658 604512
rect 248386 604500 248414 604540
rect 267826 604528 267832 604580
rect 267884 604568 267890 604580
rect 306282 604568 306288 604580
rect 267884 604540 306288 604568
rect 267884 604528 267890 604540
rect 306282 604528 306288 604540
rect 306340 604528 306346 604580
rect 347038 604528 347044 604580
rect 347096 604568 347102 604580
rect 361942 604568 361948 604580
rect 347096 604540 361948 604568
rect 347096 604528 347102 604540
rect 361942 604528 361948 604540
rect 362000 604528 362006 604580
rect 364306 604568 364334 604608
rect 379606 604596 379612 604648
rect 379664 604636 379670 604648
rect 418246 604636 418252 604648
rect 379664 604608 418252 604636
rect 379664 604596 379670 604608
rect 418246 604596 418252 604608
rect 418304 604596 418310 604648
rect 462958 604596 462964 604648
rect 463016 604636 463022 604648
rect 474274 604636 474280 604648
rect 463016 604608 474280 604636
rect 463016 604596 463022 604608
rect 474274 604596 474280 604608
rect 474332 604596 474338 604648
rect 491386 604596 491392 604648
rect 491444 604636 491450 604648
rect 529934 604636 529940 604648
rect 491444 604608 529940 604636
rect 491444 604596 491450 604608
rect 529934 604596 529940 604608
rect 529992 604596 529998 604648
rect 390278 604568 390284 604580
rect 364306 604540 390284 604568
rect 390278 604528 390284 604540
rect 390336 604528 390342 604580
rect 400950 604528 400956 604580
rect 401008 604568 401014 604580
rect 408586 604568 408592 604580
rect 401008 604540 408592 604568
rect 401008 604528 401014 604540
rect 408586 604528 408592 604540
rect 408644 604528 408650 604580
rect 429838 604528 429844 604580
rect 429896 604568 429902 604580
rect 436278 604568 436284 604580
rect 429896 604540 436284 604568
rect 429896 604528 429902 604540
rect 436278 604528 436284 604540
rect 436336 604528 436342 604580
rect 463786 604528 463792 604580
rect 463844 604568 463850 604580
rect 502242 604568 502248 604580
rect 463844 604540 502248 604568
rect 463844 604528 463850 604540
rect 502242 604528 502248 604540
rect 502300 604528 502306 604580
rect 512638 604528 512644 604580
rect 512696 604568 512702 604580
rect 520274 604568 520280 604580
rect 512696 604540 520280 604568
rect 512696 604528 512702 604540
rect 520274 604528 520280 604540
rect 520332 604528 520338 604580
rect 541618 604528 541624 604580
rect 541676 604568 541682 604580
rect 541676 604540 557534 604568
rect 541676 604528 541682 604540
rect 250254 604500 250260 604512
rect 248386 604472 250260 604500
rect 250254 604460 250260 604472
rect 250312 604460 250318 604512
rect 261478 604460 261484 604512
rect 261536 604500 261542 604512
rect 268286 604500 268292 604512
rect 261536 604472 268292 604500
rect 261536 604460 261542 604472
rect 268286 604460 268292 604472
rect 268344 604460 268350 604512
rect 289078 604460 289084 604512
rect 289136 604500 289142 604512
rect 296622 604500 296628 604512
rect 289136 604472 296628 604500
rect 289136 604460 289142 604472
rect 296622 604460 296628 604472
rect 296680 604460 296686 604512
rect 318058 604460 318064 604512
rect 318116 604500 318122 604512
rect 324590 604500 324596 604512
rect 318116 604472 324596 604500
rect 318116 604460 318122 604472
rect 324590 604460 324596 604472
rect 324648 604460 324654 604512
rect 348418 604460 348424 604512
rect 348476 604500 348482 604512
rect 352282 604500 352288 604512
rect 348476 604472 352288 604500
rect 348476 604460 348482 604472
rect 352282 604460 352288 604472
rect 352340 604460 352346 604512
rect 373258 604460 373264 604512
rect 373316 604500 373322 604512
rect 380618 604500 380624 604512
rect 373316 604472 380624 604500
rect 373316 604460 373322 604472
rect 380618 604460 380624 604472
rect 380676 604460 380682 604512
rect 428458 604460 428464 604512
rect 428516 604500 428522 604512
rect 445938 604500 445944 604512
rect 428516 604472 445944 604500
rect 428516 604460 428522 604472
rect 445938 604460 445944 604472
rect 445996 604460 446002 604512
rect 457438 604460 457444 604512
rect 457496 604500 457502 604512
rect 464614 604500 464620 604512
rect 457496 604472 464620 604500
rect 457496 604460 457502 604472
rect 464614 604460 464620 604472
rect 464672 604460 464678 604512
rect 485038 604460 485044 604512
rect 485096 604500 485102 604512
rect 492582 604500 492588 604512
rect 485096 604472 492588 604500
rect 485096 604460 485102 604472
rect 492582 604460 492588 604472
rect 492640 604460 492646 604512
rect 544378 604460 544384 604512
rect 544436 604500 544442 604512
rect 548610 604500 548616 604512
rect 544436 604472 548616 604500
rect 544436 604460 544442 604472
rect 548610 604460 548616 604472
rect 548668 604460 548674 604512
rect 557506 604500 557534 604540
rect 558270 604500 558276 604512
rect 557506 604472 558276 604500
rect 558270 604460 558276 604472
rect 558328 604460 558334 604512
rect 120166 602216 120172 602268
rect 120224 602256 120230 602268
rect 122098 602256 122104 602268
rect 120224 602228 122104 602256
rect 120224 602216 120230 602228
rect 122098 602216 122104 602228
rect 122156 602216 122162 602268
rect 124858 602216 124864 602268
rect 124916 602256 124922 602268
rect 128262 602256 128268 602268
rect 124916 602228 128268 602256
rect 124916 602216 124922 602228
rect 128262 602216 128268 602228
rect 128320 602216 128326 602268
rect 210418 602216 210424 602268
rect 210476 602256 210482 602268
rect 212350 602256 212356 602268
rect 210476 602228 212356 602256
rect 210476 602216 210482 602228
rect 212350 602216 212356 602228
rect 212408 602216 212414 602268
rect 512086 602216 512092 602268
rect 512144 602256 512150 602268
rect 514018 602256 514024 602268
rect 512144 602228 514024 602256
rect 512144 602216 512150 602228
rect 514018 602216 514024 602228
rect 514076 602216 514082 602268
rect 182082 601808 182088 601860
rect 182140 601848 182146 601860
rect 233234 601848 233240 601860
rect 182140 601820 233240 601848
rect 182140 601808 182146 601820
rect 233234 601808 233240 601820
rect 233292 601808 233298 601860
rect 350442 601808 350448 601860
rect 350500 601848 350506 601860
rect 401594 601848 401600 601860
rect 350500 601820 401600 601848
rect 350500 601808 350506 601820
rect 401594 601808 401600 601820
rect 401652 601808 401658 601860
rect 462222 601808 462228 601860
rect 462280 601848 462286 601860
rect 513374 601848 513380 601860
rect 462280 601820 513380 601848
rect 462280 601808 462286 601820
rect 513374 601808 513380 601820
rect 513432 601808 513438 601860
rect 42702 601740 42708 601792
rect 42760 601780 42766 601792
rect 93854 601780 93860 601792
rect 42760 601752 93860 601780
rect 42760 601740 42766 601752
rect 93854 601740 93860 601752
rect 93912 601740 93918 601792
rect 97902 601740 97908 601792
rect 97960 601780 97966 601792
rect 149054 601780 149060 601792
rect 97960 601752 149060 601780
rect 97960 601740 97966 601752
rect 149054 601740 149060 601752
rect 149112 601740 149118 601792
rect 154482 601740 154488 601792
rect 154540 601780 154546 601792
rect 205634 601780 205640 601792
rect 154540 601752 205640 601780
rect 154540 601740 154546 601752
rect 205634 601740 205640 601752
rect 205692 601740 205698 601792
rect 238662 601740 238668 601792
rect 238720 601780 238726 601792
rect 289814 601780 289820 601792
rect 238720 601752 289820 601780
rect 238720 601740 238726 601752
rect 289814 601740 289820 601752
rect 289872 601740 289878 601792
rect 293862 601740 293868 601792
rect 293920 601780 293926 601792
rect 345014 601780 345020 601792
rect 293920 601752 345020 601780
rect 293920 601740 293926 601752
rect 345014 601740 345020 601752
rect 345072 601740 345078 601792
rect 378042 601740 378048 601792
rect 378100 601780 378106 601792
rect 429286 601780 429292 601792
rect 378100 601752 429292 601780
rect 378100 601740 378106 601752
rect 429286 601740 429292 601752
rect 429344 601740 429350 601792
rect 434622 601740 434628 601792
rect 434680 601780 434686 601792
rect 485774 601780 485780 601792
rect 434680 601752 485780 601780
rect 434680 601740 434686 601752
rect 485774 601740 485780 601752
rect 485832 601740 485838 601792
rect 518802 601740 518808 601792
rect 518860 601780 518866 601792
rect 569954 601780 569960 601792
rect 518860 601752 569960 601780
rect 518860 601740 518866 601752
rect 569954 601740 569960 601752
rect 570012 601740 570018 601792
rect 13538 601672 13544 601724
rect 13596 601712 13602 601724
rect 66254 601712 66260 601724
rect 13596 601684 66260 601712
rect 13596 601672 13602 601684
rect 66254 601672 66260 601684
rect 66312 601672 66318 601724
rect 70302 601672 70308 601724
rect 70360 601712 70366 601724
rect 121454 601712 121460 601724
rect 70360 601684 121460 601712
rect 70360 601672 70366 601684
rect 121454 601672 121460 601684
rect 121512 601672 121518 601724
rect 126882 601672 126888 601724
rect 126940 601712 126946 601724
rect 178034 601712 178040 601724
rect 126940 601684 178040 601712
rect 126940 601672 126946 601684
rect 178034 601672 178040 601684
rect 178092 601672 178098 601724
rect 209682 601672 209688 601724
rect 209740 601712 209746 601724
rect 262214 601712 262220 601724
rect 209740 601684 262220 601712
rect 209740 601672 209746 601684
rect 262214 601672 262220 601684
rect 262272 601672 262278 601724
rect 266262 601672 266268 601724
rect 266320 601712 266326 601724
rect 317414 601712 317420 601724
rect 266320 601684 317420 601712
rect 266320 601672 266326 601684
rect 317414 601672 317420 601684
rect 317472 601672 317478 601724
rect 322842 601672 322848 601724
rect 322900 601712 322906 601724
rect 373994 601712 374000 601724
rect 322900 601684 374000 601712
rect 322900 601672 322906 601684
rect 373994 601672 374000 601684
rect 374052 601672 374058 601724
rect 405642 601672 405648 601724
rect 405700 601712 405706 601724
rect 458174 601712 458180 601724
rect 405700 601684 458180 601712
rect 405700 601672 405706 601684
rect 458174 601672 458180 601684
rect 458232 601672 458238 601724
rect 489822 601672 489828 601724
rect 489880 601712 489886 601724
rect 542354 601712 542360 601724
rect 489880 601684 542360 601712
rect 489880 601672 489886 601684
rect 542354 601672 542360 601684
rect 542412 601672 542418 601724
rect 204254 599224 204260 599276
rect 204312 599264 204318 599276
rect 204990 599264 204996 599276
rect 204312 599236 204996 599264
rect 204312 599224 204318 599236
rect 204990 599224 204996 599236
rect 205048 599224 205054 599276
rect 15194 580932 15200 580984
rect 15252 580972 15258 580984
rect 35894 580972 35900 580984
rect 15252 580944 35900 580972
rect 15252 580932 15258 580944
rect 35894 580932 35900 580944
rect 35952 580932 35958 580984
rect 36078 580932 36084 580984
rect 36136 580972 36142 580984
rect 63586 580972 63592 580984
rect 36136 580944 63592 580972
rect 36136 580932 36142 580944
rect 63586 580932 63592 580944
rect 63644 580932 63650 580984
rect 64046 580932 64052 580984
rect 64104 580972 64110 580984
rect 91922 580972 91928 580984
rect 64104 580944 91928 580972
rect 64104 580932 64110 580944
rect 91922 580932 91928 580944
rect 91980 580932 91986 580984
rect 92106 580932 92112 580984
rect 92164 580972 92170 580984
rect 119614 580972 119620 580984
rect 92164 580944 119620 580972
rect 92164 580932 92170 580944
rect 119614 580932 119620 580944
rect 119672 580932 119678 580984
rect 122098 580932 122104 580984
rect 122156 580972 122162 580984
rect 147950 580972 147956 580984
rect 122156 580944 147956 580972
rect 122156 580932 122162 580944
rect 147950 580932 147956 580944
rect 148008 580932 148014 580984
rect 148042 580932 148048 580984
rect 148100 580972 148106 580984
rect 175918 580972 175924 580984
rect 148100 580944 175924 580972
rect 148100 580932 148106 580944
rect 175918 580932 175924 580944
rect 175976 580932 175982 580984
rect 176102 580932 176108 580984
rect 176160 580972 176166 580984
rect 203610 580972 203616 580984
rect 176160 580944 203616 580972
rect 176160 580932 176166 580944
rect 203610 580932 203616 580944
rect 203668 580932 203674 580984
rect 204990 580932 204996 580984
rect 205048 580972 205054 580984
rect 231946 580972 231952 580984
rect 205048 580944 231952 580972
rect 205048 580932 205054 580944
rect 231946 580932 231952 580944
rect 232004 580932 232010 580984
rect 232038 580932 232044 580984
rect 232096 580972 232102 580984
rect 259914 580972 259920 580984
rect 232096 580944 259920 580972
rect 232096 580932 232102 580944
rect 259914 580932 259920 580944
rect 259972 580932 259978 580984
rect 260098 580932 260104 580984
rect 260156 580972 260162 580984
rect 287606 580972 287612 580984
rect 260156 580944 287612 580972
rect 260156 580932 260162 580944
rect 287606 580932 287612 580944
rect 287664 580932 287670 580984
rect 288066 580932 288072 580984
rect 288124 580972 288130 580984
rect 315942 580972 315948 580984
rect 288124 580944 315948 580972
rect 288124 580932 288130 580944
rect 315942 580932 315948 580944
rect 316000 580932 316006 580984
rect 316678 580932 316684 580984
rect 316736 580972 316742 580984
rect 343910 580972 343916 580984
rect 316736 580944 343916 580972
rect 316736 580932 316742 580944
rect 343910 580932 343916 580944
rect 343968 580932 343974 580984
rect 344094 580932 344100 580984
rect 344152 580972 344158 580984
rect 371602 580972 371608 580984
rect 344152 580944 371608 580972
rect 344152 580932 344158 580944
rect 371602 580932 371608 580944
rect 371660 580932 371666 580984
rect 372062 580932 372068 580984
rect 372120 580972 372126 580984
rect 399938 580972 399944 580984
rect 372120 580944 399944 580972
rect 372120 580932 372126 580944
rect 399938 580932 399944 580944
rect 399996 580932 400002 580984
rect 400858 580932 400864 580984
rect 400916 580972 400922 580984
rect 427906 580972 427912 580984
rect 400916 580944 427912 580972
rect 400916 580932 400922 580944
rect 427906 580932 427912 580944
rect 427964 580932 427970 580984
rect 428090 580932 428096 580984
rect 428148 580972 428154 580984
rect 455598 580972 455604 580984
rect 428148 580944 455604 580972
rect 428148 580932 428154 580944
rect 455598 580932 455604 580944
rect 455656 580932 455662 580984
rect 456058 580932 456064 580984
rect 456116 580972 456122 580984
rect 483934 580972 483940 580984
rect 456116 580944 483940 580972
rect 456116 580932 456122 580944
rect 483934 580932 483940 580944
rect 483992 580932 483998 580984
rect 484026 580932 484032 580984
rect 484084 580972 484090 580984
rect 511902 580972 511908 580984
rect 484084 580944 511908 580972
rect 484084 580932 484090 580944
rect 511902 580932 511908 580944
rect 511960 580932 511966 580984
rect 514018 580932 514024 580984
rect 514076 580972 514082 580984
rect 539594 580972 539600 580984
rect 514076 580944 539600 580972
rect 514076 580932 514082 580944
rect 539594 580932 539600 580944
rect 539652 580932 539658 580984
rect 540054 580932 540060 580984
rect 540112 580972 540118 580984
rect 567930 580972 567936 580984
rect 540112 580944 567936 580972
rect 540112 580932 540118 580944
rect 567930 580932 567936 580944
rect 567988 580932 567994 580984
rect 16574 580864 16580 580916
rect 16632 580904 16638 580916
rect 36630 580904 36636 580916
rect 16632 580876 36636 580904
rect 16632 580864 16638 580876
rect 36630 580864 36636 580876
rect 36688 580864 36694 580916
rect 44910 580864 44916 580916
rect 44968 580904 44974 580916
rect 71130 580904 71136 580916
rect 44968 580876 71136 580904
rect 44968 580864 44974 580876
rect 71130 580864 71136 580876
rect 71188 580864 71194 580916
rect 82262 580864 82268 580916
rect 82320 580904 82326 580916
rect 93118 580904 93124 580916
rect 82320 580876 93124 580904
rect 82320 580864 82326 580876
rect 93118 580864 93124 580876
rect 93176 580864 93182 580916
rect 110230 580864 110236 580916
rect 110288 580904 110294 580916
rect 124858 580904 124864 580916
rect 110288 580876 124864 580904
rect 110288 580864 110294 580876
rect 124858 580864 124864 580876
rect 124916 580864 124922 580916
rect 128630 580864 128636 580916
rect 128688 580904 128694 580916
rect 149698 580904 149704 580916
rect 128688 580876 149704 580904
rect 128688 580864 128694 580876
rect 149698 580864 149704 580876
rect 149756 580864 149762 580916
rect 156598 580864 156604 580916
rect 156656 580904 156662 580916
rect 182818 580904 182824 580916
rect 156656 580876 182824 580904
rect 156656 580864 156662 580876
rect 182818 580864 182824 580876
rect 182876 580864 182882 580916
rect 194502 580864 194508 580916
rect 194560 580904 194566 580916
rect 210418 580904 210424 580916
rect 194560 580876 210424 580904
rect 194560 580864 194566 580876
rect 210418 580864 210424 580876
rect 210476 580864 210482 580916
rect 212626 580864 212632 580916
rect 212684 580904 212690 580916
rect 232498 580904 232504 580916
rect 212684 580876 232504 580904
rect 212684 580864 212690 580876
rect 232498 580864 232504 580876
rect 232556 580864 232562 580916
rect 240594 580864 240600 580916
rect 240652 580904 240658 580916
rect 266998 580904 267004 580916
rect 240652 580876 267004 580904
rect 240652 580864 240658 580876
rect 266998 580864 267004 580876
rect 267056 580864 267062 580916
rect 278590 580864 278596 580916
rect 278648 580904 278654 580916
rect 289078 580904 289084 580916
rect 278648 580876 289084 580904
rect 278648 580864 278654 580876
rect 289078 580864 289084 580876
rect 289136 580864 289142 580916
rect 306282 580864 306288 580916
rect 306340 580904 306346 580916
rect 318058 580904 318064 580916
rect 306340 580876 318064 580904
rect 306340 580864 306346 580876
rect 318058 580864 318064 580876
rect 318116 580864 318122 580916
rect 324590 580864 324596 580916
rect 324648 580904 324654 580916
rect 347038 580904 347044 580916
rect 324648 580876 347044 580904
rect 324648 580864 324654 580876
rect 347038 580864 347044 580876
rect 347096 580864 347102 580916
rect 362586 580864 362592 580916
rect 362644 580904 362650 580916
rect 373258 580904 373264 580916
rect 362644 580876 373264 580904
rect 362644 580864 362650 580876
rect 373258 580864 373264 580876
rect 373316 580864 373322 580916
rect 390278 580864 390284 580916
rect 390336 580904 390342 580916
rect 400950 580904 400956 580916
rect 390336 580876 400956 580904
rect 390336 580864 390342 580876
rect 400950 580864 400956 580876
rect 401008 580864 401014 580916
rect 408586 580864 408592 580916
rect 408644 580904 408650 580916
rect 428458 580904 428464 580916
rect 408644 580876 428464 580904
rect 408644 580864 408650 580876
rect 428458 580864 428464 580876
rect 428516 580864 428522 580916
rect 436922 580864 436928 580916
rect 436980 580904 436986 580916
rect 462958 580904 462964 580916
rect 436980 580876 462964 580904
rect 436980 580864 436986 580876
rect 462958 580864 462964 580876
rect 463016 580864 463022 580916
rect 474274 580864 474280 580916
rect 474332 580904 474338 580916
rect 485038 580904 485044 580916
rect 474332 580876 485044 580904
rect 474332 580864 474338 580876
rect 485038 580864 485044 580876
rect 485096 580864 485102 580916
rect 502242 580864 502248 580916
rect 502300 580904 502306 580916
rect 512638 580904 512644 580916
rect 502300 580876 512644 580904
rect 502300 580864 502306 580876
rect 512638 580864 512644 580876
rect 512696 580864 512702 580916
rect 520918 580864 520924 580916
rect 520976 580904 520982 580916
rect 541618 580904 541624 580916
rect 520976 580876 541624 580904
rect 520976 580864 520982 580876
rect 541618 580864 541624 580876
rect 541676 580864 541682 580916
rect 26234 580796 26240 580848
rect 26292 580836 26298 580848
rect 43530 580836 43536 580848
rect 26292 580808 43536 580836
rect 26292 580796 26298 580808
rect 43530 580796 43536 580808
rect 43588 580796 43594 580848
rect 54570 580796 54576 580848
rect 54628 580836 54634 580848
rect 66898 580836 66904 580848
rect 54628 580808 66904 580836
rect 54628 580796 54634 580808
rect 66898 580796 66904 580808
rect 66956 580796 66962 580848
rect 138290 580796 138296 580848
rect 138348 580836 138354 580848
rect 151078 580836 151084 580848
rect 138348 580808 151084 580836
rect 138348 580796 138354 580808
rect 151078 580796 151084 580808
rect 151136 580796 151142 580848
rect 166258 580796 166264 580848
rect 166316 580836 166322 580848
rect 177298 580836 177304 580848
rect 166316 580808 177304 580836
rect 166316 580796 166322 580808
rect 177298 580796 177304 580808
rect 177356 580796 177362 580848
rect 222286 580796 222292 580848
rect 222344 580836 222350 580848
rect 233970 580836 233976 580848
rect 222344 580808 233976 580836
rect 222344 580796 222350 580808
rect 233970 580796 233976 580808
rect 234028 580796 234034 580848
rect 250254 580796 250260 580848
rect 250312 580836 250318 580848
rect 261478 580836 261484 580848
rect 250312 580808 261484 580836
rect 250312 580796 250318 580808
rect 261478 580796 261484 580808
rect 261536 580796 261542 580848
rect 334250 580796 334256 580848
rect 334308 580836 334314 580848
rect 348418 580836 348424 580848
rect 334308 580808 348424 580836
rect 334308 580796 334314 580808
rect 348418 580796 348424 580808
rect 348476 580796 348482 580848
rect 418246 580796 418252 580848
rect 418304 580836 418310 580848
rect 429838 580836 429844 580848
rect 418304 580808 429844 580836
rect 418304 580796 418310 580808
rect 429838 580796 429844 580808
rect 429896 580796 429902 580848
rect 446582 580796 446588 580848
rect 446640 580836 446646 580848
rect 457438 580836 457444 580848
rect 446640 580808 457444 580836
rect 446640 580796 446646 580808
rect 457438 580796 457444 580808
rect 457496 580796 457502 580848
rect 530578 580796 530584 580848
rect 530636 580836 530642 580848
rect 544378 580836 544384 580848
rect 530636 580808 544384 580836
rect 530636 580796 530642 580808
rect 544378 580796 544384 580808
rect 544436 580796 544442 580848
rect 558270 580252 558276 580304
rect 558328 580292 558334 580304
rect 567470 580292 567476 580304
rect 558328 580264 567476 580292
rect 558328 580252 558334 580264
rect 567470 580252 567476 580264
rect 567528 580252 567534 580304
rect 548334 578892 548340 578944
rect 548392 578932 548398 578944
rect 568022 578932 568028 578944
rect 548392 578904 568028 578932
rect 548392 578892 548398 578904
rect 568022 578892 568028 578904
rect 568080 578892 568086 578944
rect 212258 578416 212264 578468
rect 212316 578456 212322 578468
rect 232682 578456 232688 578468
rect 212316 578428 232688 578456
rect 212316 578416 212322 578428
rect 232682 578416 232688 578428
rect 232740 578416 232746 578468
rect 296346 578416 296352 578468
rect 296404 578456 296410 578468
rect 316770 578456 316776 578468
rect 296404 578428 316776 578456
rect 296404 578416 296410 578428
rect 316770 578416 316776 578428
rect 316828 578416 316834 578468
rect 408034 578416 408040 578468
rect 408092 578456 408098 578468
rect 428642 578456 428648 578468
rect 408092 578428 428648 578456
rect 408092 578416 408098 578428
rect 428642 578416 428648 578428
rect 428700 578416 428706 578468
rect 492030 578416 492036 578468
rect 492088 578456 492094 578468
rect 512730 578456 512736 578468
rect 492088 578428 512736 578456
rect 492088 578416 492094 578428
rect 512730 578416 512736 578428
rect 512788 578416 512794 578468
rect 148410 578348 148416 578400
rect 148468 578388 148474 578400
rect 165614 578388 165620 578400
rect 148468 578360 165620 578388
rect 148468 578348 148474 578360
rect 165614 578348 165620 578360
rect 165672 578348 165678 578400
rect 175458 578348 175464 578400
rect 175516 578388 175522 578400
rect 193674 578388 193680 578400
rect 175516 578360 193680 578388
rect 175516 578348 175522 578360
rect 193674 578348 193680 578360
rect 193732 578348 193738 578400
rect 203518 578348 203524 578400
rect 203576 578388 203582 578400
rect 221366 578388 221372 578400
rect 203576 578360 221372 578388
rect 203576 578348 203582 578360
rect 221366 578348 221372 578360
rect 221424 578348 221430 578400
rect 260190 578348 260196 578400
rect 260248 578388 260254 578400
rect 277670 578388 277676 578400
rect 260248 578360 277676 578388
rect 260248 578348 260254 578360
rect 277670 578348 277676 578360
rect 277728 578348 277734 578400
rect 287514 578348 287520 578400
rect 287572 578388 287578 578400
rect 305362 578388 305368 578400
rect 287572 578360 305368 578388
rect 287572 578348 287578 578360
rect 305362 578348 305368 578360
rect 305420 578348 305426 578400
rect 345658 578348 345664 578400
rect 345716 578388 345722 578400
rect 361666 578388 361672 578400
rect 345716 578360 361672 578388
rect 345716 578348 345722 578360
rect 361666 578348 361672 578360
rect 361724 578348 361730 578400
rect 371510 578348 371516 578400
rect 371568 578388 371574 578400
rect 389358 578388 389364 578400
rect 371568 578360 389364 578388
rect 371568 578348 371574 578360
rect 389358 578348 389364 578360
rect 389416 578348 389422 578400
rect 399478 578348 399484 578400
rect 399536 578388 399542 578400
rect 417694 578388 417700 578400
rect 399536 578360 417700 578388
rect 399536 578348 399542 578360
rect 417694 578348 417700 578360
rect 417752 578348 417758 578400
rect 456150 578348 456156 578400
rect 456208 578388 456214 578400
rect 473538 578388 473544 578400
rect 456208 578360 473544 578388
rect 456208 578348 456214 578360
rect 473538 578348 473544 578360
rect 473596 578348 473602 578400
rect 483474 578348 483480 578400
rect 483532 578388 483538 578400
rect 501690 578388 501696 578400
rect 483532 578360 501696 578388
rect 483532 578348 483538 578360
rect 501690 578348 501696 578360
rect 501748 578348 501754 578400
rect 36722 578280 36728 578332
rect 36780 578320 36786 578332
rect 53650 578320 53656 578332
rect 36780 578292 53656 578320
rect 36780 578280 36786 578292
rect 53650 578280 53656 578292
rect 53708 578280 53714 578332
rect 64322 578280 64328 578332
rect 64380 578320 64386 578332
rect 81434 578320 81440 578332
rect 64380 578292 81440 578320
rect 64380 578280 64386 578292
rect 81434 578280 81440 578292
rect 81492 578280 81498 578332
rect 91462 578280 91468 578332
rect 91520 578320 91526 578332
rect 109678 578320 109684 578332
rect 91520 578292 109684 578320
rect 91520 578280 91526 578292
rect 109678 578280 109684 578292
rect 109736 578280 109742 578332
rect 119430 578280 119436 578332
rect 119488 578320 119494 578332
rect 137646 578320 137652 578332
rect 119488 578292 137652 578320
rect 119488 578280 119494 578292
rect 137646 578280 137652 578292
rect 137704 578280 137710 578332
rect 156322 578280 156328 578332
rect 156380 578320 156386 578332
rect 178678 578320 178684 578332
rect 156380 578292 178684 578320
rect 156380 578280 156386 578292
rect 178678 578280 178684 578292
rect 178736 578280 178742 578332
rect 232498 578280 232504 578332
rect 232556 578320 232562 578332
rect 249702 578320 249708 578332
rect 232556 578292 249708 578320
rect 232556 578280 232562 578292
rect 249702 578280 249708 578292
rect 249760 578280 249766 578332
rect 268010 578280 268016 578332
rect 268068 578320 268074 578332
rect 287698 578320 287704 578332
rect 268068 578292 287704 578320
rect 268068 578280 268074 578292
rect 287698 578280 287704 578292
rect 287756 578280 287762 578332
rect 315482 578280 315488 578332
rect 315540 578320 315546 578332
rect 333698 578320 333704 578332
rect 315540 578292 333704 578320
rect 315540 578280 315546 578292
rect 333698 578280 333704 578292
rect 333756 578280 333762 578332
rect 352006 578280 352012 578332
rect 352064 578320 352070 578332
rect 374638 578320 374644 578332
rect 352064 578292 374644 578320
rect 352064 578280 352070 578292
rect 374638 578280 374644 578292
rect 374696 578280 374702 578332
rect 428458 578280 428464 578332
rect 428516 578320 428522 578332
rect 445662 578320 445668 578332
rect 428516 578292 445668 578320
rect 428516 578280 428522 578292
rect 445662 578280 445668 578292
rect 445720 578280 445726 578332
rect 464338 578280 464344 578332
rect 464396 578320 464402 578332
rect 483658 578320 483664 578332
rect 464396 578292 483664 578320
rect 464396 578280 464402 578292
rect 483658 578280 483664 578292
rect 483716 578280 483722 578332
rect 511442 578280 511448 578332
rect 511500 578320 511506 578332
rect 529658 578320 529664 578332
rect 511500 578292 529664 578320
rect 511500 578280 511506 578292
rect 529658 578280 529664 578292
rect 529716 578280 529722 578332
rect 541618 578280 541624 578332
rect 541676 578320 541682 578332
rect 557534 578320 557540 578332
rect 541676 578292 557540 578320
rect 541676 578280 541682 578292
rect 557534 578280 557540 578292
rect 557592 578280 557598 578332
rect 15838 578212 15844 578264
rect 15896 578252 15902 578264
rect 25682 578252 25688 578264
rect 15896 578224 25688 578252
rect 15896 578212 15902 578224
rect 25682 578212 25688 578224
rect 25740 578212 25746 578264
rect 36630 578212 36636 578264
rect 36688 578252 36694 578264
rect 63310 578252 63316 578264
rect 36688 578224 63316 578252
rect 36688 578212 36694 578224
rect 63310 578212 63316 578224
rect 63368 578212 63374 578264
rect 66898 578212 66904 578264
rect 66956 578252 66962 578264
rect 91094 578252 91100 578264
rect 66956 578224 91100 578252
rect 66956 578212 66962 578224
rect 91094 578212 91100 578224
rect 91152 578212 91158 578264
rect 93118 578212 93124 578264
rect 93176 578252 93182 578264
rect 119338 578252 119344 578264
rect 93176 578224 119344 578252
rect 93176 578212 93182 578224
rect 119338 578212 119344 578224
rect 119396 578212 119402 578264
rect 124858 578212 124864 578264
rect 124916 578252 124922 578264
rect 147306 578252 147312 578264
rect 124916 578224 147312 578252
rect 124916 578212 124922 578224
rect 147306 578212 147312 578224
rect 147364 578212 147370 578264
rect 148318 578212 148324 578264
rect 148376 578252 148382 578264
rect 175274 578252 175280 578264
rect 148376 578224 175280 578252
rect 148376 578212 148382 578224
rect 175274 578212 175280 578224
rect 175332 578212 175338 578264
rect 177298 578212 177304 578264
rect 177356 578252 177362 578264
rect 203334 578252 203340 578264
rect 177356 578224 203340 578252
rect 177356 578212 177362 578224
rect 203334 578212 203340 578224
rect 203392 578212 203398 578264
rect 204990 578212 204996 578264
rect 205048 578252 205054 578264
rect 231026 578252 231032 578264
rect 205048 578224 231032 578252
rect 205048 578212 205054 578224
rect 231026 578212 231032 578224
rect 231084 578212 231090 578264
rect 232590 578212 232596 578264
rect 232648 578252 232654 578264
rect 259362 578252 259368 578264
rect 232648 578224 259368 578252
rect 232648 578212 232654 578224
rect 259362 578212 259368 578224
rect 259420 578212 259426 578264
rect 260098 578212 260104 578264
rect 260156 578252 260162 578264
rect 287330 578252 287336 578264
rect 260156 578224 287336 578252
rect 260156 578212 260162 578224
rect 287330 578212 287336 578224
rect 287388 578212 287394 578264
rect 289078 578212 289084 578264
rect 289136 578252 289142 578264
rect 315022 578252 315028 578264
rect 289136 578224 315028 578252
rect 289136 578212 289142 578224
rect 315022 578212 315028 578224
rect 315080 578212 315086 578264
rect 316678 578212 316684 578264
rect 316736 578252 316742 578264
rect 343358 578252 343364 578264
rect 316736 578224 343364 578252
rect 316736 578212 316742 578224
rect 343358 578212 343364 578224
rect 343416 578212 343422 578264
rect 344278 578212 344284 578264
rect 344336 578252 344342 578264
rect 371326 578252 371332 578264
rect 344336 578224 371332 578252
rect 344336 578212 344342 578224
rect 371326 578212 371332 578224
rect 371384 578212 371390 578264
rect 373258 578212 373264 578264
rect 373316 578252 373322 578264
rect 399018 578252 399024 578264
rect 373316 578224 399024 578252
rect 373316 578212 373322 578224
rect 399018 578212 399024 578224
rect 399076 578212 399082 578264
rect 400858 578212 400864 578264
rect 400916 578252 400922 578264
rect 427354 578252 427360 578264
rect 400916 578224 427360 578252
rect 400916 578212 400922 578224
rect 427354 578212 427360 578224
rect 427412 578212 427418 578264
rect 428550 578212 428556 578264
rect 428608 578252 428614 578264
rect 455322 578252 455328 578264
rect 428608 578224 455328 578252
rect 428608 578212 428614 578224
rect 455322 578212 455328 578224
rect 455380 578212 455386 578264
rect 456058 578212 456064 578264
rect 456116 578252 456122 578264
rect 483198 578252 483204 578264
rect 456116 578224 483204 578252
rect 456116 578212 456122 578224
rect 483198 578212 483204 578224
rect 483256 578212 483262 578264
rect 485038 578212 485044 578264
rect 485096 578252 485102 578264
rect 511350 578252 511356 578264
rect 485096 578224 511356 578252
rect 485096 578212 485102 578224
rect 511350 578212 511356 578224
rect 511408 578212 511414 578264
rect 512638 578212 512644 578264
rect 512696 578252 512702 578264
rect 539318 578252 539324 578264
rect 512696 578224 539324 578252
rect 512696 578212 512702 578224
rect 539318 578212 539324 578224
rect 539376 578212 539382 578264
rect 540238 578212 540244 578264
rect 540296 578252 540302 578264
rect 567194 578252 567200 578264
rect 540296 578224 567200 578252
rect 540296 578212 540302 578224
rect 567194 578212 567200 578224
rect 567252 578212 567258 578264
rect 15286 575220 15292 575272
rect 15344 575260 15350 575272
rect 15930 575260 15936 575272
rect 15344 575232 15936 575260
rect 15344 575220 15350 575232
rect 15930 575220 15936 575232
rect 15988 575220 15994 575272
rect 42886 571208 42892 571260
rect 42944 571248 42950 571260
rect 43622 571248 43628 571260
rect 42944 571220 43628 571248
rect 42944 571208 42950 571220
rect 43622 571208 43628 571220
rect 43680 571208 43686 571260
rect 147674 562300 147680 562352
rect 147732 562340 147738 562352
rect 148410 562340 148416 562352
rect 147732 562312 148416 562340
rect 147732 562300 147738 562312
rect 148410 562300 148416 562312
rect 148468 562300 148474 562352
rect 259730 562300 259736 562352
rect 259788 562340 259794 562352
rect 260190 562340 260196 562352
rect 259788 562312 260196 562340
rect 259788 562300 259794 562312
rect 260190 562300 260196 562312
rect 260248 562300 260254 562352
rect 455690 562300 455696 562352
rect 455748 562340 455754 562352
rect 456150 562340 456156 562352
rect 455748 562312 456156 562340
rect 455748 562300 455754 562312
rect 456150 562300 456156 562312
rect 456208 562300 456214 562352
rect 287698 558832 287704 558884
rect 287756 558872 287762 558884
rect 295702 558872 295708 558884
rect 287756 558844 295708 558872
rect 287756 558832 287762 558844
rect 295702 558832 295708 558844
rect 295760 558832 295766 558884
rect 316770 558832 316776 558884
rect 316828 558872 316834 558884
rect 323670 558872 323676 558884
rect 316828 558844 323676 558872
rect 316828 558832 316834 558844
rect 323670 558832 323676 558844
rect 323728 558832 323734 558884
rect 63586 558288 63592 558340
rect 63644 558328 63650 558340
rect 64322 558328 64328 558340
rect 63644 558300 64328 558328
rect 63644 558288 63650 558300
rect 64322 558288 64328 558300
rect 64380 558288 64386 558340
rect 232682 558152 232688 558204
rect 232740 558192 232746 558204
rect 239766 558192 239772 558204
rect 232740 558164 239772 558192
rect 232740 558152 232746 558164
rect 239766 558152 239772 558164
rect 239824 558152 239830 558204
rect 428642 558152 428648 558204
rect 428700 558192 428706 558204
rect 435726 558192 435732 558204
rect 428700 558164 435732 558192
rect 428700 558152 428706 558164
rect 435726 558152 435732 558164
rect 435784 558152 435790 558204
rect 483658 558152 483664 558204
rect 483716 558192 483722 558204
rect 491662 558192 491668 558204
rect 483716 558164 491668 558192
rect 483716 558152 483722 558164
rect 491662 558152 491668 558164
rect 491720 558152 491726 558204
rect 512730 558152 512736 558204
rect 512788 558192 512794 558204
rect 519630 558192 519636 558204
rect 512788 558164 519636 558192
rect 512788 558152 512794 558164
rect 519630 558152 519636 558164
rect 519688 558152 519694 558204
rect 13538 557472 13544 557524
rect 13596 557512 13602 557524
rect 66254 557512 66260 557524
rect 13596 557484 66260 557512
rect 13596 557472 13602 557484
rect 66254 557472 66260 557484
rect 66312 557472 66318 557524
rect 70302 557472 70308 557524
rect 70360 557512 70366 557524
rect 121454 557512 121460 557524
rect 70360 557484 121460 557512
rect 70360 557472 70366 557484
rect 121454 557472 121460 557484
rect 121512 557472 121518 557524
rect 126882 557472 126888 557524
rect 126940 557512 126946 557524
rect 178034 557512 178040 557524
rect 126940 557484 178040 557512
rect 126940 557472 126946 557484
rect 178034 557472 178040 557484
rect 178092 557472 178098 557524
rect 209682 557472 209688 557524
rect 209740 557512 209746 557524
rect 262214 557512 262220 557524
rect 209740 557484 262220 557512
rect 209740 557472 209746 557484
rect 262214 557472 262220 557484
rect 262272 557472 262278 557524
rect 266262 557472 266268 557524
rect 266320 557512 266326 557524
rect 317414 557512 317420 557524
rect 266320 557484 317420 557512
rect 266320 557472 266326 557484
rect 317414 557472 317420 557484
rect 317472 557472 317478 557524
rect 322842 557472 322848 557524
rect 322900 557512 322906 557524
rect 373994 557512 374000 557524
rect 322900 557484 374000 557512
rect 322900 557472 322906 557484
rect 373994 557472 374000 557484
rect 374052 557472 374058 557524
rect 405642 557472 405648 557524
rect 405700 557512 405706 557524
rect 458174 557512 458180 557524
rect 405700 557484 458180 557512
rect 405700 557472 405706 557484
rect 458174 557472 458180 557484
rect 458232 557472 458238 557524
rect 489822 557472 489828 557524
rect 489880 557512 489886 557524
rect 542354 557512 542360 557524
rect 489880 557484 542360 557512
rect 489880 557472 489886 557484
rect 542354 557472 542360 557484
rect 542412 557472 542418 557524
rect 42702 557404 42708 557456
rect 42760 557444 42766 557456
rect 93854 557444 93860 557456
rect 42760 557416 93860 557444
rect 42760 557404 42766 557416
rect 93854 557404 93860 557416
rect 93912 557404 93918 557456
rect 97902 557404 97908 557456
rect 97960 557444 97966 557456
rect 149054 557444 149060 557456
rect 97960 557416 149060 557444
rect 97960 557404 97966 557416
rect 149054 557404 149060 557416
rect 149112 557404 149118 557456
rect 154482 557404 154488 557456
rect 154540 557444 154546 557456
rect 205634 557444 205640 557456
rect 154540 557416 205640 557444
rect 154540 557404 154546 557416
rect 205634 557404 205640 557416
rect 205692 557404 205698 557456
rect 238662 557404 238668 557456
rect 238720 557444 238726 557456
rect 289814 557444 289820 557456
rect 238720 557416 289820 557444
rect 238720 557404 238726 557416
rect 289814 557404 289820 557416
rect 289872 557404 289878 557456
rect 293862 557404 293868 557456
rect 293920 557444 293926 557456
rect 293920 557416 335354 557444
rect 293920 557404 293926 557416
rect 182082 557336 182088 557388
rect 182140 557376 182146 557388
rect 233234 557376 233240 557388
rect 182140 557348 233240 557376
rect 182140 557336 182146 557348
rect 233234 557336 233240 557348
rect 233292 557336 233298 557388
rect 335326 557376 335354 557416
rect 343542 557404 343548 557456
rect 343600 557444 343606 557456
rect 345658 557444 345664 557456
rect 343600 557416 345664 557444
rect 343600 557404 343606 557416
rect 345658 557404 345664 557416
rect 345716 557404 345722 557456
rect 378042 557404 378048 557456
rect 378100 557444 378106 557456
rect 429286 557444 429292 557456
rect 378100 557416 429292 557444
rect 378100 557404 378106 557416
rect 429286 557404 429292 557416
rect 429344 557404 429350 557456
rect 434622 557404 434628 557456
rect 434680 557444 434686 557456
rect 485774 557444 485780 557456
rect 434680 557416 485780 557444
rect 434680 557404 434686 557416
rect 485774 557404 485780 557416
rect 485832 557404 485838 557456
rect 518802 557404 518808 557456
rect 518860 557444 518866 557456
rect 569954 557444 569960 557456
rect 518860 557416 569960 557444
rect 518860 557404 518866 557416
rect 569954 557404 569960 557416
rect 570012 557404 570018 557456
rect 345014 557376 345020 557388
rect 335326 557348 345020 557376
rect 345014 557336 345020 557348
rect 345072 557336 345078 557388
rect 350442 557336 350448 557388
rect 350500 557376 350506 557388
rect 401594 557376 401600 557388
rect 350500 557348 401600 557376
rect 350500 557336 350506 557348
rect 401594 557336 401600 557348
rect 401652 557336 401658 557388
rect 462222 557336 462228 557388
rect 462280 557376 462286 557388
rect 513374 557376 513380 557388
rect 462280 557348 513380 557376
rect 462280 557336 462286 557348
rect 513374 557336 513380 557348
rect 513432 557336 513438 557388
rect 539502 556724 539508 556776
rect 539560 556764 539566 556776
rect 541618 556764 541624 556776
rect 539560 556736 541624 556764
rect 539560 556724 539566 556736
rect 541618 556724 541624 556736
rect 541676 556724 541682 556776
rect 35250 556656 35256 556708
rect 35308 556696 35314 556708
rect 36722 556696 36728 556708
rect 35308 556668 36728 556696
rect 35308 556656 35314 556668
rect 36722 556656 36728 556668
rect 36780 556656 36786 556708
rect 15838 556180 15844 556232
rect 15896 556220 15902 556232
rect 16574 556220 16580 556232
rect 15896 556192 16580 556220
rect 15896 556180 15902 556192
rect 16574 556180 16580 556192
rect 16632 556180 16638 556232
rect 547874 556112 547880 556164
rect 547932 556152 547938 556164
rect 548150 556152 548156 556164
rect 547932 556124 548156 556152
rect 547932 556112 547938 556124
rect 548150 556112 548156 556124
rect 548208 556112 548214 556164
rect 71866 554684 71872 554736
rect 71924 554724 71930 554736
rect 100018 554724 100024 554736
rect 71924 554696 100024 554724
rect 71924 554684 71930 554696
rect 100018 554684 100024 554696
rect 100076 554684 100082 554736
rect 127986 554724 127992 554736
rect 103486 554696 127992 554724
rect 25682 554616 25688 554668
rect 25740 554656 25746 554668
rect 36630 554656 36636 554668
rect 25740 554628 36636 554656
rect 25740 554616 25746 554628
rect 36630 554616 36636 554628
rect 36688 554616 36694 554668
rect 42886 554616 42892 554668
rect 42944 554656 42950 554668
rect 42944 554628 45554 554656
rect 42944 554616 42950 554628
rect 15286 554548 15292 554600
rect 15344 554588 15350 554600
rect 43990 554588 43996 554600
rect 15344 554560 43996 554588
rect 15344 554548 15350 554560
rect 43990 554548 43996 554560
rect 44048 554548 44054 554600
rect 45526 554588 45554 554628
rect 53650 554616 53656 554668
rect 53708 554656 53714 554668
rect 66898 554656 66904 554668
rect 53708 554628 66904 554656
rect 53708 554616 53714 554628
rect 66898 554616 66904 554628
rect 66956 554616 66962 554668
rect 81986 554616 81992 554668
rect 82044 554656 82050 554668
rect 93118 554656 93124 554668
rect 82044 554628 93124 554656
rect 82044 554616 82050 554628
rect 93118 554616 93124 554628
rect 93176 554616 93182 554668
rect 99466 554616 99472 554668
rect 99524 554656 99530 554668
rect 103486 554656 103514 554696
rect 127986 554684 127992 554696
rect 128044 554684 128050 554736
rect 165982 554684 165988 554736
rect 166040 554724 166046 554736
rect 177298 554724 177304 554736
rect 166040 554696 177304 554724
rect 166040 554684 166046 554696
rect 177298 554684 177304 554696
rect 177356 554684 177362 554736
rect 178678 554684 178684 554736
rect 178736 554724 178742 554736
rect 184014 554724 184020 554736
rect 178736 554696 184020 554724
rect 178736 554684 178742 554696
rect 184014 554684 184020 554696
rect 184072 554684 184078 554736
rect 211706 554724 211712 554736
rect 190426 554696 211712 554724
rect 99524 554628 103514 554656
rect 99524 554616 99530 554628
rect 109678 554616 109684 554668
rect 109736 554656 109742 554668
rect 124858 554656 124864 554668
rect 109736 554628 124864 554656
rect 109736 554616 109742 554628
rect 124858 554616 124864 554628
rect 124916 554616 124922 554668
rect 137646 554616 137652 554668
rect 137704 554656 137710 554668
rect 148318 554656 148324 554668
rect 137704 554628 148324 554656
rect 137704 554616 137710 554628
rect 148318 554616 148324 554628
rect 148376 554616 148382 554668
rect 183646 554616 183652 554668
rect 183704 554656 183710 554668
rect 190426 554656 190454 554696
rect 211706 554684 211712 554696
rect 211764 554684 211770 554736
rect 277670 554684 277676 554736
rect 277728 554724 277734 554736
rect 289078 554724 289084 554736
rect 277728 554696 289084 554724
rect 277728 554684 277734 554696
rect 289078 554684 289084 554696
rect 289136 554684 289142 554736
rect 306006 554684 306012 554736
rect 306064 554724 306070 554736
rect 316678 554724 316684 554736
rect 306064 554696 316684 554724
rect 306064 554684 306070 554696
rect 316678 554684 316684 554696
rect 316736 554684 316742 554736
rect 361666 554684 361672 554736
rect 361724 554724 361730 554736
rect 373258 554724 373264 554736
rect 361724 554696 373264 554724
rect 361724 554684 361730 554696
rect 373258 554684 373264 554696
rect 373316 554684 373322 554736
rect 374638 554684 374644 554736
rect 374696 554724 374702 554736
rect 379698 554724 379704 554736
rect 374696 554696 379704 554724
rect 374696 554684 374702 554696
rect 379698 554684 379704 554696
rect 379756 554684 379762 554736
rect 408034 554724 408040 554736
rect 383626 554696 408040 554724
rect 183704 554628 190454 554656
rect 183704 554616 183710 554628
rect 193674 554616 193680 554668
rect 193732 554656 193738 554668
rect 204990 554656 204996 554668
rect 193732 554628 204996 554656
rect 193732 554616 193738 554628
rect 204990 554616 204996 554628
rect 205048 554616 205054 554668
rect 222010 554616 222016 554668
rect 222068 554656 222074 554668
rect 232590 554656 232596 554668
rect 222068 554628 232596 554656
rect 222068 554616 222074 554628
rect 232590 554616 232596 554628
rect 232648 554616 232654 554668
rect 249702 554616 249708 554668
rect 249760 554656 249766 554668
rect 260098 554656 260104 554668
rect 249760 554628 260104 554656
rect 249760 554616 249766 554628
rect 260098 554616 260104 554628
rect 260156 554616 260162 554668
rect 333698 554616 333704 554668
rect 333756 554656 333762 554668
rect 344278 554656 344284 554668
rect 333756 554628 344284 554656
rect 333756 554616 333762 554628
rect 344278 554616 344284 554628
rect 344336 554616 344342 554668
rect 379606 554616 379612 554668
rect 379664 554656 379670 554668
rect 383626 554656 383654 554696
rect 408034 554684 408040 554696
rect 408092 554684 408098 554736
rect 473998 554684 474004 554736
rect 474056 554724 474062 554736
rect 485038 554724 485044 554736
rect 474056 554696 485044 554724
rect 474056 554684 474062 554696
rect 485038 554684 485044 554696
rect 485096 554684 485102 554736
rect 501690 554684 501696 554736
rect 501748 554724 501754 554736
rect 512638 554724 512644 554736
rect 501748 554696 512644 554724
rect 501748 554684 501754 554696
rect 512638 554684 512644 554696
rect 512696 554684 512702 554736
rect 548150 554684 548156 554736
rect 548208 554724 548214 554736
rect 557534 554724 557540 554736
rect 548208 554696 557540 554724
rect 548208 554684 548214 554696
rect 557534 554684 557540 554696
rect 557592 554684 557598 554736
rect 379664 554628 383654 554656
rect 379664 554616 379670 554628
rect 390002 554616 390008 554668
rect 390060 554656 390066 554668
rect 400858 554656 400864 554668
rect 390060 554628 400864 554656
rect 390060 554616 390066 554628
rect 400858 554616 400864 554628
rect 400916 554616 400922 554668
rect 417694 554616 417700 554668
rect 417752 554656 417758 554668
rect 428550 554656 428556 554668
rect 417752 554628 428556 554656
rect 417752 554616 417758 554628
rect 428550 554616 428556 554628
rect 428608 554616 428614 554668
rect 445662 554616 445668 554668
rect 445720 554656 445726 554668
rect 456058 554656 456064 554668
rect 445720 554628 456064 554656
rect 445720 554616 445726 554628
rect 456058 554616 456064 554628
rect 456116 554616 456122 554668
rect 529658 554616 529664 554668
rect 529716 554656 529722 554668
rect 540238 554656 540244 554668
rect 529716 554628 540244 554656
rect 529716 554616 529722 554628
rect 540238 554616 540244 554628
rect 540296 554616 540302 554668
rect 72050 554588 72056 554600
rect 45526 554560 72056 554588
rect 72050 554548 72056 554560
rect 72108 554548 72114 554600
rect 127066 554548 127072 554600
rect 127124 554588 127130 554600
rect 156046 554588 156052 554600
rect 127124 554560 156052 554588
rect 127124 554548 127130 554560
rect 156046 554548 156052 554560
rect 156104 554548 156110 554600
rect 238846 554548 238852 554600
rect 238904 554588 238910 554600
rect 268010 554588 268016 554600
rect 238904 554560 268016 554588
rect 238904 554548 238910 554560
rect 268010 554548 268016 554560
rect 268068 554548 268074 554600
rect 323026 554548 323032 554600
rect 323084 554588 323090 554600
rect 352006 554588 352012 554600
rect 323084 554560 352012 554588
rect 323084 554548 323090 554560
rect 352006 554548 352012 554560
rect 352064 554548 352070 554600
rect 434806 554548 434812 554600
rect 434864 554588 434870 554600
rect 463694 554588 463700 554600
rect 434864 554560 463700 554588
rect 434864 554548 434870 554560
rect 463694 554548 463700 554560
rect 463752 554548 463758 554600
rect 518986 554548 518992 554600
rect 519044 554588 519050 554600
rect 547874 554588 547880 554600
rect 519044 554560 547880 554588
rect 519044 554548 519050 554560
rect 547874 554548 547880 554560
rect 547932 554548 547938 554600
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 10318 553432 10324 553444
rect 3384 553404 10324 553432
rect 3384 553392 3390 553404
rect 10318 553392 10324 553404
rect 10376 553392 10382 553444
rect 26234 550876 26240 550928
rect 26292 550916 26298 550928
rect 35434 550916 35440 550928
rect 26292 550888 35440 550916
rect 26292 550876 26298 550888
rect 35434 550876 35440 550888
rect 35492 550876 35498 550928
rect 352006 550808 352012 550860
rect 352064 550848 352070 550860
rect 352064 550820 354674 550848
rect 352064 550808 352070 550820
rect 71130 550740 71136 550792
rect 71188 550780 71194 550792
rect 82262 550780 82268 550792
rect 71188 550752 82268 550780
rect 71188 550740 71194 550752
rect 82262 550740 82268 550752
rect 82320 550740 82326 550792
rect 99466 550740 99472 550792
rect 99524 550780 99530 550792
rect 100386 550780 100392 550792
rect 99524 550752 100392 550780
rect 99524 550740 99530 550752
rect 100386 550740 100392 550752
rect 100444 550740 100450 550792
rect 183646 550740 183652 550792
rect 183704 550780 183710 550792
rect 222286 550780 222292 550792
rect 183704 550752 222292 550780
rect 183704 550740 183710 550752
rect 222286 550740 222292 550752
rect 222344 550740 222350 550792
rect 267826 550740 267832 550792
rect 267884 550780 267890 550792
rect 267884 550752 277394 550780
rect 267884 550740 267890 550752
rect 36630 550672 36636 550724
rect 36688 550712 36694 550724
rect 53926 550712 53932 550724
rect 36688 550684 53932 550712
rect 36688 550672 36694 550684
rect 53926 550672 53932 550684
rect 53984 550672 53990 550724
rect 71866 550672 71872 550724
rect 71924 550712 71930 550724
rect 109954 550712 109960 550724
rect 71924 550684 109960 550712
rect 71924 550672 71930 550684
rect 109954 550672 109960 550684
rect 110012 550672 110018 550724
rect 151078 550672 151084 550724
rect 151136 550712 151142 550724
rect 156598 550712 156604 550724
rect 151136 550684 156604 550712
rect 151136 550672 151142 550684
rect 156598 550672 156604 550684
rect 156656 550672 156662 550724
rect 182818 550672 182824 550724
rect 182876 550712 182882 550724
rect 193950 550712 193956 550724
rect 182876 550684 193956 550712
rect 182876 550672 182882 550684
rect 193950 550672 193956 550684
rect 194008 550672 194014 550724
rect 232498 550672 232504 550724
rect 232556 550712 232562 550724
rect 232556 550684 248414 550712
rect 232556 550672 232562 550684
rect 66898 550604 66904 550656
rect 66956 550644 66962 550656
rect 72602 550644 72608 550656
rect 66956 550616 72608 550644
rect 66956 550604 66962 550616
rect 72602 550604 72608 550616
rect 72660 550604 72666 550656
rect 93118 550604 93124 550656
rect 93176 550644 93182 550656
rect 100294 550644 100300 550656
rect 93176 550616 100300 550644
rect 93176 550604 93182 550616
rect 100294 550604 100300 550616
rect 100352 550604 100358 550656
rect 100386 550604 100392 550656
rect 100444 550644 100450 550656
rect 138290 550644 138296 550656
rect 100444 550616 138296 550644
rect 100444 550604 100450 550616
rect 138290 550604 138296 550616
rect 138348 550604 138354 550656
rect 149698 550604 149704 550656
rect 149756 550644 149762 550656
rect 166258 550644 166264 550656
rect 149756 550616 166264 550644
rect 149756 550604 149762 550616
rect 166258 550604 166264 550616
rect 166316 550604 166322 550656
rect 177298 550604 177304 550656
rect 177356 550644 177362 550656
rect 184290 550644 184296 550656
rect 177356 550616 184296 550644
rect 177356 550604 177362 550616
rect 184290 550604 184296 550616
rect 184348 550604 184354 550656
rect 233970 550604 233976 550656
rect 234028 550644 234034 550656
rect 240594 550644 240600 550656
rect 234028 550616 240600 550644
rect 234028 550604 234034 550616
rect 240594 550604 240600 550616
rect 240652 550604 240658 550656
rect 248386 550644 248414 550684
rect 266998 550672 267004 550724
rect 267056 550712 267062 550724
rect 277366 550712 277394 550752
rect 295426 550740 295432 550792
rect 295484 550780 295490 550792
rect 334250 550780 334256 550792
rect 295484 550752 334256 550780
rect 295484 550740 295490 550752
rect 334250 550740 334256 550752
rect 334308 550740 334314 550792
rect 345658 550740 345664 550792
rect 345716 550780 345722 550792
rect 345716 550752 352512 550780
rect 345716 550740 345722 550752
rect 306282 550712 306288 550724
rect 267056 550684 268976 550712
rect 277366 550684 306288 550712
rect 267056 550672 267062 550684
rect 250254 550644 250260 550656
rect 248386 550616 250260 550644
rect 250254 550604 250260 550616
rect 250312 550604 250318 550656
rect 261478 550604 261484 550656
rect 261536 550644 261542 550656
rect 268286 550644 268292 550656
rect 261536 550616 268292 550644
rect 261536 550604 261542 550616
rect 268286 550604 268292 550616
rect 268344 550604 268350 550656
rect 268948 550644 268976 550684
rect 306282 550672 306288 550684
rect 306340 550672 306346 550724
rect 277946 550644 277952 550656
rect 268948 550616 277952 550644
rect 277946 550604 277952 550616
rect 278004 550604 278010 550656
rect 289078 550604 289084 550656
rect 289136 550644 289142 550656
rect 296622 550644 296628 550656
rect 289136 550616 296628 550644
rect 289136 550604 289142 550616
rect 296622 550604 296628 550616
rect 296680 550604 296686 550656
rect 318058 550604 318064 550656
rect 318116 550644 318122 550656
rect 324590 550644 324596 550656
rect 318116 550616 324596 550644
rect 318116 550604 318122 550616
rect 324590 550604 324596 550616
rect 324648 550604 324654 550656
rect 347038 550604 347044 550656
rect 347096 550644 347102 550656
rect 352282 550644 352288 550656
rect 347096 550616 352288 550644
rect 347096 550604 347102 550616
rect 352282 550604 352288 550616
rect 352340 550604 352346 550656
rect 352484 550644 352512 550752
rect 354646 550712 354674 550820
rect 463786 550808 463792 550860
rect 463844 550848 463850 550860
rect 463844 550820 470594 550848
rect 463844 550808 463850 550820
rect 379606 550740 379612 550792
rect 379664 550780 379670 550792
rect 418246 550780 418252 550792
rect 379664 550752 418252 550780
rect 379664 550740 379670 550752
rect 418246 550740 418252 550752
rect 418304 550740 418310 550792
rect 390278 550712 390284 550724
rect 354646 550684 390284 550712
rect 390278 550672 390284 550684
rect 390336 550672 390342 550724
rect 400950 550672 400956 550724
rect 401008 550712 401014 550724
rect 408586 550712 408592 550724
rect 401008 550684 408592 550712
rect 401008 550672 401014 550684
rect 408586 550672 408592 550684
rect 408644 550672 408650 550724
rect 429838 550672 429844 550724
rect 429896 550712 429902 550724
rect 436278 550712 436284 550724
rect 429896 550684 436284 550712
rect 429896 550672 429902 550684
rect 436278 550672 436284 550684
rect 436336 550672 436342 550724
rect 457438 550672 457444 550724
rect 457496 550712 457502 550724
rect 464614 550712 464620 550724
rect 457496 550684 464620 550712
rect 457496 550672 457502 550684
rect 464614 550672 464620 550684
rect 464672 550672 464678 550724
rect 470566 550712 470594 550820
rect 489886 550820 499574 550848
rect 489886 550712 489914 550820
rect 491386 550740 491392 550792
rect 491444 550780 491450 550792
rect 491444 550752 492812 550780
rect 491444 550740 491450 550752
rect 470566 550684 489914 550712
rect 361942 550644 361948 550656
rect 352484 550616 361948 550644
rect 361942 550604 361948 550616
rect 362000 550604 362006 550656
rect 373258 550604 373264 550656
rect 373316 550644 373322 550656
rect 380618 550644 380624 550656
rect 373316 550616 380624 550644
rect 373316 550604 373322 550616
rect 380618 550604 380624 550616
rect 380676 550604 380682 550656
rect 428458 550604 428464 550656
rect 428516 550644 428522 550656
rect 445938 550644 445944 550656
rect 428516 550616 445944 550644
rect 428516 550604 428522 550616
rect 445938 550604 445944 550616
rect 445996 550604 446002 550656
rect 462958 550604 462964 550656
rect 463016 550644 463022 550656
rect 474274 550644 474280 550656
rect 463016 550616 474280 550644
rect 463016 550604 463022 550616
rect 474274 550604 474280 550616
rect 474332 550604 474338 550656
rect 485038 550604 485044 550656
rect 485096 550644 485102 550656
rect 492582 550644 492588 550656
rect 485096 550616 492588 550644
rect 485096 550604 485102 550616
rect 492582 550604 492588 550616
rect 492640 550604 492646 550656
rect 492784 550644 492812 550752
rect 499546 550712 499574 550820
rect 529934 550780 529940 550792
rect 509206 550752 529940 550780
rect 502242 550712 502248 550724
rect 499546 550684 502248 550712
rect 502242 550672 502248 550684
rect 502300 550672 502306 550724
rect 509206 550644 509234 550752
rect 529934 550740 529940 550752
rect 529992 550740 529998 550792
rect 541618 550672 541624 550724
rect 541676 550712 541682 550724
rect 541676 550684 557534 550712
rect 541676 550672 541682 550684
rect 492784 550616 509234 550644
rect 514018 550604 514024 550656
rect 514076 550644 514082 550656
rect 520274 550644 520280 550656
rect 514076 550616 518894 550644
rect 514076 550604 514082 550616
rect 518866 550576 518894 550616
rect 519096 550616 520280 550644
rect 519096 550576 519124 550616
rect 520274 550604 520280 550616
rect 520332 550604 520338 550656
rect 544378 550604 544384 550656
rect 544436 550644 544442 550656
rect 548610 550644 548616 550656
rect 544436 550616 548616 550644
rect 544436 550604 544442 550616
rect 548610 550604 548616 550616
rect 548668 550604 548674 550656
rect 557506 550644 557534 550684
rect 558270 550644 558276 550656
rect 557506 550616 558276 550644
rect 558270 550604 558276 550616
rect 558328 550604 558334 550656
rect 518866 550548 519124 550576
rect 120074 548224 120080 548276
rect 120132 548264 120138 548276
rect 122098 548264 122104 548276
rect 120132 548236 122104 548264
rect 120132 548224 120138 548236
rect 122098 548224 122104 548236
rect 122156 548224 122162 548276
rect 124858 548224 124864 548276
rect 124916 548264 124922 548276
rect 128262 548264 128268 548276
rect 124916 548236 128268 548264
rect 124916 548224 124922 548236
rect 128262 548224 128268 548236
rect 128320 548224 128326 548276
rect 210418 548224 210424 548276
rect 210476 548264 210482 548276
rect 212350 548264 212356 548276
rect 210476 548236 212356 548264
rect 210476 548224 210482 548236
rect 212350 548224 212356 548236
rect 212408 548224 212414 548276
rect 204254 547068 204260 547120
rect 204312 547108 204318 547120
rect 204990 547108 204996 547120
rect 204312 547080 204996 547108
rect 204312 547068 204318 547080
rect 204990 547068 204996 547080
rect 205048 547068 205054 547120
rect 13538 529864 13544 529916
rect 13596 529904 13602 529916
rect 66254 529904 66260 529916
rect 13596 529876 66260 529904
rect 13596 529864 13602 529876
rect 66254 529864 66260 529876
rect 66312 529864 66318 529916
rect 70302 529864 70308 529916
rect 70360 529904 70366 529916
rect 121454 529904 121460 529916
rect 70360 529876 121460 529904
rect 70360 529864 70366 529876
rect 121454 529864 121460 529876
rect 121512 529864 121518 529916
rect 126882 529864 126888 529916
rect 126940 529904 126946 529916
rect 178034 529904 178040 529916
rect 126940 529876 178040 529904
rect 126940 529864 126946 529876
rect 178034 529864 178040 529876
rect 178092 529864 178098 529916
rect 209682 529864 209688 529916
rect 209740 529904 209746 529916
rect 262214 529904 262220 529916
rect 209740 529876 262220 529904
rect 209740 529864 209746 529876
rect 262214 529864 262220 529876
rect 262272 529864 262278 529916
rect 266262 529864 266268 529916
rect 266320 529904 266326 529916
rect 317414 529904 317420 529916
rect 266320 529876 317420 529904
rect 266320 529864 266326 529876
rect 317414 529864 317420 529876
rect 317472 529864 317478 529916
rect 322842 529864 322848 529916
rect 322900 529904 322906 529916
rect 373994 529904 374000 529916
rect 322900 529876 374000 529904
rect 322900 529864 322906 529876
rect 373994 529864 374000 529876
rect 374052 529864 374058 529916
rect 405642 529864 405648 529916
rect 405700 529904 405706 529916
rect 458174 529904 458180 529916
rect 405700 529876 458180 529904
rect 405700 529864 405706 529876
rect 458174 529864 458180 529876
rect 458232 529864 458238 529916
rect 489822 529864 489828 529916
rect 489880 529904 489886 529916
rect 542354 529904 542360 529916
rect 489880 529876 542360 529904
rect 489880 529864 489886 529876
rect 542354 529864 542360 529876
rect 542412 529864 542418 529916
rect 42702 529796 42708 529848
rect 42760 529836 42766 529848
rect 93854 529836 93860 529848
rect 42760 529808 93860 529836
rect 42760 529796 42766 529808
rect 93854 529796 93860 529808
rect 93912 529796 93918 529848
rect 97902 529796 97908 529848
rect 97960 529836 97966 529848
rect 149054 529836 149060 529848
rect 97960 529808 149060 529836
rect 97960 529796 97966 529808
rect 149054 529796 149060 529808
rect 149112 529796 149118 529848
rect 154482 529796 154488 529848
rect 154540 529836 154546 529848
rect 205634 529836 205640 529848
rect 154540 529808 205640 529836
rect 154540 529796 154546 529808
rect 205634 529796 205640 529808
rect 205692 529796 205698 529848
rect 238662 529796 238668 529848
rect 238720 529836 238726 529848
rect 289814 529836 289820 529848
rect 238720 529808 289820 529836
rect 238720 529796 238726 529808
rect 289814 529796 289820 529808
rect 289872 529796 289878 529848
rect 293862 529796 293868 529848
rect 293920 529836 293926 529848
rect 345014 529836 345020 529848
rect 293920 529808 345020 529836
rect 293920 529796 293926 529808
rect 345014 529796 345020 529808
rect 345072 529796 345078 529848
rect 378042 529796 378048 529848
rect 378100 529836 378106 529848
rect 429286 529836 429292 529848
rect 378100 529808 429292 529836
rect 378100 529796 378106 529808
rect 429286 529796 429292 529808
rect 429344 529796 429350 529848
rect 434622 529796 434628 529848
rect 434680 529836 434686 529848
rect 485774 529836 485780 529848
rect 434680 529808 485780 529836
rect 434680 529796 434686 529808
rect 485774 529796 485780 529808
rect 485832 529796 485838 529848
rect 518802 529796 518808 529848
rect 518860 529836 518866 529848
rect 569954 529836 569960 529848
rect 518860 529808 569960 529836
rect 518860 529796 518866 529808
rect 569954 529796 569960 529808
rect 570012 529796 570018 529848
rect 182082 529728 182088 529780
rect 182140 529768 182146 529780
rect 233234 529768 233240 529780
rect 182140 529740 233240 529768
rect 182140 529728 182146 529740
rect 233234 529728 233240 529740
rect 233292 529728 233298 529780
rect 350442 529728 350448 529780
rect 350500 529768 350506 529780
rect 401594 529768 401600 529780
rect 350500 529740 401600 529768
rect 350500 529728 350506 529740
rect 401594 529728 401600 529740
rect 401652 529728 401658 529780
rect 462222 529728 462228 529780
rect 462280 529768 462286 529780
rect 513374 529768 513380 529780
rect 462280 529740 513380 529768
rect 462280 529728 462286 529740
rect 513374 529728 513380 529740
rect 513432 529728 513438 529780
rect 2774 527144 2780 527196
rect 2832 527184 2838 527196
rect 4798 527184 4804 527196
rect 2832 527156 4804 527184
rect 2832 527144 2838 527156
rect 4798 527144 4804 527156
rect 4856 527144 4862 527196
rect 15194 527076 15200 527128
rect 15252 527116 15258 527128
rect 35894 527116 35900 527128
rect 15252 527088 35900 527116
rect 15252 527076 15258 527088
rect 35894 527076 35900 527088
rect 35952 527076 35958 527128
rect 36078 527076 36084 527128
rect 36136 527116 36142 527128
rect 63586 527116 63592 527128
rect 36136 527088 63592 527116
rect 36136 527076 36142 527088
rect 63586 527076 63592 527088
rect 63644 527076 63650 527128
rect 64046 527076 64052 527128
rect 64104 527116 64110 527128
rect 91922 527116 91928 527128
rect 64104 527088 91928 527116
rect 64104 527076 64110 527088
rect 91922 527076 91928 527088
rect 91980 527076 91986 527128
rect 92106 527076 92112 527128
rect 92164 527116 92170 527128
rect 119614 527116 119620 527128
rect 92164 527088 119620 527116
rect 92164 527076 92170 527088
rect 119614 527076 119620 527088
rect 119672 527076 119678 527128
rect 122098 527076 122104 527128
rect 122156 527116 122162 527128
rect 147950 527116 147956 527128
rect 122156 527088 147956 527116
rect 122156 527076 122162 527088
rect 147950 527076 147956 527088
rect 148008 527076 148014 527128
rect 148042 527076 148048 527128
rect 148100 527116 148106 527128
rect 175918 527116 175924 527128
rect 148100 527088 175924 527116
rect 148100 527076 148106 527088
rect 175918 527076 175924 527088
rect 175976 527076 175982 527128
rect 176102 527076 176108 527128
rect 176160 527116 176166 527128
rect 203610 527116 203616 527128
rect 176160 527088 203616 527116
rect 176160 527076 176166 527088
rect 203610 527076 203616 527088
rect 203668 527076 203674 527128
rect 204990 527076 204996 527128
rect 205048 527116 205054 527128
rect 231946 527116 231952 527128
rect 205048 527088 231952 527116
rect 205048 527076 205054 527088
rect 231946 527076 231952 527088
rect 232004 527076 232010 527128
rect 232038 527076 232044 527128
rect 232096 527116 232102 527128
rect 259914 527116 259920 527128
rect 232096 527088 259920 527116
rect 232096 527076 232102 527088
rect 259914 527076 259920 527088
rect 259972 527076 259978 527128
rect 260098 527076 260104 527128
rect 260156 527116 260162 527128
rect 287606 527116 287612 527128
rect 260156 527088 287612 527116
rect 260156 527076 260162 527088
rect 287606 527076 287612 527088
rect 287664 527076 287670 527128
rect 288066 527076 288072 527128
rect 288124 527116 288130 527128
rect 315942 527116 315948 527128
rect 288124 527088 315948 527116
rect 288124 527076 288130 527088
rect 315942 527076 315948 527088
rect 316000 527076 316006 527128
rect 316678 527076 316684 527128
rect 316736 527116 316742 527128
rect 343910 527116 343916 527128
rect 316736 527088 343916 527116
rect 316736 527076 316742 527088
rect 343910 527076 343916 527088
rect 343968 527076 343974 527128
rect 344094 527076 344100 527128
rect 344152 527116 344158 527128
rect 371602 527116 371608 527128
rect 344152 527088 371608 527116
rect 344152 527076 344158 527088
rect 371602 527076 371608 527088
rect 371660 527076 371666 527128
rect 372062 527076 372068 527128
rect 372120 527116 372126 527128
rect 399938 527116 399944 527128
rect 372120 527088 399944 527116
rect 372120 527076 372126 527088
rect 399938 527076 399944 527088
rect 399996 527076 400002 527128
rect 400858 527076 400864 527128
rect 400916 527116 400922 527128
rect 427906 527116 427912 527128
rect 400916 527088 427912 527116
rect 400916 527076 400922 527088
rect 427906 527076 427912 527088
rect 427964 527076 427970 527128
rect 428090 527076 428096 527128
rect 428148 527116 428154 527128
rect 455598 527116 455604 527128
rect 428148 527088 455604 527116
rect 428148 527076 428154 527088
rect 455598 527076 455604 527088
rect 455656 527076 455662 527128
rect 456058 527076 456064 527128
rect 456116 527116 456122 527128
rect 483934 527116 483940 527128
rect 456116 527088 483940 527116
rect 456116 527076 456122 527088
rect 483934 527076 483940 527088
rect 483992 527076 483998 527128
rect 484026 527076 484032 527128
rect 484084 527116 484090 527128
rect 511902 527116 511908 527128
rect 484084 527088 511908 527116
rect 484084 527076 484090 527088
rect 511902 527076 511908 527088
rect 511960 527076 511966 527128
rect 512086 527076 512092 527128
rect 512144 527116 512150 527128
rect 539594 527116 539600 527128
rect 512144 527088 539600 527116
rect 512144 527076 512150 527088
rect 539594 527076 539600 527088
rect 539652 527076 539658 527128
rect 540054 527076 540060 527128
rect 540112 527116 540118 527128
rect 567930 527116 567936 527128
rect 540112 527088 567936 527116
rect 540112 527076 540118 527088
rect 567930 527076 567936 527088
rect 567988 527076 567994 527128
rect 16574 527008 16580 527060
rect 16632 527048 16638 527060
rect 36630 527048 36636 527060
rect 16632 527020 36636 527048
rect 16632 527008 16638 527020
rect 36630 527008 36636 527020
rect 36688 527008 36694 527060
rect 44910 527008 44916 527060
rect 44968 527048 44974 527060
rect 71130 527048 71136 527060
rect 44968 527020 71136 527048
rect 44968 527008 44974 527020
rect 71130 527008 71136 527020
rect 71188 527008 71194 527060
rect 82262 527008 82268 527060
rect 82320 527048 82326 527060
rect 93118 527048 93124 527060
rect 82320 527020 93124 527048
rect 82320 527008 82326 527020
rect 93118 527008 93124 527020
rect 93176 527008 93182 527060
rect 110322 527008 110328 527060
rect 110380 527048 110386 527060
rect 124858 527048 124864 527060
rect 110380 527020 124864 527048
rect 110380 527008 110386 527020
rect 124858 527008 124864 527020
rect 124916 527008 124922 527060
rect 128630 527008 128636 527060
rect 128688 527048 128694 527060
rect 149698 527048 149704 527060
rect 128688 527020 149704 527048
rect 128688 527008 128694 527020
rect 149698 527008 149704 527020
rect 149756 527008 149762 527060
rect 156598 527008 156604 527060
rect 156656 527048 156662 527060
rect 182818 527048 182824 527060
rect 156656 527020 182824 527048
rect 156656 527008 156662 527020
rect 182818 527008 182824 527020
rect 182876 527008 182882 527060
rect 194502 527008 194508 527060
rect 194560 527048 194566 527060
rect 210418 527048 210424 527060
rect 194560 527020 210424 527048
rect 194560 527008 194566 527020
rect 210418 527008 210424 527020
rect 210476 527008 210482 527060
rect 212626 527008 212632 527060
rect 212684 527048 212690 527060
rect 232498 527048 232504 527060
rect 212684 527020 232504 527048
rect 212684 527008 212690 527020
rect 232498 527008 232504 527020
rect 232556 527008 232562 527060
rect 240594 527008 240600 527060
rect 240652 527048 240658 527060
rect 266998 527048 267004 527060
rect 240652 527020 267004 527048
rect 240652 527008 240658 527020
rect 266998 527008 267004 527020
rect 267056 527008 267062 527060
rect 278590 527008 278596 527060
rect 278648 527048 278654 527060
rect 289078 527048 289084 527060
rect 278648 527020 289084 527048
rect 278648 527008 278654 527020
rect 289078 527008 289084 527020
rect 289136 527008 289142 527060
rect 306282 527008 306288 527060
rect 306340 527048 306346 527060
rect 318058 527048 318064 527060
rect 306340 527020 318064 527048
rect 306340 527008 306346 527020
rect 318058 527008 318064 527020
rect 318116 527008 318122 527060
rect 324590 527008 324596 527060
rect 324648 527048 324654 527060
rect 345658 527048 345664 527060
rect 324648 527020 345664 527048
rect 324648 527008 324654 527020
rect 345658 527008 345664 527020
rect 345716 527008 345722 527060
rect 362586 527008 362592 527060
rect 362644 527048 362650 527060
rect 373258 527048 373264 527060
rect 362644 527020 373264 527048
rect 362644 527008 362650 527020
rect 373258 527008 373264 527020
rect 373316 527008 373322 527060
rect 390278 527008 390284 527060
rect 390336 527048 390342 527060
rect 400950 527048 400956 527060
rect 390336 527020 400956 527048
rect 390336 527008 390342 527020
rect 400950 527008 400956 527020
rect 401008 527008 401014 527060
rect 408586 527008 408592 527060
rect 408644 527048 408650 527060
rect 428458 527048 428464 527060
rect 408644 527020 428464 527048
rect 408644 527008 408650 527020
rect 428458 527008 428464 527020
rect 428516 527008 428522 527060
rect 436922 527008 436928 527060
rect 436980 527048 436986 527060
rect 462958 527048 462964 527060
rect 436980 527020 462964 527048
rect 436980 527008 436986 527020
rect 462958 527008 462964 527020
rect 463016 527008 463022 527060
rect 474274 527008 474280 527060
rect 474332 527048 474338 527060
rect 485038 527048 485044 527060
rect 474332 527020 485044 527048
rect 474332 527008 474338 527020
rect 485038 527008 485044 527020
rect 485096 527008 485102 527060
rect 502242 527008 502248 527060
rect 502300 527048 502306 527060
rect 514018 527048 514024 527060
rect 502300 527020 514024 527048
rect 502300 527008 502306 527020
rect 514018 527008 514024 527020
rect 514076 527008 514082 527060
rect 520918 527008 520924 527060
rect 520976 527048 520982 527060
rect 541618 527048 541624 527060
rect 520976 527020 541624 527048
rect 520976 527008 520982 527020
rect 541618 527008 541624 527020
rect 541676 527008 541682 527060
rect 26234 526940 26240 526992
rect 26292 526980 26298 526992
rect 43530 526980 43536 526992
rect 26292 526952 43536 526980
rect 26292 526940 26298 526952
rect 43530 526940 43536 526952
rect 43588 526940 43594 526992
rect 54570 526940 54576 526992
rect 54628 526980 54634 526992
rect 66898 526980 66904 526992
rect 54628 526952 66904 526980
rect 54628 526940 54634 526952
rect 66898 526940 66904 526952
rect 66956 526940 66962 526992
rect 138290 526940 138296 526992
rect 138348 526980 138354 526992
rect 151078 526980 151084 526992
rect 138348 526952 151084 526980
rect 138348 526940 138354 526952
rect 151078 526940 151084 526952
rect 151136 526940 151142 526992
rect 166258 526940 166264 526992
rect 166316 526980 166322 526992
rect 177298 526980 177304 526992
rect 166316 526952 177304 526980
rect 166316 526940 166322 526952
rect 177298 526940 177304 526952
rect 177356 526940 177362 526992
rect 222286 526940 222292 526992
rect 222344 526980 222350 526992
rect 233970 526980 233976 526992
rect 222344 526952 233976 526980
rect 222344 526940 222350 526952
rect 233970 526940 233976 526952
rect 234028 526940 234034 526992
rect 250254 526940 250260 526992
rect 250312 526980 250318 526992
rect 261478 526980 261484 526992
rect 250312 526952 261484 526980
rect 250312 526940 250318 526952
rect 261478 526940 261484 526952
rect 261536 526940 261542 526992
rect 334250 526940 334256 526992
rect 334308 526980 334314 526992
rect 347038 526980 347044 526992
rect 334308 526952 347044 526980
rect 334308 526940 334314 526952
rect 347038 526940 347044 526952
rect 347096 526940 347102 526992
rect 418246 526940 418252 526992
rect 418304 526980 418310 526992
rect 429838 526980 429844 526992
rect 418304 526952 429844 526980
rect 418304 526940 418310 526952
rect 429838 526940 429844 526952
rect 429896 526940 429902 526992
rect 446582 526940 446588 526992
rect 446640 526980 446646 526992
rect 457438 526980 457444 526992
rect 446640 526952 457444 526980
rect 446640 526940 446646 526952
rect 457438 526940 457444 526952
rect 457496 526940 457502 526992
rect 530578 526940 530584 526992
rect 530636 526980 530642 526992
rect 544378 526980 544384 526992
rect 530636 526952 544384 526980
rect 530636 526940 530642 526952
rect 544378 526940 544384 526952
rect 544436 526940 544442 526992
rect 558270 526396 558276 526448
rect 558328 526436 558334 526448
rect 567470 526436 567476 526448
rect 558328 526408 567476 526436
rect 558328 526396 558334 526408
rect 567470 526396 567476 526408
rect 567528 526396 567534 526448
rect 548334 523676 548340 523728
rect 548392 523716 548398 523728
rect 568022 523716 568028 523728
rect 548392 523688 568028 523716
rect 548392 523676 548398 523688
rect 568022 523676 568028 523688
rect 568080 523676 568086 523728
rect 212350 523200 212356 523252
rect 212408 523240 212414 523252
rect 232682 523240 232688 523252
rect 212408 523212 232688 523240
rect 212408 523200 212414 523212
rect 232682 523200 232688 523212
rect 232740 523200 232746 523252
rect 296346 523200 296352 523252
rect 296404 523240 296410 523252
rect 316770 523240 316776 523252
rect 296404 523212 316776 523240
rect 296404 523200 296410 523212
rect 316770 523200 316776 523212
rect 316828 523200 316834 523252
rect 408034 523200 408040 523252
rect 408092 523240 408098 523252
rect 428642 523240 428648 523252
rect 408092 523212 428648 523240
rect 408092 523200 408098 523212
rect 428642 523200 428648 523212
rect 428700 523200 428706 523252
rect 492030 523200 492036 523252
rect 492088 523240 492094 523252
rect 512730 523240 512736 523252
rect 492088 523212 512736 523240
rect 492088 523200 492094 523212
rect 512730 523200 512736 523212
rect 512788 523200 512794 523252
rect 148410 523132 148416 523184
rect 148468 523172 148474 523184
rect 165706 523172 165712 523184
rect 148468 523144 165712 523172
rect 148468 523132 148474 523144
rect 165706 523132 165712 523144
rect 165764 523132 165770 523184
rect 175458 523132 175464 523184
rect 175516 523172 175522 523184
rect 193674 523172 193680 523184
rect 175516 523144 193680 523172
rect 175516 523132 175522 523144
rect 193674 523132 193680 523144
rect 193732 523132 193738 523184
rect 203518 523132 203524 523184
rect 203576 523172 203582 523184
rect 221366 523172 221372 523184
rect 203576 523144 221372 523172
rect 203576 523132 203582 523144
rect 221366 523132 221372 523144
rect 221424 523132 221430 523184
rect 260190 523132 260196 523184
rect 260248 523172 260254 523184
rect 277670 523172 277676 523184
rect 260248 523144 277676 523172
rect 260248 523132 260254 523144
rect 277670 523132 277676 523144
rect 277728 523132 277734 523184
rect 287514 523132 287520 523184
rect 287572 523172 287578 523184
rect 305362 523172 305368 523184
rect 287572 523144 305368 523172
rect 287572 523132 287578 523144
rect 305362 523132 305368 523144
rect 305420 523132 305426 523184
rect 345658 523132 345664 523184
rect 345716 523172 345722 523184
rect 361666 523172 361672 523184
rect 345716 523144 361672 523172
rect 345716 523132 345722 523144
rect 361666 523132 361672 523144
rect 361724 523132 361730 523184
rect 371510 523132 371516 523184
rect 371568 523172 371574 523184
rect 389358 523172 389364 523184
rect 371568 523144 389364 523172
rect 371568 523132 371574 523144
rect 389358 523132 389364 523144
rect 389416 523132 389422 523184
rect 399478 523132 399484 523184
rect 399536 523172 399542 523184
rect 417694 523172 417700 523184
rect 399536 523144 417700 523172
rect 399536 523132 399542 523144
rect 417694 523132 417700 523144
rect 417752 523132 417758 523184
rect 456150 523132 456156 523184
rect 456208 523172 456214 523184
rect 473354 523172 473360 523184
rect 456208 523144 473360 523172
rect 456208 523132 456214 523144
rect 473354 523132 473360 523144
rect 473412 523132 473418 523184
rect 483474 523132 483480 523184
rect 483532 523172 483538 523184
rect 501690 523172 501696 523184
rect 483532 523144 501696 523172
rect 483532 523132 483538 523144
rect 501690 523132 501696 523144
rect 501748 523132 501754 523184
rect 36630 523064 36636 523116
rect 36688 523104 36694 523116
rect 53650 523104 53656 523116
rect 36688 523076 53656 523104
rect 36688 523064 36694 523076
rect 53650 523064 53656 523076
rect 53708 523064 53714 523116
rect 64322 523064 64328 523116
rect 64380 523104 64386 523116
rect 81434 523104 81440 523116
rect 64380 523076 81440 523104
rect 64380 523064 64386 523076
rect 81434 523064 81440 523076
rect 81492 523064 81498 523116
rect 91462 523064 91468 523116
rect 91520 523104 91526 523116
rect 109678 523104 109684 523116
rect 91520 523076 109684 523104
rect 91520 523064 91526 523076
rect 109678 523064 109684 523076
rect 109736 523064 109742 523116
rect 119430 523064 119436 523116
rect 119488 523104 119494 523116
rect 137646 523104 137652 523116
rect 119488 523076 137652 523104
rect 119488 523064 119494 523076
rect 137646 523064 137652 523076
rect 137704 523064 137710 523116
rect 156322 523064 156328 523116
rect 156380 523104 156386 523116
rect 178678 523104 178684 523116
rect 156380 523076 178684 523104
rect 156380 523064 156386 523076
rect 178678 523064 178684 523076
rect 178736 523064 178742 523116
rect 232498 523064 232504 523116
rect 232556 523104 232562 523116
rect 249702 523104 249708 523116
rect 232556 523076 249708 523104
rect 232556 523064 232562 523076
rect 249702 523064 249708 523076
rect 249760 523064 249766 523116
rect 268010 523064 268016 523116
rect 268068 523104 268074 523116
rect 287698 523104 287704 523116
rect 268068 523076 287704 523104
rect 268068 523064 268074 523076
rect 287698 523064 287704 523076
rect 287756 523064 287762 523116
rect 315482 523064 315488 523116
rect 315540 523104 315546 523116
rect 333698 523104 333704 523116
rect 315540 523076 333704 523104
rect 315540 523064 315546 523076
rect 333698 523064 333704 523076
rect 333756 523064 333762 523116
rect 352006 523064 352012 523116
rect 352064 523104 352070 523116
rect 374638 523104 374644 523116
rect 352064 523076 374644 523104
rect 352064 523064 352070 523076
rect 374638 523064 374644 523076
rect 374696 523064 374702 523116
rect 428458 523064 428464 523116
rect 428516 523104 428522 523116
rect 445662 523104 445668 523116
rect 428516 523076 445668 523104
rect 428516 523064 428522 523076
rect 445662 523064 445668 523076
rect 445720 523064 445726 523116
rect 464338 523064 464344 523116
rect 464396 523104 464402 523116
rect 483658 523104 483664 523116
rect 464396 523076 483664 523104
rect 464396 523064 464402 523076
rect 483658 523064 483664 523076
rect 483716 523064 483722 523116
rect 511442 523064 511448 523116
rect 511500 523104 511506 523116
rect 529658 523104 529664 523116
rect 511500 523076 529664 523104
rect 511500 523064 511506 523076
rect 529658 523064 529664 523076
rect 529716 523064 529722 523116
rect 541618 523064 541624 523116
rect 541676 523104 541682 523116
rect 557534 523104 557540 523116
rect 541676 523076 557540 523104
rect 541676 523064 541682 523076
rect 557534 523064 557540 523076
rect 557592 523064 557598 523116
rect 15102 522996 15108 523048
rect 15160 523036 15166 523048
rect 25682 523036 25688 523048
rect 15160 523008 25688 523036
rect 15160 522996 15166 523008
rect 25682 522996 25688 523008
rect 25740 522996 25746 523048
rect 36722 522996 36728 523048
rect 36780 523036 36786 523048
rect 63310 523036 63316 523048
rect 36780 523008 63316 523036
rect 36780 522996 36786 523008
rect 63310 522996 63316 523008
rect 63368 522996 63374 523048
rect 66898 522996 66904 523048
rect 66956 523036 66962 523048
rect 91094 523036 91100 523048
rect 66956 523008 91100 523036
rect 66956 522996 66962 523008
rect 91094 522996 91100 523008
rect 91152 522996 91158 523048
rect 93118 522996 93124 523048
rect 93176 523036 93182 523048
rect 119338 523036 119344 523048
rect 93176 523008 119344 523036
rect 93176 522996 93182 523008
rect 119338 522996 119344 523008
rect 119396 522996 119402 523048
rect 124858 522996 124864 523048
rect 124916 523036 124922 523048
rect 147306 523036 147312 523048
rect 124916 523008 147312 523036
rect 124916 522996 124922 523008
rect 147306 522996 147312 523008
rect 147364 522996 147370 523048
rect 148318 522996 148324 523048
rect 148376 523036 148382 523048
rect 175366 523036 175372 523048
rect 148376 523008 175372 523036
rect 148376 522996 148382 523008
rect 175366 522996 175372 523008
rect 175424 522996 175430 523048
rect 177298 522996 177304 523048
rect 177356 523036 177362 523048
rect 203334 523036 203340 523048
rect 177356 523008 203340 523036
rect 177356 522996 177362 523008
rect 203334 522996 203340 523008
rect 203392 522996 203398 523048
rect 204990 522996 204996 523048
rect 205048 523036 205054 523048
rect 231026 523036 231032 523048
rect 205048 523008 231032 523036
rect 205048 522996 205054 523008
rect 231026 522996 231032 523008
rect 231084 522996 231090 523048
rect 232590 522996 232596 523048
rect 232648 523036 232654 523048
rect 259362 523036 259368 523048
rect 232648 523008 259368 523036
rect 232648 522996 232654 523008
rect 259362 522996 259368 523008
rect 259420 522996 259426 523048
rect 260098 522996 260104 523048
rect 260156 523036 260162 523048
rect 287330 523036 287336 523048
rect 260156 523008 287336 523036
rect 260156 522996 260162 523008
rect 287330 522996 287336 523008
rect 287388 522996 287394 523048
rect 289078 522996 289084 523048
rect 289136 523036 289142 523048
rect 315022 523036 315028 523048
rect 289136 523008 315028 523036
rect 289136 522996 289142 523008
rect 315022 522996 315028 523008
rect 315080 522996 315086 523048
rect 316678 522996 316684 523048
rect 316736 523036 316742 523048
rect 343358 523036 343364 523048
rect 316736 523008 343364 523036
rect 316736 522996 316742 523008
rect 343358 522996 343364 523008
rect 343416 522996 343422 523048
rect 344278 522996 344284 523048
rect 344336 523036 344342 523048
rect 371326 523036 371332 523048
rect 344336 523008 371332 523036
rect 344336 522996 344342 523008
rect 371326 522996 371332 523008
rect 371384 522996 371390 523048
rect 373258 522996 373264 523048
rect 373316 523036 373322 523048
rect 399018 523036 399024 523048
rect 373316 523008 399024 523036
rect 373316 522996 373322 523008
rect 399018 522996 399024 523008
rect 399076 522996 399082 523048
rect 400858 522996 400864 523048
rect 400916 523036 400922 523048
rect 427354 523036 427360 523048
rect 400916 523008 427360 523036
rect 400916 522996 400922 523008
rect 427354 522996 427360 523008
rect 427412 522996 427418 523048
rect 428550 522996 428556 523048
rect 428608 523036 428614 523048
rect 455322 523036 455328 523048
rect 428608 523008 455328 523036
rect 428608 522996 428614 523008
rect 455322 522996 455328 523008
rect 455380 522996 455386 523048
rect 456058 522996 456064 523048
rect 456116 523036 456122 523048
rect 483014 523036 483020 523048
rect 456116 523008 483020 523036
rect 456116 522996 456122 523008
rect 483014 522996 483020 523008
rect 483072 522996 483078 523048
rect 485038 522996 485044 523048
rect 485096 523036 485102 523048
rect 511350 523036 511356 523048
rect 485096 523008 511356 523036
rect 485096 522996 485102 523008
rect 511350 522996 511356 523008
rect 511408 522996 511414 523048
rect 512638 522996 512644 523048
rect 512696 523036 512702 523048
rect 539318 523036 539324 523048
rect 512696 523008 539324 523036
rect 512696 522996 512702 523008
rect 539318 522996 539324 523008
rect 539376 522996 539382 523048
rect 540238 522996 540244 523048
rect 540296 523036 540302 523048
rect 567194 523036 567200 523048
rect 540296 523008 567200 523036
rect 540296 522996 540302 523008
rect 567194 522996 567200 523008
rect 567252 522996 567258 523048
rect 42702 520276 42708 520328
rect 42760 520316 42766 520328
rect 93854 520316 93860 520328
rect 42760 520288 93860 520316
rect 42760 520276 42766 520288
rect 93854 520276 93860 520288
rect 93912 520276 93918 520328
rect 97902 520276 97908 520328
rect 97960 520316 97966 520328
rect 149054 520316 149060 520328
rect 97960 520288 149060 520316
rect 97960 520276 97966 520288
rect 149054 520276 149060 520288
rect 149112 520276 149118 520328
rect 155862 520276 155868 520328
rect 155920 520316 155926 520328
rect 205634 520316 205640 520328
rect 155920 520288 205640 520316
rect 155920 520276 155926 520288
rect 205634 520276 205640 520288
rect 205692 520276 205698 520328
rect 209682 520276 209688 520328
rect 209740 520316 209746 520328
rect 262214 520316 262220 520328
rect 209740 520288 262220 520316
rect 209740 520276 209746 520288
rect 262214 520276 262220 520288
rect 262272 520276 262278 520328
rect 266262 520276 266268 520328
rect 266320 520316 266326 520328
rect 317414 520316 317420 520328
rect 266320 520288 317420 520316
rect 266320 520276 266326 520288
rect 317414 520276 317420 520288
rect 317472 520276 317478 520328
rect 322842 520276 322848 520328
rect 322900 520316 322906 520328
rect 373994 520316 374000 520328
rect 322900 520288 374000 520316
rect 322900 520276 322906 520288
rect 373994 520276 374000 520288
rect 374052 520276 374058 520328
rect 378042 520276 378048 520328
rect 378100 520316 378106 520328
rect 429286 520316 429292 520328
rect 378100 520288 429292 520316
rect 378100 520276 378106 520288
rect 429286 520276 429292 520288
rect 429344 520276 429350 520328
rect 434622 520276 434628 520328
rect 434680 520316 434686 520328
rect 485774 520316 485780 520328
rect 434680 520288 485780 520316
rect 434680 520276 434686 520288
rect 485774 520276 485780 520288
rect 485832 520276 485838 520328
rect 489822 520276 489828 520328
rect 489880 520316 489886 520328
rect 542354 520316 542360 520328
rect 489880 520288 542360 520316
rect 489880 520276 489886 520288
rect 542354 520276 542360 520288
rect 542412 520276 542418 520328
rect 154482 518848 154488 518900
rect 154540 518888 154546 518900
rect 155862 518888 155868 518900
rect 154540 518860 155868 518888
rect 154540 518848 154546 518860
rect 155862 518848 155868 518860
rect 155920 518848 155926 518900
rect 42886 514020 42892 514072
rect 42944 514060 42950 514072
rect 43622 514060 43628 514072
rect 42944 514032 43628 514060
rect 42944 514020 42950 514032
rect 43622 514020 43628 514032
rect 43680 514020 43686 514072
rect 63586 505588 63592 505640
rect 63644 505628 63650 505640
rect 64322 505628 64328 505640
rect 63644 505600 64328 505628
rect 63644 505588 63650 505600
rect 64322 505588 64328 505600
rect 64380 505588 64386 505640
rect 147674 505588 147680 505640
rect 147732 505628 147738 505640
rect 148410 505628 148416 505640
rect 147732 505600 148416 505628
rect 147732 505588 147738 505600
rect 148410 505588 148416 505600
rect 148468 505588 148474 505640
rect 259730 505588 259736 505640
rect 259788 505628 259794 505640
rect 260190 505628 260196 505640
rect 259788 505600 260196 505628
rect 259788 505588 259794 505600
rect 260190 505588 260196 505600
rect 260248 505588 260254 505640
rect 455690 505588 455696 505640
rect 455748 505628 455754 505640
rect 456150 505628 456156 505640
rect 455748 505600 456156 505628
rect 455748 505588 455754 505600
rect 456150 505588 456156 505600
rect 456208 505588 456214 505640
rect 287698 504568 287704 504620
rect 287756 504608 287762 504620
rect 295702 504608 295708 504620
rect 287756 504580 295708 504608
rect 287756 504568 287762 504580
rect 295702 504568 295708 504580
rect 295760 504568 295766 504620
rect 428642 504364 428648 504416
rect 428700 504404 428706 504416
rect 435726 504404 435732 504416
rect 428700 504376 435732 504404
rect 428700 504364 428706 504376
rect 435726 504364 435732 504376
rect 435784 504364 435790 504416
rect 483658 504296 483664 504348
rect 483716 504336 483722 504348
rect 491662 504336 491668 504348
rect 483716 504308 491668 504336
rect 483716 504296 483722 504308
rect 491662 504296 491668 504308
rect 491720 504296 491726 504348
rect 512730 504296 512736 504348
rect 512788 504336 512794 504348
rect 519630 504336 519636 504348
rect 512788 504308 519636 504336
rect 512788 504296 512794 504308
rect 519630 504296 519636 504308
rect 519688 504296 519694 504348
rect 232682 504228 232688 504280
rect 232740 504268 232746 504280
rect 239766 504268 239772 504280
rect 232740 504240 239772 504268
rect 232740 504228 232746 504240
rect 239766 504228 239772 504240
rect 239824 504228 239830 504280
rect 316770 503752 316776 503804
rect 316828 503792 316834 503804
rect 323670 503792 323676 503804
rect 316828 503764 323676 503792
rect 316828 503752 316834 503764
rect 323670 503752 323676 503764
rect 323728 503752 323734 503804
rect 13538 503616 13544 503668
rect 13596 503656 13602 503668
rect 66254 503656 66260 503668
rect 13596 503628 66260 503656
rect 13596 503616 13602 503628
rect 66254 503616 66260 503628
rect 66312 503616 66318 503668
rect 70302 503616 70308 503668
rect 70360 503656 70366 503668
rect 121454 503656 121460 503668
rect 70360 503628 121460 503656
rect 70360 503616 70366 503628
rect 121454 503616 121460 503628
rect 121512 503616 121518 503668
rect 126882 503616 126888 503668
rect 126940 503656 126946 503668
rect 178034 503656 178040 503668
rect 126940 503628 178040 503656
rect 126940 503616 126946 503628
rect 178034 503616 178040 503628
rect 178092 503616 178098 503668
rect 182082 503616 182088 503668
rect 182140 503656 182146 503668
rect 233234 503656 233240 503668
rect 182140 503628 233240 503656
rect 182140 503616 182146 503628
rect 233234 503616 233240 503628
rect 233292 503616 233298 503668
rect 238662 503616 238668 503668
rect 238720 503656 238726 503668
rect 289814 503656 289820 503668
rect 238720 503628 289820 503656
rect 238720 503616 238726 503628
rect 289814 503616 289820 503628
rect 289872 503616 289878 503668
rect 293862 503616 293868 503668
rect 293920 503656 293926 503668
rect 345014 503656 345020 503668
rect 293920 503628 345020 503656
rect 293920 503616 293926 503628
rect 345014 503616 345020 503628
rect 345072 503616 345078 503668
rect 350442 503616 350448 503668
rect 350500 503656 350506 503668
rect 401594 503656 401600 503668
rect 350500 503628 401600 503656
rect 350500 503616 350506 503628
rect 401594 503616 401600 503628
rect 401652 503616 401658 503668
rect 405642 503616 405648 503668
rect 405700 503656 405706 503668
rect 458174 503656 458180 503668
rect 405700 503628 458180 503656
rect 405700 503616 405706 503628
rect 458174 503616 458180 503628
rect 458232 503616 458238 503668
rect 462222 503616 462228 503668
rect 462280 503656 462286 503668
rect 513374 503656 513380 503668
rect 462280 503628 513380 503656
rect 462280 503616 462286 503628
rect 513374 503616 513380 503628
rect 513432 503616 513438 503668
rect 518802 503616 518808 503668
rect 518860 503656 518866 503668
rect 569954 503656 569960 503668
rect 518860 503628 569960 503656
rect 518860 503616 518866 503628
rect 569954 503616 569960 503628
rect 570012 503616 570018 503668
rect 539502 503548 539508 503600
rect 539560 503588 539566 503600
rect 541618 503588 541624 503600
rect 539560 503560 541624 503588
rect 539560 503548 539566 503560
rect 541618 503548 541624 503560
rect 541676 503548 541682 503600
rect 15102 502664 15108 502716
rect 15160 502704 15166 502716
rect 16574 502704 16580 502716
rect 15160 502676 16580 502704
rect 15160 502664 15166 502676
rect 16574 502664 16580 502676
rect 16632 502664 16638 502716
rect 547874 502664 547880 502716
rect 547932 502704 547938 502716
rect 548150 502704 548156 502716
rect 547932 502676 548156 502704
rect 547932 502664 547938 502676
rect 548150 502664 548156 502676
rect 548208 502664 548214 502716
rect 35250 502256 35256 502308
rect 35308 502296 35314 502308
rect 36630 502296 36636 502308
rect 35308 502268 36636 502296
rect 35308 502256 35314 502268
rect 36630 502256 36636 502268
rect 36688 502256 36694 502308
rect 71866 500896 71872 500948
rect 71924 500936 71930 500948
rect 100018 500936 100024 500948
rect 71924 500908 100024 500936
rect 71924 500896 71930 500908
rect 100018 500896 100024 500908
rect 100076 500896 100082 500948
rect 127986 500936 127992 500948
rect 103486 500908 127992 500936
rect 25682 500828 25688 500880
rect 25740 500868 25746 500880
rect 36722 500868 36728 500880
rect 25740 500840 36728 500868
rect 25740 500828 25746 500840
rect 36722 500828 36728 500840
rect 36780 500828 36786 500880
rect 42886 500828 42892 500880
rect 42944 500868 42950 500880
rect 42944 500840 45554 500868
rect 42944 500828 42950 500840
rect 15286 500760 15292 500812
rect 15344 500800 15350 500812
rect 43990 500800 43996 500812
rect 15344 500772 43996 500800
rect 15344 500760 15350 500772
rect 43990 500760 43996 500772
rect 44048 500760 44054 500812
rect 45526 500800 45554 500840
rect 53650 500828 53656 500880
rect 53708 500868 53714 500880
rect 66898 500868 66904 500880
rect 53708 500840 66904 500868
rect 53708 500828 53714 500840
rect 66898 500828 66904 500840
rect 66956 500828 66962 500880
rect 81986 500828 81992 500880
rect 82044 500868 82050 500880
rect 93118 500868 93124 500880
rect 82044 500840 93124 500868
rect 82044 500828 82050 500840
rect 93118 500828 93124 500840
rect 93176 500828 93182 500880
rect 99466 500828 99472 500880
rect 99524 500868 99530 500880
rect 103486 500868 103514 500908
rect 127986 500896 127992 500908
rect 128044 500896 128050 500948
rect 165982 500896 165988 500948
rect 166040 500936 166046 500948
rect 177298 500936 177304 500948
rect 166040 500908 177304 500936
rect 166040 500896 166046 500908
rect 177298 500896 177304 500908
rect 177356 500896 177362 500948
rect 178678 500896 178684 500948
rect 178736 500936 178742 500948
rect 184014 500936 184020 500948
rect 178736 500908 184020 500936
rect 178736 500896 178742 500908
rect 184014 500896 184020 500908
rect 184072 500896 184078 500948
rect 211706 500936 211712 500948
rect 190426 500908 211712 500936
rect 99524 500840 103514 500868
rect 99524 500828 99530 500840
rect 109678 500828 109684 500880
rect 109736 500868 109742 500880
rect 124858 500868 124864 500880
rect 109736 500840 124864 500868
rect 109736 500828 109742 500840
rect 124858 500828 124864 500840
rect 124916 500828 124922 500880
rect 137646 500828 137652 500880
rect 137704 500868 137710 500880
rect 148318 500868 148324 500880
rect 137704 500840 148324 500868
rect 137704 500828 137710 500840
rect 148318 500828 148324 500840
rect 148376 500828 148382 500880
rect 183646 500828 183652 500880
rect 183704 500868 183710 500880
rect 190426 500868 190454 500908
rect 211706 500896 211712 500908
rect 211764 500896 211770 500948
rect 277670 500896 277676 500948
rect 277728 500936 277734 500948
rect 289078 500936 289084 500948
rect 277728 500908 289084 500936
rect 277728 500896 277734 500908
rect 289078 500896 289084 500908
rect 289136 500896 289142 500948
rect 306006 500896 306012 500948
rect 306064 500936 306070 500948
rect 316678 500936 316684 500948
rect 306064 500908 316684 500936
rect 306064 500896 306070 500908
rect 316678 500896 316684 500908
rect 316736 500896 316742 500948
rect 343358 500896 343364 500948
rect 343416 500936 343422 500948
rect 345658 500936 345664 500948
rect 343416 500908 345664 500936
rect 343416 500896 343422 500908
rect 345658 500896 345664 500908
rect 345716 500896 345722 500948
rect 361666 500896 361672 500948
rect 361724 500936 361730 500948
rect 373258 500936 373264 500948
rect 361724 500908 373264 500936
rect 361724 500896 361730 500908
rect 373258 500896 373264 500908
rect 373316 500896 373322 500948
rect 379606 500896 379612 500948
rect 379664 500936 379670 500948
rect 408034 500936 408040 500948
rect 379664 500908 408040 500936
rect 379664 500896 379670 500908
rect 408034 500896 408040 500908
rect 408092 500896 408098 500948
rect 473998 500896 474004 500948
rect 474056 500936 474062 500948
rect 485038 500936 485044 500948
rect 474056 500908 485044 500936
rect 474056 500896 474062 500908
rect 485038 500896 485044 500908
rect 485096 500896 485102 500948
rect 501690 500896 501696 500948
rect 501748 500936 501754 500948
rect 512638 500936 512644 500948
rect 501748 500908 512644 500936
rect 501748 500896 501754 500908
rect 512638 500896 512644 500908
rect 512696 500896 512702 500948
rect 548150 500896 548156 500948
rect 548208 500936 548214 500948
rect 557534 500936 557540 500948
rect 548208 500908 557540 500936
rect 548208 500896 548214 500908
rect 557534 500896 557540 500908
rect 557592 500896 557598 500948
rect 183704 500840 190454 500868
rect 183704 500828 183710 500840
rect 193674 500828 193680 500880
rect 193732 500868 193738 500880
rect 204990 500868 204996 500880
rect 193732 500840 204996 500868
rect 193732 500828 193738 500840
rect 204990 500828 204996 500840
rect 205048 500828 205054 500880
rect 222010 500828 222016 500880
rect 222068 500868 222074 500880
rect 232590 500868 232596 500880
rect 222068 500840 232596 500868
rect 222068 500828 222074 500840
rect 232590 500828 232596 500840
rect 232648 500828 232654 500880
rect 249702 500828 249708 500880
rect 249760 500868 249766 500880
rect 260098 500868 260104 500880
rect 249760 500840 260104 500868
rect 249760 500828 249766 500840
rect 260098 500828 260104 500840
rect 260156 500828 260162 500880
rect 333698 500828 333704 500880
rect 333756 500868 333762 500880
rect 344278 500868 344284 500880
rect 333756 500840 344284 500868
rect 333756 500828 333762 500840
rect 344278 500828 344284 500840
rect 344336 500828 344342 500880
rect 374638 500828 374644 500880
rect 374696 500868 374702 500880
rect 379698 500868 379704 500880
rect 374696 500840 379704 500868
rect 374696 500828 374702 500840
rect 379698 500828 379704 500840
rect 379756 500828 379762 500880
rect 390002 500828 390008 500880
rect 390060 500868 390066 500880
rect 400858 500868 400864 500880
rect 390060 500840 400864 500868
rect 390060 500828 390066 500840
rect 400858 500828 400864 500840
rect 400916 500828 400922 500880
rect 417694 500828 417700 500880
rect 417752 500868 417758 500880
rect 428550 500868 428556 500880
rect 417752 500840 428556 500868
rect 417752 500828 417758 500840
rect 428550 500828 428556 500840
rect 428608 500828 428614 500880
rect 445662 500828 445668 500880
rect 445720 500868 445726 500880
rect 456058 500868 456064 500880
rect 445720 500840 456064 500868
rect 445720 500828 445726 500840
rect 456058 500828 456064 500840
rect 456116 500828 456122 500880
rect 529658 500828 529664 500880
rect 529716 500868 529722 500880
rect 540238 500868 540244 500880
rect 529716 500840 540244 500868
rect 529716 500828 529722 500840
rect 540238 500828 540244 500840
rect 540296 500828 540302 500880
rect 72050 500800 72056 500812
rect 45526 500772 72056 500800
rect 72050 500760 72056 500772
rect 72108 500760 72114 500812
rect 127066 500760 127072 500812
rect 127124 500800 127130 500812
rect 156046 500800 156052 500812
rect 127124 500772 156052 500800
rect 127124 500760 127130 500772
rect 156046 500760 156052 500772
rect 156104 500760 156110 500812
rect 238846 500760 238852 500812
rect 238904 500800 238910 500812
rect 268010 500800 268016 500812
rect 238904 500772 268016 500800
rect 238904 500760 238910 500772
rect 268010 500760 268016 500772
rect 268068 500760 268074 500812
rect 323026 500760 323032 500812
rect 323084 500800 323090 500812
rect 352006 500800 352012 500812
rect 323084 500772 352012 500800
rect 323084 500760 323090 500772
rect 352006 500760 352012 500772
rect 352064 500760 352070 500812
rect 434806 500760 434812 500812
rect 434864 500800 434870 500812
rect 463694 500800 463700 500812
rect 434864 500772 463700 500800
rect 434864 500760 434870 500772
rect 463694 500760 463700 500772
rect 463752 500760 463758 500812
rect 518986 500760 518992 500812
rect 519044 500800 519050 500812
rect 547874 500800 547880 500812
rect 519044 500772 547880 500800
rect 519044 500760 519050 500772
rect 547874 500760 547880 500772
rect 547932 500760 547938 500812
rect 71130 496952 71136 497004
rect 71188 496992 71194 497004
rect 82262 496992 82268 497004
rect 71188 496964 82268 496992
rect 71188 496952 71194 496964
rect 82262 496952 82268 496964
rect 82320 496952 82326 497004
rect 184198 496952 184204 497004
rect 184256 496992 184262 497004
rect 222286 496992 222292 497004
rect 184256 496964 222292 496992
rect 184256 496952 184262 496964
rect 222286 496952 222292 496964
rect 222344 496952 222350 497004
rect 266998 496952 267004 497004
rect 267056 496992 267062 497004
rect 277946 496992 277952 497004
rect 267056 496964 277952 496992
rect 267056 496952 267062 496964
rect 277946 496952 277952 496964
rect 278004 496952 278010 497004
rect 296162 496952 296168 497004
rect 296220 496992 296226 497004
rect 334250 496992 334256 497004
rect 296220 496964 334256 496992
rect 296220 496952 296226 496964
rect 334250 496952 334256 496964
rect 334308 496952 334314 497004
rect 352190 496952 352196 497004
rect 352248 496992 352254 497004
rect 352248 496964 364334 496992
rect 352248 496952 352254 496964
rect 26234 496884 26240 496936
rect 26292 496924 26298 496936
rect 35434 496924 35440 496936
rect 26292 496896 35440 496924
rect 26292 496884 26298 496896
rect 35434 496884 35440 496896
rect 35492 496884 35498 496936
rect 36630 496884 36636 496936
rect 36688 496924 36694 496936
rect 53926 496924 53932 496936
rect 36688 496896 53932 496924
rect 36688 496884 36694 496896
rect 53926 496884 53932 496896
rect 53984 496884 53990 496936
rect 72234 496884 72240 496936
rect 72292 496924 72298 496936
rect 109954 496924 109960 496936
rect 72292 496896 109960 496924
rect 72292 496884 72298 496896
rect 109954 496884 109960 496896
rect 110012 496884 110018 496936
rect 151078 496884 151084 496936
rect 151136 496924 151142 496936
rect 156598 496924 156604 496936
rect 151136 496896 156604 496924
rect 151136 496884 151142 496896
rect 156598 496884 156604 496896
rect 156656 496884 156662 496936
rect 182818 496884 182824 496936
rect 182876 496924 182882 496936
rect 193950 496924 193956 496936
rect 182876 496896 193956 496924
rect 182876 496884 182882 496896
rect 193950 496884 193956 496896
rect 194008 496884 194014 496936
rect 232498 496884 232504 496936
rect 232556 496924 232562 496936
rect 232556 496896 248414 496924
rect 232556 496884 232562 496896
rect 66898 496816 66904 496868
rect 66956 496856 66962 496868
rect 72602 496856 72608 496868
rect 66956 496828 72608 496856
rect 66956 496816 66962 496828
rect 72602 496816 72608 496828
rect 72660 496816 72666 496868
rect 93118 496816 93124 496868
rect 93176 496856 93182 496868
rect 100294 496856 100300 496868
rect 93176 496828 100300 496856
rect 93176 496816 93182 496828
rect 100294 496816 100300 496828
rect 100352 496816 100358 496868
rect 138290 496856 138296 496868
rect 100404 496828 138296 496856
rect 100202 496748 100208 496800
rect 100260 496788 100266 496800
rect 100404 496788 100432 496828
rect 138290 496816 138296 496828
rect 138348 496816 138354 496868
rect 149698 496816 149704 496868
rect 149756 496856 149762 496868
rect 166258 496856 166264 496868
rect 149756 496828 166264 496856
rect 149756 496816 149762 496828
rect 166258 496816 166264 496828
rect 166316 496816 166322 496868
rect 177298 496816 177304 496868
rect 177356 496856 177362 496868
rect 184290 496856 184296 496868
rect 177356 496828 184296 496856
rect 177356 496816 177362 496828
rect 184290 496816 184296 496828
rect 184348 496816 184354 496868
rect 233970 496816 233976 496868
rect 234028 496856 234034 496868
rect 240594 496856 240600 496868
rect 234028 496828 240600 496856
rect 234028 496816 234034 496828
rect 240594 496816 240600 496828
rect 240652 496816 240658 496868
rect 248386 496856 248414 496896
rect 268194 496884 268200 496936
rect 268252 496924 268258 496936
rect 306282 496924 306288 496936
rect 268252 496896 306288 496924
rect 268252 496884 268258 496896
rect 306282 496884 306288 496896
rect 306340 496884 306346 496936
rect 345658 496884 345664 496936
rect 345716 496924 345722 496936
rect 361942 496924 361948 496936
rect 345716 496896 361948 496924
rect 345716 496884 345722 496896
rect 361942 496884 361948 496896
rect 362000 496884 362006 496936
rect 364306 496924 364334 496964
rect 380250 496952 380256 497004
rect 380308 496992 380314 497004
rect 418246 496992 418252 497004
rect 380308 496964 418252 496992
rect 380308 496952 380314 496964
rect 418246 496952 418252 496964
rect 418304 496952 418310 497004
rect 464154 496952 464160 497004
rect 464212 496992 464218 497004
rect 464212 496964 470594 496992
rect 464212 496952 464218 496964
rect 390278 496924 390284 496936
rect 364306 496896 390284 496924
rect 390278 496884 390284 496896
rect 390336 496884 390342 496936
rect 400950 496884 400956 496936
rect 401008 496924 401014 496936
rect 408586 496924 408592 496936
rect 401008 496896 408592 496924
rect 401008 496884 401014 496896
rect 408586 496884 408592 496896
rect 408644 496884 408650 496936
rect 429838 496884 429844 496936
rect 429896 496924 429902 496936
rect 436278 496924 436284 496936
rect 429896 496896 436284 496924
rect 429896 496884 429902 496896
rect 436278 496884 436284 496896
rect 436336 496884 436342 496936
rect 457438 496884 457444 496936
rect 457496 496924 457502 496936
rect 464614 496924 464620 496936
rect 457496 496896 464620 496924
rect 457496 496884 457502 496896
rect 464614 496884 464620 496896
rect 464672 496884 464678 496936
rect 470566 496924 470594 496964
rect 485038 496952 485044 497004
rect 485096 496992 485102 497004
rect 492582 496992 492588 497004
rect 485096 496964 492588 496992
rect 485096 496952 485102 496964
rect 492582 496952 492588 496964
rect 492640 496952 492646 497004
rect 502242 496924 502248 496936
rect 470566 496896 502248 496924
rect 502242 496884 502248 496896
rect 502300 496884 502306 496936
rect 514018 496884 514024 496936
rect 514076 496924 514082 496936
rect 520274 496924 520280 496936
rect 514076 496896 520280 496924
rect 514076 496884 514082 496896
rect 520274 496884 520280 496896
rect 520332 496884 520338 496936
rect 250254 496856 250260 496868
rect 248386 496828 250260 496856
rect 250254 496816 250260 496828
rect 250312 496816 250318 496868
rect 261478 496816 261484 496868
rect 261536 496856 261542 496868
rect 268286 496856 268292 496868
rect 261536 496828 268292 496856
rect 261536 496816 261542 496828
rect 268286 496816 268292 496828
rect 268344 496816 268350 496868
rect 289078 496816 289084 496868
rect 289136 496856 289142 496868
rect 296622 496856 296628 496868
rect 289136 496828 296628 496856
rect 289136 496816 289142 496828
rect 296622 496816 296628 496828
rect 296680 496816 296686 496868
rect 318058 496816 318064 496868
rect 318116 496856 318122 496868
rect 324590 496856 324596 496868
rect 318116 496828 324596 496856
rect 318116 496816 318122 496828
rect 324590 496816 324596 496828
rect 324648 496816 324654 496868
rect 347038 496816 347044 496868
rect 347096 496856 347102 496868
rect 352282 496856 352288 496868
rect 347096 496828 352288 496856
rect 347096 496816 347102 496828
rect 352282 496816 352288 496828
rect 352340 496816 352346 496868
rect 373258 496816 373264 496868
rect 373316 496856 373322 496868
rect 380618 496856 380624 496868
rect 373316 496828 380624 496856
rect 373316 496816 373322 496828
rect 380618 496816 380624 496828
rect 380676 496816 380682 496868
rect 428458 496816 428464 496868
rect 428516 496856 428522 496868
rect 445938 496856 445944 496868
rect 428516 496828 445944 496856
rect 428516 496816 428522 496828
rect 445938 496816 445944 496828
rect 445996 496816 446002 496868
rect 462958 496816 462964 496868
rect 463016 496856 463022 496868
rect 474274 496856 474280 496868
rect 463016 496828 474280 496856
rect 463016 496816 463022 496828
rect 474274 496816 474280 496828
rect 474332 496816 474338 496868
rect 492122 496816 492128 496868
rect 492180 496856 492186 496868
rect 529934 496856 529940 496868
rect 492180 496828 529940 496856
rect 492180 496816 492186 496828
rect 529934 496816 529940 496828
rect 529992 496816 529998 496868
rect 541618 496816 541624 496868
rect 541676 496856 541682 496868
rect 558270 496856 558276 496868
rect 541676 496828 558276 496856
rect 541676 496816 541682 496828
rect 558270 496816 558276 496828
rect 558328 496816 558334 496868
rect 100260 496760 100432 496788
rect 100260 496748 100266 496760
rect 120166 494232 120172 494284
rect 120224 494272 120230 494284
rect 122098 494272 122104 494284
rect 120224 494244 122104 494272
rect 120224 494232 120230 494244
rect 122098 494232 122104 494244
rect 122156 494232 122162 494284
rect 124858 494232 124864 494284
rect 124916 494272 124922 494284
rect 128262 494272 128268 494284
rect 124916 494244 128268 494272
rect 124916 494232 124922 494244
rect 128262 494232 128268 494244
rect 128320 494232 128326 494284
rect 210418 494232 210424 494284
rect 210476 494272 210482 494284
rect 212350 494272 212356 494284
rect 210476 494244 212356 494272
rect 210476 494232 210482 494244
rect 212350 494232 212356 494244
rect 212408 494232 212414 494284
rect 544378 494028 544384 494080
rect 544436 494068 544442 494080
rect 548334 494068 548340 494080
rect 544436 494040 548340 494068
rect 544436 494028 544442 494040
rect 548334 494028 548340 494040
rect 548392 494028 548398 494080
rect 204254 492056 204260 492108
rect 204312 492096 204318 492108
rect 204990 492096 204996 492108
rect 204312 492068 204996 492096
rect 204312 492056 204318 492068
rect 204990 492056 204996 492068
rect 205048 492056 205054 492108
rect 13538 476008 13544 476060
rect 13596 476048 13602 476060
rect 66254 476048 66260 476060
rect 13596 476020 66260 476048
rect 13596 476008 13602 476020
rect 66254 476008 66260 476020
rect 66312 476008 66318 476060
rect 70302 476008 70308 476060
rect 70360 476048 70366 476060
rect 121454 476048 121460 476060
rect 70360 476020 121460 476048
rect 70360 476008 70366 476020
rect 121454 476008 121460 476020
rect 121512 476008 121518 476060
rect 126882 476008 126888 476060
rect 126940 476048 126946 476060
rect 178034 476048 178040 476060
rect 126940 476020 178040 476048
rect 126940 476008 126946 476020
rect 178034 476008 178040 476020
rect 178092 476008 178098 476060
rect 209682 476008 209688 476060
rect 209740 476048 209746 476060
rect 262214 476048 262220 476060
rect 209740 476020 262220 476048
rect 209740 476008 209746 476020
rect 262214 476008 262220 476020
rect 262272 476008 262278 476060
rect 266262 476008 266268 476060
rect 266320 476048 266326 476060
rect 317414 476048 317420 476060
rect 266320 476020 317420 476048
rect 266320 476008 266326 476020
rect 317414 476008 317420 476020
rect 317472 476008 317478 476060
rect 322842 476008 322848 476060
rect 322900 476048 322906 476060
rect 373994 476048 374000 476060
rect 322900 476020 374000 476048
rect 322900 476008 322906 476020
rect 373994 476008 374000 476020
rect 374052 476008 374058 476060
rect 405642 476008 405648 476060
rect 405700 476048 405706 476060
rect 458174 476048 458180 476060
rect 405700 476020 458180 476048
rect 405700 476008 405706 476020
rect 458174 476008 458180 476020
rect 458232 476008 458238 476060
rect 489822 476008 489828 476060
rect 489880 476048 489886 476060
rect 542354 476048 542360 476060
rect 489880 476020 542360 476048
rect 489880 476008 489886 476020
rect 542354 476008 542360 476020
rect 542412 476008 542418 476060
rect 42702 475940 42708 475992
rect 42760 475980 42766 475992
rect 93854 475980 93860 475992
rect 42760 475952 93860 475980
rect 42760 475940 42766 475952
rect 93854 475940 93860 475952
rect 93912 475940 93918 475992
rect 97902 475940 97908 475992
rect 97960 475980 97966 475992
rect 149054 475980 149060 475992
rect 97960 475952 149060 475980
rect 97960 475940 97966 475952
rect 149054 475940 149060 475952
rect 149112 475940 149118 475992
rect 154482 475940 154488 475992
rect 154540 475980 154546 475992
rect 205634 475980 205640 475992
rect 154540 475952 205640 475980
rect 154540 475940 154546 475952
rect 205634 475940 205640 475952
rect 205692 475940 205698 475992
rect 238662 475940 238668 475992
rect 238720 475980 238726 475992
rect 289814 475980 289820 475992
rect 238720 475952 289820 475980
rect 238720 475940 238726 475952
rect 289814 475940 289820 475952
rect 289872 475940 289878 475992
rect 293862 475940 293868 475992
rect 293920 475980 293926 475992
rect 345014 475980 345020 475992
rect 293920 475952 345020 475980
rect 293920 475940 293926 475952
rect 345014 475940 345020 475952
rect 345072 475940 345078 475992
rect 378042 475940 378048 475992
rect 378100 475980 378106 475992
rect 429286 475980 429292 475992
rect 378100 475952 429292 475980
rect 378100 475940 378106 475952
rect 429286 475940 429292 475952
rect 429344 475940 429350 475992
rect 462222 475940 462228 475992
rect 462280 475980 462286 475992
rect 513374 475980 513380 475992
rect 462280 475952 513380 475980
rect 462280 475940 462286 475952
rect 513374 475940 513380 475952
rect 513432 475940 513438 475992
rect 518802 475940 518808 475992
rect 518860 475980 518866 475992
rect 569954 475980 569960 475992
rect 518860 475952 569960 475980
rect 518860 475940 518866 475952
rect 569954 475940 569960 475952
rect 570012 475940 570018 475992
rect 182082 475872 182088 475924
rect 182140 475912 182146 475924
rect 233234 475912 233240 475924
rect 182140 475884 233240 475912
rect 182140 475872 182146 475884
rect 233234 475872 233240 475884
rect 233292 475872 233298 475924
rect 350442 475872 350448 475924
rect 350500 475912 350506 475924
rect 401594 475912 401600 475924
rect 350500 475884 401600 475912
rect 350500 475872 350506 475884
rect 401594 475872 401600 475884
rect 401652 475872 401658 475924
rect 434622 475872 434628 475924
rect 434680 475912 434686 475924
rect 485774 475912 485780 475924
rect 434680 475884 485780 475912
rect 434680 475872 434686 475884
rect 485774 475872 485780 475884
rect 485832 475872 485838 475924
rect 15194 473288 15200 473340
rect 15252 473328 15258 473340
rect 35894 473328 35900 473340
rect 15252 473300 35900 473328
rect 15252 473288 15258 473300
rect 35894 473288 35900 473300
rect 35952 473288 35958 473340
rect 36078 473288 36084 473340
rect 36136 473328 36142 473340
rect 63586 473328 63592 473340
rect 36136 473300 63592 473328
rect 36136 473288 36142 473300
rect 63586 473288 63592 473300
rect 63644 473288 63650 473340
rect 64046 473288 64052 473340
rect 64104 473328 64110 473340
rect 91922 473328 91928 473340
rect 64104 473300 91928 473328
rect 64104 473288 64110 473300
rect 91922 473288 91928 473300
rect 91980 473288 91986 473340
rect 92106 473288 92112 473340
rect 92164 473328 92170 473340
rect 119614 473328 119620 473340
rect 92164 473300 119620 473328
rect 92164 473288 92170 473300
rect 119614 473288 119620 473300
rect 119672 473288 119678 473340
rect 122098 473288 122104 473340
rect 122156 473328 122162 473340
rect 147950 473328 147956 473340
rect 122156 473300 147956 473328
rect 122156 473288 122162 473300
rect 147950 473288 147956 473300
rect 148008 473288 148014 473340
rect 148042 473288 148048 473340
rect 148100 473328 148106 473340
rect 175918 473328 175924 473340
rect 148100 473300 175924 473328
rect 148100 473288 148106 473300
rect 175918 473288 175924 473300
rect 175976 473288 175982 473340
rect 176102 473288 176108 473340
rect 176160 473328 176166 473340
rect 203610 473328 203616 473340
rect 176160 473300 203616 473328
rect 176160 473288 176166 473300
rect 203610 473288 203616 473300
rect 203668 473288 203674 473340
rect 204990 473288 204996 473340
rect 205048 473328 205054 473340
rect 231946 473328 231952 473340
rect 205048 473300 231952 473328
rect 205048 473288 205054 473300
rect 231946 473288 231952 473300
rect 232004 473288 232010 473340
rect 232038 473288 232044 473340
rect 232096 473328 232102 473340
rect 259914 473328 259920 473340
rect 232096 473300 259920 473328
rect 232096 473288 232102 473300
rect 259914 473288 259920 473300
rect 259972 473288 259978 473340
rect 260098 473288 260104 473340
rect 260156 473328 260162 473340
rect 287606 473328 287612 473340
rect 260156 473300 287612 473328
rect 260156 473288 260162 473300
rect 287606 473288 287612 473300
rect 287664 473288 287670 473340
rect 288066 473288 288072 473340
rect 288124 473328 288130 473340
rect 315942 473328 315948 473340
rect 288124 473300 315948 473328
rect 288124 473288 288130 473300
rect 315942 473288 315948 473300
rect 316000 473288 316006 473340
rect 316678 473288 316684 473340
rect 316736 473328 316742 473340
rect 343910 473328 343916 473340
rect 316736 473300 343916 473328
rect 316736 473288 316742 473300
rect 343910 473288 343916 473300
rect 343968 473288 343974 473340
rect 344094 473288 344100 473340
rect 344152 473328 344158 473340
rect 371602 473328 371608 473340
rect 344152 473300 371608 473328
rect 344152 473288 344158 473300
rect 371602 473288 371608 473300
rect 371660 473288 371666 473340
rect 372062 473288 372068 473340
rect 372120 473328 372126 473340
rect 399938 473328 399944 473340
rect 372120 473300 399944 473328
rect 372120 473288 372126 473300
rect 399938 473288 399944 473300
rect 399996 473288 400002 473340
rect 400858 473288 400864 473340
rect 400916 473328 400922 473340
rect 427906 473328 427912 473340
rect 400916 473300 427912 473328
rect 400916 473288 400922 473300
rect 427906 473288 427912 473300
rect 427964 473288 427970 473340
rect 428090 473288 428096 473340
rect 428148 473328 428154 473340
rect 455598 473328 455604 473340
rect 428148 473300 455604 473328
rect 428148 473288 428154 473300
rect 455598 473288 455604 473300
rect 455656 473288 455662 473340
rect 456058 473288 456064 473340
rect 456116 473328 456122 473340
rect 483934 473328 483940 473340
rect 456116 473300 483940 473328
rect 456116 473288 456122 473300
rect 483934 473288 483940 473300
rect 483992 473288 483998 473340
rect 484026 473288 484032 473340
rect 484084 473328 484090 473340
rect 511902 473328 511908 473340
rect 484084 473300 511908 473328
rect 484084 473288 484090 473300
rect 511902 473288 511908 473300
rect 511960 473288 511966 473340
rect 512086 473288 512092 473340
rect 512144 473328 512150 473340
rect 539594 473328 539600 473340
rect 512144 473300 539600 473328
rect 512144 473288 512150 473300
rect 539594 473288 539600 473300
rect 539652 473288 539658 473340
rect 540054 473288 540060 473340
rect 540112 473328 540118 473340
rect 567930 473328 567936 473340
rect 540112 473300 567936 473328
rect 540112 473288 540118 473300
rect 567930 473288 567936 473300
rect 567988 473288 567994 473340
rect 16574 473220 16580 473272
rect 16632 473260 16638 473272
rect 36630 473260 36636 473272
rect 16632 473232 36636 473260
rect 16632 473220 16638 473232
rect 36630 473220 36636 473232
rect 36688 473220 36694 473272
rect 44910 473220 44916 473272
rect 44968 473260 44974 473272
rect 71130 473260 71136 473272
rect 44968 473232 71136 473260
rect 44968 473220 44974 473232
rect 71130 473220 71136 473232
rect 71188 473220 71194 473272
rect 82262 473220 82268 473272
rect 82320 473260 82326 473272
rect 93118 473260 93124 473272
rect 82320 473232 93124 473260
rect 82320 473220 82326 473232
rect 93118 473220 93124 473232
rect 93176 473220 93182 473272
rect 110230 473220 110236 473272
rect 110288 473260 110294 473272
rect 124858 473260 124864 473272
rect 110288 473232 124864 473260
rect 110288 473220 110294 473232
rect 124858 473220 124864 473232
rect 124916 473220 124922 473272
rect 128630 473220 128636 473272
rect 128688 473260 128694 473272
rect 149698 473260 149704 473272
rect 128688 473232 149704 473260
rect 128688 473220 128694 473232
rect 149698 473220 149704 473232
rect 149756 473220 149762 473272
rect 156598 473220 156604 473272
rect 156656 473260 156662 473272
rect 182818 473260 182824 473272
rect 156656 473232 182824 473260
rect 156656 473220 156662 473232
rect 182818 473220 182824 473232
rect 182876 473220 182882 473272
rect 194502 473220 194508 473272
rect 194560 473260 194566 473272
rect 210418 473260 210424 473272
rect 194560 473232 210424 473260
rect 194560 473220 194566 473232
rect 210418 473220 210424 473232
rect 210476 473220 210482 473272
rect 212626 473220 212632 473272
rect 212684 473260 212690 473272
rect 232498 473260 232504 473272
rect 212684 473232 232504 473260
rect 212684 473220 212690 473232
rect 232498 473220 232504 473232
rect 232556 473220 232562 473272
rect 240594 473220 240600 473272
rect 240652 473260 240658 473272
rect 266998 473260 267004 473272
rect 240652 473232 267004 473260
rect 240652 473220 240658 473232
rect 266998 473220 267004 473232
rect 267056 473220 267062 473272
rect 278590 473220 278596 473272
rect 278648 473260 278654 473272
rect 289078 473260 289084 473272
rect 278648 473232 289084 473260
rect 278648 473220 278654 473232
rect 289078 473220 289084 473232
rect 289136 473220 289142 473272
rect 306282 473220 306288 473272
rect 306340 473260 306346 473272
rect 318058 473260 318064 473272
rect 306340 473232 318064 473260
rect 306340 473220 306346 473232
rect 318058 473220 318064 473232
rect 318116 473220 318122 473272
rect 324590 473220 324596 473272
rect 324648 473260 324654 473272
rect 345658 473260 345664 473272
rect 324648 473232 345664 473260
rect 324648 473220 324654 473232
rect 345658 473220 345664 473232
rect 345716 473220 345722 473272
rect 362586 473220 362592 473272
rect 362644 473260 362650 473272
rect 373258 473260 373264 473272
rect 362644 473232 373264 473260
rect 362644 473220 362650 473232
rect 373258 473220 373264 473232
rect 373316 473220 373322 473272
rect 390278 473220 390284 473272
rect 390336 473260 390342 473272
rect 400950 473260 400956 473272
rect 390336 473232 400956 473260
rect 390336 473220 390342 473232
rect 400950 473220 400956 473232
rect 401008 473220 401014 473272
rect 408586 473220 408592 473272
rect 408644 473260 408650 473272
rect 428458 473260 428464 473272
rect 408644 473232 428464 473260
rect 408644 473220 408650 473232
rect 428458 473220 428464 473232
rect 428516 473220 428522 473272
rect 436922 473220 436928 473272
rect 436980 473260 436986 473272
rect 462958 473260 462964 473272
rect 436980 473232 462964 473260
rect 436980 473220 436986 473232
rect 462958 473220 462964 473232
rect 463016 473220 463022 473272
rect 474274 473220 474280 473272
rect 474332 473260 474338 473272
rect 485038 473260 485044 473272
rect 474332 473232 485044 473260
rect 474332 473220 474338 473232
rect 485038 473220 485044 473232
rect 485096 473220 485102 473272
rect 502242 473220 502248 473272
rect 502300 473260 502306 473272
rect 514018 473260 514024 473272
rect 502300 473232 514024 473260
rect 502300 473220 502306 473232
rect 514018 473220 514024 473232
rect 514076 473220 514082 473272
rect 520918 473220 520924 473272
rect 520976 473260 520982 473272
rect 541618 473260 541624 473272
rect 520976 473232 541624 473260
rect 520976 473220 520982 473232
rect 541618 473220 541624 473232
rect 541676 473220 541682 473272
rect 26234 473152 26240 473204
rect 26292 473192 26298 473204
rect 43530 473192 43536 473204
rect 26292 473164 43536 473192
rect 26292 473152 26298 473164
rect 43530 473152 43536 473164
rect 43588 473152 43594 473204
rect 54570 473152 54576 473204
rect 54628 473192 54634 473204
rect 66898 473192 66904 473204
rect 54628 473164 66904 473192
rect 54628 473152 54634 473164
rect 66898 473152 66904 473164
rect 66956 473152 66962 473204
rect 138290 473152 138296 473204
rect 138348 473192 138354 473204
rect 151078 473192 151084 473204
rect 138348 473164 151084 473192
rect 138348 473152 138354 473164
rect 151078 473152 151084 473164
rect 151136 473152 151142 473204
rect 166258 473152 166264 473204
rect 166316 473192 166322 473204
rect 177298 473192 177304 473204
rect 166316 473164 177304 473192
rect 166316 473152 166322 473164
rect 177298 473152 177304 473164
rect 177356 473152 177362 473204
rect 222286 473152 222292 473204
rect 222344 473192 222350 473204
rect 233970 473192 233976 473204
rect 222344 473164 233976 473192
rect 222344 473152 222350 473164
rect 233970 473152 233976 473164
rect 234028 473152 234034 473204
rect 250254 473152 250260 473204
rect 250312 473192 250318 473204
rect 261478 473192 261484 473204
rect 250312 473164 261484 473192
rect 250312 473152 250318 473164
rect 261478 473152 261484 473164
rect 261536 473152 261542 473204
rect 334250 473152 334256 473204
rect 334308 473192 334314 473204
rect 347038 473192 347044 473204
rect 334308 473164 347044 473192
rect 334308 473152 334314 473164
rect 347038 473152 347044 473164
rect 347096 473152 347102 473204
rect 418246 473152 418252 473204
rect 418304 473192 418310 473204
rect 429838 473192 429844 473204
rect 418304 473164 429844 473192
rect 418304 473152 418310 473164
rect 429838 473152 429844 473164
rect 429896 473152 429902 473204
rect 446582 473152 446588 473204
rect 446640 473192 446646 473204
rect 457438 473192 457444 473204
rect 446640 473164 457444 473192
rect 446640 473152 446646 473164
rect 457438 473152 457444 473164
rect 457496 473152 457502 473204
rect 530578 473152 530584 473204
rect 530636 473192 530642 473204
rect 544378 473192 544384 473204
rect 530636 473164 544384 473192
rect 530636 473152 530642 473164
rect 544378 473152 544384 473164
rect 544436 473152 544442 473204
rect 558270 472608 558276 472660
rect 558328 472648 558334 472660
rect 567470 472648 567476 472660
rect 558328 472620 567476 472648
rect 558328 472608 558334 472620
rect 567470 472608 567476 472620
rect 567528 472608 567534 472660
rect 64322 470568 64328 470620
rect 64380 470608 64386 470620
rect 579982 470608 579988 470620
rect 64380 470580 579988 470608
rect 64380 470568 64386 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 548334 469820 548340 469872
rect 548392 469860 548398 469872
rect 568022 469860 568028 469872
rect 548392 469832 568028 469860
rect 548392 469820 548398 469832
rect 568022 469820 568028 469832
rect 568080 469820 568086 469872
rect 212350 469412 212356 469464
rect 212408 469452 212414 469464
rect 232682 469452 232688 469464
rect 212408 469424 232688 469452
rect 212408 469412 212414 469424
rect 232682 469412 232688 469424
rect 232740 469412 232746 469464
rect 296346 469412 296352 469464
rect 296404 469452 296410 469464
rect 316770 469452 316776 469464
rect 296404 469424 316776 469452
rect 296404 469412 296410 469424
rect 316770 469412 316776 469424
rect 316828 469412 316834 469464
rect 408034 469412 408040 469464
rect 408092 469452 408098 469464
rect 428642 469452 428648 469464
rect 408092 469424 428648 469452
rect 408092 469412 408098 469424
rect 428642 469412 428648 469424
rect 428700 469412 428706 469464
rect 148318 469344 148324 469396
rect 148376 469384 148382 469396
rect 165706 469384 165712 469396
rect 148376 469356 165712 469384
rect 148376 469344 148382 469356
rect 165706 469344 165712 469356
rect 165764 469344 165770 469396
rect 175458 469344 175464 469396
rect 175516 469384 175522 469396
rect 193674 469384 193680 469396
rect 175516 469356 193680 469384
rect 175516 469344 175522 469356
rect 193674 469344 193680 469356
rect 193732 469344 193738 469396
rect 203518 469344 203524 469396
rect 203576 469384 203582 469396
rect 221366 469384 221372 469396
rect 203576 469356 221372 469384
rect 203576 469344 203582 469356
rect 221366 469344 221372 469356
rect 221424 469344 221430 469396
rect 260098 469344 260104 469396
rect 260156 469384 260162 469396
rect 277670 469384 277676 469396
rect 260156 469356 277676 469384
rect 260156 469344 260162 469356
rect 277670 469344 277676 469356
rect 277728 469344 277734 469396
rect 287514 469344 287520 469396
rect 287572 469384 287578 469396
rect 305362 469384 305368 469396
rect 287572 469356 305368 469384
rect 287572 469344 287578 469356
rect 305362 469344 305368 469356
rect 305420 469344 305426 469396
rect 345658 469344 345664 469396
rect 345716 469384 345722 469396
rect 361666 469384 361672 469396
rect 345716 469356 361672 469384
rect 345716 469344 345722 469356
rect 361666 469344 361672 469356
rect 361724 469344 361730 469396
rect 371510 469344 371516 469396
rect 371568 469384 371574 469396
rect 389358 469384 389364 469396
rect 371568 469356 389364 469384
rect 371568 469344 371574 469356
rect 389358 469344 389364 469356
rect 389416 469344 389422 469396
rect 399478 469344 399484 469396
rect 399536 469384 399542 469396
rect 417694 469384 417700 469396
rect 399536 469356 417700 469384
rect 399536 469344 399542 469356
rect 417694 469344 417700 469356
rect 417752 469344 417758 469396
rect 456150 469344 456156 469396
rect 456208 469384 456214 469396
rect 473354 469384 473360 469396
rect 456208 469356 473360 469384
rect 456208 469344 456214 469356
rect 473354 469344 473360 469356
rect 473412 469344 473418 469396
rect 483474 469344 483480 469396
rect 483532 469384 483538 469396
rect 501690 469384 501696 469396
rect 483532 469356 501696 469384
rect 483532 469344 483538 469356
rect 501690 469344 501696 469356
rect 501748 469344 501754 469396
rect 511442 469344 511448 469396
rect 511500 469384 511506 469396
rect 529658 469384 529664 469396
rect 511500 469356 529664 469384
rect 511500 469344 511506 469356
rect 529658 469344 529664 469356
rect 529716 469344 529722 469396
rect 36722 469276 36728 469328
rect 36780 469316 36786 469328
rect 53650 469316 53656 469328
rect 36780 469288 53656 469316
rect 36780 469276 36786 469288
rect 53650 469276 53656 469288
rect 53708 469276 53714 469328
rect 64414 469276 64420 469328
rect 64472 469316 64478 469328
rect 81434 469316 81440 469328
rect 64472 469288 81440 469316
rect 64472 469276 64478 469288
rect 81434 469276 81440 469288
rect 81492 469276 81498 469328
rect 91462 469276 91468 469328
rect 91520 469316 91526 469328
rect 109678 469316 109684 469328
rect 91520 469288 109684 469316
rect 91520 469276 91526 469288
rect 109678 469276 109684 469288
rect 109736 469276 109742 469328
rect 119430 469276 119436 469328
rect 119488 469316 119494 469328
rect 137646 469316 137652 469328
rect 119488 469288 137652 469316
rect 119488 469276 119494 469288
rect 137646 469276 137652 469288
rect 137704 469276 137710 469328
rect 156322 469276 156328 469328
rect 156380 469316 156386 469328
rect 178678 469316 178684 469328
rect 156380 469288 178684 469316
rect 156380 469276 156386 469288
rect 178678 469276 178684 469288
rect 178736 469276 178742 469328
rect 232590 469276 232596 469328
rect 232648 469316 232654 469328
rect 249702 469316 249708 469328
rect 232648 469288 249708 469316
rect 232648 469276 232654 469288
rect 249702 469276 249708 469288
rect 249760 469276 249766 469328
rect 268010 469276 268016 469328
rect 268068 469316 268074 469328
rect 287698 469316 287704 469328
rect 268068 469288 287704 469316
rect 268068 469276 268074 469288
rect 287698 469276 287704 469288
rect 287756 469276 287762 469328
rect 315482 469276 315488 469328
rect 315540 469316 315546 469328
rect 333698 469316 333704 469328
rect 315540 469288 333704 469316
rect 315540 469276 315546 469288
rect 333698 469276 333704 469288
rect 333756 469276 333762 469328
rect 352006 469276 352012 469328
rect 352064 469316 352070 469328
rect 374638 469316 374644 469328
rect 352064 469288 374644 469316
rect 352064 469276 352070 469288
rect 374638 469276 374644 469288
rect 374696 469276 374702 469328
rect 428458 469276 428464 469328
rect 428516 469316 428522 469328
rect 445662 469316 445668 469328
rect 428516 469288 445668 469316
rect 428516 469276 428522 469288
rect 445662 469276 445668 469288
rect 445720 469276 445726 469328
rect 464338 469276 464344 469328
rect 464396 469316 464402 469328
rect 483658 469316 483664 469328
rect 464396 469288 483664 469316
rect 464396 469276 464402 469288
rect 483658 469276 483664 469288
rect 483716 469276 483722 469328
rect 492030 469276 492036 469328
rect 492088 469316 492094 469328
rect 512730 469316 512736 469328
rect 492088 469288 512736 469316
rect 492088 469276 492094 469288
rect 512730 469276 512736 469288
rect 512788 469276 512794 469328
rect 541618 469276 541624 469328
rect 541676 469316 541682 469328
rect 557534 469316 557540 469328
rect 541676 469288 557540 469316
rect 541676 469276 541682 469288
rect 557534 469276 557540 469288
rect 557592 469276 557598 469328
rect 15654 469208 15660 469260
rect 15712 469248 15718 469260
rect 25682 469248 25688 469260
rect 15712 469220 25688 469248
rect 15712 469208 15718 469220
rect 25682 469208 25688 469220
rect 25740 469208 25746 469260
rect 36630 469208 36636 469260
rect 36688 469248 36694 469260
rect 63310 469248 63316 469260
rect 36688 469220 63316 469248
rect 36688 469208 36694 469220
rect 63310 469208 63316 469220
rect 63368 469208 63374 469260
rect 66898 469208 66904 469260
rect 66956 469248 66962 469260
rect 91094 469248 91100 469260
rect 66956 469220 91100 469248
rect 66956 469208 66962 469220
rect 91094 469208 91100 469220
rect 91152 469208 91158 469260
rect 93118 469208 93124 469260
rect 93176 469248 93182 469260
rect 119338 469248 119344 469260
rect 93176 469220 119344 469248
rect 93176 469208 93182 469220
rect 119338 469208 119344 469220
rect 119396 469208 119402 469260
rect 124858 469208 124864 469260
rect 124916 469248 124922 469260
rect 147306 469248 147312 469260
rect 124916 469220 147312 469248
rect 124916 469208 124922 469220
rect 147306 469208 147312 469220
rect 147364 469208 147370 469260
rect 148410 469208 148416 469260
rect 148468 469248 148474 469260
rect 175366 469248 175372 469260
rect 148468 469220 175372 469248
rect 148468 469208 148474 469220
rect 175366 469208 175372 469220
rect 175424 469208 175430 469260
rect 177298 469208 177304 469260
rect 177356 469248 177362 469260
rect 203334 469248 203340 469260
rect 177356 469220 203340 469248
rect 177356 469208 177362 469220
rect 203334 469208 203340 469220
rect 203392 469208 203398 469260
rect 204990 469208 204996 469260
rect 205048 469248 205054 469260
rect 231026 469248 231032 469260
rect 205048 469220 231032 469248
rect 205048 469208 205054 469220
rect 231026 469208 231032 469220
rect 231084 469208 231090 469260
rect 232498 469208 232504 469260
rect 232556 469248 232562 469260
rect 259362 469248 259368 469260
rect 232556 469220 259368 469248
rect 232556 469208 232562 469220
rect 259362 469208 259368 469220
rect 259420 469208 259426 469260
rect 260190 469208 260196 469260
rect 260248 469248 260254 469260
rect 287330 469248 287336 469260
rect 260248 469220 287336 469248
rect 260248 469208 260254 469220
rect 287330 469208 287336 469220
rect 287388 469208 287394 469260
rect 289078 469208 289084 469260
rect 289136 469248 289142 469260
rect 315022 469248 315028 469260
rect 289136 469220 315028 469248
rect 289136 469208 289142 469220
rect 315022 469208 315028 469220
rect 315080 469208 315086 469260
rect 316678 469208 316684 469260
rect 316736 469248 316742 469260
rect 343358 469248 343364 469260
rect 316736 469220 343364 469248
rect 316736 469208 316742 469220
rect 343358 469208 343364 469220
rect 343416 469208 343422 469260
rect 344278 469208 344284 469260
rect 344336 469248 344342 469260
rect 371326 469248 371332 469260
rect 344336 469220 371332 469248
rect 344336 469208 344342 469220
rect 371326 469208 371332 469220
rect 371384 469208 371390 469260
rect 373258 469208 373264 469260
rect 373316 469248 373322 469260
rect 399018 469248 399024 469260
rect 373316 469220 399024 469248
rect 373316 469208 373322 469220
rect 399018 469208 399024 469220
rect 399076 469208 399082 469260
rect 400858 469208 400864 469260
rect 400916 469248 400922 469260
rect 427354 469248 427360 469260
rect 400916 469220 427360 469248
rect 400916 469208 400922 469220
rect 427354 469208 427360 469220
rect 427412 469208 427418 469260
rect 428550 469208 428556 469260
rect 428608 469248 428614 469260
rect 455322 469248 455328 469260
rect 428608 469220 455328 469248
rect 428608 469208 428614 469220
rect 455322 469208 455328 469220
rect 455380 469208 455386 469260
rect 456058 469208 456064 469260
rect 456116 469248 456122 469260
rect 483014 469248 483020 469260
rect 456116 469220 483020 469248
rect 456116 469208 456122 469220
rect 483014 469208 483020 469220
rect 483072 469208 483078 469260
rect 485038 469208 485044 469260
rect 485096 469248 485102 469260
rect 511350 469248 511356 469260
rect 485096 469220 511356 469248
rect 485096 469208 485102 469220
rect 511350 469208 511356 469220
rect 511408 469208 511414 469260
rect 512638 469208 512644 469260
rect 512696 469248 512702 469260
rect 539318 469248 539324 469260
rect 512696 469220 539324 469248
rect 512696 469208 512702 469220
rect 539318 469208 539324 469220
rect 539376 469208 539382 469260
rect 540238 469208 540244 469260
rect 540296 469248 540302 469260
rect 567194 469248 567200 469260
rect 540296 469220 567200 469248
rect 540296 469208 540302 469220
rect 567194 469208 567200 469220
rect 567252 469208 567258 469260
rect 15286 467236 15292 467288
rect 15344 467276 15350 467288
rect 15930 467276 15936 467288
rect 15344 467248 15936 467276
rect 15344 467236 15350 467248
rect 15930 467236 15936 467248
rect 15988 467236 15994 467288
rect 182082 466556 182088 466608
rect 182140 466596 182146 466608
rect 233234 466596 233240 466608
rect 182140 466568 233240 466596
rect 182140 466556 182146 466568
rect 233234 466556 233240 466568
rect 233292 466556 233298 466608
rect 350442 466556 350448 466608
rect 350500 466596 350506 466608
rect 401594 466596 401600 466608
rect 350500 466568 401600 466596
rect 350500 466556 350506 466568
rect 401594 466556 401600 466568
rect 401652 466556 401658 466608
rect 462222 466556 462228 466608
rect 462280 466596 462286 466608
rect 513374 466596 513380 466608
rect 462280 466568 513380 466596
rect 462280 466556 462286 466568
rect 513374 466556 513380 466568
rect 513432 466556 513438 466608
rect 42702 466488 42708 466540
rect 42760 466528 42766 466540
rect 93854 466528 93860 466540
rect 42760 466500 93860 466528
rect 42760 466488 42766 466500
rect 93854 466488 93860 466500
rect 93912 466488 93918 466540
rect 97902 466488 97908 466540
rect 97960 466528 97966 466540
rect 149054 466528 149060 466540
rect 97960 466500 149060 466528
rect 97960 466488 97966 466500
rect 149054 466488 149060 466500
rect 149112 466488 149118 466540
rect 154482 466488 154488 466540
rect 154540 466528 154546 466540
rect 205634 466528 205640 466540
rect 154540 466500 205640 466528
rect 154540 466488 154546 466500
rect 205634 466488 205640 466500
rect 205692 466488 205698 466540
rect 238662 466488 238668 466540
rect 238720 466528 238726 466540
rect 289814 466528 289820 466540
rect 238720 466500 289820 466528
rect 238720 466488 238726 466500
rect 289814 466488 289820 466500
rect 289872 466488 289878 466540
rect 293862 466488 293868 466540
rect 293920 466528 293926 466540
rect 345014 466528 345020 466540
rect 293920 466500 345020 466528
rect 293920 466488 293926 466500
rect 345014 466488 345020 466500
rect 345072 466488 345078 466540
rect 378042 466488 378048 466540
rect 378100 466528 378106 466540
rect 429286 466528 429292 466540
rect 378100 466500 429292 466528
rect 378100 466488 378106 466500
rect 429286 466488 429292 466500
rect 429344 466488 429350 466540
rect 434622 466488 434628 466540
rect 434680 466528 434686 466540
rect 485774 466528 485780 466540
rect 434680 466500 485780 466528
rect 434680 466488 434686 466500
rect 485774 466488 485780 466500
rect 485832 466488 485838 466540
rect 518802 466488 518808 466540
rect 518860 466528 518866 466540
rect 569954 466528 569960 466540
rect 518860 466500 569960 466528
rect 518860 466488 518866 466500
rect 569954 466488 569960 466500
rect 570012 466488 570018 466540
rect 13538 466420 13544 466472
rect 13596 466460 13602 466472
rect 66254 466460 66260 466472
rect 13596 466432 66260 466460
rect 13596 466420 13602 466432
rect 66254 466420 66260 466432
rect 66312 466420 66318 466472
rect 70302 466420 70308 466472
rect 70360 466460 70366 466472
rect 121454 466460 121460 466472
rect 70360 466432 121460 466460
rect 70360 466420 70366 466432
rect 121454 466420 121460 466432
rect 121512 466420 121518 466472
rect 126882 466420 126888 466472
rect 126940 466460 126946 466472
rect 178034 466460 178040 466472
rect 126940 466432 178040 466460
rect 126940 466420 126946 466432
rect 178034 466420 178040 466432
rect 178092 466420 178098 466472
rect 209682 466420 209688 466472
rect 209740 466460 209746 466472
rect 262214 466460 262220 466472
rect 209740 466432 262220 466460
rect 209740 466420 209746 466432
rect 262214 466420 262220 466432
rect 262272 466420 262278 466472
rect 266262 466420 266268 466472
rect 266320 466460 266326 466472
rect 317414 466460 317420 466472
rect 266320 466432 317420 466460
rect 266320 466420 266326 466432
rect 317414 466420 317420 466432
rect 317472 466420 317478 466472
rect 322842 466420 322848 466472
rect 322900 466460 322906 466472
rect 373994 466460 374000 466472
rect 322900 466432 374000 466460
rect 322900 466420 322906 466432
rect 373994 466420 374000 466432
rect 374052 466420 374058 466472
rect 405642 466420 405648 466472
rect 405700 466460 405706 466472
rect 458174 466460 458180 466472
rect 405700 466432 458180 466460
rect 405700 466420 405706 466432
rect 458174 466420 458180 466432
rect 458232 466420 458238 466472
rect 489822 466420 489828 466472
rect 489880 466460 489886 466472
rect 542354 466460 542360 466472
rect 489880 466432 542360 466460
rect 489880 466420 489886 466432
rect 542354 466420 542360 466432
rect 542412 466420 542418 466472
rect 42886 464040 42892 464092
rect 42944 464080 42950 464092
rect 43622 464080 43628 464092
rect 42944 464052 43628 464080
rect 42944 464040 42950 464052
rect 43622 464040 43628 464052
rect 43680 464040 43686 464092
rect 428642 450508 428648 450560
rect 428700 450548 428706 450560
rect 435726 450548 435732 450560
rect 428700 450520 435732 450548
rect 428700 450508 428706 450520
rect 435726 450508 435732 450520
rect 435784 450508 435790 450560
rect 512730 450440 512736 450492
rect 512788 450480 512794 450492
rect 519630 450480 519636 450492
rect 512788 450452 519636 450480
rect 512788 450440 512794 450452
rect 519630 450440 519636 450452
rect 519688 450440 519694 450492
rect 483658 450304 483664 450356
rect 483716 450344 483722 450356
rect 491662 450344 491668 450356
rect 483716 450316 491668 450344
rect 483716 450304 483722 450316
rect 491662 450304 491668 450316
rect 491720 450304 491726 450356
rect 232682 449896 232688 449948
rect 232740 449936 232746 449948
rect 239766 449936 239772 449948
rect 232740 449908 239772 449936
rect 232740 449896 232746 449908
rect 239766 449896 239772 449908
rect 239824 449896 239830 449948
rect 287698 449896 287704 449948
rect 287756 449936 287762 449948
rect 295702 449936 295708 449948
rect 287756 449908 295708 449936
rect 287756 449896 287762 449908
rect 295702 449896 295708 449908
rect 295760 449896 295766 449948
rect 316770 449896 316776 449948
rect 316828 449936 316834 449948
rect 323670 449936 323676 449948
rect 316828 449908 323676 449936
rect 316828 449896 316834 449908
rect 323670 449896 323676 449908
rect 323728 449896 323734 449948
rect 63586 449624 63592 449676
rect 63644 449664 63650 449676
rect 64414 449664 64420 449676
rect 63644 449636 64420 449664
rect 63644 449624 63650 449636
rect 64414 449624 64420 449636
rect 64472 449624 64478 449676
rect 455690 449624 455696 449676
rect 455748 449664 455754 449676
rect 456150 449664 456156 449676
rect 455748 449636 456156 449664
rect 455748 449624 455754 449636
rect 456150 449624 456156 449636
rect 456208 449624 456214 449676
rect 15838 448672 15844 448724
rect 15896 448712 15902 448724
rect 16666 448712 16672 448724
rect 15896 448684 16672 448712
rect 15896 448672 15902 448684
rect 16666 448672 16672 448684
rect 16724 448672 16730 448724
rect 2774 448604 2780 448656
rect 2832 448644 2838 448656
rect 4890 448644 4896 448656
rect 2832 448616 4896 448644
rect 2832 448604 2838 448616
rect 4890 448604 4896 448616
rect 4948 448604 4954 448656
rect 35250 448468 35256 448520
rect 35308 448508 35314 448520
rect 36722 448508 36728 448520
rect 35308 448480 36728 448508
rect 35308 448468 35314 448480
rect 36722 448468 36728 448480
rect 36780 448468 36786 448520
rect 231670 448468 231676 448520
rect 231728 448508 231734 448520
rect 232590 448508 232596 448520
rect 231728 448480 232596 448508
rect 231728 448468 231734 448480
rect 232590 448468 232596 448480
rect 232648 448468 232654 448520
rect 343634 448468 343640 448520
rect 343692 448508 343698 448520
rect 345658 448508 345664 448520
rect 343692 448480 345664 448508
rect 343692 448468 343698 448480
rect 345658 448468 345664 448480
rect 345716 448468 345722 448520
rect 539502 448468 539508 448520
rect 539560 448508 539566 448520
rect 541618 448508 541624 448520
rect 539560 448480 541624 448508
rect 539560 448468 539566 448480
rect 541618 448468 541624 448480
rect 541676 448468 541682 448520
rect 547874 448468 547880 448520
rect 547932 448508 547938 448520
rect 548150 448508 548156 448520
rect 547932 448480 548156 448508
rect 547932 448468 547938 448480
rect 548150 448468 548156 448480
rect 548208 448468 548214 448520
rect 71866 445680 71872 445732
rect 71924 445720 71930 445732
rect 100018 445720 100024 445732
rect 71924 445692 100024 445720
rect 71924 445680 71930 445692
rect 100018 445680 100024 445692
rect 100076 445680 100082 445732
rect 127986 445720 127992 445732
rect 103486 445692 127992 445720
rect 25682 445612 25688 445664
rect 25740 445652 25746 445664
rect 36630 445652 36636 445664
rect 25740 445624 36636 445652
rect 25740 445612 25746 445624
rect 36630 445612 36636 445624
rect 36688 445612 36694 445664
rect 42886 445612 42892 445664
rect 42944 445652 42950 445664
rect 42944 445624 45554 445652
rect 42944 445612 42950 445624
rect 15286 445544 15292 445596
rect 15344 445584 15350 445596
rect 43990 445584 43996 445596
rect 15344 445556 43996 445584
rect 15344 445544 15350 445556
rect 43990 445544 43996 445556
rect 44048 445544 44054 445596
rect 45526 445584 45554 445624
rect 53650 445612 53656 445664
rect 53708 445652 53714 445664
rect 66898 445652 66904 445664
rect 53708 445624 66904 445652
rect 53708 445612 53714 445624
rect 66898 445612 66904 445624
rect 66956 445612 66962 445664
rect 81986 445612 81992 445664
rect 82044 445652 82050 445664
rect 93118 445652 93124 445664
rect 82044 445624 93124 445652
rect 82044 445612 82050 445624
rect 93118 445612 93124 445624
rect 93176 445612 93182 445664
rect 99466 445612 99472 445664
rect 99524 445652 99530 445664
rect 103486 445652 103514 445692
rect 127986 445680 127992 445692
rect 128044 445680 128050 445732
rect 165982 445680 165988 445732
rect 166040 445720 166046 445732
rect 177298 445720 177304 445732
rect 166040 445692 177304 445720
rect 166040 445680 166046 445692
rect 177298 445680 177304 445692
rect 177356 445680 177362 445732
rect 178678 445680 178684 445732
rect 178736 445720 178742 445732
rect 184014 445720 184020 445732
rect 178736 445692 184020 445720
rect 178736 445680 178742 445692
rect 184014 445680 184020 445692
rect 184072 445680 184078 445732
rect 211706 445720 211712 445732
rect 190426 445692 211712 445720
rect 99524 445624 103514 445652
rect 99524 445612 99530 445624
rect 109678 445612 109684 445664
rect 109736 445652 109742 445664
rect 124858 445652 124864 445664
rect 109736 445624 124864 445652
rect 109736 445612 109742 445624
rect 124858 445612 124864 445624
rect 124916 445612 124922 445664
rect 137646 445612 137652 445664
rect 137704 445652 137710 445664
rect 148410 445652 148416 445664
rect 137704 445624 148416 445652
rect 137704 445612 137710 445624
rect 148410 445612 148416 445624
rect 148468 445612 148474 445664
rect 183646 445612 183652 445664
rect 183704 445652 183710 445664
rect 190426 445652 190454 445692
rect 211706 445680 211712 445692
rect 211764 445680 211770 445732
rect 222010 445680 222016 445732
rect 222068 445720 222074 445732
rect 232498 445720 232504 445732
rect 222068 445692 232504 445720
rect 222068 445680 222074 445692
rect 232498 445680 232504 445692
rect 232556 445680 232562 445732
rect 277670 445680 277676 445732
rect 277728 445720 277734 445732
rect 289078 445720 289084 445732
rect 277728 445692 289084 445720
rect 277728 445680 277734 445692
rect 289078 445680 289084 445692
rect 289136 445680 289142 445732
rect 306006 445680 306012 445732
rect 306064 445720 306070 445732
rect 316678 445720 316684 445732
rect 306064 445692 316684 445720
rect 306064 445680 306070 445692
rect 316678 445680 316684 445692
rect 316736 445680 316742 445732
rect 361666 445680 361672 445732
rect 361724 445720 361730 445732
rect 373258 445720 373264 445732
rect 361724 445692 373264 445720
rect 361724 445680 361730 445692
rect 373258 445680 373264 445692
rect 373316 445680 373322 445732
rect 379606 445680 379612 445732
rect 379664 445720 379670 445732
rect 408034 445720 408040 445732
rect 379664 445692 408040 445720
rect 379664 445680 379670 445692
rect 408034 445680 408040 445692
rect 408092 445680 408098 445732
rect 473998 445680 474004 445732
rect 474056 445720 474062 445732
rect 485038 445720 485044 445732
rect 474056 445692 485044 445720
rect 474056 445680 474062 445692
rect 485038 445680 485044 445692
rect 485096 445680 485102 445732
rect 501690 445680 501696 445732
rect 501748 445720 501754 445732
rect 512638 445720 512644 445732
rect 501748 445692 512644 445720
rect 501748 445680 501754 445692
rect 512638 445680 512644 445692
rect 512696 445680 512702 445732
rect 548150 445680 548156 445732
rect 548208 445720 548214 445732
rect 557534 445720 557540 445732
rect 548208 445692 557540 445720
rect 548208 445680 548214 445692
rect 557534 445680 557540 445692
rect 557592 445680 557598 445732
rect 183704 445624 190454 445652
rect 183704 445612 183710 445624
rect 193674 445612 193680 445664
rect 193732 445652 193738 445664
rect 204990 445652 204996 445664
rect 193732 445624 204996 445652
rect 193732 445612 193738 445624
rect 204990 445612 204996 445624
rect 205048 445612 205054 445664
rect 249702 445612 249708 445664
rect 249760 445652 249766 445664
rect 260190 445652 260196 445664
rect 249760 445624 260196 445652
rect 249760 445612 249766 445624
rect 260190 445612 260196 445624
rect 260248 445612 260254 445664
rect 333698 445612 333704 445664
rect 333756 445652 333762 445664
rect 344278 445652 344284 445664
rect 333756 445624 344284 445652
rect 333756 445612 333762 445624
rect 344278 445612 344284 445624
rect 344336 445612 344342 445664
rect 374638 445612 374644 445664
rect 374696 445652 374702 445664
rect 379698 445652 379704 445664
rect 374696 445624 379704 445652
rect 374696 445612 374702 445624
rect 379698 445612 379704 445624
rect 379756 445612 379762 445664
rect 390002 445612 390008 445664
rect 390060 445652 390066 445664
rect 400858 445652 400864 445664
rect 390060 445624 400864 445652
rect 390060 445612 390066 445624
rect 400858 445612 400864 445624
rect 400916 445612 400922 445664
rect 417694 445612 417700 445664
rect 417752 445652 417758 445664
rect 428550 445652 428556 445664
rect 417752 445624 428556 445652
rect 417752 445612 417758 445624
rect 428550 445612 428556 445624
rect 428608 445612 428614 445664
rect 445662 445612 445668 445664
rect 445720 445652 445726 445664
rect 456058 445652 456064 445664
rect 445720 445624 456064 445652
rect 445720 445612 445726 445624
rect 456058 445612 456064 445624
rect 456116 445612 456122 445664
rect 529658 445612 529664 445664
rect 529716 445652 529722 445664
rect 540238 445652 540244 445664
rect 529716 445624 540244 445652
rect 529716 445612 529722 445624
rect 540238 445612 540244 445624
rect 540296 445612 540302 445664
rect 72050 445584 72056 445596
rect 45526 445556 72056 445584
rect 72050 445544 72056 445556
rect 72108 445544 72114 445596
rect 127066 445544 127072 445596
rect 127124 445584 127130 445596
rect 156046 445584 156052 445596
rect 127124 445556 156052 445584
rect 127124 445544 127130 445556
rect 156046 445544 156052 445556
rect 156104 445544 156110 445596
rect 238846 445544 238852 445596
rect 238904 445584 238910 445596
rect 268010 445584 268016 445596
rect 238904 445556 268016 445584
rect 238904 445544 238910 445556
rect 268010 445544 268016 445556
rect 268068 445544 268074 445596
rect 323026 445544 323032 445596
rect 323084 445584 323090 445596
rect 352006 445584 352012 445596
rect 323084 445556 352012 445584
rect 323084 445544 323090 445556
rect 352006 445544 352012 445556
rect 352064 445544 352070 445596
rect 434806 445544 434812 445596
rect 434864 445584 434870 445596
rect 463694 445584 463700 445596
rect 434864 445556 463700 445584
rect 434864 445544 434870 445556
rect 463694 445544 463700 445556
rect 463752 445544 463758 445596
rect 518986 445544 518992 445596
rect 519044 445584 519050 445596
rect 547874 445584 547880 445596
rect 519044 445556 547880 445584
rect 519044 445544 519050 445556
rect 547874 445544 547880 445556
rect 547932 445544 547938 445596
rect 26602 443368 26608 443420
rect 26660 443408 26666 443420
rect 35434 443408 35440 443420
rect 26660 443380 35440 443408
rect 26660 443368 26666 443380
rect 35434 443368 35440 443380
rect 35492 443368 35498 443420
rect 71130 443096 71136 443148
rect 71188 443136 71194 443148
rect 82262 443136 82268 443148
rect 71188 443108 82268 443136
rect 71188 443096 71194 443108
rect 82262 443096 82268 443108
rect 82320 443096 82326 443148
rect 99374 443096 99380 443148
rect 99432 443136 99438 443148
rect 100294 443136 100300 443148
rect 99432 443108 100300 443136
rect 99432 443096 99438 443108
rect 100294 443096 100300 443108
rect 100352 443096 100358 443148
rect 183646 443096 183652 443148
rect 183704 443136 183710 443148
rect 222194 443136 222200 443148
rect 183704 443108 222200 443136
rect 183704 443096 183710 443108
rect 222194 443096 222200 443108
rect 222252 443096 222258 443148
rect 266998 443096 267004 443148
rect 267056 443136 267062 443148
rect 277946 443136 277952 443148
rect 267056 443108 277952 443136
rect 267056 443096 267062 443108
rect 277946 443096 277952 443108
rect 278004 443096 278010 443148
rect 295426 443096 295432 443148
rect 295484 443136 295490 443148
rect 334250 443136 334256 443148
rect 295484 443108 334256 443136
rect 295484 443096 295490 443108
rect 334250 443096 334256 443108
rect 334308 443096 334314 443148
rect 352006 443096 352012 443148
rect 352064 443136 352070 443148
rect 352064 443108 364334 443136
rect 352064 443096 352070 443108
rect 36630 443028 36636 443080
rect 36688 443068 36694 443080
rect 53926 443068 53932 443080
rect 36688 443040 53932 443068
rect 36688 443028 36694 443040
rect 53926 443028 53932 443040
rect 53984 443028 53990 443080
rect 71866 443028 71872 443080
rect 71924 443068 71930 443080
rect 109954 443068 109960 443080
rect 71924 443040 109960 443068
rect 71924 443028 71930 443040
rect 109954 443028 109960 443040
rect 110012 443028 110018 443080
rect 124858 443028 124864 443080
rect 124916 443068 124922 443080
rect 128354 443068 128360 443080
rect 124916 443040 128360 443068
rect 124916 443028 124922 443040
rect 128354 443028 128360 443040
rect 128412 443028 128418 443080
rect 151078 443028 151084 443080
rect 151136 443068 151142 443080
rect 156598 443068 156604 443080
rect 151136 443040 156604 443068
rect 151136 443028 151142 443040
rect 156598 443028 156604 443040
rect 156656 443028 156662 443080
rect 182818 443028 182824 443080
rect 182876 443068 182882 443080
rect 193950 443068 193956 443080
rect 182876 443040 193956 443068
rect 182876 443028 182882 443040
rect 193950 443028 193956 443040
rect 194008 443028 194014 443080
rect 232498 443028 232504 443080
rect 232556 443068 232562 443080
rect 232556 443040 248414 443068
rect 232556 443028 232562 443040
rect 66898 442960 66904 443012
rect 66956 443000 66962 443012
rect 72602 443000 72608 443012
rect 66956 442972 72608 443000
rect 66956 442960 66962 442972
rect 72602 442960 72608 442972
rect 72660 442960 72666 443012
rect 93118 442960 93124 443012
rect 93176 443000 93182 443012
rect 99374 443000 99380 443012
rect 93176 442972 99380 443000
rect 93176 442960 93182 442972
rect 99374 442960 99380 442972
rect 99432 442960 99438 443012
rect 99466 442960 99472 443012
rect 99524 443000 99530 443012
rect 138014 443000 138020 443012
rect 99524 442972 138020 443000
rect 99524 442960 99530 442972
rect 138014 442960 138020 442972
rect 138072 442960 138078 443012
rect 149698 442960 149704 443012
rect 149756 443000 149762 443012
rect 166258 443000 166264 443012
rect 149756 442972 166264 443000
rect 149756 442960 149762 442972
rect 166258 442960 166264 442972
rect 166316 442960 166322 443012
rect 177298 442960 177304 443012
rect 177356 443000 177362 443012
rect 184290 443000 184296 443012
rect 177356 442972 184296 443000
rect 177356 442960 177362 442972
rect 184290 442960 184296 442972
rect 184348 442960 184354 443012
rect 233970 442960 233976 443012
rect 234028 443000 234034 443012
rect 240594 443000 240600 443012
rect 234028 442972 240600 443000
rect 234028 442960 234034 442972
rect 240594 442960 240600 442972
rect 240652 442960 240658 443012
rect 248386 443000 248414 443040
rect 267826 443028 267832 443080
rect 267884 443068 267890 443080
rect 306282 443068 306288 443080
rect 267884 443040 306288 443068
rect 267884 443028 267890 443040
rect 306282 443028 306288 443040
rect 306340 443028 306346 443080
rect 345658 443028 345664 443080
rect 345716 443068 345722 443080
rect 361942 443068 361948 443080
rect 345716 443040 361948 443068
rect 345716 443028 345722 443040
rect 361942 443028 361948 443040
rect 362000 443028 362006 443080
rect 364306 443068 364334 443108
rect 379606 443096 379612 443148
rect 379664 443136 379670 443148
rect 418246 443136 418252 443148
rect 379664 443108 418252 443136
rect 379664 443096 379670 443108
rect 418246 443096 418252 443108
rect 418304 443096 418310 443148
rect 462958 443096 462964 443148
rect 463016 443136 463022 443148
rect 474274 443136 474280 443148
rect 463016 443108 474280 443136
rect 463016 443096 463022 443108
rect 474274 443096 474280 443108
rect 474332 443096 474338 443148
rect 485038 443096 485044 443148
rect 485096 443136 485102 443148
rect 492582 443136 492588 443148
rect 485096 443108 492588 443136
rect 485096 443096 485102 443108
rect 492582 443096 492588 443108
rect 492640 443096 492646 443148
rect 390278 443068 390284 443080
rect 364306 443040 390284 443068
rect 390278 443028 390284 443040
rect 390336 443028 390342 443080
rect 400858 443028 400864 443080
rect 400916 443068 400922 443080
rect 408586 443068 408592 443080
rect 400916 443040 408592 443068
rect 400916 443028 400922 443040
rect 408586 443028 408592 443040
rect 408644 443028 408650 443080
rect 429838 443028 429844 443080
rect 429896 443068 429902 443080
rect 436278 443068 436284 443080
rect 429896 443040 436284 443068
rect 429896 443028 429902 443040
rect 436278 443028 436284 443040
rect 436336 443028 436342 443080
rect 463786 443028 463792 443080
rect 463844 443068 463850 443080
rect 502242 443068 502248 443080
rect 463844 443040 502248 443068
rect 463844 443028 463850 443040
rect 502242 443028 502248 443040
rect 502300 443028 502306 443080
rect 514018 443028 514024 443080
rect 514076 443068 514082 443080
rect 520274 443068 520280 443080
rect 514076 443040 520280 443068
rect 514076 443028 514082 443040
rect 520274 443028 520280 443040
rect 520332 443028 520338 443080
rect 250254 443000 250260 443012
rect 248386 442972 250260 443000
rect 250254 442960 250260 442972
rect 250312 442960 250318 443012
rect 261478 442960 261484 443012
rect 261536 443000 261542 443012
rect 268286 443000 268292 443012
rect 261536 442972 268292 443000
rect 261536 442960 261542 442972
rect 268286 442960 268292 442972
rect 268344 442960 268350 443012
rect 289078 442960 289084 443012
rect 289136 443000 289142 443012
rect 296622 443000 296628 443012
rect 289136 442972 296628 443000
rect 289136 442960 289142 442972
rect 296622 442960 296628 442972
rect 296680 442960 296686 443012
rect 318058 442960 318064 443012
rect 318116 443000 318122 443012
rect 324590 443000 324596 443012
rect 318116 442972 324596 443000
rect 318116 442960 318122 442972
rect 324590 442960 324596 442972
rect 324648 442960 324654 443012
rect 347038 442960 347044 443012
rect 347096 443000 347102 443012
rect 352282 443000 352288 443012
rect 347096 442972 352288 443000
rect 347096 442960 347102 442972
rect 352282 442960 352288 442972
rect 352340 442960 352346 443012
rect 373258 442960 373264 443012
rect 373316 443000 373322 443012
rect 380618 443000 380624 443012
rect 373316 442972 380624 443000
rect 373316 442960 373322 442972
rect 380618 442960 380624 442972
rect 380676 442960 380682 443012
rect 428458 442960 428464 443012
rect 428516 443000 428522 443012
rect 445938 443000 445944 443012
rect 428516 442972 445944 443000
rect 428516 442960 428522 442972
rect 445938 442960 445944 442972
rect 445996 442960 446002 443012
rect 457438 442960 457444 443012
rect 457496 443000 457502 443012
rect 464614 443000 464620 443012
rect 457496 442972 464620 443000
rect 457496 442960 457502 442972
rect 464614 442960 464620 442972
rect 464672 442960 464678 443012
rect 491386 442960 491392 443012
rect 491444 443000 491450 443012
rect 529934 443000 529940 443012
rect 491444 442972 529940 443000
rect 491444 442960 491450 442972
rect 529934 442960 529940 442972
rect 529992 442960 529998 443012
rect 541618 442960 541624 443012
rect 541676 443000 541682 443012
rect 558270 443000 558276 443012
rect 541676 442972 558276 443000
rect 541676 442960 541682 442972
rect 558270 442960 558276 442972
rect 558328 442960 558334 443012
rect 210418 441600 210424 441652
rect 210476 441640 210482 441652
rect 212534 441640 212540 441652
rect 210476 441612 212540 441640
rect 210476 441600 210482 441612
rect 212534 441600 212540 441612
rect 212592 441600 212598 441652
rect 42702 440240 42708 440292
rect 42760 440280 42766 440292
rect 93854 440280 93860 440292
rect 42760 440252 93860 440280
rect 42760 440240 42766 440252
rect 93854 440240 93860 440252
rect 93912 440240 93918 440292
rect 97902 440240 97908 440292
rect 97960 440280 97966 440292
rect 149054 440280 149060 440292
rect 97960 440252 149060 440280
rect 97960 440240 97966 440252
rect 149054 440240 149060 440252
rect 149112 440240 149118 440292
rect 154482 440240 154488 440292
rect 154540 440280 154546 440292
rect 205634 440280 205640 440292
rect 154540 440252 205640 440280
rect 154540 440240 154546 440252
rect 205634 440240 205640 440252
rect 205692 440240 205698 440292
rect 209682 440240 209688 440292
rect 209740 440280 209746 440292
rect 262214 440280 262220 440292
rect 209740 440252 262220 440280
rect 209740 440240 209746 440252
rect 262214 440240 262220 440252
rect 262272 440240 262278 440292
rect 266262 440240 266268 440292
rect 266320 440280 266326 440292
rect 317414 440280 317420 440292
rect 266320 440252 317420 440280
rect 266320 440240 266326 440252
rect 317414 440240 317420 440252
rect 317472 440240 317478 440292
rect 322842 440240 322848 440292
rect 322900 440280 322906 440292
rect 373994 440280 374000 440292
rect 322900 440252 374000 440280
rect 322900 440240 322906 440252
rect 373994 440240 374000 440252
rect 374052 440240 374058 440292
rect 378042 440240 378048 440292
rect 378100 440280 378106 440292
rect 429286 440280 429292 440292
rect 378100 440252 429292 440280
rect 378100 440240 378106 440252
rect 429286 440240 429292 440252
rect 429344 440240 429350 440292
rect 434622 440240 434628 440292
rect 434680 440280 434686 440292
rect 485774 440280 485780 440292
rect 434680 440252 485780 440280
rect 434680 440240 434686 440252
rect 485774 440240 485780 440252
rect 485832 440240 485838 440292
rect 489822 440240 489828 440292
rect 489880 440280 489886 440292
rect 542354 440280 542360 440292
rect 489880 440252 542360 440280
rect 489880 440240 489886 440252
rect 542354 440240 542360 440252
rect 542412 440240 542418 440292
rect 544378 440240 544384 440292
rect 544436 440280 544442 440292
rect 548334 440280 548340 440292
rect 544436 440252 548340 440280
rect 544436 440240 544442 440252
rect 548334 440240 548340 440252
rect 548392 440240 548398 440292
rect 120258 440172 120264 440224
rect 120316 440212 120322 440224
rect 122098 440212 122104 440224
rect 120316 440184 122104 440212
rect 120316 440172 120322 440184
rect 122098 440172 122104 440184
rect 122156 440172 122162 440224
rect 204254 436092 204260 436144
rect 204312 436132 204318 436144
rect 204990 436132 204996 436144
rect 204312 436104 204996 436132
rect 204312 436092 204318 436104
rect 204990 436092 204996 436104
rect 205048 436092 205054 436144
rect 400306 436092 400312 436144
rect 400364 436132 400370 436144
rect 400950 436132 400956 436144
rect 400364 436104 400956 436132
rect 400364 436092 400370 436104
rect 400950 436092 400956 436104
rect 401008 436092 401014 436144
rect 13538 422220 13544 422272
rect 13596 422260 13602 422272
rect 66254 422260 66260 422272
rect 13596 422232 66260 422260
rect 13596 422220 13602 422232
rect 66254 422220 66260 422232
rect 66312 422220 66318 422272
rect 70302 422220 70308 422272
rect 70360 422260 70366 422272
rect 121454 422260 121460 422272
rect 70360 422232 121460 422260
rect 70360 422220 70366 422232
rect 121454 422220 121460 422232
rect 121512 422220 121518 422272
rect 126882 422220 126888 422272
rect 126940 422260 126946 422272
rect 178034 422260 178040 422272
rect 126940 422232 178040 422260
rect 126940 422220 126946 422232
rect 178034 422220 178040 422232
rect 178092 422220 178098 422272
rect 182082 422220 182088 422272
rect 182140 422260 182146 422272
rect 233234 422260 233240 422272
rect 182140 422232 233240 422260
rect 182140 422220 182146 422232
rect 233234 422220 233240 422232
rect 233292 422220 233298 422272
rect 238662 422220 238668 422272
rect 238720 422260 238726 422272
rect 289814 422260 289820 422272
rect 238720 422232 289820 422260
rect 238720 422220 238726 422232
rect 289814 422220 289820 422232
rect 289872 422220 289878 422272
rect 293862 422220 293868 422272
rect 293920 422260 293926 422272
rect 345014 422260 345020 422272
rect 293920 422232 345020 422260
rect 293920 422220 293926 422232
rect 345014 422220 345020 422232
rect 345072 422220 345078 422272
rect 350442 422220 350448 422272
rect 350500 422260 350506 422272
rect 401594 422260 401600 422272
rect 350500 422232 401600 422260
rect 350500 422220 350506 422232
rect 401594 422220 401600 422232
rect 401652 422220 401658 422272
rect 405642 422220 405648 422272
rect 405700 422260 405706 422272
rect 458174 422260 458180 422272
rect 405700 422232 458180 422260
rect 405700 422220 405706 422232
rect 458174 422220 458180 422232
rect 458232 422220 458238 422272
rect 462222 422220 462228 422272
rect 462280 422260 462286 422272
rect 513374 422260 513380 422272
rect 462280 422232 513380 422260
rect 462280 422220 462286 422232
rect 513374 422220 513380 422232
rect 513432 422220 513438 422272
rect 518802 422220 518808 422272
rect 518860 422260 518866 422272
rect 569954 422260 569960 422272
rect 518860 422232 569960 422260
rect 518860 422220 518866 422232
rect 569954 422220 569960 422232
rect 570012 422220 570018 422272
rect 15194 419432 15200 419484
rect 15252 419472 15258 419484
rect 35894 419472 35900 419484
rect 15252 419444 35900 419472
rect 15252 419432 15258 419444
rect 35894 419432 35900 419444
rect 35952 419432 35958 419484
rect 36078 419432 36084 419484
rect 36136 419472 36142 419484
rect 63586 419472 63592 419484
rect 36136 419444 63592 419472
rect 36136 419432 36142 419444
rect 63586 419432 63592 419444
rect 63644 419432 63650 419484
rect 64046 419432 64052 419484
rect 64104 419472 64110 419484
rect 91922 419472 91928 419484
rect 64104 419444 91928 419472
rect 64104 419432 64110 419444
rect 91922 419432 91928 419444
rect 91980 419432 91986 419484
rect 92106 419432 92112 419484
rect 92164 419472 92170 419484
rect 119614 419472 119620 419484
rect 92164 419444 119620 419472
rect 92164 419432 92170 419444
rect 119614 419432 119620 419444
rect 119672 419432 119678 419484
rect 122098 419432 122104 419484
rect 122156 419472 122162 419484
rect 147950 419472 147956 419484
rect 122156 419444 147956 419472
rect 122156 419432 122162 419444
rect 147950 419432 147956 419444
rect 148008 419432 148014 419484
rect 148042 419432 148048 419484
rect 148100 419472 148106 419484
rect 175918 419472 175924 419484
rect 148100 419444 175924 419472
rect 148100 419432 148106 419444
rect 175918 419432 175924 419444
rect 175976 419432 175982 419484
rect 176102 419432 176108 419484
rect 176160 419472 176166 419484
rect 203610 419472 203616 419484
rect 176160 419444 203616 419472
rect 176160 419432 176166 419444
rect 203610 419432 203616 419444
rect 203668 419432 203674 419484
rect 204990 419432 204996 419484
rect 205048 419472 205054 419484
rect 231946 419472 231952 419484
rect 205048 419444 231952 419472
rect 205048 419432 205054 419444
rect 231946 419432 231952 419444
rect 232004 419432 232010 419484
rect 232038 419432 232044 419484
rect 232096 419472 232102 419484
rect 259914 419472 259920 419484
rect 232096 419444 259920 419472
rect 232096 419432 232102 419444
rect 259914 419432 259920 419444
rect 259972 419432 259978 419484
rect 260098 419432 260104 419484
rect 260156 419472 260162 419484
rect 287606 419472 287612 419484
rect 260156 419444 287612 419472
rect 260156 419432 260162 419444
rect 287606 419432 287612 419444
rect 287664 419432 287670 419484
rect 288066 419432 288072 419484
rect 288124 419472 288130 419484
rect 315942 419472 315948 419484
rect 288124 419444 315948 419472
rect 288124 419432 288130 419444
rect 315942 419432 315948 419444
rect 316000 419432 316006 419484
rect 316678 419432 316684 419484
rect 316736 419472 316742 419484
rect 343910 419472 343916 419484
rect 316736 419444 343916 419472
rect 316736 419432 316742 419444
rect 343910 419432 343916 419444
rect 343968 419432 343974 419484
rect 344094 419432 344100 419484
rect 344152 419472 344158 419484
rect 371602 419472 371608 419484
rect 344152 419444 371608 419472
rect 344152 419432 344158 419444
rect 371602 419432 371608 419444
rect 371660 419432 371666 419484
rect 372062 419432 372068 419484
rect 372120 419472 372126 419484
rect 399938 419472 399944 419484
rect 372120 419444 399944 419472
rect 372120 419432 372126 419444
rect 399938 419432 399944 419444
rect 399996 419432 400002 419484
rect 400950 419432 400956 419484
rect 401008 419472 401014 419484
rect 427906 419472 427912 419484
rect 401008 419444 427912 419472
rect 401008 419432 401014 419444
rect 427906 419432 427912 419444
rect 427964 419432 427970 419484
rect 428090 419432 428096 419484
rect 428148 419472 428154 419484
rect 455598 419472 455604 419484
rect 428148 419444 455604 419472
rect 428148 419432 428154 419444
rect 455598 419432 455604 419444
rect 455656 419432 455662 419484
rect 456058 419432 456064 419484
rect 456116 419472 456122 419484
rect 483934 419472 483940 419484
rect 456116 419444 483940 419472
rect 456116 419432 456122 419444
rect 483934 419432 483940 419444
rect 483992 419432 483998 419484
rect 484026 419432 484032 419484
rect 484084 419472 484090 419484
rect 511902 419472 511908 419484
rect 484084 419444 511908 419472
rect 484084 419432 484090 419444
rect 511902 419432 511908 419444
rect 511960 419432 511966 419484
rect 512086 419432 512092 419484
rect 512144 419472 512150 419484
rect 539594 419472 539600 419484
rect 512144 419444 539600 419472
rect 512144 419432 512150 419444
rect 539594 419432 539600 419444
rect 539652 419432 539658 419484
rect 540054 419432 540060 419484
rect 540112 419472 540118 419484
rect 567930 419472 567936 419484
rect 540112 419444 567936 419472
rect 540112 419432 540118 419444
rect 567930 419432 567936 419444
rect 567988 419432 567994 419484
rect 16574 419364 16580 419416
rect 16632 419404 16638 419416
rect 36630 419404 36636 419416
rect 16632 419376 36636 419404
rect 16632 419364 16638 419376
rect 36630 419364 36636 419376
rect 36688 419364 36694 419416
rect 44910 419364 44916 419416
rect 44968 419404 44974 419416
rect 71130 419404 71136 419416
rect 44968 419376 71136 419404
rect 44968 419364 44974 419376
rect 71130 419364 71136 419376
rect 71188 419364 71194 419416
rect 82262 419364 82268 419416
rect 82320 419404 82326 419416
rect 93118 419404 93124 419416
rect 82320 419376 93124 419404
rect 82320 419364 82326 419376
rect 93118 419364 93124 419376
rect 93176 419364 93182 419416
rect 110230 419364 110236 419416
rect 110288 419404 110294 419416
rect 124858 419404 124864 419416
rect 110288 419376 124864 419404
rect 110288 419364 110294 419376
rect 124858 419364 124864 419376
rect 124916 419364 124922 419416
rect 128630 419364 128636 419416
rect 128688 419404 128694 419416
rect 149698 419404 149704 419416
rect 128688 419376 149704 419404
rect 128688 419364 128694 419376
rect 149698 419364 149704 419376
rect 149756 419364 149762 419416
rect 156598 419364 156604 419416
rect 156656 419404 156662 419416
rect 182818 419404 182824 419416
rect 156656 419376 182824 419404
rect 156656 419364 156662 419376
rect 182818 419364 182824 419376
rect 182876 419364 182882 419416
rect 194502 419364 194508 419416
rect 194560 419404 194566 419416
rect 210418 419404 210424 419416
rect 194560 419376 210424 419404
rect 194560 419364 194566 419376
rect 210418 419364 210424 419376
rect 210476 419364 210482 419416
rect 212626 419364 212632 419416
rect 212684 419404 212690 419416
rect 232498 419404 232504 419416
rect 212684 419376 232504 419404
rect 212684 419364 212690 419376
rect 232498 419364 232504 419376
rect 232556 419364 232562 419416
rect 240594 419364 240600 419416
rect 240652 419404 240658 419416
rect 266998 419404 267004 419416
rect 240652 419376 267004 419404
rect 240652 419364 240658 419376
rect 266998 419364 267004 419376
rect 267056 419364 267062 419416
rect 278590 419364 278596 419416
rect 278648 419404 278654 419416
rect 289078 419404 289084 419416
rect 278648 419376 289084 419404
rect 278648 419364 278654 419376
rect 289078 419364 289084 419376
rect 289136 419364 289142 419416
rect 306282 419364 306288 419416
rect 306340 419404 306346 419416
rect 318058 419404 318064 419416
rect 306340 419376 318064 419404
rect 306340 419364 306346 419376
rect 318058 419364 318064 419376
rect 318116 419364 318122 419416
rect 324590 419364 324596 419416
rect 324648 419404 324654 419416
rect 345658 419404 345664 419416
rect 324648 419376 345664 419404
rect 324648 419364 324654 419376
rect 345658 419364 345664 419376
rect 345716 419364 345722 419416
rect 362586 419364 362592 419416
rect 362644 419404 362650 419416
rect 373258 419404 373264 419416
rect 362644 419376 373264 419404
rect 362644 419364 362650 419376
rect 373258 419364 373264 419376
rect 373316 419364 373322 419416
rect 390278 419364 390284 419416
rect 390336 419404 390342 419416
rect 400858 419404 400864 419416
rect 390336 419376 400864 419404
rect 390336 419364 390342 419376
rect 400858 419364 400864 419376
rect 400916 419364 400922 419416
rect 408586 419364 408592 419416
rect 408644 419404 408650 419416
rect 428458 419404 428464 419416
rect 408644 419376 428464 419404
rect 408644 419364 408650 419376
rect 428458 419364 428464 419376
rect 428516 419364 428522 419416
rect 436922 419364 436928 419416
rect 436980 419404 436986 419416
rect 462958 419404 462964 419416
rect 436980 419376 462964 419404
rect 436980 419364 436986 419376
rect 462958 419364 462964 419376
rect 463016 419364 463022 419416
rect 474274 419364 474280 419416
rect 474332 419404 474338 419416
rect 485038 419404 485044 419416
rect 474332 419376 485044 419404
rect 474332 419364 474338 419376
rect 485038 419364 485044 419376
rect 485096 419364 485102 419416
rect 502242 419364 502248 419416
rect 502300 419404 502306 419416
rect 514018 419404 514024 419416
rect 502300 419376 514024 419404
rect 502300 419364 502306 419376
rect 514018 419364 514024 419376
rect 514076 419364 514082 419416
rect 520918 419364 520924 419416
rect 520976 419404 520982 419416
rect 541618 419404 541624 419416
rect 520976 419376 541624 419404
rect 520976 419364 520982 419376
rect 541618 419364 541624 419376
rect 541676 419364 541682 419416
rect 26234 419296 26240 419348
rect 26292 419336 26298 419348
rect 43530 419336 43536 419348
rect 26292 419308 43536 419336
rect 26292 419296 26298 419308
rect 43530 419296 43536 419308
rect 43588 419296 43594 419348
rect 54570 419296 54576 419348
rect 54628 419336 54634 419348
rect 66898 419336 66904 419348
rect 54628 419308 66904 419336
rect 54628 419296 54634 419308
rect 66898 419296 66904 419308
rect 66956 419296 66962 419348
rect 138290 419296 138296 419348
rect 138348 419336 138354 419348
rect 151078 419336 151084 419348
rect 138348 419308 151084 419336
rect 138348 419296 138354 419308
rect 151078 419296 151084 419308
rect 151136 419296 151142 419348
rect 166258 419296 166264 419348
rect 166316 419336 166322 419348
rect 177298 419336 177304 419348
rect 166316 419308 177304 419336
rect 166316 419296 166322 419308
rect 177298 419296 177304 419308
rect 177356 419296 177362 419348
rect 222286 419296 222292 419348
rect 222344 419336 222350 419348
rect 233970 419336 233976 419348
rect 222344 419308 233976 419336
rect 222344 419296 222350 419308
rect 233970 419296 233976 419308
rect 234028 419296 234034 419348
rect 250254 419296 250260 419348
rect 250312 419336 250318 419348
rect 261478 419336 261484 419348
rect 250312 419308 261484 419336
rect 250312 419296 250318 419308
rect 261478 419296 261484 419308
rect 261536 419296 261542 419348
rect 334250 419296 334256 419348
rect 334308 419336 334314 419348
rect 347038 419336 347044 419348
rect 334308 419308 347044 419336
rect 334308 419296 334314 419308
rect 347038 419296 347044 419308
rect 347096 419296 347102 419348
rect 418246 419296 418252 419348
rect 418304 419336 418310 419348
rect 429838 419336 429844 419348
rect 418304 419308 429844 419336
rect 418304 419296 418310 419308
rect 429838 419296 429844 419308
rect 429896 419296 429902 419348
rect 446582 419296 446588 419348
rect 446640 419336 446646 419348
rect 457438 419336 457444 419348
rect 446640 419308 457444 419336
rect 446640 419296 446646 419308
rect 457438 419296 457444 419308
rect 457496 419296 457502 419348
rect 530578 419296 530584 419348
rect 530636 419336 530642 419348
rect 544378 419336 544384 419348
rect 530636 419308 544384 419336
rect 530636 419296 530642 419308
rect 544378 419296 544384 419308
rect 544436 419296 544442 419348
rect 558270 418752 558276 418804
rect 558328 418792 558334 418804
rect 567470 418792 567476 418804
rect 558328 418764 567476 418792
rect 558328 418752 558334 418764
rect 567470 418752 567476 418764
rect 567528 418752 567534 418804
rect 548334 416032 548340 416084
rect 548392 416072 548398 416084
rect 568022 416072 568028 416084
rect 548392 416044 568028 416072
rect 548392 416032 548398 416044
rect 568022 416032 568028 416044
rect 568080 416032 568086 416084
rect 212350 415624 212356 415676
rect 212408 415664 212414 415676
rect 232682 415664 232688 415676
rect 212408 415636 232688 415664
rect 212408 415624 212414 415636
rect 232682 415624 232688 415636
rect 232740 415624 232746 415676
rect 296346 415624 296352 415676
rect 296404 415664 296410 415676
rect 316770 415664 316776 415676
rect 296404 415636 316776 415664
rect 296404 415624 296410 415636
rect 316770 415624 316776 415636
rect 316828 415624 316834 415676
rect 408034 415624 408040 415676
rect 408092 415664 408098 415676
rect 428642 415664 428648 415676
rect 408092 415636 428648 415664
rect 408092 415624 408098 415636
rect 428642 415624 428648 415636
rect 428700 415624 428706 415676
rect 119430 415556 119436 415608
rect 119488 415596 119494 415608
rect 137646 415596 137652 415608
rect 119488 415568 137652 415596
rect 119488 415556 119494 415568
rect 137646 415556 137652 415568
rect 137704 415556 137710 415608
rect 148318 415556 148324 415608
rect 148376 415596 148382 415608
rect 165706 415596 165712 415608
rect 148376 415568 165712 415596
rect 148376 415556 148382 415568
rect 165706 415556 165712 415568
rect 165764 415556 165770 415608
rect 175458 415556 175464 415608
rect 175516 415596 175522 415608
rect 193674 415596 193680 415608
rect 175516 415568 193680 415596
rect 175516 415556 175522 415568
rect 193674 415556 193680 415568
rect 193732 415556 193738 415608
rect 203518 415556 203524 415608
rect 203576 415596 203582 415608
rect 221366 415596 221372 415608
rect 203576 415568 221372 415596
rect 203576 415556 203582 415568
rect 221366 415556 221372 415568
rect 221424 415556 221430 415608
rect 260098 415556 260104 415608
rect 260156 415596 260162 415608
rect 277670 415596 277676 415608
rect 260156 415568 277676 415596
rect 260156 415556 260162 415568
rect 277670 415556 277676 415568
rect 277728 415556 277734 415608
rect 287514 415556 287520 415608
rect 287572 415596 287578 415608
rect 305362 415596 305368 415608
rect 287572 415568 305368 415596
rect 287572 415556 287578 415568
rect 305362 415556 305368 415568
rect 305420 415556 305426 415608
rect 345658 415556 345664 415608
rect 345716 415596 345722 415608
rect 361666 415596 361672 415608
rect 345716 415568 361672 415596
rect 345716 415556 345722 415568
rect 361666 415556 361672 415568
rect 361724 415556 361730 415608
rect 371510 415556 371516 415608
rect 371568 415596 371574 415608
rect 389358 415596 389364 415608
rect 371568 415568 389364 415596
rect 371568 415556 371574 415568
rect 389358 415556 389364 415568
rect 389416 415556 389422 415608
rect 399478 415556 399484 415608
rect 399536 415596 399542 415608
rect 417694 415596 417700 415608
rect 399536 415568 417700 415596
rect 399536 415556 399542 415568
rect 417694 415556 417700 415568
rect 417752 415556 417758 415608
rect 456058 415556 456064 415608
rect 456116 415596 456122 415608
rect 473354 415596 473360 415608
rect 456116 415568 473360 415596
rect 456116 415556 456122 415568
rect 473354 415556 473360 415568
rect 473412 415556 473418 415608
rect 483474 415556 483480 415608
rect 483532 415596 483538 415608
rect 501690 415596 501696 415608
rect 483532 415568 501696 415596
rect 483532 415556 483538 415568
rect 501690 415556 501696 415568
rect 501748 415556 501754 415608
rect 511442 415556 511448 415608
rect 511500 415596 511506 415608
rect 529658 415596 529664 415608
rect 511500 415568 529664 415596
rect 511500 415556 511506 415568
rect 529658 415556 529664 415568
rect 529716 415556 529722 415608
rect 36722 415488 36728 415540
rect 36780 415528 36786 415540
rect 53650 415528 53656 415540
rect 36780 415500 53656 415528
rect 36780 415488 36786 415500
rect 53650 415488 53656 415500
rect 53708 415488 53714 415540
rect 64414 415488 64420 415540
rect 64472 415528 64478 415540
rect 81434 415528 81440 415540
rect 64472 415500 81440 415528
rect 64472 415488 64478 415500
rect 81434 415488 81440 415500
rect 81492 415488 81498 415540
rect 91462 415488 91468 415540
rect 91520 415528 91526 415540
rect 109678 415528 109684 415540
rect 91520 415500 109684 415528
rect 91520 415488 91526 415500
rect 109678 415488 109684 415500
rect 109736 415488 109742 415540
rect 127986 415488 127992 415540
rect 128044 415528 128050 415540
rect 148502 415528 148508 415540
rect 128044 415500 148508 415528
rect 128044 415488 128050 415500
rect 148502 415488 148508 415500
rect 148560 415488 148566 415540
rect 156322 415488 156328 415540
rect 156380 415528 156386 415540
rect 178678 415528 178684 415540
rect 156380 415500 178684 415528
rect 156380 415488 156386 415500
rect 178678 415488 178684 415500
rect 178736 415488 178742 415540
rect 232590 415488 232596 415540
rect 232648 415528 232654 415540
rect 249702 415528 249708 415540
rect 232648 415500 249708 415528
rect 232648 415488 232654 415500
rect 249702 415488 249708 415500
rect 249760 415488 249766 415540
rect 268010 415488 268016 415540
rect 268068 415528 268074 415540
rect 287698 415528 287704 415540
rect 268068 415500 287704 415528
rect 268068 415488 268074 415500
rect 287698 415488 287704 415500
rect 287756 415488 287762 415540
rect 315482 415488 315488 415540
rect 315540 415528 315546 415540
rect 333698 415528 333704 415540
rect 315540 415500 333704 415528
rect 315540 415488 315546 415500
rect 333698 415488 333704 415500
rect 333756 415488 333762 415540
rect 352006 415488 352012 415540
rect 352064 415528 352070 415540
rect 374638 415528 374644 415540
rect 352064 415500 374644 415528
rect 352064 415488 352070 415500
rect 374638 415488 374644 415500
rect 374696 415488 374702 415540
rect 428458 415488 428464 415540
rect 428516 415528 428522 415540
rect 445662 415528 445668 415540
rect 428516 415500 445668 415528
rect 428516 415488 428522 415500
rect 445662 415488 445668 415500
rect 445720 415488 445726 415540
rect 464338 415488 464344 415540
rect 464396 415528 464402 415540
rect 483658 415528 483664 415540
rect 464396 415500 483664 415528
rect 464396 415488 464402 415500
rect 483658 415488 483664 415500
rect 483716 415488 483722 415540
rect 492030 415488 492036 415540
rect 492088 415528 492094 415540
rect 512730 415528 512736 415540
rect 492088 415500 512736 415528
rect 492088 415488 492094 415500
rect 512730 415488 512736 415500
rect 512788 415488 512794 415540
rect 541618 415488 541624 415540
rect 541676 415528 541682 415540
rect 557534 415528 557540 415540
rect 541676 415500 557540 415528
rect 541676 415488 541682 415500
rect 557534 415488 557540 415500
rect 557592 415488 557598 415540
rect 15102 415420 15108 415472
rect 15160 415460 15166 415472
rect 25682 415460 25688 415472
rect 15160 415432 25688 415460
rect 15160 415420 15166 415432
rect 25682 415420 25688 415432
rect 25740 415420 25746 415472
rect 36630 415420 36636 415472
rect 36688 415460 36694 415472
rect 63310 415460 63316 415472
rect 36688 415432 63316 415460
rect 36688 415420 36694 415432
rect 63310 415420 63316 415432
rect 63368 415420 63374 415472
rect 66898 415420 66904 415472
rect 66956 415460 66962 415472
rect 91094 415460 91100 415472
rect 66956 415432 91100 415460
rect 66956 415420 66962 415432
rect 91094 415420 91100 415432
rect 91152 415420 91158 415472
rect 93118 415420 93124 415472
rect 93176 415460 93182 415472
rect 119338 415460 119344 415472
rect 93176 415432 119344 415460
rect 93176 415420 93182 415432
rect 119338 415420 119344 415432
rect 119396 415420 119402 415472
rect 122098 415420 122104 415472
rect 122156 415460 122162 415472
rect 147306 415460 147312 415472
rect 122156 415432 147312 415460
rect 122156 415420 122162 415432
rect 147306 415420 147312 415432
rect 147364 415420 147370 415472
rect 148410 415420 148416 415472
rect 148468 415460 148474 415472
rect 175366 415460 175372 415472
rect 148468 415432 175372 415460
rect 148468 415420 148474 415432
rect 175366 415420 175372 415432
rect 175424 415420 175430 415472
rect 177298 415420 177304 415472
rect 177356 415460 177362 415472
rect 203334 415460 203340 415472
rect 177356 415432 203340 415460
rect 177356 415420 177362 415432
rect 203334 415420 203340 415432
rect 203392 415420 203398 415472
rect 204990 415420 204996 415472
rect 205048 415460 205054 415472
rect 231026 415460 231032 415472
rect 205048 415432 231032 415460
rect 205048 415420 205054 415432
rect 231026 415420 231032 415432
rect 231084 415420 231090 415472
rect 232498 415420 232504 415472
rect 232556 415460 232562 415472
rect 259362 415460 259368 415472
rect 232556 415432 259368 415460
rect 232556 415420 232562 415432
rect 259362 415420 259368 415432
rect 259420 415420 259426 415472
rect 260190 415420 260196 415472
rect 260248 415460 260254 415472
rect 287330 415460 287336 415472
rect 260248 415432 287336 415460
rect 260248 415420 260254 415432
rect 287330 415420 287336 415432
rect 287388 415420 287394 415472
rect 289078 415420 289084 415472
rect 289136 415460 289142 415472
rect 315022 415460 315028 415472
rect 289136 415432 315028 415460
rect 289136 415420 289142 415432
rect 315022 415420 315028 415432
rect 315080 415420 315086 415472
rect 316678 415420 316684 415472
rect 316736 415460 316742 415472
rect 343358 415460 343364 415472
rect 316736 415432 343364 415460
rect 316736 415420 316742 415432
rect 343358 415420 343364 415432
rect 343416 415420 343422 415472
rect 344278 415420 344284 415472
rect 344336 415460 344342 415472
rect 371326 415460 371332 415472
rect 344336 415432 371332 415460
rect 344336 415420 344342 415432
rect 371326 415420 371332 415432
rect 371384 415420 371390 415472
rect 373258 415420 373264 415472
rect 373316 415460 373322 415472
rect 399018 415460 399024 415472
rect 373316 415432 399024 415460
rect 373316 415420 373322 415432
rect 399018 415420 399024 415432
rect 399076 415420 399082 415472
rect 400858 415420 400864 415472
rect 400916 415460 400922 415472
rect 427354 415460 427360 415472
rect 400916 415432 427360 415460
rect 400916 415420 400922 415432
rect 427354 415420 427360 415432
rect 427412 415420 427418 415472
rect 428550 415420 428556 415472
rect 428608 415460 428614 415472
rect 455322 415460 455328 415472
rect 428608 415432 455328 415460
rect 428608 415420 428614 415432
rect 455322 415420 455328 415432
rect 455380 415420 455386 415472
rect 456150 415420 456156 415472
rect 456208 415460 456214 415472
rect 483014 415460 483020 415472
rect 456208 415432 483020 415460
rect 456208 415420 456214 415432
rect 483014 415420 483020 415432
rect 483072 415420 483078 415472
rect 485038 415420 485044 415472
rect 485096 415460 485102 415472
rect 511350 415460 511356 415472
rect 485096 415432 511356 415460
rect 485096 415420 485102 415432
rect 511350 415420 511356 415432
rect 511408 415420 511414 415472
rect 512638 415420 512644 415472
rect 512696 415460 512702 415472
rect 539318 415460 539324 415472
rect 512696 415432 539324 415460
rect 512696 415420 512702 415432
rect 539318 415420 539324 415432
rect 539376 415420 539382 415472
rect 540238 415420 540244 415472
rect 540296 415460 540302 415472
rect 567194 415460 567200 415472
rect 540296 415432 567200 415460
rect 540296 415420 540302 415432
rect 567194 415420 567200 415432
rect 567252 415420 567258 415472
rect 3142 410320 3148 410372
rect 3200 410360 3206 410372
rect 8938 410360 8944 410372
rect 3200 410332 8944 410360
rect 3200 410320 3206 410332
rect 8938 410320 8944 410332
rect 8996 410320 9002 410372
rect 42886 405900 42892 405952
rect 42944 405940 42950 405952
rect 43622 405940 43628 405952
rect 42944 405912 43628 405940
rect 42944 405900 42950 405912
rect 43622 405900 43628 405912
rect 43680 405900 43686 405952
rect 148502 395292 148508 395344
rect 148560 395332 148566 395344
rect 155862 395332 155868 395344
rect 148560 395304 155868 395332
rect 148560 395292 148566 395304
rect 155862 395292 155868 395304
rect 155920 395292 155926 395344
rect 428642 395292 428648 395344
rect 428700 395332 428706 395344
rect 435726 395332 435732 395344
rect 428700 395304 435732 395332
rect 428700 395292 428706 395304
rect 435726 395292 435732 395304
rect 435784 395292 435790 395344
rect 287698 395088 287704 395140
rect 287756 395128 287762 395140
rect 295794 395128 295800 395140
rect 287756 395100 295800 395128
rect 287756 395088 287762 395100
rect 295794 395088 295800 395100
rect 295852 395088 295858 395140
rect 316770 395088 316776 395140
rect 316828 395128 316834 395140
rect 323670 395128 323676 395140
rect 316828 395100 323676 395128
rect 316828 395088 316834 395100
rect 323670 395088 323676 395100
rect 323728 395088 323734 395140
rect 232682 395020 232688 395072
rect 232740 395060 232746 395072
rect 239766 395060 239772 395072
rect 232740 395032 239772 395060
rect 232740 395020 232746 395032
rect 239766 395020 239772 395032
rect 239824 395020 239830 395072
rect 483658 395020 483664 395072
rect 483716 395060 483722 395072
rect 491662 395060 491668 395072
rect 483716 395032 491668 395060
rect 483716 395020 483722 395032
rect 491662 395020 491668 395032
rect 491720 395020 491726 395072
rect 512730 395020 512736 395072
rect 512788 395060 512794 395072
rect 519630 395060 519636 395072
rect 512788 395032 519636 395060
rect 512788 395020 512794 395032
rect 519630 395020 519636 395032
rect 519688 395020 519694 395072
rect 547874 394680 547880 394732
rect 547932 394720 547938 394732
rect 548150 394720 548156 394732
rect 547932 394692 548156 394720
rect 547932 394680 547938 394692
rect 548150 394680 548156 394692
rect 548208 394680 548214 394732
rect 13538 394612 13544 394664
rect 13596 394652 13602 394664
rect 13596 394624 59952 394652
rect 13596 394612 13602 394624
rect 35250 394544 35256 394596
rect 35308 394584 35314 394596
rect 36722 394584 36728 394596
rect 35308 394556 36728 394584
rect 35308 394544 35314 394556
rect 36722 394544 36728 394556
rect 36780 394544 36786 394596
rect 42702 394544 42708 394596
rect 42760 394584 42766 394596
rect 42760 394556 45554 394584
rect 42760 394544 42766 394556
rect 45526 394448 45554 394556
rect 59924 394516 59952 394624
rect 63586 394612 63592 394664
rect 63644 394652 63650 394664
rect 64414 394652 64420 394664
rect 63644 394624 64420 394652
rect 63644 394612 63650 394624
rect 64414 394612 64420 394624
rect 64472 394612 64478 394664
rect 70302 394612 70308 394664
rect 70360 394652 70366 394664
rect 121454 394652 121460 394664
rect 70360 394624 121460 394652
rect 70360 394612 70366 394624
rect 121454 394612 121460 394624
rect 121512 394612 121518 394664
rect 126882 394612 126888 394664
rect 126940 394652 126946 394664
rect 178034 394652 178040 394664
rect 126940 394624 178040 394652
rect 126940 394612 126946 394624
rect 178034 394612 178040 394624
rect 178092 394612 178098 394664
rect 209682 394612 209688 394664
rect 209740 394652 209746 394664
rect 262214 394652 262220 394664
rect 209740 394624 262220 394652
rect 209740 394612 209746 394624
rect 262214 394612 262220 394624
rect 262272 394612 262278 394664
rect 266262 394612 266268 394664
rect 266320 394652 266326 394664
rect 317414 394652 317420 394664
rect 266320 394624 317420 394652
rect 266320 394612 266326 394624
rect 317414 394612 317420 394624
rect 317472 394612 317478 394664
rect 322842 394612 322848 394664
rect 322900 394652 322906 394664
rect 373994 394652 374000 394664
rect 322900 394624 374000 394652
rect 322900 394612 322906 394624
rect 373994 394612 374000 394624
rect 374052 394612 374058 394664
rect 405642 394612 405648 394664
rect 405700 394652 405706 394664
rect 458174 394652 458180 394664
rect 405700 394624 458180 394652
rect 405700 394612 405706 394624
rect 458174 394612 458180 394624
rect 458232 394612 458238 394664
rect 489822 394612 489828 394664
rect 489880 394652 489886 394664
rect 542354 394652 542360 394664
rect 489880 394624 542360 394652
rect 489880 394612 489886 394624
rect 542354 394612 542360 394624
rect 542412 394612 542418 394664
rect 93854 394584 93860 394596
rect 74506 394556 93860 394584
rect 66254 394516 66260 394528
rect 59924 394488 66260 394516
rect 66254 394476 66260 394488
rect 66312 394476 66318 394528
rect 74506 394448 74534 394556
rect 93854 394544 93860 394556
rect 93912 394544 93918 394596
rect 97902 394544 97908 394596
rect 97960 394584 97966 394596
rect 149054 394584 149060 394596
rect 97960 394556 149060 394584
rect 97960 394544 97966 394556
rect 149054 394544 149060 394556
rect 149112 394544 149118 394596
rect 182082 394544 182088 394596
rect 182140 394584 182146 394596
rect 233234 394584 233240 394596
rect 182140 394556 233240 394584
rect 182140 394544 182146 394556
rect 233234 394544 233240 394556
rect 233292 394544 233298 394596
rect 238662 394544 238668 394596
rect 238720 394584 238726 394596
rect 289814 394584 289820 394596
rect 238720 394556 289820 394584
rect 238720 394544 238726 394556
rect 289814 394544 289820 394556
rect 289872 394544 289878 394596
rect 293862 394544 293868 394596
rect 293920 394584 293926 394596
rect 293920 394556 335354 394584
rect 293920 394544 293926 394556
rect 154482 394476 154488 394528
rect 154540 394516 154546 394528
rect 205634 394516 205640 394528
rect 154540 394488 205640 394516
rect 154540 394476 154546 394488
rect 205634 394476 205640 394488
rect 205692 394476 205698 394528
rect 335326 394516 335354 394556
rect 343634 394544 343640 394596
rect 343692 394584 343698 394596
rect 345658 394584 345664 394596
rect 343692 394556 345664 394584
rect 343692 394544 343698 394556
rect 345658 394544 345664 394556
rect 345716 394544 345722 394596
rect 378042 394544 378048 394596
rect 378100 394584 378106 394596
rect 429286 394584 429292 394596
rect 378100 394556 429292 394584
rect 378100 394544 378106 394556
rect 429286 394544 429292 394556
rect 429344 394544 429350 394596
rect 462222 394544 462228 394596
rect 462280 394584 462286 394596
rect 513374 394584 513380 394596
rect 462280 394556 513380 394584
rect 462280 394544 462286 394556
rect 513374 394544 513380 394556
rect 513432 394544 513438 394596
rect 518802 394544 518808 394596
rect 518860 394584 518866 394596
rect 569954 394584 569960 394596
rect 518860 394556 569960 394584
rect 518860 394544 518866 394556
rect 569954 394544 569960 394556
rect 570012 394544 570018 394596
rect 345014 394516 345020 394528
rect 335326 394488 345020 394516
rect 345014 394476 345020 394488
rect 345072 394476 345078 394528
rect 350442 394476 350448 394528
rect 350500 394516 350506 394528
rect 401594 394516 401600 394528
rect 350500 394488 401600 394516
rect 350500 394476 350506 394488
rect 401594 394476 401600 394488
rect 401652 394476 401658 394528
rect 434622 394476 434628 394528
rect 434680 394516 434686 394528
rect 485774 394516 485780 394528
rect 434680 394488 485780 394516
rect 434680 394476 434686 394488
rect 485774 394476 485780 394488
rect 485832 394476 485838 394528
rect 45526 394420 74534 394448
rect 231578 393252 231584 393304
rect 231636 393292 231642 393304
rect 232590 393292 232596 393304
rect 231636 393264 232596 393292
rect 231636 393252 231642 393264
rect 232590 393252 232596 393264
rect 232648 393252 232654 393304
rect 539318 393252 539324 393304
rect 539376 393292 539382 393304
rect 541618 393292 541624 393304
rect 539376 393264 541624 393292
rect 539376 393252 539382 393264
rect 541618 393252 541624 393264
rect 541676 393252 541682 393304
rect 71866 391892 71872 391944
rect 71924 391932 71930 391944
rect 100018 391932 100024 391944
rect 71924 391904 100024 391932
rect 71924 391892 71930 391904
rect 100018 391892 100024 391904
rect 100076 391892 100082 391944
rect 127986 391932 127992 391944
rect 103486 391904 127992 391932
rect 25682 391824 25688 391876
rect 25740 391864 25746 391876
rect 36630 391864 36636 391876
rect 25740 391836 36636 391864
rect 25740 391824 25746 391836
rect 36630 391824 36636 391836
rect 36688 391824 36694 391876
rect 42886 391824 42892 391876
rect 42944 391864 42950 391876
rect 42944 391836 45554 391864
rect 42944 391824 42950 391836
rect 15286 391756 15292 391808
rect 15344 391796 15350 391808
rect 43990 391796 43996 391808
rect 15344 391768 43996 391796
rect 15344 391756 15350 391768
rect 43990 391756 43996 391768
rect 44048 391756 44054 391808
rect 45526 391796 45554 391836
rect 53650 391824 53656 391876
rect 53708 391864 53714 391876
rect 66898 391864 66904 391876
rect 53708 391836 66904 391864
rect 53708 391824 53714 391836
rect 66898 391824 66904 391836
rect 66956 391824 66962 391876
rect 81986 391824 81992 391876
rect 82044 391864 82050 391876
rect 93118 391864 93124 391876
rect 82044 391836 93124 391864
rect 82044 391824 82050 391836
rect 93118 391824 93124 391836
rect 93176 391824 93182 391876
rect 99466 391824 99472 391876
rect 99524 391864 99530 391876
rect 103486 391864 103514 391904
rect 127986 391892 127992 391904
rect 128044 391892 128050 391944
rect 165982 391892 165988 391944
rect 166040 391932 166046 391944
rect 177298 391932 177304 391944
rect 166040 391904 177304 391932
rect 166040 391892 166046 391904
rect 177298 391892 177304 391904
rect 177356 391892 177362 391944
rect 178678 391892 178684 391944
rect 178736 391932 178742 391944
rect 184014 391932 184020 391944
rect 178736 391904 184020 391932
rect 178736 391892 178742 391904
rect 184014 391892 184020 391904
rect 184072 391892 184078 391944
rect 211706 391932 211712 391944
rect 190426 391904 211712 391932
rect 99524 391836 103514 391864
rect 99524 391824 99530 391836
rect 109678 391824 109684 391876
rect 109736 391864 109742 391876
rect 122098 391864 122104 391876
rect 109736 391836 122104 391864
rect 109736 391824 109742 391836
rect 122098 391824 122104 391836
rect 122156 391824 122162 391876
rect 137646 391824 137652 391876
rect 137704 391864 137710 391876
rect 148410 391864 148416 391876
rect 137704 391836 148416 391864
rect 137704 391824 137710 391836
rect 148410 391824 148416 391836
rect 148468 391824 148474 391876
rect 183646 391824 183652 391876
rect 183704 391864 183710 391876
rect 190426 391864 190454 391904
rect 211706 391892 211712 391904
rect 211764 391892 211770 391944
rect 221918 391892 221924 391944
rect 221976 391932 221982 391944
rect 232498 391932 232504 391944
rect 221976 391904 232504 391932
rect 221976 391892 221982 391904
rect 232498 391892 232504 391904
rect 232556 391892 232562 391944
rect 277670 391892 277676 391944
rect 277728 391932 277734 391944
rect 289078 391932 289084 391944
rect 277728 391904 289084 391932
rect 277728 391892 277734 391904
rect 289078 391892 289084 391904
rect 289136 391892 289142 391944
rect 306006 391892 306012 391944
rect 306064 391932 306070 391944
rect 316678 391932 316684 391944
rect 306064 391904 316684 391932
rect 306064 391892 306070 391904
rect 316678 391892 316684 391904
rect 316736 391892 316742 391944
rect 361666 391892 361672 391944
rect 361724 391932 361730 391944
rect 373258 391932 373264 391944
rect 361724 391904 373264 391932
rect 361724 391892 361730 391904
rect 373258 391892 373264 391904
rect 373316 391892 373322 391944
rect 379606 391892 379612 391944
rect 379664 391932 379670 391944
rect 408034 391932 408040 391944
rect 379664 391904 408040 391932
rect 379664 391892 379670 391904
rect 408034 391892 408040 391904
rect 408092 391892 408098 391944
rect 473998 391892 474004 391944
rect 474056 391932 474062 391944
rect 485038 391932 485044 391944
rect 474056 391904 485044 391932
rect 474056 391892 474062 391904
rect 485038 391892 485044 391904
rect 485096 391892 485102 391944
rect 501690 391892 501696 391944
rect 501748 391932 501754 391944
rect 512638 391932 512644 391944
rect 501748 391904 512644 391932
rect 501748 391892 501754 391904
rect 512638 391892 512644 391904
rect 512696 391892 512702 391944
rect 548150 391892 548156 391944
rect 548208 391932 548214 391944
rect 557534 391932 557540 391944
rect 548208 391904 557540 391932
rect 548208 391892 548214 391904
rect 557534 391892 557540 391904
rect 557592 391892 557598 391944
rect 183704 391836 190454 391864
rect 183704 391824 183710 391836
rect 193674 391824 193680 391876
rect 193732 391864 193738 391876
rect 204990 391864 204996 391876
rect 193732 391836 204996 391864
rect 193732 391824 193738 391836
rect 204990 391824 204996 391836
rect 205048 391824 205054 391876
rect 249702 391824 249708 391876
rect 249760 391864 249766 391876
rect 260190 391864 260196 391876
rect 249760 391836 260196 391864
rect 249760 391824 249766 391836
rect 260190 391824 260196 391836
rect 260248 391824 260254 391876
rect 333698 391824 333704 391876
rect 333756 391864 333762 391876
rect 344278 391864 344284 391876
rect 333756 391836 344284 391864
rect 333756 391824 333762 391836
rect 344278 391824 344284 391836
rect 344336 391824 344342 391876
rect 374638 391824 374644 391876
rect 374696 391864 374702 391876
rect 379698 391864 379704 391876
rect 374696 391836 379704 391864
rect 374696 391824 374702 391836
rect 379698 391824 379704 391836
rect 379756 391824 379762 391876
rect 390002 391824 390008 391876
rect 390060 391864 390066 391876
rect 400858 391864 400864 391876
rect 390060 391836 400864 391864
rect 390060 391824 390066 391836
rect 400858 391824 400864 391836
rect 400916 391824 400922 391876
rect 417694 391824 417700 391876
rect 417752 391864 417758 391876
rect 428550 391864 428556 391876
rect 417752 391836 428556 391864
rect 417752 391824 417758 391836
rect 428550 391824 428556 391836
rect 428608 391824 428614 391876
rect 445662 391824 445668 391876
rect 445720 391864 445726 391876
rect 456150 391864 456156 391876
rect 445720 391836 456156 391864
rect 445720 391824 445726 391836
rect 456150 391824 456156 391836
rect 456208 391824 456214 391876
rect 529658 391824 529664 391876
rect 529716 391864 529722 391876
rect 540238 391864 540244 391876
rect 529716 391836 540244 391864
rect 529716 391824 529722 391836
rect 540238 391824 540244 391836
rect 540296 391824 540302 391876
rect 71958 391796 71964 391808
rect 45526 391768 71964 391796
rect 71958 391756 71964 391768
rect 72016 391756 72022 391808
rect 238846 391756 238852 391808
rect 238904 391796 238910 391808
rect 268010 391796 268016 391808
rect 238904 391768 268016 391796
rect 238904 391756 238910 391768
rect 268010 391756 268016 391768
rect 268068 391756 268074 391808
rect 323026 391756 323032 391808
rect 323084 391796 323090 391808
rect 352006 391796 352012 391808
rect 323084 391768 352012 391796
rect 323084 391756 323090 391768
rect 352006 391756 352012 391768
rect 352064 391756 352070 391808
rect 434806 391756 434812 391808
rect 434864 391796 434870 391808
rect 463786 391796 463792 391808
rect 434864 391768 463792 391796
rect 434864 391756 434870 391768
rect 463786 391756 463792 391768
rect 463844 391756 463850 391808
rect 518986 391756 518992 391808
rect 519044 391796 519050 391808
rect 547874 391796 547880 391808
rect 519044 391768 547880 391796
rect 519044 391756 519050 391768
rect 547874 391756 547880 391768
rect 547932 391756 547938 391808
rect 15102 390396 15108 390448
rect 15160 390436 15166 390448
rect 16574 390436 16580 390448
rect 15160 390408 16580 390436
rect 15160 390396 15166 390408
rect 16574 390396 16580 390408
rect 16632 390396 16638 390448
rect 26234 389784 26240 389836
rect 26292 389824 26298 389836
rect 35434 389824 35440 389836
rect 26292 389796 35440 389824
rect 26292 389784 26298 389796
rect 35434 389784 35440 389796
rect 35492 389784 35498 389836
rect 489886 389388 499574 389416
rect 71130 389308 71136 389360
rect 71188 389348 71194 389360
rect 82262 389348 82268 389360
rect 71188 389320 82268 389348
rect 71188 389308 71194 389320
rect 82262 389308 82268 389320
rect 82320 389308 82326 389360
rect 99466 389308 99472 389360
rect 99524 389348 99530 389360
rect 100386 389348 100392 389360
rect 99524 389320 100392 389348
rect 99524 389308 99530 389320
rect 100386 389308 100392 389320
rect 100444 389308 100450 389360
rect 183646 389308 183652 389360
rect 183704 389348 183710 389360
rect 222286 389348 222292 389360
rect 183704 389320 222292 389348
rect 183704 389308 183710 389320
rect 222286 389308 222292 389320
rect 222344 389308 222350 389360
rect 266998 389308 267004 389360
rect 267056 389348 267062 389360
rect 277946 389348 277952 389360
rect 267056 389320 277952 389348
rect 267056 389308 267062 389320
rect 277946 389308 277952 389320
rect 278004 389308 278010 389360
rect 295426 389308 295432 389360
rect 295484 389348 295490 389360
rect 334250 389348 334256 389360
rect 295484 389320 334256 389348
rect 295484 389308 295490 389320
rect 334250 389308 334256 389320
rect 334308 389308 334314 389360
rect 352006 389308 352012 389360
rect 352064 389348 352070 389360
rect 352064 389320 364334 389348
rect 352064 389308 352070 389320
rect 36630 389240 36636 389292
rect 36688 389280 36694 389292
rect 53926 389280 53932 389292
rect 36688 389252 53932 389280
rect 36688 389240 36694 389252
rect 53926 389240 53932 389252
rect 53984 389240 53990 389292
rect 71866 389240 71872 389292
rect 71924 389280 71930 389292
rect 109954 389280 109960 389292
rect 71924 389252 109960 389280
rect 71924 389240 71930 389252
rect 109954 389240 109960 389252
rect 110012 389240 110018 389292
rect 151078 389240 151084 389292
rect 151136 389280 151142 389292
rect 156598 389280 156604 389292
rect 151136 389252 156604 389280
rect 151136 389240 151142 389252
rect 156598 389240 156604 389252
rect 156656 389240 156662 389292
rect 182818 389240 182824 389292
rect 182876 389280 182882 389292
rect 193950 389280 193956 389292
rect 182876 389252 193956 389280
rect 182876 389240 182882 389252
rect 193950 389240 193956 389252
rect 194008 389240 194014 389292
rect 232498 389240 232504 389292
rect 232556 389280 232562 389292
rect 232556 389252 248414 389280
rect 232556 389240 232562 389252
rect 66898 389172 66904 389224
rect 66956 389212 66962 389224
rect 72602 389212 72608 389224
rect 66956 389184 72608 389212
rect 66956 389172 66962 389184
rect 72602 389172 72608 389184
rect 72660 389172 72666 389224
rect 93118 389172 93124 389224
rect 93176 389212 93182 389224
rect 100294 389212 100300 389224
rect 93176 389184 100300 389212
rect 93176 389172 93182 389184
rect 100294 389172 100300 389184
rect 100352 389172 100358 389224
rect 100386 389172 100392 389224
rect 100444 389212 100450 389224
rect 138290 389212 138296 389224
rect 100444 389184 138296 389212
rect 100444 389172 100450 389184
rect 138290 389172 138296 389184
rect 138348 389172 138354 389224
rect 149698 389172 149704 389224
rect 149756 389212 149762 389224
rect 166258 389212 166264 389224
rect 149756 389184 166264 389212
rect 149756 389172 149762 389184
rect 166258 389172 166264 389184
rect 166316 389172 166322 389224
rect 177298 389172 177304 389224
rect 177356 389212 177362 389224
rect 184290 389212 184296 389224
rect 177356 389184 184296 389212
rect 177356 389172 177362 389184
rect 184290 389172 184296 389184
rect 184348 389172 184354 389224
rect 233970 389172 233976 389224
rect 234028 389212 234034 389224
rect 240594 389212 240600 389224
rect 234028 389184 240600 389212
rect 234028 389172 234034 389184
rect 240594 389172 240600 389184
rect 240652 389172 240658 389224
rect 248386 389212 248414 389252
rect 267826 389240 267832 389292
rect 267884 389280 267890 389292
rect 306282 389280 306288 389292
rect 267884 389252 306288 389280
rect 267884 389240 267890 389252
rect 306282 389240 306288 389252
rect 306340 389240 306346 389292
rect 345658 389240 345664 389292
rect 345716 389280 345722 389292
rect 361942 389280 361948 389292
rect 345716 389252 361948 389280
rect 345716 389240 345722 389252
rect 361942 389240 361948 389252
rect 362000 389240 362006 389292
rect 364306 389280 364334 389320
rect 379606 389308 379612 389360
rect 379664 389348 379670 389360
rect 418246 389348 418252 389360
rect 379664 389320 418252 389348
rect 379664 389308 379670 389320
rect 418246 389308 418252 389320
rect 418304 389308 418310 389360
rect 463786 389308 463792 389360
rect 463844 389348 463850 389360
rect 463844 389320 470594 389348
rect 463844 389308 463850 389320
rect 390278 389280 390284 389292
rect 364306 389252 390284 389280
rect 390278 389240 390284 389252
rect 390336 389240 390342 389292
rect 400950 389240 400956 389292
rect 401008 389280 401014 389292
rect 408586 389280 408592 389292
rect 401008 389252 408592 389280
rect 401008 389240 401014 389252
rect 408586 389240 408592 389252
rect 408644 389240 408650 389292
rect 429838 389240 429844 389292
rect 429896 389280 429902 389292
rect 436278 389280 436284 389292
rect 429896 389252 436284 389280
rect 429896 389240 429902 389252
rect 436278 389240 436284 389252
rect 436336 389240 436342 389292
rect 457438 389240 457444 389292
rect 457496 389280 457502 389292
rect 464614 389280 464620 389292
rect 457496 389252 464620 389280
rect 457496 389240 457502 389252
rect 464614 389240 464620 389252
rect 464672 389240 464678 389292
rect 470566 389280 470594 389320
rect 489886 389280 489914 389388
rect 491386 389308 491392 389360
rect 491444 389348 491450 389360
rect 491444 389320 492812 389348
rect 491444 389308 491450 389320
rect 470566 389252 489914 389280
rect 250254 389212 250260 389224
rect 248386 389184 250260 389212
rect 250254 389172 250260 389184
rect 250312 389172 250318 389224
rect 261478 389172 261484 389224
rect 261536 389212 261542 389224
rect 268286 389212 268292 389224
rect 261536 389184 268292 389212
rect 261536 389172 261542 389184
rect 268286 389172 268292 389184
rect 268344 389172 268350 389224
rect 289078 389172 289084 389224
rect 289136 389212 289142 389224
rect 296622 389212 296628 389224
rect 289136 389184 296628 389212
rect 289136 389172 289142 389184
rect 296622 389172 296628 389184
rect 296680 389172 296686 389224
rect 318058 389172 318064 389224
rect 318116 389212 318122 389224
rect 324590 389212 324596 389224
rect 318116 389184 324596 389212
rect 318116 389172 318122 389184
rect 324590 389172 324596 389184
rect 324648 389172 324654 389224
rect 347038 389172 347044 389224
rect 347096 389212 347102 389224
rect 352282 389212 352288 389224
rect 347096 389184 352288 389212
rect 347096 389172 347102 389184
rect 352282 389172 352288 389184
rect 352340 389172 352346 389224
rect 373258 389172 373264 389224
rect 373316 389212 373322 389224
rect 380618 389212 380624 389224
rect 373316 389184 380624 389212
rect 373316 389172 373322 389184
rect 380618 389172 380624 389184
rect 380676 389172 380682 389224
rect 428458 389172 428464 389224
rect 428516 389212 428522 389224
rect 445938 389212 445944 389224
rect 428516 389184 445944 389212
rect 428516 389172 428522 389184
rect 445938 389172 445944 389184
rect 445996 389172 446002 389224
rect 462958 389172 462964 389224
rect 463016 389212 463022 389224
rect 474274 389212 474280 389224
rect 463016 389184 474280 389212
rect 463016 389172 463022 389184
rect 474274 389172 474280 389184
rect 474332 389172 474338 389224
rect 485038 389172 485044 389224
rect 485096 389212 485102 389224
rect 492582 389212 492588 389224
rect 485096 389184 492588 389212
rect 485096 389172 485102 389184
rect 492582 389172 492588 389184
rect 492640 389172 492646 389224
rect 492784 389212 492812 389320
rect 499546 389280 499574 389388
rect 502242 389280 502248 389292
rect 499546 389252 502248 389280
rect 502242 389240 502248 389252
rect 502300 389240 502306 389292
rect 514018 389240 514024 389292
rect 514076 389280 514082 389292
rect 520274 389280 520280 389292
rect 514076 389252 520280 389280
rect 514076 389240 514082 389252
rect 520274 389240 520280 389252
rect 520332 389240 520338 389292
rect 529934 389212 529940 389224
rect 492784 389184 529940 389212
rect 529934 389172 529940 389184
rect 529992 389172 529998 389224
rect 541618 389172 541624 389224
rect 541676 389212 541682 389224
rect 558270 389212 558276 389224
rect 541676 389184 558276 389212
rect 541676 389172 541682 389184
rect 558270 389172 558276 389184
rect 558328 389172 558334 389224
rect 122806 386600 132494 386628
rect 42702 386452 42708 386504
rect 42760 386492 42766 386504
rect 93854 386492 93860 386504
rect 42760 386464 93860 386492
rect 42760 386452 42766 386464
rect 93854 386452 93860 386464
rect 93912 386452 93918 386504
rect 97902 386452 97908 386504
rect 97960 386492 97966 386504
rect 122806 386492 122834 386600
rect 126882 386520 126888 386572
rect 126940 386560 126946 386572
rect 126940 386532 128492 386560
rect 126940 386520 126946 386532
rect 97960 386464 122834 386492
rect 97960 386452 97966 386464
rect 13538 386384 13544 386436
rect 13596 386424 13602 386436
rect 66254 386424 66260 386436
rect 13596 386396 66260 386424
rect 13596 386384 13602 386396
rect 66254 386384 66260 386396
rect 66312 386384 66318 386436
rect 70302 386384 70308 386436
rect 70360 386424 70366 386436
rect 121454 386424 121460 386436
rect 70360 386396 121460 386424
rect 70360 386384 70366 386396
rect 121454 386384 121460 386396
rect 121512 386384 121518 386436
rect 124858 386384 124864 386436
rect 124916 386424 124922 386436
rect 128262 386424 128268 386436
rect 124916 386396 128268 386424
rect 124916 386384 124922 386396
rect 128262 386384 128268 386396
rect 128320 386384 128326 386436
rect 128464 386424 128492 386532
rect 132466 386492 132494 386600
rect 182082 386520 182088 386572
rect 182140 386560 182146 386572
rect 233234 386560 233240 386572
rect 182140 386532 233240 386560
rect 182140 386520 182146 386532
rect 233234 386520 233240 386532
rect 233292 386520 233298 386572
rect 350442 386520 350448 386572
rect 350500 386560 350506 386572
rect 401594 386560 401600 386572
rect 350500 386532 401600 386560
rect 350500 386520 350506 386532
rect 401594 386520 401600 386532
rect 401652 386520 401658 386572
rect 462222 386520 462228 386572
rect 462280 386560 462286 386572
rect 513374 386560 513380 386572
rect 462280 386532 513380 386560
rect 462280 386520 462286 386532
rect 513374 386520 513380 386532
rect 513432 386520 513438 386572
rect 149054 386492 149060 386504
rect 132466 386464 149060 386492
rect 149054 386452 149060 386464
rect 149112 386452 149118 386504
rect 154482 386452 154488 386504
rect 154540 386492 154546 386504
rect 205634 386492 205640 386504
rect 154540 386464 205640 386492
rect 154540 386452 154546 386464
rect 205634 386452 205640 386464
rect 205692 386452 205698 386504
rect 238662 386452 238668 386504
rect 238720 386492 238726 386504
rect 289814 386492 289820 386504
rect 238720 386464 289820 386492
rect 238720 386452 238726 386464
rect 289814 386452 289820 386464
rect 289872 386452 289878 386504
rect 293862 386452 293868 386504
rect 293920 386492 293926 386504
rect 345014 386492 345020 386504
rect 293920 386464 345020 386492
rect 293920 386452 293926 386464
rect 345014 386452 345020 386464
rect 345072 386452 345078 386504
rect 378042 386452 378048 386504
rect 378100 386492 378106 386504
rect 429286 386492 429292 386504
rect 378100 386464 429292 386492
rect 378100 386452 378106 386464
rect 429286 386452 429292 386464
rect 429344 386452 429350 386504
rect 434622 386452 434628 386504
rect 434680 386492 434686 386504
rect 485774 386492 485780 386504
rect 434680 386464 485780 386492
rect 434680 386452 434686 386464
rect 485774 386452 485780 386464
rect 485832 386452 485838 386504
rect 518802 386452 518808 386504
rect 518860 386492 518866 386504
rect 569954 386492 569960 386504
rect 518860 386464 569960 386492
rect 518860 386452 518866 386464
rect 569954 386452 569960 386464
rect 570012 386452 570018 386504
rect 178034 386424 178040 386436
rect 128464 386396 178040 386424
rect 178034 386384 178040 386396
rect 178092 386384 178098 386436
rect 209682 386384 209688 386436
rect 209740 386424 209746 386436
rect 262214 386424 262220 386436
rect 209740 386396 262220 386424
rect 209740 386384 209746 386396
rect 262214 386384 262220 386396
rect 262272 386384 262278 386436
rect 266262 386384 266268 386436
rect 266320 386424 266326 386436
rect 317414 386424 317420 386436
rect 266320 386396 317420 386424
rect 266320 386384 266326 386396
rect 317414 386384 317420 386396
rect 317472 386384 317478 386436
rect 322842 386384 322848 386436
rect 322900 386424 322906 386436
rect 373994 386424 374000 386436
rect 322900 386396 374000 386424
rect 322900 386384 322906 386396
rect 373994 386384 374000 386396
rect 374052 386384 374058 386436
rect 405642 386384 405648 386436
rect 405700 386424 405706 386436
rect 458174 386424 458180 386436
rect 405700 386396 458180 386424
rect 405700 386384 405706 386396
rect 458174 386384 458180 386396
rect 458232 386384 458238 386436
rect 489822 386384 489828 386436
rect 489880 386424 489886 386436
rect 542354 386424 542360 386436
rect 489880 386396 542360 386424
rect 489880 386384 489886 386396
rect 542354 386384 542360 386396
rect 542412 386384 542418 386436
rect 544378 386384 544384 386436
rect 544436 386424 544442 386436
rect 548334 386424 548340 386436
rect 544436 386396 548340 386424
rect 544436 386384 544442 386396
rect 548334 386384 548340 386396
rect 548392 386384 548398 386436
rect 120258 386248 120264 386300
rect 120316 386288 120322 386300
rect 122098 386288 122104 386300
rect 120316 386260 122104 386288
rect 120316 386248 120322 386260
rect 122098 386248 122104 386260
rect 122156 386248 122162 386300
rect 204070 385024 204076 385076
rect 204128 385064 204134 385076
rect 212442 385064 212448 385076
rect 204128 385036 212448 385064
rect 204128 385024 204134 385036
rect 212442 385024 212448 385036
rect 212500 385024 212506 385076
rect 204254 384956 204260 385008
rect 204312 384996 204318 385008
rect 204990 384996 204996 385008
rect 204312 384968 204996 384996
rect 204312 384956 204318 384968
rect 204990 384956 204996 384968
rect 205048 384956 205054 385008
rect 568114 378156 568120 378208
rect 568172 378196 568178 378208
rect 580166 378196 580172 378208
rect 568172 378168 580172 378196
rect 568172 378156 568178 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 15194 365644 15200 365696
rect 15252 365684 15258 365696
rect 35894 365684 35900 365696
rect 15252 365656 35900 365684
rect 15252 365644 15258 365656
rect 35894 365644 35900 365656
rect 35952 365644 35958 365696
rect 36078 365644 36084 365696
rect 36136 365684 36142 365696
rect 63586 365684 63592 365696
rect 36136 365656 63592 365684
rect 36136 365644 36142 365656
rect 63586 365644 63592 365656
rect 63644 365644 63650 365696
rect 64046 365644 64052 365696
rect 64104 365684 64110 365696
rect 91922 365684 91928 365696
rect 64104 365656 91928 365684
rect 64104 365644 64110 365656
rect 91922 365644 91928 365656
rect 91980 365644 91986 365696
rect 92106 365644 92112 365696
rect 92164 365684 92170 365696
rect 119614 365684 119620 365696
rect 92164 365656 119620 365684
rect 92164 365644 92170 365656
rect 119614 365644 119620 365656
rect 119672 365644 119678 365696
rect 122098 365644 122104 365696
rect 122156 365684 122162 365696
rect 147950 365684 147956 365696
rect 122156 365656 147956 365684
rect 122156 365644 122162 365656
rect 147950 365644 147956 365656
rect 148008 365644 148014 365696
rect 148042 365644 148048 365696
rect 148100 365684 148106 365696
rect 175918 365684 175924 365696
rect 148100 365656 175924 365684
rect 148100 365644 148106 365656
rect 175918 365644 175924 365656
rect 175976 365644 175982 365696
rect 176102 365644 176108 365696
rect 176160 365684 176166 365696
rect 203610 365684 203616 365696
rect 176160 365656 203616 365684
rect 176160 365644 176166 365656
rect 203610 365644 203616 365656
rect 203668 365644 203674 365696
rect 204990 365644 204996 365696
rect 205048 365684 205054 365696
rect 231946 365684 231952 365696
rect 205048 365656 231952 365684
rect 205048 365644 205054 365656
rect 231946 365644 231952 365656
rect 232004 365644 232010 365696
rect 232038 365644 232044 365696
rect 232096 365684 232102 365696
rect 259914 365684 259920 365696
rect 232096 365656 259920 365684
rect 232096 365644 232102 365656
rect 259914 365644 259920 365656
rect 259972 365644 259978 365696
rect 260098 365644 260104 365696
rect 260156 365684 260162 365696
rect 287606 365684 287612 365696
rect 260156 365656 287612 365684
rect 260156 365644 260162 365656
rect 287606 365644 287612 365656
rect 287664 365644 287670 365696
rect 288066 365644 288072 365696
rect 288124 365684 288130 365696
rect 315942 365684 315948 365696
rect 288124 365656 315948 365684
rect 288124 365644 288130 365656
rect 315942 365644 315948 365656
rect 316000 365644 316006 365696
rect 316678 365644 316684 365696
rect 316736 365684 316742 365696
rect 343910 365684 343916 365696
rect 316736 365656 343916 365684
rect 316736 365644 316742 365656
rect 343910 365644 343916 365656
rect 343968 365644 343974 365696
rect 344094 365644 344100 365696
rect 344152 365684 344158 365696
rect 371602 365684 371608 365696
rect 344152 365656 371608 365684
rect 344152 365644 344158 365656
rect 371602 365644 371608 365656
rect 371660 365644 371666 365696
rect 372062 365644 372068 365696
rect 372120 365684 372126 365696
rect 399938 365684 399944 365696
rect 372120 365656 399944 365684
rect 372120 365644 372126 365656
rect 399938 365644 399944 365656
rect 399996 365644 400002 365696
rect 400858 365644 400864 365696
rect 400916 365684 400922 365696
rect 427906 365684 427912 365696
rect 400916 365656 427912 365684
rect 400916 365644 400922 365656
rect 427906 365644 427912 365656
rect 427964 365644 427970 365696
rect 428090 365644 428096 365696
rect 428148 365684 428154 365696
rect 455598 365684 455604 365696
rect 428148 365656 455604 365684
rect 428148 365644 428154 365656
rect 455598 365644 455604 365656
rect 455656 365644 455662 365696
rect 456058 365644 456064 365696
rect 456116 365684 456122 365696
rect 483934 365684 483940 365696
rect 456116 365656 483940 365684
rect 456116 365644 456122 365656
rect 483934 365644 483940 365656
rect 483992 365644 483998 365696
rect 484026 365644 484032 365696
rect 484084 365684 484090 365696
rect 511902 365684 511908 365696
rect 484084 365656 511908 365684
rect 484084 365644 484090 365656
rect 511902 365644 511908 365656
rect 511960 365644 511966 365696
rect 512086 365644 512092 365696
rect 512144 365684 512150 365696
rect 539594 365684 539600 365696
rect 512144 365656 539600 365684
rect 512144 365644 512150 365656
rect 539594 365644 539600 365656
rect 539652 365644 539658 365696
rect 540054 365644 540060 365696
rect 540112 365684 540118 365696
rect 567930 365684 567936 365696
rect 540112 365656 567936 365684
rect 540112 365644 540118 365656
rect 567930 365644 567936 365656
rect 567988 365644 567994 365696
rect 16574 365576 16580 365628
rect 16632 365616 16638 365628
rect 36630 365616 36636 365628
rect 16632 365588 36636 365616
rect 16632 365576 16638 365588
rect 36630 365576 36636 365588
rect 36688 365576 36694 365628
rect 44910 365576 44916 365628
rect 44968 365616 44974 365628
rect 71130 365616 71136 365628
rect 44968 365588 71136 365616
rect 44968 365576 44974 365588
rect 71130 365576 71136 365588
rect 71188 365576 71194 365628
rect 82262 365576 82268 365628
rect 82320 365616 82326 365628
rect 93118 365616 93124 365628
rect 82320 365588 93124 365616
rect 82320 365576 82326 365588
rect 93118 365576 93124 365588
rect 93176 365576 93182 365628
rect 110230 365576 110236 365628
rect 110288 365616 110294 365628
rect 124858 365616 124864 365628
rect 110288 365588 124864 365616
rect 110288 365576 110294 365588
rect 124858 365576 124864 365588
rect 124916 365576 124922 365628
rect 128630 365576 128636 365628
rect 128688 365616 128694 365628
rect 149698 365616 149704 365628
rect 128688 365588 149704 365616
rect 128688 365576 128694 365588
rect 149698 365576 149704 365588
rect 149756 365576 149762 365628
rect 156598 365576 156604 365628
rect 156656 365616 156662 365628
rect 182818 365616 182824 365628
rect 156656 365588 182824 365616
rect 156656 365576 156662 365588
rect 182818 365576 182824 365588
rect 182876 365576 182882 365628
rect 194502 365576 194508 365628
rect 194560 365616 194566 365628
rect 204070 365616 204076 365628
rect 194560 365588 204076 365616
rect 194560 365576 194566 365588
rect 204070 365576 204076 365588
rect 204128 365576 204134 365628
rect 212626 365576 212632 365628
rect 212684 365616 212690 365628
rect 232498 365616 232504 365628
rect 212684 365588 232504 365616
rect 212684 365576 212690 365588
rect 232498 365576 232504 365588
rect 232556 365576 232562 365628
rect 240594 365576 240600 365628
rect 240652 365616 240658 365628
rect 266998 365616 267004 365628
rect 240652 365588 267004 365616
rect 240652 365576 240658 365588
rect 266998 365576 267004 365588
rect 267056 365576 267062 365628
rect 278590 365576 278596 365628
rect 278648 365616 278654 365628
rect 289078 365616 289084 365628
rect 278648 365588 289084 365616
rect 278648 365576 278654 365588
rect 289078 365576 289084 365588
rect 289136 365576 289142 365628
rect 306282 365576 306288 365628
rect 306340 365616 306346 365628
rect 318058 365616 318064 365628
rect 306340 365588 318064 365616
rect 306340 365576 306346 365588
rect 318058 365576 318064 365588
rect 318116 365576 318122 365628
rect 324590 365576 324596 365628
rect 324648 365616 324654 365628
rect 345658 365616 345664 365628
rect 324648 365588 345664 365616
rect 324648 365576 324654 365588
rect 345658 365576 345664 365588
rect 345716 365576 345722 365628
rect 362586 365576 362592 365628
rect 362644 365616 362650 365628
rect 373258 365616 373264 365628
rect 362644 365588 373264 365616
rect 362644 365576 362650 365588
rect 373258 365576 373264 365588
rect 373316 365576 373322 365628
rect 390278 365576 390284 365628
rect 390336 365616 390342 365628
rect 400950 365616 400956 365628
rect 390336 365588 400956 365616
rect 390336 365576 390342 365588
rect 400950 365576 400956 365588
rect 401008 365576 401014 365628
rect 408586 365576 408592 365628
rect 408644 365616 408650 365628
rect 428458 365616 428464 365628
rect 408644 365588 428464 365616
rect 408644 365576 408650 365588
rect 428458 365576 428464 365588
rect 428516 365576 428522 365628
rect 436922 365576 436928 365628
rect 436980 365616 436986 365628
rect 462958 365616 462964 365628
rect 436980 365588 462964 365616
rect 436980 365576 436986 365588
rect 462958 365576 462964 365588
rect 463016 365576 463022 365628
rect 474274 365576 474280 365628
rect 474332 365616 474338 365628
rect 485038 365616 485044 365628
rect 474332 365588 485044 365616
rect 474332 365576 474338 365588
rect 485038 365576 485044 365588
rect 485096 365576 485102 365628
rect 502242 365576 502248 365628
rect 502300 365616 502306 365628
rect 514018 365616 514024 365628
rect 502300 365588 514024 365616
rect 502300 365576 502306 365588
rect 514018 365576 514024 365588
rect 514076 365576 514082 365628
rect 520918 365576 520924 365628
rect 520976 365616 520982 365628
rect 541618 365616 541624 365628
rect 520976 365588 541624 365616
rect 520976 365576 520982 365588
rect 541618 365576 541624 365588
rect 541676 365576 541682 365628
rect 26234 365508 26240 365560
rect 26292 365548 26298 365560
rect 43530 365548 43536 365560
rect 26292 365520 43536 365548
rect 26292 365508 26298 365520
rect 43530 365508 43536 365520
rect 43588 365508 43594 365560
rect 54570 365508 54576 365560
rect 54628 365548 54634 365560
rect 66898 365548 66904 365560
rect 54628 365520 66904 365548
rect 54628 365508 54634 365520
rect 66898 365508 66904 365520
rect 66956 365508 66962 365560
rect 138290 365508 138296 365560
rect 138348 365548 138354 365560
rect 151078 365548 151084 365560
rect 138348 365520 151084 365548
rect 138348 365508 138354 365520
rect 151078 365508 151084 365520
rect 151136 365508 151142 365560
rect 166258 365508 166264 365560
rect 166316 365548 166322 365560
rect 177298 365548 177304 365560
rect 166316 365520 177304 365548
rect 166316 365508 166322 365520
rect 177298 365508 177304 365520
rect 177356 365508 177362 365560
rect 222286 365508 222292 365560
rect 222344 365548 222350 365560
rect 233970 365548 233976 365560
rect 222344 365520 233976 365548
rect 222344 365508 222350 365520
rect 233970 365508 233976 365520
rect 234028 365508 234034 365560
rect 250254 365508 250260 365560
rect 250312 365548 250318 365560
rect 261478 365548 261484 365560
rect 250312 365520 261484 365548
rect 250312 365508 250318 365520
rect 261478 365508 261484 365520
rect 261536 365508 261542 365560
rect 334250 365508 334256 365560
rect 334308 365548 334314 365560
rect 347038 365548 347044 365560
rect 334308 365520 347044 365548
rect 334308 365508 334314 365520
rect 347038 365508 347044 365520
rect 347096 365508 347102 365560
rect 418246 365508 418252 365560
rect 418304 365548 418310 365560
rect 429838 365548 429844 365560
rect 418304 365520 429844 365548
rect 418304 365508 418310 365520
rect 429838 365508 429844 365520
rect 429896 365508 429902 365560
rect 446582 365508 446588 365560
rect 446640 365548 446646 365560
rect 457438 365548 457444 365560
rect 446640 365520 457444 365548
rect 446640 365508 446646 365520
rect 457438 365508 457444 365520
rect 457496 365508 457502 365560
rect 530578 365508 530584 365560
rect 530636 365548 530642 365560
rect 544378 365548 544384 365560
rect 530636 365520 544384 365548
rect 530636 365508 530642 365520
rect 544378 365508 544384 365520
rect 544436 365508 544442 365560
rect 558270 364964 558276 365016
rect 558328 365004 558334 365016
rect 567470 365004 567476 365016
rect 558328 364976 567476 365004
rect 558328 364964 558334 364976
rect 567470 364964 567476 364976
rect 567528 364964 567534 365016
rect 548334 362176 548340 362228
rect 548392 362216 548398 362228
rect 568114 362216 568120 362228
rect 548392 362188 568120 362216
rect 548392 362176 548398 362188
rect 568114 362176 568120 362188
rect 568172 362176 568178 362228
rect 148410 361700 148416 361752
rect 148468 361740 148474 361752
rect 165706 361740 165712 361752
rect 148468 361712 165712 361740
rect 148468 361700 148474 361712
rect 165706 361700 165712 361712
rect 165764 361700 165770 361752
rect 175458 361700 175464 361752
rect 175516 361740 175522 361752
rect 193674 361740 193680 361752
rect 175516 361712 193680 361740
rect 175516 361700 175522 361712
rect 193674 361700 193680 361712
rect 193732 361700 193738 361752
rect 203518 361700 203524 361752
rect 203576 361740 203582 361752
rect 221366 361740 221372 361752
rect 203576 361712 221372 361740
rect 203576 361700 203582 361712
rect 221366 361700 221372 361712
rect 221424 361700 221430 361752
rect 232590 361700 232596 361752
rect 232648 361740 232654 361752
rect 249702 361740 249708 361752
rect 232648 361712 249708 361740
rect 232648 361700 232654 361712
rect 249702 361700 249708 361712
rect 249760 361700 249766 361752
rect 260098 361700 260104 361752
rect 260156 361740 260162 361752
rect 277670 361740 277676 361752
rect 260156 361712 277676 361740
rect 260156 361700 260162 361712
rect 277670 361700 277676 361712
rect 277728 361700 277734 361752
rect 296346 361700 296352 361752
rect 296404 361740 296410 361752
rect 316770 361740 316776 361752
rect 296404 361712 316776 361740
rect 296404 361700 296410 361712
rect 316770 361700 316776 361712
rect 316828 361700 316834 361752
rect 345658 361700 345664 361752
rect 345716 361740 345722 361752
rect 361666 361740 361672 361752
rect 345716 361712 361672 361740
rect 345716 361700 345722 361712
rect 361666 361700 361672 361712
rect 361724 361700 361730 361752
rect 371510 361700 371516 361752
rect 371568 361740 371574 361752
rect 389358 361740 389364 361752
rect 371568 361712 389364 361740
rect 371568 361700 371574 361712
rect 389358 361700 389364 361712
rect 389416 361700 389422 361752
rect 399478 361700 399484 361752
rect 399536 361740 399542 361752
rect 417694 361740 417700 361752
rect 399536 361712 417700 361740
rect 399536 361700 399542 361712
rect 417694 361700 417700 361712
rect 417752 361700 417758 361752
rect 428458 361700 428464 361752
rect 428516 361740 428522 361752
rect 445662 361740 445668 361752
rect 428516 361712 445668 361740
rect 428516 361700 428522 361712
rect 445662 361700 445668 361712
rect 445720 361700 445726 361752
rect 456058 361700 456064 361752
rect 456116 361740 456122 361752
rect 473354 361740 473360 361752
rect 456116 361712 473360 361740
rect 456116 361700 456122 361712
rect 473354 361700 473360 361712
rect 473412 361700 473418 361752
rect 483474 361700 483480 361752
rect 483532 361740 483538 361752
rect 501690 361740 501696 361752
rect 483532 361712 501696 361740
rect 483532 361700 483538 361712
rect 501690 361700 501696 361712
rect 501748 361700 501754 361752
rect 511442 361700 511448 361752
rect 511500 361740 511506 361752
rect 529658 361740 529664 361752
rect 511500 361712 529664 361740
rect 511500 361700 511506 361712
rect 529658 361700 529664 361712
rect 529716 361700 529722 361752
rect 36630 361632 36636 361684
rect 36688 361672 36694 361684
rect 53650 361672 53656 361684
rect 36688 361644 53656 361672
rect 36688 361632 36694 361644
rect 53650 361632 53656 361644
rect 53708 361632 53714 361684
rect 64414 361632 64420 361684
rect 64472 361672 64478 361684
rect 81434 361672 81440 361684
rect 64472 361644 81440 361672
rect 64472 361632 64478 361644
rect 81434 361632 81440 361644
rect 81492 361632 81498 361684
rect 119430 361632 119436 361684
rect 119488 361672 119494 361684
rect 137646 361672 137652 361684
rect 119488 361644 137652 361672
rect 119488 361632 119494 361644
rect 137646 361632 137652 361644
rect 137704 361632 137710 361684
rect 156322 361632 156328 361684
rect 156380 361672 156386 361684
rect 178678 361672 178684 361684
rect 156380 361644 178684 361672
rect 156380 361632 156386 361644
rect 178678 361632 178684 361644
rect 178736 361632 178742 361684
rect 212350 361632 212356 361684
rect 212408 361672 212414 361684
rect 232682 361672 232688 361684
rect 212408 361644 232688 361672
rect 212408 361632 212414 361644
rect 232682 361632 232688 361644
rect 232740 361632 232746 361684
rect 268010 361632 268016 361684
rect 268068 361672 268074 361684
rect 287698 361672 287704 361684
rect 268068 361644 287704 361672
rect 268068 361632 268074 361644
rect 287698 361632 287704 361644
rect 287756 361632 287762 361684
rect 315482 361632 315488 361684
rect 315540 361672 315546 361684
rect 333698 361672 333704 361684
rect 315540 361644 333704 361672
rect 315540 361632 315546 361644
rect 333698 361632 333704 361644
rect 333756 361632 333762 361684
rect 352006 361632 352012 361684
rect 352064 361672 352070 361684
rect 374638 361672 374644 361684
rect 352064 361644 374644 361672
rect 352064 361632 352070 361644
rect 374638 361632 374644 361644
rect 374696 361632 374702 361684
rect 408034 361632 408040 361684
rect 408092 361672 408098 361684
rect 428642 361672 428648 361684
rect 408092 361644 428648 361672
rect 408092 361632 408098 361644
rect 428642 361632 428648 361644
rect 428700 361632 428706 361684
rect 464338 361632 464344 361684
rect 464396 361672 464402 361684
rect 483658 361672 483664 361684
rect 464396 361644 483664 361672
rect 464396 361632 464402 361644
rect 483658 361632 483664 361644
rect 483716 361632 483722 361684
rect 492030 361632 492036 361684
rect 492088 361672 492094 361684
rect 512730 361672 512736 361684
rect 492088 361644 512736 361672
rect 492088 361632 492094 361644
rect 512730 361632 512736 361644
rect 512788 361632 512794 361684
rect 541618 361632 541624 361684
rect 541676 361672 541682 361684
rect 557534 361672 557540 361684
rect 541676 361644 557540 361672
rect 541676 361632 541682 361644
rect 557534 361632 557540 361644
rect 557592 361632 557598 361684
rect 15102 361564 15108 361616
rect 15160 361604 15166 361616
rect 25682 361604 25688 361616
rect 15160 361576 25688 361604
rect 15160 361564 15166 361576
rect 25682 361564 25688 361576
rect 25740 361564 25746 361616
rect 36722 361564 36728 361616
rect 36780 361604 36786 361616
rect 63310 361604 63316 361616
rect 36780 361576 63316 361604
rect 36780 361564 36786 361576
rect 63310 361564 63316 361576
rect 63368 361564 63374 361616
rect 66898 361564 66904 361616
rect 66956 361604 66962 361616
rect 91094 361604 91100 361616
rect 66956 361576 91100 361604
rect 66956 361564 66962 361576
rect 91094 361564 91100 361576
rect 91152 361564 91158 361616
rect 93118 361564 93124 361616
rect 93176 361604 93182 361616
rect 119338 361604 119344 361616
rect 93176 361576 119344 361604
rect 93176 361564 93182 361576
rect 119338 361564 119344 361576
rect 119396 361564 119402 361616
rect 122098 361564 122104 361616
rect 122156 361604 122162 361616
rect 147306 361604 147312 361616
rect 122156 361576 147312 361604
rect 122156 361564 122162 361576
rect 147306 361564 147312 361576
rect 147364 361564 147370 361616
rect 148318 361564 148324 361616
rect 148376 361604 148382 361616
rect 175366 361604 175372 361616
rect 148376 361576 175372 361604
rect 148376 361564 148382 361576
rect 175366 361564 175372 361576
rect 175424 361564 175430 361616
rect 177298 361564 177304 361616
rect 177356 361604 177362 361616
rect 203334 361604 203340 361616
rect 177356 361576 203340 361604
rect 177356 361564 177362 361576
rect 203334 361564 203340 361576
rect 203392 361564 203398 361616
rect 204990 361564 204996 361616
rect 205048 361604 205054 361616
rect 231026 361604 231032 361616
rect 205048 361576 231032 361604
rect 205048 361564 205054 361576
rect 231026 361564 231032 361576
rect 231084 361564 231090 361616
rect 232498 361564 232504 361616
rect 232556 361604 232562 361616
rect 259362 361604 259368 361616
rect 232556 361576 259368 361604
rect 232556 361564 232562 361576
rect 259362 361564 259368 361576
rect 259420 361564 259426 361616
rect 260190 361564 260196 361616
rect 260248 361604 260254 361616
rect 287330 361604 287336 361616
rect 260248 361576 287336 361604
rect 260248 361564 260254 361576
rect 287330 361564 287336 361576
rect 287388 361564 287394 361616
rect 289078 361564 289084 361616
rect 289136 361604 289142 361616
rect 315022 361604 315028 361616
rect 289136 361576 315028 361604
rect 289136 361564 289142 361576
rect 315022 361564 315028 361576
rect 315080 361564 315086 361616
rect 316678 361564 316684 361616
rect 316736 361604 316742 361616
rect 343358 361604 343364 361616
rect 316736 361576 343364 361604
rect 316736 361564 316742 361576
rect 343358 361564 343364 361576
rect 343416 361564 343422 361616
rect 344278 361564 344284 361616
rect 344336 361604 344342 361616
rect 371326 361604 371332 361616
rect 344336 361576 371332 361604
rect 344336 361564 344342 361576
rect 371326 361564 371332 361576
rect 371384 361564 371390 361616
rect 373258 361564 373264 361616
rect 373316 361604 373322 361616
rect 399018 361604 399024 361616
rect 373316 361576 399024 361604
rect 373316 361564 373322 361576
rect 399018 361564 399024 361576
rect 399076 361564 399082 361616
rect 400858 361564 400864 361616
rect 400916 361604 400922 361616
rect 427354 361604 427360 361616
rect 400916 361576 427360 361604
rect 400916 361564 400922 361576
rect 427354 361564 427360 361576
rect 427412 361564 427418 361616
rect 428550 361564 428556 361616
rect 428608 361604 428614 361616
rect 455322 361604 455328 361616
rect 428608 361576 455328 361604
rect 428608 361564 428614 361576
rect 455322 361564 455328 361576
rect 455380 361564 455386 361616
rect 456150 361564 456156 361616
rect 456208 361604 456214 361616
rect 483014 361604 483020 361616
rect 456208 361576 483020 361604
rect 456208 361564 456214 361576
rect 483014 361564 483020 361576
rect 483072 361564 483078 361616
rect 485038 361564 485044 361616
rect 485096 361604 485102 361616
rect 511350 361604 511356 361616
rect 485096 361576 511356 361604
rect 485096 361564 485102 361576
rect 511350 361564 511356 361576
rect 511408 361564 511414 361616
rect 512638 361564 512644 361616
rect 512696 361604 512702 361616
rect 539318 361604 539324 361616
rect 512696 361576 539324 361604
rect 512696 361564 512702 361576
rect 539318 361564 539324 361576
rect 539376 361564 539382 361616
rect 540238 361564 540244 361616
rect 540296 361604 540302 361616
rect 567194 361604 567200 361616
rect 540296 361576 567200 361604
rect 540296 361564 540302 361576
rect 567194 361564 567200 361576
rect 567252 361564 567258 361616
rect 109310 359252 109316 359304
rect 109368 359252 109374 359304
rect 305362 359292 305368 359304
rect 296686 359264 305368 359292
rect 91462 358776 91468 358828
rect 91520 358816 91526 358828
rect 109328 358816 109356 359252
rect 91520 358788 109356 358816
rect 91520 358776 91526 358788
rect 287514 358776 287520 358828
rect 287572 358816 287578 358828
rect 296686 358816 296714 359264
rect 305362 359252 305368 359264
rect 305420 359252 305426 359304
rect 287572 358788 296714 358816
rect 287572 358776 287578 358788
rect 42886 356940 42892 356992
rect 42944 356980 42950 356992
rect 43622 356980 43628 356992
rect 42944 356952 43628 356980
rect 42944 356940 42950 356952
rect 43622 356940 43628 356952
rect 43680 356940 43686 356992
rect 2774 345176 2780 345228
rect 2832 345216 2838 345228
rect 4982 345216 4988 345228
rect 2832 345188 4988 345216
rect 2832 345176 2838 345188
rect 4982 345176 4988 345188
rect 5040 345176 5046 345228
rect 63586 342524 63592 342576
rect 63644 342564 63650 342576
rect 64414 342564 64420 342576
rect 63644 342536 64420 342564
rect 63644 342524 63650 342536
rect 64414 342524 64420 342536
rect 64472 342524 64478 342576
rect 147674 342524 147680 342576
rect 147732 342564 147738 342576
rect 148410 342564 148416 342576
rect 147732 342536 148416 342564
rect 147732 342524 147738 342536
rect 148410 342524 148416 342536
rect 148468 342524 148474 342576
rect 512730 341912 512736 341964
rect 512788 341952 512794 341964
rect 519630 341952 519636 341964
rect 512788 341924 519636 341952
rect 512788 341912 512794 341924
rect 519630 341912 519636 341924
rect 519688 341912 519694 341964
rect 287698 341504 287704 341556
rect 287756 341544 287762 341556
rect 295702 341544 295708 341556
rect 287756 341516 295708 341544
rect 287756 341504 287762 341516
rect 295702 341504 295708 341516
rect 295760 341504 295766 341556
rect 428642 341504 428648 341556
rect 428700 341544 428706 341556
rect 435726 341544 435732 341556
rect 428700 341516 435732 341544
rect 428700 341504 428706 341516
rect 435726 341504 435732 341516
rect 435784 341504 435790 341556
rect 232682 341368 232688 341420
rect 232740 341408 232746 341420
rect 239766 341408 239772 341420
rect 232740 341380 239772 341408
rect 232740 341368 232746 341380
rect 239766 341368 239772 341380
rect 239824 341368 239830 341420
rect 483658 341368 483664 341420
rect 483716 341408 483722 341420
rect 491662 341408 491668 341420
rect 483716 341380 491668 341408
rect 483716 341368 483722 341380
rect 491662 341368 491668 341380
rect 491720 341368 491726 341420
rect 316770 341232 316776 341284
rect 316828 341272 316834 341284
rect 323670 341272 323676 341284
rect 316828 341244 323676 341272
rect 316828 341232 316834 341244
rect 323670 341232 323676 341244
rect 323728 341232 323734 341284
rect 13538 340824 13544 340876
rect 13596 340864 13602 340876
rect 66254 340864 66260 340876
rect 13596 340836 66260 340864
rect 13596 340824 13602 340836
rect 66254 340824 66260 340836
rect 66312 340824 66318 340876
rect 70302 340824 70308 340876
rect 70360 340864 70366 340876
rect 121454 340864 121460 340876
rect 70360 340836 121460 340864
rect 70360 340824 70366 340836
rect 121454 340824 121460 340836
rect 121512 340824 121518 340876
rect 126882 340824 126888 340876
rect 126940 340864 126946 340876
rect 178034 340864 178040 340876
rect 126940 340836 178040 340864
rect 126940 340824 126946 340836
rect 178034 340824 178040 340836
rect 178092 340824 178098 340876
rect 209682 340824 209688 340876
rect 209740 340864 209746 340876
rect 262214 340864 262220 340876
rect 209740 340836 262220 340864
rect 209740 340824 209746 340836
rect 262214 340824 262220 340836
rect 262272 340824 262278 340876
rect 266262 340824 266268 340876
rect 266320 340864 266326 340876
rect 317414 340864 317420 340876
rect 266320 340836 317420 340864
rect 266320 340824 266326 340836
rect 317414 340824 317420 340836
rect 317472 340824 317478 340876
rect 322842 340824 322848 340876
rect 322900 340864 322906 340876
rect 373994 340864 374000 340876
rect 322900 340836 374000 340864
rect 322900 340824 322906 340836
rect 373994 340824 374000 340836
rect 374052 340824 374058 340876
rect 405642 340824 405648 340876
rect 405700 340864 405706 340876
rect 458174 340864 458180 340876
rect 405700 340836 458180 340864
rect 405700 340824 405706 340836
rect 458174 340824 458180 340836
rect 458232 340824 458238 340876
rect 489822 340824 489828 340876
rect 489880 340864 489886 340876
rect 489880 340836 539364 340864
rect 489880 340824 489886 340836
rect 42702 340756 42708 340808
rect 42760 340796 42766 340808
rect 93854 340796 93860 340808
rect 42760 340768 93860 340796
rect 42760 340756 42766 340768
rect 93854 340756 93860 340768
rect 93912 340756 93918 340808
rect 97902 340756 97908 340808
rect 97960 340796 97966 340808
rect 149054 340796 149060 340808
rect 97960 340768 149060 340796
rect 97960 340756 97966 340768
rect 149054 340756 149060 340768
rect 149112 340756 149118 340808
rect 154482 340756 154488 340808
rect 154540 340796 154546 340808
rect 205634 340796 205640 340808
rect 154540 340768 205640 340796
rect 154540 340756 154546 340768
rect 205634 340756 205640 340768
rect 205692 340756 205698 340808
rect 231670 340756 231676 340808
rect 231728 340796 231734 340808
rect 232590 340796 232596 340808
rect 231728 340768 232596 340796
rect 231728 340756 231734 340768
rect 232590 340756 232596 340768
rect 232648 340756 232654 340808
rect 238662 340756 238668 340808
rect 238720 340796 238726 340808
rect 289814 340796 289820 340808
rect 238720 340768 289820 340796
rect 238720 340756 238726 340768
rect 289814 340756 289820 340768
rect 289872 340756 289878 340808
rect 293862 340756 293868 340808
rect 293920 340796 293926 340808
rect 345014 340796 345020 340808
rect 293920 340768 345020 340796
rect 293920 340756 293926 340768
rect 345014 340756 345020 340768
rect 345072 340756 345078 340808
rect 378042 340756 378048 340808
rect 378100 340796 378106 340808
rect 429286 340796 429292 340808
rect 378100 340768 429292 340796
rect 378100 340756 378106 340768
rect 429286 340756 429292 340768
rect 429344 340756 429350 340808
rect 434622 340756 434628 340808
rect 434680 340796 434686 340808
rect 485774 340796 485780 340808
rect 434680 340768 485780 340796
rect 434680 340756 434686 340768
rect 485774 340756 485780 340768
rect 485832 340756 485838 340808
rect 518802 340756 518808 340808
rect 518860 340796 518866 340808
rect 518860 340768 528554 340796
rect 518860 340756 518866 340768
rect 35250 340688 35256 340740
rect 35308 340728 35314 340740
rect 36630 340728 36636 340740
rect 35308 340700 36636 340728
rect 35308 340688 35314 340700
rect 36630 340688 36636 340700
rect 36688 340688 36694 340740
rect 182082 340688 182088 340740
rect 182140 340728 182146 340740
rect 233234 340728 233240 340740
rect 182140 340700 233240 340728
rect 182140 340688 182146 340700
rect 233234 340688 233240 340700
rect 233292 340688 233298 340740
rect 343634 340688 343640 340740
rect 343692 340728 343698 340740
rect 345658 340728 345664 340740
rect 343692 340700 345664 340728
rect 343692 340688 343698 340700
rect 345658 340688 345664 340700
rect 345716 340688 345722 340740
rect 350442 340688 350448 340740
rect 350500 340728 350506 340740
rect 401594 340728 401600 340740
rect 350500 340700 401600 340728
rect 350500 340688 350506 340700
rect 401594 340688 401600 340700
rect 401652 340688 401658 340740
rect 462222 340688 462228 340740
rect 462280 340728 462286 340740
rect 513374 340728 513380 340740
rect 462280 340700 513380 340728
rect 462280 340688 462286 340700
rect 513374 340688 513380 340700
rect 513432 340688 513438 340740
rect 528526 340660 528554 340768
rect 539336 340728 539364 340836
rect 539502 340824 539508 340876
rect 539560 340864 539566 340876
rect 541618 340864 541624 340876
rect 539560 340836 541624 340864
rect 539560 340824 539566 340836
rect 541618 340824 541624 340836
rect 541676 340824 541682 340876
rect 569954 340796 569960 340808
rect 547846 340768 569960 340796
rect 542354 340728 542360 340740
rect 539336 340700 542360 340728
rect 542354 340688 542360 340700
rect 542412 340688 542418 340740
rect 547846 340660 547874 340768
rect 569954 340756 569960 340768
rect 570012 340756 570018 340808
rect 528526 340632 547874 340660
rect 547874 340552 547880 340604
rect 547932 340592 547938 340604
rect 548150 340592 548156 340604
rect 547932 340564 548156 340592
rect 547932 340552 547938 340564
rect 548150 340552 548156 340564
rect 548208 340552 548214 340604
rect 71866 338036 71872 338088
rect 71924 338076 71930 338088
rect 100018 338076 100024 338088
rect 71924 338048 100024 338076
rect 71924 338036 71930 338048
rect 100018 338036 100024 338048
rect 100076 338036 100082 338088
rect 127986 338076 127992 338088
rect 103486 338048 127992 338076
rect 25682 337968 25688 338020
rect 25740 338008 25746 338020
rect 36722 338008 36728 338020
rect 25740 337980 36728 338008
rect 25740 337968 25746 337980
rect 36722 337968 36728 337980
rect 36780 337968 36786 338020
rect 42886 337968 42892 338020
rect 42944 338008 42950 338020
rect 42944 337980 45554 338008
rect 42944 337968 42950 337980
rect 15286 337900 15292 337952
rect 15344 337940 15350 337952
rect 43990 337940 43996 337952
rect 15344 337912 43996 337940
rect 15344 337900 15350 337912
rect 43990 337900 43996 337912
rect 44048 337900 44054 337952
rect 45526 337940 45554 337980
rect 53650 337968 53656 338020
rect 53708 338008 53714 338020
rect 66898 338008 66904 338020
rect 53708 337980 66904 338008
rect 53708 337968 53714 337980
rect 66898 337968 66904 337980
rect 66956 337968 66962 338020
rect 81986 337968 81992 338020
rect 82044 338008 82050 338020
rect 93118 338008 93124 338020
rect 82044 337980 93124 338008
rect 82044 337968 82050 337980
rect 93118 337968 93124 337980
rect 93176 337968 93182 338020
rect 99466 337968 99472 338020
rect 99524 338008 99530 338020
rect 103486 338008 103514 338048
rect 127986 338036 127992 338048
rect 128044 338036 128050 338088
rect 165982 338036 165988 338088
rect 166040 338076 166046 338088
rect 177298 338076 177304 338088
rect 166040 338048 177304 338076
rect 166040 338036 166046 338048
rect 177298 338036 177304 338048
rect 177356 338036 177362 338088
rect 178678 338036 178684 338088
rect 178736 338076 178742 338088
rect 184014 338076 184020 338088
rect 178736 338048 184020 338076
rect 178736 338036 178742 338048
rect 184014 338036 184020 338048
rect 184072 338036 184078 338088
rect 211706 338076 211712 338088
rect 190426 338048 211712 338076
rect 99524 337980 103514 338008
rect 99524 337968 99530 337980
rect 109678 337968 109684 338020
rect 109736 338008 109742 338020
rect 122098 338008 122104 338020
rect 109736 337980 122104 338008
rect 109736 337968 109742 337980
rect 122098 337968 122104 337980
rect 122156 337968 122162 338020
rect 137646 337968 137652 338020
rect 137704 338008 137710 338020
rect 148318 338008 148324 338020
rect 137704 337980 148324 338008
rect 137704 337968 137710 337980
rect 148318 337968 148324 337980
rect 148376 337968 148382 338020
rect 183646 337968 183652 338020
rect 183704 338008 183710 338020
rect 190426 338008 190454 338048
rect 211706 338036 211712 338048
rect 211764 338036 211770 338088
rect 277670 338036 277676 338088
rect 277728 338076 277734 338088
rect 289078 338076 289084 338088
rect 277728 338048 289084 338076
rect 277728 338036 277734 338048
rect 289078 338036 289084 338048
rect 289136 338036 289142 338088
rect 306006 338036 306012 338088
rect 306064 338076 306070 338088
rect 316678 338076 316684 338088
rect 306064 338048 316684 338076
rect 306064 338036 306070 338048
rect 316678 338036 316684 338048
rect 316736 338036 316742 338088
rect 361666 338036 361672 338088
rect 361724 338076 361730 338088
rect 373258 338076 373264 338088
rect 361724 338048 373264 338076
rect 361724 338036 361730 338048
rect 373258 338036 373264 338048
rect 373316 338036 373322 338088
rect 374638 338036 374644 338088
rect 374696 338076 374702 338088
rect 379698 338076 379704 338088
rect 374696 338048 379704 338076
rect 374696 338036 374702 338048
rect 379698 338036 379704 338048
rect 379756 338036 379762 338088
rect 408034 338076 408040 338088
rect 383626 338048 408040 338076
rect 183704 337980 190454 338008
rect 183704 337968 183710 337980
rect 193674 337968 193680 338020
rect 193732 338008 193738 338020
rect 204990 338008 204996 338020
rect 193732 337980 204996 338008
rect 193732 337968 193738 337980
rect 204990 337968 204996 337980
rect 205048 337968 205054 338020
rect 222010 337968 222016 338020
rect 222068 338008 222074 338020
rect 232498 338008 232504 338020
rect 222068 337980 232504 338008
rect 222068 337968 222074 337980
rect 232498 337968 232504 337980
rect 232556 337968 232562 338020
rect 249702 337968 249708 338020
rect 249760 338008 249766 338020
rect 260190 338008 260196 338020
rect 249760 337980 260196 338008
rect 249760 337968 249766 337980
rect 260190 337968 260196 337980
rect 260248 337968 260254 338020
rect 333698 337968 333704 338020
rect 333756 338008 333762 338020
rect 344278 338008 344284 338020
rect 333756 337980 344284 338008
rect 333756 337968 333762 337980
rect 344278 337968 344284 337980
rect 344336 337968 344342 338020
rect 379606 337968 379612 338020
rect 379664 338008 379670 338020
rect 383626 338008 383654 338048
rect 408034 338036 408040 338048
rect 408092 338036 408098 338088
rect 473998 338036 474004 338088
rect 474056 338076 474062 338088
rect 485038 338076 485044 338088
rect 474056 338048 485044 338076
rect 474056 338036 474062 338048
rect 485038 338036 485044 338048
rect 485096 338036 485102 338088
rect 501690 338036 501696 338088
rect 501748 338076 501754 338088
rect 512638 338076 512644 338088
rect 501748 338048 512644 338076
rect 501748 338036 501754 338048
rect 512638 338036 512644 338048
rect 512696 338036 512702 338088
rect 548150 338036 548156 338088
rect 548208 338076 548214 338088
rect 557534 338076 557540 338088
rect 548208 338048 557540 338076
rect 548208 338036 548214 338048
rect 557534 338036 557540 338048
rect 557592 338036 557598 338088
rect 379664 337980 383654 338008
rect 379664 337968 379670 337980
rect 390002 337968 390008 338020
rect 390060 338008 390066 338020
rect 400858 338008 400864 338020
rect 390060 337980 400864 338008
rect 390060 337968 390066 337980
rect 400858 337968 400864 337980
rect 400916 337968 400922 338020
rect 417694 337968 417700 338020
rect 417752 338008 417758 338020
rect 428550 338008 428556 338020
rect 417752 337980 428556 338008
rect 417752 337968 417758 337980
rect 428550 337968 428556 337980
rect 428608 337968 428614 338020
rect 445662 337968 445668 338020
rect 445720 338008 445726 338020
rect 456150 338008 456156 338020
rect 445720 337980 456156 338008
rect 445720 337968 445726 337980
rect 456150 337968 456156 337980
rect 456208 337968 456214 338020
rect 529658 337968 529664 338020
rect 529716 338008 529722 338020
rect 540238 338008 540244 338020
rect 529716 337980 540244 338008
rect 529716 337968 529722 337980
rect 540238 337968 540244 337980
rect 540296 337968 540302 338020
rect 72050 337940 72056 337952
rect 45526 337912 72056 337940
rect 72050 337900 72056 337912
rect 72108 337900 72114 337952
rect 127066 337900 127072 337952
rect 127124 337940 127130 337952
rect 156046 337940 156052 337952
rect 127124 337912 156052 337940
rect 127124 337900 127130 337912
rect 156046 337900 156052 337912
rect 156104 337900 156110 337952
rect 238846 337900 238852 337952
rect 238904 337940 238910 337952
rect 268010 337940 268016 337952
rect 238904 337912 268016 337940
rect 238904 337900 238910 337912
rect 268010 337900 268016 337912
rect 268068 337900 268074 337952
rect 323026 337900 323032 337952
rect 323084 337940 323090 337952
rect 352006 337940 352012 337952
rect 323084 337912 352012 337940
rect 323084 337900 323090 337912
rect 352006 337900 352012 337912
rect 352064 337900 352070 337952
rect 434806 337900 434812 337952
rect 434864 337940 434870 337952
rect 463694 337940 463700 337952
rect 434864 337912 463700 337940
rect 434864 337900 434870 337912
rect 463694 337900 463700 337912
rect 463752 337900 463758 337952
rect 518986 337900 518992 337952
rect 519044 337940 519050 337952
rect 547874 337940 547880 337952
rect 519044 337912 547880 337940
rect 519044 337900 519050 337912
rect 547874 337900 547880 337912
rect 547932 337900 547938 337952
rect 26234 335724 26240 335776
rect 26292 335764 26298 335776
rect 35434 335764 35440 335776
rect 26292 335736 35440 335764
rect 26292 335724 26298 335736
rect 35434 335724 35440 335736
rect 35492 335724 35498 335776
rect 71130 335452 71136 335504
rect 71188 335492 71194 335504
rect 82262 335492 82268 335504
rect 71188 335464 82268 335492
rect 71188 335452 71194 335464
rect 82262 335452 82268 335464
rect 82320 335452 82326 335504
rect 99374 335452 99380 335504
rect 99432 335492 99438 335504
rect 100294 335492 100300 335504
rect 99432 335464 100300 335492
rect 99432 335452 99438 335464
rect 100294 335452 100300 335464
rect 100352 335452 100358 335504
rect 183646 335452 183652 335504
rect 183704 335492 183710 335504
rect 222286 335492 222292 335504
rect 183704 335464 222292 335492
rect 183704 335452 183710 335464
rect 222286 335452 222292 335464
rect 222344 335452 222350 335504
rect 261478 335452 261484 335504
rect 261536 335492 261542 335504
rect 268286 335492 268292 335504
rect 261536 335464 268292 335492
rect 261536 335452 261542 335464
rect 268286 335452 268292 335464
rect 268344 335452 268350 335504
rect 295426 335452 295432 335504
rect 295484 335492 295490 335504
rect 334250 335492 334256 335504
rect 295484 335464 334256 335492
rect 295484 335452 295490 335464
rect 334250 335452 334256 335464
rect 334308 335452 334314 335504
rect 379606 335452 379612 335504
rect 379664 335492 379670 335504
rect 418246 335492 418252 335504
rect 379664 335464 418252 335492
rect 379664 335452 379670 335464
rect 418246 335452 418252 335464
rect 418304 335452 418310 335504
rect 463786 335452 463792 335504
rect 463844 335492 463850 335504
rect 463844 335464 470594 335492
rect 463844 335452 463850 335464
rect 36630 335384 36636 335436
rect 36688 335424 36694 335436
rect 53926 335424 53932 335436
rect 36688 335396 53932 335424
rect 36688 335384 36694 335396
rect 53926 335384 53932 335396
rect 53984 335384 53990 335436
rect 71866 335384 71872 335436
rect 71924 335424 71930 335436
rect 109954 335424 109960 335436
rect 71924 335396 109960 335424
rect 71924 335384 71930 335396
rect 109954 335384 109960 335396
rect 110012 335384 110018 335436
rect 124858 335384 124864 335436
rect 124916 335424 124922 335436
rect 128630 335424 128636 335436
rect 124916 335396 128636 335424
rect 124916 335384 124922 335396
rect 128630 335384 128636 335396
rect 128688 335384 128694 335436
rect 151078 335384 151084 335436
rect 151136 335424 151142 335436
rect 156598 335424 156604 335436
rect 151136 335396 156604 335424
rect 151136 335384 151142 335396
rect 156598 335384 156604 335396
rect 156656 335384 156662 335436
rect 182818 335384 182824 335436
rect 182876 335424 182882 335436
rect 193950 335424 193956 335436
rect 182876 335396 193956 335424
rect 182876 335384 182882 335396
rect 193950 335384 193956 335396
rect 194008 335384 194014 335436
rect 232498 335384 232504 335436
rect 232556 335424 232562 335436
rect 232556 335396 248414 335424
rect 232556 335384 232562 335396
rect 15102 335316 15108 335368
rect 15160 335356 15166 335368
rect 16574 335356 16580 335368
rect 15160 335328 16580 335356
rect 15160 335316 15166 335328
rect 16574 335316 16580 335328
rect 16632 335316 16638 335368
rect 66898 335316 66904 335368
rect 66956 335356 66962 335368
rect 72602 335356 72608 335368
rect 66956 335328 72608 335356
rect 66956 335316 66962 335328
rect 72602 335316 72608 335328
rect 72660 335316 72666 335368
rect 93118 335316 93124 335368
rect 93176 335356 93182 335368
rect 99374 335356 99380 335368
rect 93176 335328 99380 335356
rect 93176 335316 93182 335328
rect 99374 335316 99380 335328
rect 99432 335316 99438 335368
rect 99466 335316 99472 335368
rect 99524 335356 99530 335368
rect 138290 335356 138296 335368
rect 99524 335328 138296 335356
rect 99524 335316 99530 335328
rect 138290 335316 138296 335328
rect 138348 335316 138354 335368
rect 149698 335316 149704 335368
rect 149756 335356 149762 335368
rect 166258 335356 166264 335368
rect 149756 335328 166264 335356
rect 149756 335316 149762 335328
rect 166258 335316 166264 335328
rect 166316 335316 166322 335368
rect 177298 335316 177304 335368
rect 177356 335356 177362 335368
rect 184290 335356 184296 335368
rect 177356 335328 184296 335356
rect 177356 335316 177362 335328
rect 184290 335316 184296 335328
rect 184348 335316 184354 335368
rect 233970 335316 233976 335368
rect 234028 335356 234034 335368
rect 240594 335356 240600 335368
rect 234028 335328 240600 335356
rect 234028 335316 234034 335328
rect 240594 335316 240600 335328
rect 240652 335316 240658 335368
rect 248386 335356 248414 335396
rect 267826 335384 267832 335436
rect 267884 335424 267890 335436
rect 306282 335424 306288 335436
rect 267884 335396 306288 335424
rect 267884 335384 267890 335396
rect 306282 335384 306288 335396
rect 306340 335384 306346 335436
rect 352006 335384 352012 335436
rect 352064 335424 352070 335436
rect 390278 335424 390284 335436
rect 352064 335396 390284 335424
rect 352064 335384 352070 335396
rect 390278 335384 390284 335396
rect 390336 335384 390342 335436
rect 400858 335384 400864 335436
rect 400916 335424 400922 335436
rect 408586 335424 408592 335436
rect 400916 335396 408592 335424
rect 400916 335384 400922 335396
rect 408586 335384 408592 335396
rect 408644 335384 408650 335436
rect 429838 335384 429844 335436
rect 429896 335424 429902 335436
rect 436278 335424 436284 335436
rect 429896 335396 436284 335424
rect 429896 335384 429902 335396
rect 436278 335384 436284 335396
rect 436336 335384 436342 335436
rect 457438 335384 457444 335436
rect 457496 335424 457502 335436
rect 464614 335424 464620 335436
rect 457496 335396 464620 335424
rect 457496 335384 457502 335396
rect 464614 335384 464620 335396
rect 464672 335384 464678 335436
rect 470566 335424 470594 335464
rect 491386 335452 491392 335504
rect 491444 335492 491450 335504
rect 529934 335492 529940 335504
rect 491444 335464 529940 335492
rect 491444 335452 491450 335464
rect 529934 335452 529940 335464
rect 529992 335452 529998 335504
rect 502242 335424 502248 335436
rect 470566 335396 502248 335424
rect 502242 335384 502248 335396
rect 502300 335384 502306 335436
rect 512638 335384 512644 335436
rect 512696 335424 512702 335436
rect 520274 335424 520280 335436
rect 512696 335396 520280 335424
rect 512696 335384 512702 335396
rect 520274 335384 520280 335396
rect 520332 335384 520338 335436
rect 250254 335356 250260 335368
rect 248386 335328 250260 335356
rect 250254 335316 250260 335328
rect 250312 335316 250318 335368
rect 266998 335316 267004 335368
rect 267056 335356 267062 335368
rect 277946 335356 277952 335368
rect 267056 335328 277952 335356
rect 267056 335316 267062 335328
rect 277946 335316 277952 335328
rect 278004 335316 278010 335368
rect 289078 335316 289084 335368
rect 289136 335356 289142 335368
rect 296530 335356 296536 335368
rect 289136 335328 296536 335356
rect 289136 335316 289142 335328
rect 296530 335316 296536 335328
rect 296588 335316 296594 335368
rect 318058 335316 318064 335368
rect 318116 335356 318122 335368
rect 324590 335356 324596 335368
rect 318116 335328 324596 335356
rect 318116 335316 318122 335328
rect 324590 335316 324596 335328
rect 324648 335316 324654 335368
rect 347038 335316 347044 335368
rect 347096 335356 347102 335368
rect 361942 335356 361948 335368
rect 347096 335328 361948 335356
rect 347096 335316 347102 335328
rect 361942 335316 361948 335328
rect 362000 335316 362006 335368
rect 373258 335316 373264 335368
rect 373316 335356 373322 335368
rect 380618 335356 380624 335368
rect 373316 335328 380624 335356
rect 373316 335316 373322 335328
rect 380618 335316 380624 335328
rect 380676 335316 380682 335368
rect 428458 335316 428464 335368
rect 428516 335356 428522 335368
rect 445938 335356 445944 335368
rect 428516 335328 445944 335356
rect 428516 335316 428522 335328
rect 445938 335316 445944 335328
rect 445996 335316 446002 335368
rect 462958 335316 462964 335368
rect 463016 335356 463022 335368
rect 474274 335356 474280 335368
rect 463016 335328 474280 335356
rect 463016 335316 463022 335328
rect 474274 335316 474280 335328
rect 474332 335316 474338 335368
rect 485038 335316 485044 335368
rect 485096 335356 485102 335368
rect 492582 335356 492588 335368
rect 485096 335328 492588 335356
rect 485096 335316 485102 335328
rect 492582 335316 492588 335328
rect 492640 335316 492646 335368
rect 511810 335316 511816 335368
rect 511868 335356 511874 335368
rect 514018 335356 514024 335368
rect 511868 335328 514024 335356
rect 511868 335316 511874 335328
rect 514018 335316 514024 335328
rect 514076 335316 514082 335368
rect 541618 335316 541624 335368
rect 541676 335356 541682 335368
rect 558270 335356 558276 335368
rect 541676 335328 558276 335356
rect 541676 335316 541682 335328
rect 558270 335316 558276 335328
rect 558328 335316 558334 335368
rect 348418 332528 348424 332580
rect 348476 332568 348482 332580
rect 352282 332568 352288 332580
rect 348476 332540 352288 332568
rect 348476 332528 348482 332540
rect 352282 332528 352288 332540
rect 352340 332528 352346 332580
rect 544378 332528 544384 332580
rect 544436 332568 544442 332580
rect 548334 332568 548340 332580
rect 544436 332540 548340 332568
rect 544436 332528 544442 332540
rect 548334 332528 548340 332540
rect 548392 332528 548398 332580
rect 568022 332392 568028 332444
rect 568080 332392 568086 332444
rect 120166 332256 120172 332308
rect 120224 332296 120230 332308
rect 122098 332296 122104 332308
rect 120224 332268 122104 332296
rect 120224 332256 120230 332268
rect 122098 332256 122104 332268
rect 122156 332256 122162 332308
rect 568040 332240 568068 332392
rect 568022 332188 568028 332240
rect 568080 332188 568086 332240
rect 209682 331304 209688 331356
rect 209740 331344 209746 331356
rect 262214 331344 262220 331356
rect 209740 331316 262220 331344
rect 209740 331304 209746 331316
rect 262214 331304 262220 331316
rect 262272 331304 262278 331356
rect 204070 331236 204076 331288
rect 204128 331276 204134 331288
rect 212442 331276 212448 331288
rect 204128 331248 212448 331276
rect 204128 331236 204134 331248
rect 212442 331236 212448 331248
rect 212500 331236 212506 331288
rect 293862 331236 293868 331288
rect 293920 331276 293926 331288
rect 345014 331276 345020 331288
rect 293920 331248 345020 331276
rect 293920 331236 293926 331248
rect 345014 331236 345020 331248
rect 345072 331236 345078 331288
rect 405642 331236 405648 331288
rect 405700 331276 405706 331288
rect 458174 331276 458180 331288
rect 405700 331248 458180 331276
rect 405700 331236 405706 331248
rect 458174 331236 458180 331248
rect 458232 331236 458238 331288
rect 489822 331236 489828 331288
rect 489880 331276 489886 331288
rect 542354 331276 542360 331288
rect 489880 331248 542360 331276
rect 489880 331236 489886 331248
rect 542354 331236 542360 331248
rect 542412 331236 542418 331288
rect 204254 328992 204260 329044
rect 204312 329032 204318 329044
rect 204990 329032 204996 329044
rect 204312 329004 204996 329032
rect 204312 328992 204318 329004
rect 204990 328992 204996 329004
rect 205048 328992 205054 329044
rect 400306 328992 400312 329044
rect 400364 329032 400370 329044
rect 400950 329032 400956 329044
rect 400364 329004 400956 329032
rect 400364 328992 400370 329004
rect 400950 328992 400956 329004
rect 401008 328992 401014 329044
rect 570598 324300 570604 324352
rect 570656 324340 570662 324352
rect 579982 324340 579988 324352
rect 570656 324312 579988 324340
rect 570656 324300 570662 324312
rect 579982 324300 579988 324312
rect 580040 324300 580046 324352
rect 13538 314576 13544 314628
rect 13596 314616 13602 314628
rect 66254 314616 66260 314628
rect 13596 314588 66260 314616
rect 13596 314576 13602 314588
rect 66254 314576 66260 314588
rect 66312 314576 66318 314628
rect 70302 314576 70308 314628
rect 70360 314616 70366 314628
rect 121454 314616 121460 314628
rect 70360 314588 121460 314616
rect 70360 314576 70366 314588
rect 121454 314576 121460 314588
rect 121512 314576 121518 314628
rect 126882 314576 126888 314628
rect 126940 314616 126946 314628
rect 178034 314616 178040 314628
rect 126940 314588 178040 314616
rect 126940 314576 126946 314588
rect 178034 314576 178040 314588
rect 178092 314576 178098 314628
rect 182082 314576 182088 314628
rect 182140 314616 182146 314628
rect 233234 314616 233240 314628
rect 182140 314588 233240 314616
rect 182140 314576 182146 314588
rect 233234 314576 233240 314588
rect 233292 314576 233298 314628
rect 238662 314576 238668 314628
rect 238720 314616 238726 314628
rect 289814 314616 289820 314628
rect 238720 314588 289820 314616
rect 238720 314576 238726 314588
rect 289814 314576 289820 314588
rect 289872 314576 289878 314628
rect 322842 314576 322848 314628
rect 322900 314616 322906 314628
rect 373994 314616 374000 314628
rect 322900 314588 374000 314616
rect 322900 314576 322906 314588
rect 373994 314576 374000 314588
rect 374052 314576 374058 314628
rect 378042 314576 378048 314628
rect 378100 314616 378106 314628
rect 429286 314616 429292 314628
rect 378100 314588 429292 314616
rect 378100 314576 378106 314588
rect 429286 314576 429292 314588
rect 429344 314576 429350 314628
rect 434622 314576 434628 314628
rect 434680 314616 434686 314628
rect 485774 314616 485780 314628
rect 434680 314588 485780 314616
rect 434680 314576 434686 314588
rect 485774 314576 485780 314588
rect 485832 314576 485838 314628
rect 518802 314576 518808 314628
rect 518860 314616 518866 314628
rect 569954 314616 569960 314628
rect 518860 314588 569960 314616
rect 518860 314576 518866 314588
rect 569954 314576 569960 314588
rect 570012 314576 570018 314628
rect 42702 314508 42708 314560
rect 42760 314548 42766 314560
rect 93854 314548 93860 314560
rect 42760 314520 93860 314548
rect 42760 314508 42766 314520
rect 93854 314508 93860 314520
rect 93912 314508 93918 314560
rect 97902 314508 97908 314560
rect 97960 314548 97966 314560
rect 149054 314548 149060 314560
rect 97960 314520 149060 314548
rect 97960 314508 97966 314520
rect 149054 314508 149060 314520
rect 149112 314508 149118 314560
rect 154482 314508 154488 314560
rect 154540 314548 154546 314560
rect 205634 314548 205640 314560
rect 154540 314520 205640 314548
rect 154540 314508 154546 314520
rect 205634 314508 205640 314520
rect 205692 314508 205698 314560
rect 266262 314508 266268 314560
rect 266320 314548 266326 314560
rect 317414 314548 317420 314560
rect 266320 314520 317420 314548
rect 266320 314508 266326 314520
rect 317414 314508 317420 314520
rect 317472 314508 317478 314560
rect 350442 314508 350448 314560
rect 350500 314548 350506 314560
rect 401594 314548 401600 314560
rect 350500 314520 401600 314548
rect 350500 314508 350506 314520
rect 401594 314508 401600 314520
rect 401652 314508 401658 314560
rect 462222 314508 462228 314560
rect 462280 314548 462286 314560
rect 513374 314548 513380 314560
rect 462280 314520 513380 314548
rect 462280 314508 462286 314520
rect 513374 314508 513380 314520
rect 513432 314508 513438 314560
rect 15194 311788 15200 311840
rect 15252 311828 15258 311840
rect 35894 311828 35900 311840
rect 15252 311800 35900 311828
rect 15252 311788 15258 311800
rect 35894 311788 35900 311800
rect 35952 311788 35958 311840
rect 36078 311788 36084 311840
rect 36136 311828 36142 311840
rect 63586 311828 63592 311840
rect 36136 311800 63592 311828
rect 36136 311788 36142 311800
rect 63586 311788 63592 311800
rect 63644 311788 63650 311840
rect 64046 311788 64052 311840
rect 64104 311828 64110 311840
rect 91922 311828 91928 311840
rect 64104 311800 91928 311828
rect 64104 311788 64110 311800
rect 91922 311788 91928 311800
rect 91980 311788 91986 311840
rect 92106 311788 92112 311840
rect 92164 311828 92170 311840
rect 119614 311828 119620 311840
rect 92164 311800 119620 311828
rect 92164 311788 92170 311800
rect 119614 311788 119620 311800
rect 119672 311788 119678 311840
rect 122098 311788 122104 311840
rect 122156 311828 122162 311840
rect 147950 311828 147956 311840
rect 122156 311800 147956 311828
rect 122156 311788 122162 311800
rect 147950 311788 147956 311800
rect 148008 311788 148014 311840
rect 148042 311788 148048 311840
rect 148100 311828 148106 311840
rect 175918 311828 175924 311840
rect 148100 311800 175924 311828
rect 148100 311788 148106 311800
rect 175918 311788 175924 311800
rect 175976 311788 175982 311840
rect 176102 311788 176108 311840
rect 176160 311828 176166 311840
rect 203610 311828 203616 311840
rect 176160 311800 203616 311828
rect 176160 311788 176166 311800
rect 203610 311788 203616 311800
rect 203668 311788 203674 311840
rect 204990 311788 204996 311840
rect 205048 311828 205054 311840
rect 231946 311828 231952 311840
rect 205048 311800 231952 311828
rect 205048 311788 205054 311800
rect 231946 311788 231952 311800
rect 232004 311788 232010 311840
rect 232038 311788 232044 311840
rect 232096 311828 232102 311840
rect 259914 311828 259920 311840
rect 232096 311800 259920 311828
rect 232096 311788 232102 311800
rect 259914 311788 259920 311800
rect 259972 311788 259978 311840
rect 260098 311788 260104 311840
rect 260156 311828 260162 311840
rect 287606 311828 287612 311840
rect 260156 311800 287612 311828
rect 260156 311788 260162 311800
rect 287606 311788 287612 311800
rect 287664 311788 287670 311840
rect 288066 311788 288072 311840
rect 288124 311828 288130 311840
rect 315942 311828 315948 311840
rect 288124 311800 315948 311828
rect 288124 311788 288130 311800
rect 315942 311788 315948 311800
rect 316000 311788 316006 311840
rect 316678 311788 316684 311840
rect 316736 311828 316742 311840
rect 343910 311828 343916 311840
rect 316736 311800 343916 311828
rect 316736 311788 316742 311800
rect 343910 311788 343916 311800
rect 343968 311788 343974 311840
rect 344094 311788 344100 311840
rect 344152 311828 344158 311840
rect 371602 311828 371608 311840
rect 344152 311800 371608 311828
rect 344152 311788 344158 311800
rect 371602 311788 371608 311800
rect 371660 311788 371666 311840
rect 372062 311788 372068 311840
rect 372120 311828 372126 311840
rect 399938 311828 399944 311840
rect 372120 311800 399944 311828
rect 372120 311788 372126 311800
rect 399938 311788 399944 311800
rect 399996 311788 400002 311840
rect 400950 311788 400956 311840
rect 401008 311828 401014 311840
rect 427906 311828 427912 311840
rect 401008 311800 427912 311828
rect 401008 311788 401014 311800
rect 427906 311788 427912 311800
rect 427964 311788 427970 311840
rect 428090 311788 428096 311840
rect 428148 311828 428154 311840
rect 455598 311828 455604 311840
rect 428148 311800 455604 311828
rect 428148 311788 428154 311800
rect 455598 311788 455604 311800
rect 455656 311788 455662 311840
rect 456058 311788 456064 311840
rect 456116 311828 456122 311840
rect 483934 311828 483940 311840
rect 456116 311800 483940 311828
rect 456116 311788 456122 311800
rect 483934 311788 483940 311800
rect 483992 311788 483998 311840
rect 484026 311788 484032 311840
rect 484084 311828 484090 311840
rect 511902 311828 511908 311840
rect 484084 311800 511908 311828
rect 484084 311788 484090 311800
rect 511902 311788 511908 311800
rect 511960 311788 511966 311840
rect 514018 311788 514024 311840
rect 514076 311828 514082 311840
rect 539594 311828 539600 311840
rect 514076 311800 539600 311828
rect 514076 311788 514082 311800
rect 539594 311788 539600 311800
rect 539652 311788 539658 311840
rect 540054 311788 540060 311840
rect 540112 311828 540118 311840
rect 567930 311828 567936 311840
rect 540112 311800 567936 311828
rect 540112 311788 540118 311800
rect 567930 311788 567936 311800
rect 567988 311788 567994 311840
rect 16574 311720 16580 311772
rect 16632 311760 16638 311772
rect 36630 311760 36636 311772
rect 16632 311732 36636 311760
rect 16632 311720 16638 311732
rect 36630 311720 36636 311732
rect 36688 311720 36694 311772
rect 44910 311720 44916 311772
rect 44968 311760 44974 311772
rect 71130 311760 71136 311772
rect 44968 311732 71136 311760
rect 44968 311720 44974 311732
rect 71130 311720 71136 311732
rect 71188 311720 71194 311772
rect 82262 311720 82268 311772
rect 82320 311760 82326 311772
rect 93118 311760 93124 311772
rect 82320 311732 93124 311760
rect 82320 311720 82326 311732
rect 93118 311720 93124 311732
rect 93176 311720 93182 311772
rect 110230 311720 110236 311772
rect 110288 311760 110294 311772
rect 124858 311760 124864 311772
rect 110288 311732 124864 311760
rect 110288 311720 110294 311732
rect 124858 311720 124864 311732
rect 124916 311720 124922 311772
rect 128630 311720 128636 311772
rect 128688 311760 128694 311772
rect 149698 311760 149704 311772
rect 128688 311732 149704 311760
rect 128688 311720 128694 311732
rect 149698 311720 149704 311732
rect 149756 311720 149762 311772
rect 156598 311720 156604 311772
rect 156656 311760 156662 311772
rect 182818 311760 182824 311772
rect 156656 311732 182824 311760
rect 156656 311720 156662 311732
rect 182818 311720 182824 311732
rect 182876 311720 182882 311772
rect 194502 311720 194508 311772
rect 194560 311760 194566 311772
rect 204070 311760 204076 311772
rect 194560 311732 204076 311760
rect 194560 311720 194566 311732
rect 204070 311720 204076 311732
rect 204128 311720 204134 311772
rect 212626 311720 212632 311772
rect 212684 311760 212690 311772
rect 232498 311760 232504 311772
rect 212684 311732 232504 311760
rect 212684 311720 212690 311732
rect 232498 311720 232504 311732
rect 232556 311720 232562 311772
rect 240594 311720 240600 311772
rect 240652 311760 240658 311772
rect 266998 311760 267004 311772
rect 240652 311732 267004 311760
rect 240652 311720 240658 311732
rect 266998 311720 267004 311732
rect 267056 311720 267062 311772
rect 278590 311720 278596 311772
rect 278648 311760 278654 311772
rect 289078 311760 289084 311772
rect 278648 311732 289084 311760
rect 278648 311720 278654 311732
rect 289078 311720 289084 311732
rect 289136 311720 289142 311772
rect 306282 311720 306288 311772
rect 306340 311760 306346 311772
rect 318058 311760 318064 311772
rect 306340 311732 318064 311760
rect 306340 311720 306346 311732
rect 318058 311720 318064 311732
rect 318116 311720 318122 311772
rect 324590 311720 324596 311772
rect 324648 311760 324654 311772
rect 347038 311760 347044 311772
rect 324648 311732 347044 311760
rect 324648 311720 324654 311732
rect 347038 311720 347044 311732
rect 347096 311720 347102 311772
rect 362586 311720 362592 311772
rect 362644 311760 362650 311772
rect 373258 311760 373264 311772
rect 362644 311732 373264 311760
rect 362644 311720 362650 311732
rect 373258 311720 373264 311732
rect 373316 311720 373322 311772
rect 390278 311720 390284 311772
rect 390336 311760 390342 311772
rect 400858 311760 400864 311772
rect 390336 311732 400864 311760
rect 390336 311720 390342 311732
rect 400858 311720 400864 311732
rect 400916 311720 400922 311772
rect 408586 311720 408592 311772
rect 408644 311760 408650 311772
rect 428458 311760 428464 311772
rect 408644 311732 428464 311760
rect 408644 311720 408650 311732
rect 428458 311720 428464 311732
rect 428516 311720 428522 311772
rect 436922 311720 436928 311772
rect 436980 311760 436986 311772
rect 462958 311760 462964 311772
rect 436980 311732 462964 311760
rect 436980 311720 436986 311732
rect 462958 311720 462964 311732
rect 463016 311720 463022 311772
rect 474274 311720 474280 311772
rect 474332 311760 474338 311772
rect 485038 311760 485044 311772
rect 474332 311732 485044 311760
rect 474332 311720 474338 311732
rect 485038 311720 485044 311732
rect 485096 311720 485102 311772
rect 502242 311720 502248 311772
rect 502300 311760 502306 311772
rect 512638 311760 512644 311772
rect 502300 311732 512644 311760
rect 502300 311720 502306 311732
rect 512638 311720 512644 311732
rect 512696 311720 512702 311772
rect 520918 311720 520924 311772
rect 520976 311760 520982 311772
rect 541618 311760 541624 311772
rect 520976 311732 541624 311760
rect 520976 311720 520982 311732
rect 541618 311720 541624 311732
rect 541676 311720 541682 311772
rect 26234 311652 26240 311704
rect 26292 311692 26298 311704
rect 43530 311692 43536 311704
rect 26292 311664 43536 311692
rect 26292 311652 26298 311664
rect 43530 311652 43536 311664
rect 43588 311652 43594 311704
rect 54570 311652 54576 311704
rect 54628 311692 54634 311704
rect 66898 311692 66904 311704
rect 54628 311664 66904 311692
rect 54628 311652 54634 311664
rect 66898 311652 66904 311664
rect 66956 311652 66962 311704
rect 138290 311652 138296 311704
rect 138348 311692 138354 311704
rect 151078 311692 151084 311704
rect 138348 311664 151084 311692
rect 138348 311652 138354 311664
rect 151078 311652 151084 311664
rect 151136 311652 151142 311704
rect 166258 311652 166264 311704
rect 166316 311692 166322 311704
rect 177298 311692 177304 311704
rect 166316 311664 177304 311692
rect 166316 311652 166322 311664
rect 177298 311652 177304 311664
rect 177356 311652 177362 311704
rect 222286 311652 222292 311704
rect 222344 311692 222350 311704
rect 233970 311692 233976 311704
rect 222344 311664 233976 311692
rect 222344 311652 222350 311664
rect 233970 311652 233976 311664
rect 234028 311652 234034 311704
rect 250254 311652 250260 311704
rect 250312 311692 250318 311704
rect 261478 311692 261484 311704
rect 250312 311664 261484 311692
rect 250312 311652 250318 311664
rect 261478 311652 261484 311664
rect 261536 311652 261542 311704
rect 334250 311652 334256 311704
rect 334308 311692 334314 311704
rect 348418 311692 348424 311704
rect 334308 311664 348424 311692
rect 334308 311652 334314 311664
rect 348418 311652 348424 311664
rect 348476 311652 348482 311704
rect 418246 311652 418252 311704
rect 418304 311692 418310 311704
rect 429838 311692 429844 311704
rect 418304 311664 429844 311692
rect 418304 311652 418310 311664
rect 429838 311652 429844 311664
rect 429896 311652 429902 311704
rect 446582 311652 446588 311704
rect 446640 311692 446646 311704
rect 457438 311692 457444 311704
rect 446640 311664 457444 311692
rect 446640 311652 446646 311664
rect 457438 311652 457444 311664
rect 457496 311652 457502 311704
rect 530578 311652 530584 311704
rect 530636 311692 530642 311704
rect 544378 311692 544384 311704
rect 530636 311664 544384 311692
rect 530636 311652 530642 311664
rect 544378 311652 544384 311664
rect 544436 311652 544442 311704
rect 558270 311108 558276 311160
rect 558328 311148 558334 311160
rect 567470 311148 567476 311160
rect 558328 311120 567476 311148
rect 558328 311108 558334 311120
rect 567470 311108 567476 311120
rect 567528 311108 567534 311160
rect 548334 308388 548340 308440
rect 548392 308428 548398 308440
rect 568114 308428 568120 308440
rect 548392 308400 568120 308428
rect 548392 308388 548398 308400
rect 568114 308388 568120 308400
rect 568172 308388 568178 308440
rect 212258 307980 212264 308032
rect 212316 308020 212322 308032
rect 232682 308020 232688 308032
rect 212316 307992 232688 308020
rect 212316 307980 212322 307992
rect 232682 307980 232688 307992
rect 232740 307980 232746 308032
rect 296346 307980 296352 308032
rect 296404 308020 296410 308032
rect 316770 308020 316776 308032
rect 296404 307992 316776 308020
rect 296404 307980 296410 307992
rect 316770 307980 316776 307992
rect 316828 307980 316834 308032
rect 408034 307980 408040 308032
rect 408092 308020 408098 308032
rect 428642 308020 428648 308032
rect 408092 307992 428648 308020
rect 408092 307980 408098 307992
rect 428642 307980 428648 307992
rect 428700 307980 428706 308032
rect 148318 307912 148324 307964
rect 148376 307952 148382 307964
rect 165614 307952 165620 307964
rect 148376 307924 165620 307952
rect 148376 307912 148382 307924
rect 165614 307912 165620 307924
rect 165672 307912 165678 307964
rect 175458 307912 175464 307964
rect 175516 307952 175522 307964
rect 193674 307952 193680 307964
rect 175516 307924 193680 307952
rect 175516 307912 175522 307924
rect 193674 307912 193680 307924
rect 193732 307912 193738 307964
rect 203518 307912 203524 307964
rect 203576 307952 203582 307964
rect 221366 307952 221372 307964
rect 203576 307924 221372 307952
rect 203576 307912 203582 307924
rect 221366 307912 221372 307924
rect 221424 307912 221430 307964
rect 260190 307912 260196 307964
rect 260248 307952 260254 307964
rect 277670 307952 277676 307964
rect 260248 307924 277676 307952
rect 260248 307912 260254 307924
rect 277670 307912 277676 307924
rect 277728 307912 277734 307964
rect 287514 307912 287520 307964
rect 287572 307952 287578 307964
rect 305362 307952 305368 307964
rect 287572 307924 305368 307952
rect 287572 307912 287578 307924
rect 305362 307912 305368 307924
rect 305420 307912 305426 307964
rect 345658 307912 345664 307964
rect 345716 307952 345722 307964
rect 361666 307952 361672 307964
rect 345716 307924 361672 307952
rect 345716 307912 345722 307924
rect 361666 307912 361672 307924
rect 361724 307912 361730 307964
rect 371510 307912 371516 307964
rect 371568 307952 371574 307964
rect 389358 307952 389364 307964
rect 371568 307924 389364 307952
rect 371568 307912 371574 307924
rect 389358 307912 389364 307924
rect 389416 307912 389422 307964
rect 399478 307912 399484 307964
rect 399536 307952 399542 307964
rect 417694 307952 417700 307964
rect 399536 307924 417700 307952
rect 399536 307912 399542 307924
rect 417694 307912 417700 307924
rect 417752 307912 417758 307964
rect 456150 307912 456156 307964
rect 456208 307952 456214 307964
rect 473538 307952 473544 307964
rect 456208 307924 473544 307952
rect 456208 307912 456214 307924
rect 473538 307912 473544 307924
rect 473596 307912 473602 307964
rect 483474 307912 483480 307964
rect 483532 307952 483538 307964
rect 501690 307952 501696 307964
rect 483532 307924 501696 307952
rect 483532 307912 483538 307924
rect 501690 307912 501696 307924
rect 501748 307912 501754 307964
rect 511442 307912 511448 307964
rect 511500 307952 511506 307964
rect 529658 307952 529664 307964
rect 511500 307924 529664 307952
rect 511500 307912 511506 307924
rect 529658 307912 529664 307924
rect 529716 307912 529722 307964
rect 36722 307844 36728 307896
rect 36780 307884 36786 307896
rect 53650 307884 53656 307896
rect 36780 307856 53656 307884
rect 36780 307844 36786 307856
rect 53650 307844 53656 307856
rect 53708 307844 53714 307896
rect 64414 307844 64420 307896
rect 64472 307884 64478 307896
rect 81434 307884 81440 307896
rect 64472 307856 81440 307884
rect 64472 307844 64478 307856
rect 81434 307844 81440 307856
rect 81492 307844 81498 307896
rect 91462 307844 91468 307896
rect 91520 307884 91526 307896
rect 109678 307884 109684 307896
rect 91520 307856 109684 307884
rect 91520 307844 91526 307856
rect 109678 307844 109684 307856
rect 109736 307844 109742 307896
rect 119430 307844 119436 307896
rect 119488 307884 119494 307896
rect 137646 307884 137652 307896
rect 119488 307856 137652 307884
rect 119488 307844 119494 307856
rect 137646 307844 137652 307856
rect 137704 307844 137710 307896
rect 156322 307844 156328 307896
rect 156380 307884 156386 307896
rect 178678 307884 178684 307896
rect 156380 307856 178684 307884
rect 156380 307844 156386 307856
rect 178678 307844 178684 307856
rect 178736 307844 178742 307896
rect 232498 307844 232504 307896
rect 232556 307884 232562 307896
rect 249702 307884 249708 307896
rect 232556 307856 249708 307884
rect 232556 307844 232562 307856
rect 249702 307844 249708 307856
rect 249760 307844 249766 307896
rect 268010 307844 268016 307896
rect 268068 307884 268074 307896
rect 287698 307884 287704 307896
rect 268068 307856 287704 307884
rect 268068 307844 268074 307856
rect 287698 307844 287704 307856
rect 287756 307844 287762 307896
rect 315482 307844 315488 307896
rect 315540 307884 315546 307896
rect 333698 307884 333704 307896
rect 315540 307856 333704 307884
rect 315540 307844 315546 307856
rect 333698 307844 333704 307856
rect 333756 307844 333762 307896
rect 352006 307844 352012 307896
rect 352064 307884 352070 307896
rect 374638 307884 374644 307896
rect 352064 307856 374644 307884
rect 352064 307844 352070 307856
rect 374638 307844 374644 307856
rect 374696 307844 374702 307896
rect 428550 307844 428556 307896
rect 428608 307884 428614 307896
rect 445662 307884 445668 307896
rect 428608 307856 445668 307884
rect 428608 307844 428614 307856
rect 445662 307844 445668 307856
rect 445720 307844 445726 307896
rect 464338 307844 464344 307896
rect 464396 307884 464402 307896
rect 483658 307884 483664 307896
rect 464396 307856 483664 307884
rect 464396 307844 464402 307856
rect 483658 307844 483664 307856
rect 483716 307844 483722 307896
rect 492030 307844 492036 307896
rect 492088 307884 492094 307896
rect 512730 307884 512736 307896
rect 492088 307856 512736 307884
rect 492088 307844 492094 307856
rect 512730 307844 512736 307856
rect 512788 307844 512794 307896
rect 541618 307844 541624 307896
rect 541676 307884 541682 307896
rect 557534 307884 557540 307896
rect 541676 307856 557540 307884
rect 541676 307844 541682 307856
rect 557534 307844 557540 307856
rect 557592 307844 557598 307896
rect 15102 307776 15108 307828
rect 15160 307816 15166 307828
rect 25682 307816 25688 307828
rect 15160 307788 25688 307816
rect 15160 307776 15166 307788
rect 25682 307776 25688 307788
rect 25740 307776 25746 307828
rect 36630 307776 36636 307828
rect 36688 307816 36694 307828
rect 63310 307816 63316 307828
rect 36688 307788 63316 307816
rect 36688 307776 36694 307788
rect 63310 307776 63316 307788
rect 63368 307776 63374 307828
rect 66898 307776 66904 307828
rect 66956 307816 66962 307828
rect 91094 307816 91100 307828
rect 66956 307788 91100 307816
rect 66956 307776 66962 307788
rect 91094 307776 91100 307788
rect 91152 307776 91158 307828
rect 93118 307776 93124 307828
rect 93176 307816 93182 307828
rect 119338 307816 119344 307828
rect 93176 307788 119344 307816
rect 93176 307776 93182 307788
rect 119338 307776 119344 307788
rect 119396 307776 119402 307828
rect 122098 307776 122104 307828
rect 122156 307816 122162 307828
rect 147306 307816 147312 307828
rect 122156 307788 147312 307816
rect 122156 307776 122162 307788
rect 147306 307776 147312 307788
rect 147364 307776 147370 307828
rect 148410 307776 148416 307828
rect 148468 307816 148474 307828
rect 175274 307816 175280 307828
rect 148468 307788 175280 307816
rect 148468 307776 148474 307788
rect 175274 307776 175280 307788
rect 175332 307776 175338 307828
rect 177298 307776 177304 307828
rect 177356 307816 177362 307828
rect 203334 307816 203340 307828
rect 177356 307788 203340 307816
rect 177356 307776 177362 307788
rect 203334 307776 203340 307788
rect 203392 307776 203398 307828
rect 204990 307776 204996 307828
rect 205048 307816 205054 307828
rect 231026 307816 231032 307828
rect 205048 307788 231032 307816
rect 205048 307776 205054 307788
rect 231026 307776 231032 307788
rect 231084 307776 231090 307828
rect 232590 307776 232596 307828
rect 232648 307816 232654 307828
rect 259362 307816 259368 307828
rect 232648 307788 259368 307816
rect 232648 307776 232654 307788
rect 259362 307776 259368 307788
rect 259420 307776 259426 307828
rect 260098 307776 260104 307828
rect 260156 307816 260162 307828
rect 287330 307816 287336 307828
rect 260156 307788 287336 307816
rect 260156 307776 260162 307788
rect 287330 307776 287336 307788
rect 287388 307776 287394 307828
rect 289078 307776 289084 307828
rect 289136 307816 289142 307828
rect 315022 307816 315028 307828
rect 289136 307788 315028 307816
rect 289136 307776 289142 307788
rect 315022 307776 315028 307788
rect 315080 307776 315086 307828
rect 316678 307776 316684 307828
rect 316736 307816 316742 307828
rect 343358 307816 343364 307828
rect 316736 307788 343364 307816
rect 316736 307776 316742 307788
rect 343358 307776 343364 307788
rect 343416 307776 343422 307828
rect 344278 307776 344284 307828
rect 344336 307816 344342 307828
rect 371326 307816 371332 307828
rect 344336 307788 371332 307816
rect 344336 307776 344342 307788
rect 371326 307776 371332 307788
rect 371384 307776 371390 307828
rect 373258 307776 373264 307828
rect 373316 307816 373322 307828
rect 399018 307816 399024 307828
rect 373316 307788 399024 307816
rect 373316 307776 373322 307788
rect 399018 307776 399024 307788
rect 399076 307776 399082 307828
rect 400858 307776 400864 307828
rect 400916 307816 400922 307828
rect 427354 307816 427360 307828
rect 400916 307788 427360 307816
rect 400916 307776 400922 307788
rect 427354 307776 427360 307788
rect 427412 307776 427418 307828
rect 428458 307776 428464 307828
rect 428516 307816 428522 307828
rect 455322 307816 455328 307828
rect 428516 307788 455328 307816
rect 428516 307776 428522 307788
rect 455322 307776 455328 307788
rect 455380 307776 455386 307828
rect 456058 307776 456064 307828
rect 456116 307816 456122 307828
rect 483198 307816 483204 307828
rect 456116 307788 483204 307816
rect 456116 307776 456122 307788
rect 483198 307776 483204 307788
rect 483256 307776 483262 307828
rect 485038 307776 485044 307828
rect 485096 307816 485102 307828
rect 511350 307816 511356 307828
rect 485096 307788 511356 307816
rect 485096 307776 485102 307788
rect 511350 307776 511356 307788
rect 511408 307776 511414 307828
rect 512638 307776 512644 307828
rect 512696 307816 512702 307828
rect 539318 307816 539324 307828
rect 512696 307788 539324 307816
rect 512696 307776 512702 307788
rect 539318 307776 539324 307788
rect 539376 307776 539382 307828
rect 540238 307776 540244 307828
rect 540296 307816 540302 307828
rect 567194 307816 567200 307828
rect 540296 307788 567200 307816
rect 540296 307776 540302 307788
rect 567194 307776 567200 307788
rect 567252 307776 567258 307828
rect 42886 300976 42892 301028
rect 42944 301016 42950 301028
rect 43622 301016 43628 301028
rect 42944 300988 43628 301016
rect 42944 300976 42950 300988
rect 43622 300976 43628 300988
rect 43680 300976 43686 301028
rect 3326 293088 3332 293140
rect 3384 293128 3390 293140
rect 7558 293128 7564 293140
rect 3384 293100 7564 293128
rect 3384 293088 3390 293100
rect 7558 293088 7564 293100
rect 7616 293088 7622 293140
rect 63586 291864 63592 291916
rect 63644 291904 63650 291916
rect 64414 291904 64420 291916
rect 63644 291876 64420 291904
rect 63644 291864 63650 291876
rect 64414 291864 64420 291876
rect 64472 291864 64478 291916
rect 259730 291864 259736 291916
rect 259788 291904 259794 291916
rect 260190 291904 260196 291916
rect 259788 291876 260196 291904
rect 259788 291864 259794 291876
rect 260190 291864 260196 291876
rect 260248 291864 260254 291916
rect 455690 291864 455696 291916
rect 455748 291904 455754 291916
rect 456150 291904 456156 291916
rect 455748 291876 456156 291904
rect 455748 291864 455754 291876
rect 456150 291864 456156 291876
rect 456208 291864 456214 291916
rect 287698 288328 287704 288380
rect 287756 288368 287762 288380
rect 295702 288368 295708 288380
rect 287756 288340 295708 288368
rect 287756 288328 287762 288340
rect 295702 288328 295708 288340
rect 295760 288328 295766 288380
rect 316770 288328 316776 288380
rect 316828 288368 316834 288380
rect 323670 288368 323676 288380
rect 316828 288340 323676 288368
rect 316828 288328 316834 288340
rect 323670 288328 323676 288340
rect 323728 288328 323734 288380
rect 232682 287920 232688 287972
rect 232740 287960 232746 287972
rect 239766 287960 239772 287972
rect 232740 287932 239772 287960
rect 232740 287920 232746 287932
rect 239766 287920 239772 287932
rect 239824 287920 239830 287972
rect 428642 287648 428648 287700
rect 428700 287688 428706 287700
rect 435726 287688 435732 287700
rect 428700 287660 435732 287688
rect 428700 287648 428706 287660
rect 435726 287648 435732 287660
rect 435784 287648 435790 287700
rect 512730 287512 512736 287564
rect 512788 287552 512794 287564
rect 519630 287552 519636 287564
rect 512788 287524 519636 287552
rect 512788 287512 512794 287524
rect 519630 287512 519636 287524
rect 519688 287512 519694 287564
rect 483658 287376 483664 287428
rect 483716 287416 483722 287428
rect 491662 287416 491668 287428
rect 483716 287388 491668 287416
rect 483716 287376 483722 287388
rect 491662 287376 491668 287388
rect 491720 287376 491726 287428
rect 13538 286968 13544 287020
rect 13596 287008 13602 287020
rect 66254 287008 66260 287020
rect 13596 286980 66260 287008
rect 13596 286968 13602 286980
rect 66254 286968 66260 286980
rect 66312 286968 66318 287020
rect 70302 286968 70308 287020
rect 70360 287008 70366 287020
rect 121454 287008 121460 287020
rect 70360 286980 121460 287008
rect 70360 286968 70366 286980
rect 121454 286968 121460 286980
rect 121512 286968 121518 287020
rect 154482 286968 154488 287020
rect 154540 287008 154546 287020
rect 205634 287008 205640 287020
rect 154540 286980 205640 287008
rect 154540 286968 154546 286980
rect 205634 286968 205640 286980
rect 205692 286968 205698 287020
rect 209682 286968 209688 287020
rect 209740 287008 209746 287020
rect 262214 287008 262220 287020
rect 209740 286980 262220 287008
rect 209740 286968 209746 286980
rect 262214 286968 262220 286980
rect 262272 286968 262278 287020
rect 266262 286968 266268 287020
rect 266320 287008 266326 287020
rect 317414 287008 317420 287020
rect 266320 286980 317420 287008
rect 266320 286968 266326 286980
rect 317414 286968 317420 286980
rect 317472 286968 317478 287020
rect 322842 286968 322848 287020
rect 322900 287008 322906 287020
rect 373994 287008 374000 287020
rect 322900 286980 374000 287008
rect 322900 286968 322906 286980
rect 373994 286968 374000 286980
rect 374052 286968 374058 287020
rect 405642 286968 405648 287020
rect 405700 287008 405706 287020
rect 458174 287008 458180 287020
rect 405700 286980 458180 287008
rect 405700 286968 405706 286980
rect 458174 286968 458180 286980
rect 458232 286968 458238 287020
rect 489822 286968 489828 287020
rect 489880 287008 489886 287020
rect 542354 287008 542360 287020
rect 489880 286980 542360 287008
rect 489880 286968 489886 286980
rect 542354 286968 542360 286980
rect 542412 286968 542418 287020
rect 42702 286900 42708 286952
rect 42760 286940 42766 286952
rect 93854 286940 93860 286952
rect 42760 286912 93860 286940
rect 42760 286900 42766 286912
rect 93854 286900 93860 286912
rect 93912 286900 93918 286952
rect 97902 286900 97908 286952
rect 97960 286940 97966 286952
rect 149054 286940 149060 286952
rect 97960 286912 149060 286940
rect 97960 286900 97966 286912
rect 149054 286900 149060 286912
rect 149112 286900 149118 286952
rect 182082 286900 182088 286952
rect 182140 286940 182146 286952
rect 233234 286940 233240 286952
rect 182140 286912 233240 286940
rect 182140 286900 182146 286912
rect 233234 286900 233240 286912
rect 233292 286900 233298 286952
rect 238662 286900 238668 286952
rect 238720 286940 238726 286952
rect 289814 286940 289820 286952
rect 238720 286912 289820 286940
rect 238720 286900 238726 286912
rect 289814 286900 289820 286912
rect 289872 286900 289878 286952
rect 293862 286900 293868 286952
rect 293920 286940 293926 286952
rect 293920 286912 335354 286940
rect 293920 286900 293926 286912
rect 126882 286832 126888 286884
rect 126940 286872 126946 286884
rect 178034 286872 178040 286884
rect 126940 286844 178040 286872
rect 126940 286832 126946 286844
rect 178034 286832 178040 286844
rect 178092 286832 178098 286884
rect 335326 286872 335354 286912
rect 343542 286900 343548 286952
rect 343600 286940 343606 286952
rect 345658 286940 345664 286952
rect 343600 286912 345664 286940
rect 343600 286900 343606 286912
rect 345658 286900 345664 286912
rect 345716 286900 345722 286952
rect 378042 286900 378048 286952
rect 378100 286940 378106 286952
rect 429286 286940 429292 286952
rect 378100 286912 429292 286940
rect 378100 286900 378106 286912
rect 429286 286900 429292 286912
rect 429344 286900 429350 286952
rect 434622 286900 434628 286952
rect 434680 286940 434686 286952
rect 485774 286940 485780 286952
rect 434680 286912 485780 286940
rect 434680 286900 434686 286912
rect 485774 286900 485780 286912
rect 485832 286900 485838 286952
rect 518802 286900 518808 286952
rect 518860 286940 518866 286952
rect 569954 286940 569960 286952
rect 518860 286912 569960 286940
rect 518860 286900 518866 286912
rect 569954 286900 569960 286912
rect 570012 286900 570018 286952
rect 345014 286872 345020 286884
rect 335326 286844 345020 286872
rect 345014 286832 345020 286844
rect 345072 286832 345078 286884
rect 350442 286832 350448 286884
rect 350500 286872 350506 286884
rect 401594 286872 401600 286884
rect 350500 286844 401600 286872
rect 350500 286832 350506 286844
rect 401594 286832 401600 286844
rect 401652 286832 401658 286884
rect 462222 286832 462228 286884
rect 462280 286872 462286 286884
rect 513374 286872 513380 286884
rect 462280 286844 513380 286872
rect 462280 286832 462286 286844
rect 513374 286832 513380 286844
rect 513432 286832 513438 286884
rect 427722 286764 427728 286816
rect 427780 286804 427786 286816
rect 428550 286804 428556 286816
rect 427780 286776 428556 286804
rect 427780 286764 427786 286776
rect 428550 286764 428556 286776
rect 428608 286764 428614 286816
rect 539502 286764 539508 286816
rect 539560 286804 539566 286816
rect 541618 286804 541624 286816
rect 539560 286776 541624 286804
rect 539560 286764 539566 286776
rect 541618 286764 541624 286776
rect 541676 286764 541682 286816
rect 35250 286696 35256 286748
rect 35308 286736 35314 286748
rect 36722 286736 36728 286748
rect 35308 286708 36728 286736
rect 35308 286696 35314 286708
rect 36722 286696 36728 286708
rect 36780 286696 36786 286748
rect 547874 286152 547880 286204
rect 547932 286192 547938 286204
rect 548150 286192 548156 286204
rect 547932 286164 548156 286192
rect 547932 286152 547938 286164
rect 548150 286152 548156 286164
rect 548208 286152 548214 286204
rect 15102 285676 15108 285728
rect 15160 285716 15166 285728
rect 16574 285716 16580 285728
rect 15160 285688 16580 285716
rect 15160 285676 15166 285688
rect 16574 285676 16580 285688
rect 16632 285676 16638 285728
rect 71866 284248 71872 284300
rect 71924 284288 71930 284300
rect 100018 284288 100024 284300
rect 71924 284260 100024 284288
rect 71924 284248 71930 284260
rect 100018 284248 100024 284260
rect 100076 284248 100082 284300
rect 127986 284288 127992 284300
rect 103486 284260 127992 284288
rect 25682 284180 25688 284232
rect 25740 284220 25746 284232
rect 36630 284220 36636 284232
rect 25740 284192 36636 284220
rect 25740 284180 25746 284192
rect 36630 284180 36636 284192
rect 36688 284180 36694 284232
rect 42886 284180 42892 284232
rect 42944 284220 42950 284232
rect 42944 284192 45554 284220
rect 42944 284180 42950 284192
rect 15286 284112 15292 284164
rect 15344 284152 15350 284164
rect 43990 284152 43996 284164
rect 15344 284124 43996 284152
rect 15344 284112 15350 284124
rect 43990 284112 43996 284124
rect 44048 284112 44054 284164
rect 45526 284152 45554 284192
rect 53650 284180 53656 284232
rect 53708 284220 53714 284232
rect 66898 284220 66904 284232
rect 53708 284192 66904 284220
rect 53708 284180 53714 284192
rect 66898 284180 66904 284192
rect 66956 284180 66962 284232
rect 81986 284180 81992 284232
rect 82044 284220 82050 284232
rect 93118 284220 93124 284232
rect 82044 284192 93124 284220
rect 82044 284180 82050 284192
rect 93118 284180 93124 284192
rect 93176 284180 93182 284232
rect 99466 284180 99472 284232
rect 99524 284220 99530 284232
rect 103486 284220 103514 284260
rect 127986 284248 127992 284260
rect 128044 284248 128050 284300
rect 165982 284248 165988 284300
rect 166040 284288 166046 284300
rect 177298 284288 177304 284300
rect 166040 284260 177304 284288
rect 166040 284248 166046 284260
rect 177298 284248 177304 284260
rect 177356 284248 177362 284300
rect 178678 284248 178684 284300
rect 178736 284288 178742 284300
rect 184014 284288 184020 284300
rect 178736 284260 184020 284288
rect 178736 284248 178742 284260
rect 184014 284248 184020 284260
rect 184072 284248 184078 284300
rect 211706 284288 211712 284300
rect 190426 284260 211712 284288
rect 99524 284192 103514 284220
rect 99524 284180 99530 284192
rect 109678 284180 109684 284232
rect 109736 284220 109742 284232
rect 122098 284220 122104 284232
rect 109736 284192 122104 284220
rect 109736 284180 109742 284192
rect 122098 284180 122104 284192
rect 122156 284180 122162 284232
rect 137646 284180 137652 284232
rect 137704 284220 137710 284232
rect 148410 284220 148416 284232
rect 137704 284192 148416 284220
rect 137704 284180 137710 284192
rect 148410 284180 148416 284192
rect 148468 284180 148474 284232
rect 183646 284180 183652 284232
rect 183704 284220 183710 284232
rect 190426 284220 190454 284260
rect 211706 284248 211712 284260
rect 211764 284248 211770 284300
rect 277670 284248 277676 284300
rect 277728 284288 277734 284300
rect 289078 284288 289084 284300
rect 277728 284260 289084 284288
rect 277728 284248 277734 284260
rect 289078 284248 289084 284260
rect 289136 284248 289142 284300
rect 306006 284248 306012 284300
rect 306064 284288 306070 284300
rect 316678 284288 316684 284300
rect 306064 284260 316684 284288
rect 306064 284248 306070 284260
rect 316678 284248 316684 284260
rect 316736 284248 316742 284300
rect 361666 284248 361672 284300
rect 361724 284288 361730 284300
rect 373258 284288 373264 284300
rect 361724 284260 373264 284288
rect 361724 284248 361730 284260
rect 373258 284248 373264 284260
rect 373316 284248 373322 284300
rect 374638 284248 374644 284300
rect 374696 284288 374702 284300
rect 379698 284288 379704 284300
rect 374696 284260 379704 284288
rect 374696 284248 374702 284260
rect 379698 284248 379704 284260
rect 379756 284248 379762 284300
rect 408034 284288 408040 284300
rect 383626 284260 408040 284288
rect 183704 284192 190454 284220
rect 183704 284180 183710 284192
rect 193674 284180 193680 284232
rect 193732 284220 193738 284232
rect 204990 284220 204996 284232
rect 193732 284192 204996 284220
rect 193732 284180 193738 284192
rect 204990 284180 204996 284192
rect 205048 284180 205054 284232
rect 222010 284180 222016 284232
rect 222068 284220 222074 284232
rect 232590 284220 232596 284232
rect 222068 284192 232596 284220
rect 222068 284180 222074 284192
rect 232590 284180 232596 284192
rect 232648 284180 232654 284232
rect 249702 284180 249708 284232
rect 249760 284220 249766 284232
rect 260098 284220 260104 284232
rect 249760 284192 260104 284220
rect 249760 284180 249766 284192
rect 260098 284180 260104 284192
rect 260156 284180 260162 284232
rect 333698 284180 333704 284232
rect 333756 284220 333762 284232
rect 344278 284220 344284 284232
rect 333756 284192 344284 284220
rect 333756 284180 333762 284192
rect 344278 284180 344284 284192
rect 344336 284180 344342 284232
rect 379606 284180 379612 284232
rect 379664 284220 379670 284232
rect 383626 284220 383654 284260
rect 408034 284248 408040 284260
rect 408092 284248 408098 284300
rect 473998 284248 474004 284300
rect 474056 284288 474062 284300
rect 485038 284288 485044 284300
rect 474056 284260 485044 284288
rect 474056 284248 474062 284260
rect 485038 284248 485044 284260
rect 485096 284248 485102 284300
rect 501690 284248 501696 284300
rect 501748 284288 501754 284300
rect 512638 284288 512644 284300
rect 501748 284260 512644 284288
rect 501748 284248 501754 284260
rect 512638 284248 512644 284260
rect 512696 284248 512702 284300
rect 548150 284248 548156 284300
rect 548208 284288 548214 284300
rect 557534 284288 557540 284300
rect 548208 284260 557540 284288
rect 548208 284248 548214 284260
rect 557534 284248 557540 284260
rect 557592 284248 557598 284300
rect 379664 284192 383654 284220
rect 379664 284180 379670 284192
rect 390002 284180 390008 284232
rect 390060 284220 390066 284232
rect 400858 284220 400864 284232
rect 390060 284192 400864 284220
rect 390060 284180 390066 284192
rect 400858 284180 400864 284192
rect 400916 284180 400922 284232
rect 417694 284180 417700 284232
rect 417752 284220 417758 284232
rect 428458 284220 428464 284232
rect 417752 284192 428464 284220
rect 417752 284180 417758 284192
rect 428458 284180 428464 284192
rect 428516 284180 428522 284232
rect 445662 284180 445668 284232
rect 445720 284220 445726 284232
rect 456058 284220 456064 284232
rect 445720 284192 456064 284220
rect 445720 284180 445726 284192
rect 456058 284180 456064 284192
rect 456116 284180 456122 284232
rect 529658 284180 529664 284232
rect 529716 284220 529722 284232
rect 540238 284220 540244 284232
rect 529716 284192 540244 284220
rect 529716 284180 529722 284192
rect 540238 284180 540244 284192
rect 540296 284180 540302 284232
rect 72050 284152 72056 284164
rect 45526 284124 72056 284152
rect 72050 284112 72056 284124
rect 72108 284112 72114 284164
rect 127066 284112 127072 284164
rect 127124 284152 127130 284164
rect 156046 284152 156052 284164
rect 127124 284124 156052 284152
rect 127124 284112 127130 284124
rect 156046 284112 156052 284124
rect 156104 284112 156110 284164
rect 238846 284112 238852 284164
rect 238904 284152 238910 284164
rect 268010 284152 268016 284164
rect 238904 284124 268016 284152
rect 238904 284112 238910 284124
rect 268010 284112 268016 284124
rect 268068 284112 268074 284164
rect 323026 284112 323032 284164
rect 323084 284152 323090 284164
rect 352006 284152 352012 284164
rect 323084 284124 352012 284152
rect 323084 284112 323090 284124
rect 352006 284112 352012 284124
rect 352064 284112 352070 284164
rect 434806 284112 434812 284164
rect 434864 284152 434870 284164
rect 463694 284152 463700 284164
rect 434864 284124 463700 284152
rect 434864 284112 434870 284124
rect 463694 284112 463700 284124
rect 463752 284112 463758 284164
rect 518986 284112 518992 284164
rect 519044 284152 519050 284164
rect 547874 284152 547880 284164
rect 519044 284124 547880 284152
rect 519044 284112 519050 284124
rect 547874 284112 547880 284124
rect 547932 284112 547938 284164
rect 26234 280372 26240 280424
rect 26292 280412 26298 280424
rect 35434 280412 35440 280424
rect 26292 280384 35440 280412
rect 26292 280372 26298 280384
rect 35434 280372 35440 280384
rect 35492 280372 35498 280424
rect 71866 280372 71872 280424
rect 71924 280412 71930 280424
rect 71924 280384 74534 280412
rect 71924 280372 71930 280384
rect 71130 280304 71136 280356
rect 71188 280344 71194 280356
rect 71188 280316 72832 280344
rect 71188 280304 71194 280316
rect 36630 280236 36636 280288
rect 36688 280276 36694 280288
rect 53926 280276 53932 280288
rect 36688 280248 53932 280276
rect 36688 280236 36694 280248
rect 53926 280236 53932 280248
rect 53984 280236 53990 280288
rect 39298 280168 39304 280220
rect 39356 280208 39362 280220
rect 44266 280208 44272 280220
rect 39356 280180 44272 280208
rect 39356 280168 39362 280180
rect 44266 280168 44272 280180
rect 44324 280168 44330 280220
rect 66898 280168 66904 280220
rect 66956 280208 66962 280220
rect 72602 280208 72608 280220
rect 66956 280180 72608 280208
rect 66956 280168 66962 280180
rect 72602 280168 72608 280180
rect 72660 280168 72666 280220
rect 72804 280208 72832 280316
rect 74506 280276 74534 280384
rect 352006 280372 352012 280424
rect 352064 280412 352070 280424
rect 352064 280384 354674 280412
rect 352064 280372 352070 280384
rect 99466 280304 99472 280356
rect 99524 280344 99530 280356
rect 100386 280344 100392 280356
rect 99524 280316 100392 280344
rect 99524 280304 99530 280316
rect 100386 280304 100392 280316
rect 100444 280304 100450 280356
rect 183646 280304 183652 280356
rect 183704 280344 183710 280356
rect 222286 280344 222292 280356
rect 183704 280316 222292 280344
rect 183704 280304 183710 280316
rect 222286 280304 222292 280316
rect 222344 280304 222350 280356
rect 266998 280304 267004 280356
rect 267056 280344 267062 280356
rect 277946 280344 277952 280356
rect 267056 280316 277952 280344
rect 267056 280304 267062 280316
rect 277946 280304 277952 280316
rect 278004 280304 278010 280356
rect 295426 280304 295432 280356
rect 295484 280344 295490 280356
rect 334250 280344 334256 280356
rect 295484 280316 334256 280344
rect 295484 280304 295490 280316
rect 334250 280304 334256 280316
rect 334308 280304 334314 280356
rect 347038 280304 347044 280356
rect 347096 280344 347102 280356
rect 347096 280316 352512 280344
rect 347096 280304 347102 280316
rect 109954 280276 109960 280288
rect 74506 280248 109960 280276
rect 109954 280236 109960 280248
rect 110012 280236 110018 280288
rect 124858 280236 124864 280288
rect 124916 280276 124922 280288
rect 128630 280276 128636 280288
rect 124916 280248 128636 280276
rect 124916 280236 124922 280248
rect 128630 280236 128636 280248
rect 128688 280236 128694 280288
rect 151078 280236 151084 280288
rect 151136 280276 151142 280288
rect 156598 280276 156604 280288
rect 151136 280248 156604 280276
rect 151136 280236 151142 280248
rect 156598 280236 156604 280248
rect 156656 280236 156662 280288
rect 182818 280236 182824 280288
rect 182876 280276 182882 280288
rect 193950 280276 193956 280288
rect 182876 280248 193956 280276
rect 182876 280236 182882 280248
rect 193950 280236 193956 280248
rect 194008 280236 194014 280288
rect 232498 280236 232504 280288
rect 232556 280276 232562 280288
rect 232556 280248 248414 280276
rect 232556 280236 232562 280248
rect 82262 280208 82268 280220
rect 72804 280180 82268 280208
rect 82262 280168 82268 280180
rect 82320 280168 82326 280220
rect 93118 280168 93124 280220
rect 93176 280208 93182 280220
rect 100294 280208 100300 280220
rect 93176 280180 100300 280208
rect 93176 280168 93182 280180
rect 100294 280168 100300 280180
rect 100352 280168 100358 280220
rect 100386 280168 100392 280220
rect 100444 280208 100450 280220
rect 138290 280208 138296 280220
rect 100444 280180 138296 280208
rect 100444 280168 100450 280180
rect 138290 280168 138296 280180
rect 138348 280168 138354 280220
rect 149698 280168 149704 280220
rect 149756 280208 149762 280220
rect 166258 280208 166264 280220
rect 149756 280180 166264 280208
rect 149756 280168 149762 280180
rect 166258 280168 166264 280180
rect 166316 280168 166322 280220
rect 177298 280168 177304 280220
rect 177356 280208 177362 280220
rect 184290 280208 184296 280220
rect 177356 280180 184296 280208
rect 177356 280168 177362 280180
rect 184290 280168 184296 280180
rect 184348 280168 184354 280220
rect 233970 280168 233976 280220
rect 234028 280208 234034 280220
rect 240594 280208 240600 280220
rect 234028 280180 240600 280208
rect 234028 280168 234034 280180
rect 240594 280168 240600 280180
rect 240652 280168 240658 280220
rect 248386 280208 248414 280248
rect 267826 280236 267832 280288
rect 267884 280276 267890 280288
rect 306282 280276 306288 280288
rect 267884 280248 306288 280276
rect 267884 280236 267890 280248
rect 306282 280236 306288 280248
rect 306340 280236 306346 280288
rect 250254 280208 250260 280220
rect 248386 280180 250260 280208
rect 250254 280168 250260 280180
rect 250312 280168 250318 280220
rect 261478 280168 261484 280220
rect 261536 280208 261542 280220
rect 268286 280208 268292 280220
rect 261536 280180 268292 280208
rect 261536 280168 261542 280180
rect 268286 280168 268292 280180
rect 268344 280168 268350 280220
rect 289078 280168 289084 280220
rect 289136 280208 289142 280220
rect 296622 280208 296628 280220
rect 289136 280180 296628 280208
rect 289136 280168 289142 280180
rect 296622 280168 296628 280180
rect 296680 280168 296686 280220
rect 318058 280168 318064 280220
rect 318116 280208 318122 280220
rect 324590 280208 324596 280220
rect 318116 280180 324596 280208
rect 318116 280168 318122 280180
rect 324590 280168 324596 280180
rect 324648 280168 324654 280220
rect 348418 280168 348424 280220
rect 348476 280208 348482 280220
rect 352282 280208 352288 280220
rect 348476 280180 352288 280208
rect 348476 280168 348482 280180
rect 352282 280168 352288 280180
rect 352340 280168 352346 280220
rect 352484 280208 352512 280316
rect 354646 280276 354674 280384
rect 463786 280372 463792 280424
rect 463844 280412 463850 280424
rect 463844 280384 470594 280412
rect 463844 280372 463850 280384
rect 379606 280304 379612 280356
rect 379664 280344 379670 280356
rect 418246 280344 418252 280356
rect 379664 280316 418252 280344
rect 379664 280304 379670 280316
rect 418246 280304 418252 280316
rect 418304 280304 418310 280356
rect 390278 280276 390284 280288
rect 354646 280248 390284 280276
rect 390278 280236 390284 280248
rect 390336 280236 390342 280288
rect 400858 280236 400864 280288
rect 400916 280276 400922 280288
rect 408586 280276 408592 280288
rect 400916 280248 408592 280276
rect 400916 280236 400922 280248
rect 408586 280236 408592 280248
rect 408644 280236 408650 280288
rect 429838 280236 429844 280288
rect 429896 280276 429902 280288
rect 436278 280276 436284 280288
rect 429896 280248 436284 280276
rect 429896 280236 429902 280248
rect 436278 280236 436284 280248
rect 436336 280236 436342 280288
rect 457438 280236 457444 280288
rect 457496 280276 457502 280288
rect 464614 280276 464620 280288
rect 457496 280248 464620 280276
rect 457496 280236 457502 280248
rect 464614 280236 464620 280248
rect 464672 280236 464678 280288
rect 470566 280276 470594 280384
rect 491386 280304 491392 280356
rect 491444 280344 491450 280356
rect 529934 280344 529940 280356
rect 491444 280316 529940 280344
rect 491444 280304 491450 280316
rect 529934 280304 529940 280316
rect 529992 280304 529998 280356
rect 502242 280276 502248 280288
rect 470566 280248 502248 280276
rect 502242 280236 502248 280248
rect 502300 280236 502306 280288
rect 541618 280236 541624 280288
rect 541676 280276 541682 280288
rect 541676 280248 557534 280276
rect 541676 280236 541682 280248
rect 361942 280208 361948 280220
rect 352484 280180 361948 280208
rect 361942 280168 361948 280180
rect 362000 280168 362006 280220
rect 373258 280168 373264 280220
rect 373316 280208 373322 280220
rect 380618 280208 380624 280220
rect 373316 280180 380624 280208
rect 373316 280168 373322 280180
rect 380618 280168 380624 280180
rect 380676 280168 380682 280220
rect 428458 280168 428464 280220
rect 428516 280208 428522 280220
rect 445938 280208 445944 280220
rect 428516 280180 445944 280208
rect 428516 280168 428522 280180
rect 445938 280168 445944 280180
rect 445996 280168 446002 280220
rect 462958 280168 462964 280220
rect 463016 280208 463022 280220
rect 474274 280208 474280 280220
rect 463016 280180 474280 280208
rect 463016 280168 463022 280180
rect 474274 280168 474280 280180
rect 474332 280168 474338 280220
rect 485038 280168 485044 280220
rect 485096 280208 485102 280220
rect 492582 280208 492588 280220
rect 485096 280180 492588 280208
rect 485096 280168 485102 280180
rect 492582 280168 492588 280180
rect 492640 280168 492646 280220
rect 512638 280168 512644 280220
rect 512696 280208 512702 280220
rect 520274 280208 520280 280220
rect 512696 280180 520280 280208
rect 512696 280168 512702 280180
rect 520274 280168 520280 280180
rect 520332 280168 520338 280220
rect 544378 280168 544384 280220
rect 544436 280208 544442 280220
rect 548610 280208 548616 280220
rect 544436 280180 548616 280208
rect 544436 280168 544442 280180
rect 548610 280168 548616 280180
rect 548668 280168 548674 280220
rect 557506 280208 557534 280248
rect 558270 280208 558276 280220
rect 557506 280180 558276 280208
rect 558270 280168 558276 280180
rect 558328 280168 558334 280220
rect 568022 278400 568028 278452
rect 568080 278400 568086 278452
rect 120166 278264 120172 278316
rect 120224 278304 120230 278316
rect 122098 278304 122104 278316
rect 120224 278276 122104 278304
rect 120224 278264 120230 278276
rect 122098 278264 122104 278276
rect 122156 278264 122162 278316
rect 512086 278264 512092 278316
rect 512144 278304 512150 278316
rect 514018 278304 514024 278316
rect 512144 278276 514024 278304
rect 512144 278264 512150 278276
rect 514018 278264 514024 278276
rect 514076 278264 514082 278316
rect 568040 278248 568068 278400
rect 568022 278196 568028 278248
rect 568080 278196 568086 278248
rect 126882 277516 126888 277568
rect 126940 277556 126946 277568
rect 178034 277556 178040 277568
rect 126940 277528 178040 277556
rect 126940 277516 126946 277528
rect 178034 277516 178040 277528
rect 178092 277516 178098 277568
rect 182082 277516 182088 277568
rect 182140 277556 182146 277568
rect 233234 277556 233240 277568
rect 182140 277528 233240 277556
rect 182140 277516 182146 277528
rect 233234 277516 233240 277528
rect 233292 277516 233298 277568
rect 462222 277516 462228 277568
rect 462280 277556 462286 277568
rect 513374 277556 513380 277568
rect 462280 277528 513380 277556
rect 462280 277516 462286 277528
rect 513374 277516 513380 277528
rect 513432 277516 513438 277568
rect 42702 277448 42708 277500
rect 42760 277488 42766 277500
rect 93854 277488 93860 277500
rect 42760 277460 93860 277488
rect 42760 277448 42766 277460
rect 93854 277448 93860 277460
rect 93912 277448 93918 277500
rect 97902 277448 97908 277500
rect 97960 277488 97966 277500
rect 149054 277488 149060 277500
rect 97960 277460 149060 277488
rect 97960 277448 97966 277460
rect 149054 277448 149060 277460
rect 149112 277448 149118 277500
rect 154482 277448 154488 277500
rect 154540 277488 154546 277500
rect 205634 277488 205640 277500
rect 154540 277460 205640 277488
rect 154540 277448 154546 277460
rect 205634 277448 205640 277460
rect 205692 277448 205698 277500
rect 209682 277448 209688 277500
rect 209740 277488 209746 277500
rect 262214 277488 262220 277500
rect 209740 277460 262220 277488
rect 209740 277448 209746 277460
rect 262214 277448 262220 277460
rect 262272 277448 262278 277500
rect 266262 277448 266268 277500
rect 266320 277488 266326 277500
rect 317414 277488 317420 277500
rect 266320 277460 317420 277488
rect 266320 277448 266326 277460
rect 317414 277448 317420 277460
rect 317472 277448 317478 277500
rect 322842 277448 322848 277500
rect 322900 277488 322906 277500
rect 373994 277488 374000 277500
rect 322900 277460 374000 277488
rect 322900 277448 322906 277460
rect 373994 277448 374000 277460
rect 374052 277448 374058 277500
rect 378042 277448 378048 277500
rect 378100 277488 378106 277500
rect 429286 277488 429292 277500
rect 378100 277460 429292 277488
rect 378100 277448 378106 277460
rect 429286 277448 429292 277460
rect 429344 277448 429350 277500
rect 434622 277448 434628 277500
rect 434680 277488 434686 277500
rect 485774 277488 485780 277500
rect 434680 277460 485780 277488
rect 434680 277448 434686 277460
rect 485774 277448 485780 277460
rect 485832 277448 485838 277500
rect 518802 277448 518808 277500
rect 518860 277488 518866 277500
rect 569954 277488 569960 277500
rect 518860 277460 569960 277488
rect 518860 277448 518866 277460
rect 569954 277448 569960 277460
rect 570012 277448 570018 277500
rect 13538 277380 13544 277432
rect 13596 277420 13602 277432
rect 66254 277420 66260 277432
rect 13596 277392 66260 277420
rect 13596 277380 13602 277392
rect 66254 277380 66260 277392
rect 66312 277380 66318 277432
rect 70302 277380 70308 277432
rect 70360 277420 70366 277432
rect 121454 277420 121460 277432
rect 70360 277392 121460 277420
rect 70360 277380 70366 277392
rect 121454 277380 121460 277392
rect 121512 277380 121518 277432
rect 204070 277380 204076 277432
rect 204128 277420 204134 277432
rect 212442 277420 212448 277432
rect 204128 277392 212448 277420
rect 204128 277380 204134 277392
rect 212442 277380 212448 277392
rect 212500 277380 212506 277432
rect 238662 277380 238668 277432
rect 238720 277420 238726 277432
rect 289814 277420 289820 277432
rect 238720 277392 289820 277420
rect 238720 277380 238726 277392
rect 289814 277380 289820 277392
rect 289872 277380 289878 277432
rect 293862 277380 293868 277432
rect 293920 277420 293926 277432
rect 345014 277420 345020 277432
rect 293920 277392 345020 277420
rect 293920 277380 293926 277392
rect 345014 277380 345020 277392
rect 345072 277380 345078 277432
rect 350442 277380 350448 277432
rect 350500 277420 350506 277432
rect 401594 277420 401600 277432
rect 350500 277392 401600 277420
rect 350500 277380 350506 277392
rect 401594 277380 401600 277392
rect 401652 277380 401658 277432
rect 405642 277380 405648 277432
rect 405700 277420 405706 277432
rect 458174 277420 458180 277432
rect 405700 277392 458180 277420
rect 405700 277380 405706 277392
rect 458174 277380 458180 277392
rect 458232 277380 458238 277432
rect 489822 277380 489828 277432
rect 489880 277420 489886 277432
rect 542354 277420 542360 277432
rect 489880 277392 542360 277420
rect 489880 277380 489886 277392
rect 542354 277380 542360 277392
rect 542412 277380 542418 277432
rect 204254 272552 204260 272604
rect 204312 272592 204318 272604
rect 204990 272592 204996 272604
rect 204312 272564 204996 272592
rect 204312 272552 204318 272564
rect 204990 272552 204996 272564
rect 205048 272552 205054 272604
rect 400306 272552 400312 272604
rect 400364 272592 400370 272604
rect 400950 272592 400956 272604
rect 400364 272564 400956 272592
rect 400364 272552 400370 272564
rect 400950 272552 400956 272564
rect 401008 272552 401014 272604
rect 15194 256640 15200 256692
rect 15252 256680 15258 256692
rect 35894 256680 35900 256692
rect 15252 256652 35900 256680
rect 15252 256640 15258 256652
rect 35894 256640 35900 256652
rect 35952 256640 35958 256692
rect 36078 256640 36084 256692
rect 36136 256680 36142 256692
rect 63586 256680 63592 256692
rect 36136 256652 63592 256680
rect 36136 256640 36142 256652
rect 63586 256640 63592 256652
rect 63644 256640 63650 256692
rect 64046 256640 64052 256692
rect 64104 256680 64110 256692
rect 91922 256680 91928 256692
rect 64104 256652 91928 256680
rect 64104 256640 64110 256652
rect 91922 256640 91928 256652
rect 91980 256640 91986 256692
rect 92106 256640 92112 256692
rect 92164 256680 92170 256692
rect 119614 256680 119620 256692
rect 92164 256652 119620 256680
rect 92164 256640 92170 256652
rect 119614 256640 119620 256652
rect 119672 256640 119678 256692
rect 122098 256640 122104 256692
rect 122156 256680 122162 256692
rect 147950 256680 147956 256692
rect 122156 256652 147956 256680
rect 122156 256640 122162 256652
rect 147950 256640 147956 256652
rect 148008 256640 148014 256692
rect 148042 256640 148048 256692
rect 148100 256680 148106 256692
rect 175918 256680 175924 256692
rect 148100 256652 175924 256680
rect 148100 256640 148106 256652
rect 175918 256640 175924 256652
rect 175976 256640 175982 256692
rect 176102 256640 176108 256692
rect 176160 256680 176166 256692
rect 203610 256680 203616 256692
rect 176160 256652 203616 256680
rect 176160 256640 176166 256652
rect 203610 256640 203616 256652
rect 203668 256640 203674 256692
rect 204990 256640 204996 256692
rect 205048 256680 205054 256692
rect 231946 256680 231952 256692
rect 205048 256652 231952 256680
rect 205048 256640 205054 256652
rect 231946 256640 231952 256652
rect 232004 256640 232010 256692
rect 232038 256640 232044 256692
rect 232096 256680 232102 256692
rect 259914 256680 259920 256692
rect 232096 256652 259920 256680
rect 232096 256640 232102 256652
rect 259914 256640 259920 256652
rect 259972 256640 259978 256692
rect 260098 256640 260104 256692
rect 260156 256680 260162 256692
rect 287606 256680 287612 256692
rect 260156 256652 287612 256680
rect 260156 256640 260162 256652
rect 287606 256640 287612 256652
rect 287664 256640 287670 256692
rect 288066 256640 288072 256692
rect 288124 256680 288130 256692
rect 315942 256680 315948 256692
rect 288124 256652 315948 256680
rect 288124 256640 288130 256652
rect 315942 256640 315948 256652
rect 316000 256640 316006 256692
rect 316678 256640 316684 256692
rect 316736 256680 316742 256692
rect 343910 256680 343916 256692
rect 316736 256652 343916 256680
rect 316736 256640 316742 256652
rect 343910 256640 343916 256652
rect 343968 256640 343974 256692
rect 344094 256640 344100 256692
rect 344152 256680 344158 256692
rect 371602 256680 371608 256692
rect 344152 256652 371608 256680
rect 344152 256640 344158 256652
rect 371602 256640 371608 256652
rect 371660 256640 371666 256692
rect 372062 256640 372068 256692
rect 372120 256680 372126 256692
rect 399938 256680 399944 256692
rect 372120 256652 399944 256680
rect 372120 256640 372126 256652
rect 399938 256640 399944 256652
rect 399996 256640 400002 256692
rect 400950 256640 400956 256692
rect 401008 256680 401014 256692
rect 427906 256680 427912 256692
rect 401008 256652 427912 256680
rect 401008 256640 401014 256652
rect 427906 256640 427912 256652
rect 427964 256640 427970 256692
rect 428090 256640 428096 256692
rect 428148 256680 428154 256692
rect 455598 256680 455604 256692
rect 428148 256652 455604 256680
rect 428148 256640 428154 256652
rect 455598 256640 455604 256652
rect 455656 256640 455662 256692
rect 456058 256640 456064 256692
rect 456116 256680 456122 256692
rect 483934 256680 483940 256692
rect 456116 256652 483940 256680
rect 456116 256640 456122 256652
rect 483934 256640 483940 256652
rect 483992 256640 483998 256692
rect 484026 256640 484032 256692
rect 484084 256680 484090 256692
rect 511902 256680 511908 256692
rect 484084 256652 511908 256680
rect 484084 256640 484090 256652
rect 511902 256640 511908 256652
rect 511960 256640 511966 256692
rect 514018 256640 514024 256692
rect 514076 256680 514082 256692
rect 539594 256680 539600 256692
rect 514076 256652 539600 256680
rect 514076 256640 514082 256652
rect 539594 256640 539600 256652
rect 539652 256640 539658 256692
rect 540054 256640 540060 256692
rect 540112 256680 540118 256692
rect 567930 256680 567936 256692
rect 540112 256652 567936 256680
rect 540112 256640 540118 256652
rect 567930 256640 567936 256652
rect 567988 256640 567994 256692
rect 16574 256572 16580 256624
rect 16632 256612 16638 256624
rect 36630 256612 36636 256624
rect 16632 256584 36636 256612
rect 16632 256572 16638 256584
rect 36630 256572 36636 256584
rect 36688 256572 36694 256624
rect 44910 256572 44916 256624
rect 44968 256612 44974 256624
rect 71130 256612 71136 256624
rect 44968 256584 71136 256612
rect 44968 256572 44974 256584
rect 71130 256572 71136 256584
rect 71188 256572 71194 256624
rect 82262 256572 82268 256624
rect 82320 256612 82326 256624
rect 93118 256612 93124 256624
rect 82320 256584 93124 256612
rect 82320 256572 82326 256584
rect 93118 256572 93124 256584
rect 93176 256572 93182 256624
rect 110322 256572 110328 256624
rect 110380 256612 110386 256624
rect 124858 256612 124864 256624
rect 110380 256584 124864 256612
rect 110380 256572 110386 256584
rect 124858 256572 124864 256584
rect 124916 256572 124922 256624
rect 128630 256572 128636 256624
rect 128688 256612 128694 256624
rect 149698 256612 149704 256624
rect 128688 256584 149704 256612
rect 128688 256572 128694 256584
rect 149698 256572 149704 256584
rect 149756 256572 149762 256624
rect 156598 256572 156604 256624
rect 156656 256612 156662 256624
rect 182818 256612 182824 256624
rect 156656 256584 182824 256612
rect 156656 256572 156662 256584
rect 182818 256572 182824 256584
rect 182876 256572 182882 256624
rect 194502 256572 194508 256624
rect 194560 256612 194566 256624
rect 204070 256612 204076 256624
rect 194560 256584 204076 256612
rect 194560 256572 194566 256584
rect 204070 256572 204076 256584
rect 204128 256572 204134 256624
rect 212626 256572 212632 256624
rect 212684 256612 212690 256624
rect 232498 256612 232504 256624
rect 212684 256584 232504 256612
rect 212684 256572 212690 256584
rect 232498 256572 232504 256584
rect 232556 256572 232562 256624
rect 240594 256572 240600 256624
rect 240652 256612 240658 256624
rect 266998 256612 267004 256624
rect 240652 256584 267004 256612
rect 240652 256572 240658 256584
rect 266998 256572 267004 256584
rect 267056 256572 267062 256624
rect 278590 256572 278596 256624
rect 278648 256612 278654 256624
rect 289078 256612 289084 256624
rect 278648 256584 289084 256612
rect 278648 256572 278654 256584
rect 289078 256572 289084 256584
rect 289136 256572 289142 256624
rect 306282 256572 306288 256624
rect 306340 256612 306346 256624
rect 318058 256612 318064 256624
rect 306340 256584 318064 256612
rect 306340 256572 306346 256584
rect 318058 256572 318064 256584
rect 318116 256572 318122 256624
rect 324590 256572 324596 256624
rect 324648 256612 324654 256624
rect 347038 256612 347044 256624
rect 324648 256584 347044 256612
rect 324648 256572 324654 256584
rect 347038 256572 347044 256584
rect 347096 256572 347102 256624
rect 362586 256572 362592 256624
rect 362644 256612 362650 256624
rect 373258 256612 373264 256624
rect 362644 256584 373264 256612
rect 362644 256572 362650 256584
rect 373258 256572 373264 256584
rect 373316 256572 373322 256624
rect 390278 256572 390284 256624
rect 390336 256612 390342 256624
rect 400858 256612 400864 256624
rect 390336 256584 400864 256612
rect 390336 256572 390342 256584
rect 400858 256572 400864 256584
rect 400916 256572 400922 256624
rect 408586 256572 408592 256624
rect 408644 256612 408650 256624
rect 428458 256612 428464 256624
rect 408644 256584 428464 256612
rect 408644 256572 408650 256584
rect 428458 256572 428464 256584
rect 428516 256572 428522 256624
rect 436922 256572 436928 256624
rect 436980 256612 436986 256624
rect 462958 256612 462964 256624
rect 436980 256584 462964 256612
rect 436980 256572 436986 256584
rect 462958 256572 462964 256584
rect 463016 256572 463022 256624
rect 474274 256572 474280 256624
rect 474332 256612 474338 256624
rect 485038 256612 485044 256624
rect 474332 256584 485044 256612
rect 474332 256572 474338 256584
rect 485038 256572 485044 256584
rect 485096 256572 485102 256624
rect 502242 256572 502248 256624
rect 502300 256612 502306 256624
rect 512638 256612 512644 256624
rect 502300 256584 512644 256612
rect 502300 256572 502306 256584
rect 512638 256572 512644 256584
rect 512696 256572 512702 256624
rect 520918 256572 520924 256624
rect 520976 256612 520982 256624
rect 541618 256612 541624 256624
rect 520976 256584 541624 256612
rect 520976 256572 520982 256584
rect 541618 256572 541624 256584
rect 541676 256572 541682 256624
rect 26234 256504 26240 256556
rect 26292 256544 26298 256556
rect 39298 256544 39304 256556
rect 26292 256516 39304 256544
rect 26292 256504 26298 256516
rect 39298 256504 39304 256516
rect 39356 256504 39362 256556
rect 54570 256504 54576 256556
rect 54628 256544 54634 256556
rect 66898 256544 66904 256556
rect 54628 256516 66904 256544
rect 54628 256504 54634 256516
rect 66898 256504 66904 256516
rect 66956 256504 66962 256556
rect 138290 256504 138296 256556
rect 138348 256544 138354 256556
rect 151078 256544 151084 256556
rect 138348 256516 151084 256544
rect 138348 256504 138354 256516
rect 151078 256504 151084 256516
rect 151136 256504 151142 256556
rect 166258 256504 166264 256556
rect 166316 256544 166322 256556
rect 177298 256544 177304 256556
rect 166316 256516 177304 256544
rect 166316 256504 166322 256516
rect 177298 256504 177304 256516
rect 177356 256504 177362 256556
rect 222286 256504 222292 256556
rect 222344 256544 222350 256556
rect 233970 256544 233976 256556
rect 222344 256516 233976 256544
rect 222344 256504 222350 256516
rect 233970 256504 233976 256516
rect 234028 256504 234034 256556
rect 250254 256504 250260 256556
rect 250312 256544 250318 256556
rect 261478 256544 261484 256556
rect 250312 256516 261484 256544
rect 250312 256504 250318 256516
rect 261478 256504 261484 256516
rect 261536 256504 261542 256556
rect 334250 256504 334256 256556
rect 334308 256544 334314 256556
rect 348418 256544 348424 256556
rect 334308 256516 348424 256544
rect 334308 256504 334314 256516
rect 348418 256504 348424 256516
rect 348476 256504 348482 256556
rect 418246 256504 418252 256556
rect 418304 256544 418310 256556
rect 429838 256544 429844 256556
rect 418304 256516 429844 256544
rect 418304 256504 418310 256516
rect 429838 256504 429844 256516
rect 429896 256504 429902 256556
rect 446582 256504 446588 256556
rect 446640 256544 446646 256556
rect 457438 256544 457444 256556
rect 446640 256516 457444 256544
rect 446640 256504 446646 256516
rect 457438 256504 457444 256516
rect 457496 256504 457502 256556
rect 530578 256504 530584 256556
rect 530636 256544 530642 256556
rect 544378 256544 544384 256556
rect 530636 256516 544384 256544
rect 530636 256504 530642 256516
rect 544378 256504 544384 256516
rect 544436 256504 544442 256556
rect 558270 255960 558276 256012
rect 558328 256000 558334 256012
rect 567470 256000 567476 256012
rect 558328 255972 567476 256000
rect 558328 255960 558334 255972
rect 567470 255960 567476 255972
rect 567528 255960 567534 256012
rect 548334 254532 548340 254584
rect 548392 254572 548398 254584
rect 568114 254572 568120 254584
rect 548392 254544 568120 254572
rect 548392 254532 548398 254544
rect 568114 254532 568120 254544
rect 568172 254532 568178 254584
rect 212350 254124 212356 254176
rect 212408 254164 212414 254176
rect 232682 254164 232688 254176
rect 212408 254136 232688 254164
rect 212408 254124 212414 254136
rect 232682 254124 232688 254136
rect 232740 254124 232746 254176
rect 296346 254124 296352 254176
rect 296404 254164 296410 254176
rect 316770 254164 316776 254176
rect 296404 254136 316776 254164
rect 296404 254124 296410 254136
rect 316770 254124 316776 254136
rect 316828 254124 316834 254176
rect 408034 254124 408040 254176
rect 408092 254164 408098 254176
rect 428642 254164 428648 254176
rect 408092 254136 428648 254164
rect 408092 254124 408098 254136
rect 428642 254124 428648 254136
rect 428700 254124 428706 254176
rect 492030 254124 492036 254176
rect 492088 254164 492094 254176
rect 512730 254164 512736 254176
rect 492088 254136 512736 254164
rect 492088 254124 492094 254136
rect 512730 254124 512736 254136
rect 512788 254124 512794 254176
rect 2774 254056 2780 254108
rect 2832 254096 2838 254108
rect 5074 254096 5080 254108
rect 2832 254068 5080 254096
rect 2832 254056 2838 254068
rect 5074 254056 5080 254068
rect 5132 254056 5138 254108
rect 148410 254056 148416 254108
rect 148468 254096 148474 254108
rect 165706 254096 165712 254108
rect 148468 254068 165712 254096
rect 148468 254056 148474 254068
rect 165706 254056 165712 254068
rect 165764 254056 165770 254108
rect 175458 254056 175464 254108
rect 175516 254096 175522 254108
rect 193674 254096 193680 254108
rect 175516 254068 193680 254096
rect 175516 254056 175522 254068
rect 193674 254056 193680 254068
rect 193732 254056 193738 254108
rect 203518 254056 203524 254108
rect 203576 254096 203582 254108
rect 221366 254096 221372 254108
rect 203576 254068 221372 254096
rect 203576 254056 203582 254068
rect 221366 254056 221372 254068
rect 221424 254056 221430 254108
rect 260098 254056 260104 254108
rect 260156 254096 260162 254108
rect 277670 254096 277676 254108
rect 260156 254068 277676 254096
rect 260156 254056 260162 254068
rect 277670 254056 277676 254068
rect 277728 254056 277734 254108
rect 287514 254056 287520 254108
rect 287572 254096 287578 254108
rect 305362 254096 305368 254108
rect 287572 254068 305368 254096
rect 287572 254056 287578 254068
rect 305362 254056 305368 254068
rect 305420 254056 305426 254108
rect 345658 254056 345664 254108
rect 345716 254096 345722 254108
rect 361666 254096 361672 254108
rect 345716 254068 361672 254096
rect 345716 254056 345722 254068
rect 361666 254056 361672 254068
rect 361724 254056 361730 254108
rect 371510 254056 371516 254108
rect 371568 254096 371574 254108
rect 389358 254096 389364 254108
rect 371568 254068 389364 254096
rect 371568 254056 371574 254068
rect 389358 254056 389364 254068
rect 389416 254056 389422 254108
rect 399478 254056 399484 254108
rect 399536 254096 399542 254108
rect 417694 254096 417700 254108
rect 399536 254068 417700 254096
rect 399536 254056 399542 254068
rect 417694 254056 417700 254068
rect 417752 254056 417758 254108
rect 456058 254056 456064 254108
rect 456116 254096 456122 254108
rect 473354 254096 473360 254108
rect 456116 254068 473360 254096
rect 456116 254056 456122 254068
rect 473354 254056 473360 254068
rect 473412 254056 473418 254108
rect 483474 254056 483480 254108
rect 483532 254096 483538 254108
rect 501690 254096 501696 254108
rect 483532 254068 501696 254096
rect 483532 254056 483538 254068
rect 501690 254056 501696 254068
rect 501748 254056 501754 254108
rect 36722 253988 36728 254040
rect 36780 254028 36786 254040
rect 53650 254028 53656 254040
rect 36780 254000 53656 254028
rect 36780 253988 36786 254000
rect 53650 253988 53656 254000
rect 53708 253988 53714 254040
rect 64414 253988 64420 254040
rect 64472 254028 64478 254040
rect 81434 254028 81440 254040
rect 64472 254000 81440 254028
rect 64472 253988 64478 254000
rect 81434 253988 81440 254000
rect 81492 253988 81498 254040
rect 91462 253988 91468 254040
rect 91520 254028 91526 254040
rect 109678 254028 109684 254040
rect 91520 254000 109684 254028
rect 91520 253988 91526 254000
rect 109678 253988 109684 254000
rect 109736 253988 109742 254040
rect 119430 253988 119436 254040
rect 119488 254028 119494 254040
rect 137646 254028 137652 254040
rect 119488 254000 137652 254028
rect 119488 253988 119494 254000
rect 137646 253988 137652 254000
rect 137704 253988 137710 254040
rect 156322 253988 156328 254040
rect 156380 254028 156386 254040
rect 178678 254028 178684 254040
rect 156380 254000 178684 254028
rect 156380 253988 156386 254000
rect 178678 253988 178684 254000
rect 178736 253988 178742 254040
rect 232498 253988 232504 254040
rect 232556 254028 232562 254040
rect 249702 254028 249708 254040
rect 232556 254000 249708 254028
rect 232556 253988 232562 254000
rect 249702 253988 249708 254000
rect 249760 253988 249766 254040
rect 268010 253988 268016 254040
rect 268068 254028 268074 254040
rect 287698 254028 287704 254040
rect 268068 254000 287704 254028
rect 268068 253988 268074 254000
rect 287698 253988 287704 254000
rect 287756 253988 287762 254040
rect 315482 253988 315488 254040
rect 315540 254028 315546 254040
rect 333698 254028 333704 254040
rect 315540 254000 333704 254028
rect 315540 253988 315546 254000
rect 333698 253988 333704 254000
rect 333756 253988 333762 254040
rect 352006 253988 352012 254040
rect 352064 254028 352070 254040
rect 374638 254028 374644 254040
rect 352064 254000 374644 254028
rect 352064 253988 352070 254000
rect 374638 253988 374644 254000
rect 374696 253988 374702 254040
rect 428550 253988 428556 254040
rect 428608 254028 428614 254040
rect 445662 254028 445668 254040
rect 428608 254000 445668 254028
rect 428608 253988 428614 254000
rect 445662 253988 445668 254000
rect 445720 253988 445726 254040
rect 464338 253988 464344 254040
rect 464396 254028 464402 254040
rect 483658 254028 483664 254040
rect 464396 254000 483664 254028
rect 464396 253988 464402 254000
rect 483658 253988 483664 254000
rect 483716 253988 483722 254040
rect 511442 253988 511448 254040
rect 511500 254028 511506 254040
rect 529658 254028 529664 254040
rect 511500 254000 529664 254028
rect 511500 253988 511506 254000
rect 529658 253988 529664 254000
rect 529716 253988 529722 254040
rect 541618 253988 541624 254040
rect 541676 254028 541682 254040
rect 557534 254028 557540 254040
rect 541676 254000 557540 254028
rect 541676 253988 541682 254000
rect 557534 253988 557540 254000
rect 557592 253988 557598 254040
rect 15102 253920 15108 253972
rect 15160 253960 15166 253972
rect 25682 253960 25688 253972
rect 15160 253932 25688 253960
rect 15160 253920 15166 253932
rect 25682 253920 25688 253932
rect 25740 253920 25746 253972
rect 36630 253920 36636 253972
rect 36688 253960 36694 253972
rect 63310 253960 63316 253972
rect 36688 253932 63316 253960
rect 36688 253920 36694 253932
rect 63310 253920 63316 253932
rect 63368 253920 63374 253972
rect 66898 253920 66904 253972
rect 66956 253960 66962 253972
rect 91094 253960 91100 253972
rect 66956 253932 91100 253960
rect 66956 253920 66962 253932
rect 91094 253920 91100 253932
rect 91152 253920 91158 253972
rect 93118 253920 93124 253972
rect 93176 253960 93182 253972
rect 119338 253960 119344 253972
rect 93176 253932 119344 253960
rect 93176 253920 93182 253932
rect 119338 253920 119344 253932
rect 119396 253920 119402 253972
rect 122098 253920 122104 253972
rect 122156 253960 122162 253972
rect 147306 253960 147312 253972
rect 122156 253932 147312 253960
rect 122156 253920 122162 253932
rect 147306 253920 147312 253932
rect 147364 253920 147370 253972
rect 148318 253920 148324 253972
rect 148376 253960 148382 253972
rect 175366 253960 175372 253972
rect 148376 253932 175372 253960
rect 148376 253920 148382 253932
rect 175366 253920 175372 253932
rect 175424 253920 175430 253972
rect 177298 253920 177304 253972
rect 177356 253960 177362 253972
rect 203334 253960 203340 253972
rect 177356 253932 203340 253960
rect 177356 253920 177362 253932
rect 203334 253920 203340 253932
rect 203392 253920 203398 253972
rect 204990 253920 204996 253972
rect 205048 253960 205054 253972
rect 231026 253960 231032 253972
rect 205048 253932 231032 253960
rect 205048 253920 205054 253932
rect 231026 253920 231032 253932
rect 231084 253920 231090 253972
rect 232590 253920 232596 253972
rect 232648 253960 232654 253972
rect 259362 253960 259368 253972
rect 232648 253932 259368 253960
rect 232648 253920 232654 253932
rect 259362 253920 259368 253932
rect 259420 253920 259426 253972
rect 260190 253920 260196 253972
rect 260248 253960 260254 253972
rect 287330 253960 287336 253972
rect 260248 253932 287336 253960
rect 260248 253920 260254 253932
rect 287330 253920 287336 253932
rect 287388 253920 287394 253972
rect 289078 253920 289084 253972
rect 289136 253960 289142 253972
rect 315022 253960 315028 253972
rect 289136 253932 315028 253960
rect 289136 253920 289142 253932
rect 315022 253920 315028 253932
rect 315080 253920 315086 253972
rect 316678 253920 316684 253972
rect 316736 253960 316742 253972
rect 343358 253960 343364 253972
rect 316736 253932 343364 253960
rect 316736 253920 316742 253932
rect 343358 253920 343364 253932
rect 343416 253920 343422 253972
rect 344278 253920 344284 253972
rect 344336 253960 344342 253972
rect 371326 253960 371332 253972
rect 344336 253932 371332 253960
rect 344336 253920 344342 253932
rect 371326 253920 371332 253932
rect 371384 253920 371390 253972
rect 373258 253920 373264 253972
rect 373316 253960 373322 253972
rect 399018 253960 399024 253972
rect 373316 253932 399024 253960
rect 373316 253920 373322 253932
rect 399018 253920 399024 253932
rect 399076 253920 399082 253972
rect 400858 253920 400864 253972
rect 400916 253960 400922 253972
rect 427354 253960 427360 253972
rect 400916 253932 427360 253960
rect 400916 253920 400922 253932
rect 427354 253920 427360 253932
rect 427412 253920 427418 253972
rect 428458 253920 428464 253972
rect 428516 253960 428522 253972
rect 455322 253960 455328 253972
rect 428516 253932 455328 253960
rect 428516 253920 428522 253932
rect 455322 253920 455328 253932
rect 455380 253920 455386 253972
rect 456150 253920 456156 253972
rect 456208 253960 456214 253972
rect 483014 253960 483020 253972
rect 456208 253932 483020 253960
rect 456208 253920 456214 253932
rect 483014 253920 483020 253932
rect 483072 253920 483078 253972
rect 485038 253920 485044 253972
rect 485096 253960 485102 253972
rect 511350 253960 511356 253972
rect 485096 253932 511356 253960
rect 485096 253920 485102 253932
rect 511350 253920 511356 253932
rect 511408 253920 511414 253972
rect 512638 253920 512644 253972
rect 512696 253960 512702 253972
rect 539318 253960 539324 253972
rect 512696 253932 539324 253960
rect 512696 253920 512702 253932
rect 539318 253920 539324 253932
rect 539376 253920 539382 253972
rect 540238 253920 540244 253972
rect 540296 253960 540302 253972
rect 567194 253960 567200 253972
rect 540296 253932 567200 253960
rect 540296 253920 540302 253932
rect 567194 253920 567200 253932
rect 567252 253920 567258 253972
rect 350442 251336 350448 251388
rect 350500 251376 350506 251388
rect 401594 251376 401600 251388
rect 350500 251348 401600 251376
rect 350500 251336 350506 251348
rect 401594 251336 401600 251348
rect 401652 251336 401658 251388
rect 462222 251336 462228 251388
rect 462280 251376 462286 251388
rect 513374 251376 513380 251388
rect 462280 251348 513380 251376
rect 462280 251336 462286 251348
rect 513374 251336 513380 251348
rect 513432 251336 513438 251388
rect 42702 251268 42708 251320
rect 42760 251308 42766 251320
rect 42760 251280 45554 251308
rect 42760 251268 42766 251280
rect 45526 251240 45554 251280
rect 126882 251268 126888 251320
rect 126940 251308 126946 251320
rect 178034 251308 178040 251320
rect 126940 251280 178040 251308
rect 126940 251268 126946 251280
rect 178034 251268 178040 251280
rect 178092 251268 178098 251320
rect 182082 251268 182088 251320
rect 182140 251308 182146 251320
rect 233234 251308 233240 251320
rect 182140 251280 233240 251308
rect 182140 251268 182146 251280
rect 233234 251268 233240 251280
rect 233292 251268 233298 251320
rect 238662 251268 238668 251320
rect 238720 251308 238726 251320
rect 289814 251308 289820 251320
rect 238720 251280 289820 251308
rect 238720 251268 238726 251280
rect 289814 251268 289820 251280
rect 289872 251268 289878 251320
rect 293862 251268 293868 251320
rect 293920 251308 293926 251320
rect 345014 251308 345020 251320
rect 293920 251280 345020 251308
rect 293920 251268 293926 251280
rect 345014 251268 345020 251280
rect 345072 251268 345078 251320
rect 378042 251268 378048 251320
rect 378100 251308 378106 251320
rect 429286 251308 429292 251320
rect 378100 251280 429292 251308
rect 378100 251268 378106 251280
rect 429286 251268 429292 251280
rect 429344 251268 429350 251320
rect 434622 251268 434628 251320
rect 434680 251308 434686 251320
rect 485774 251308 485780 251320
rect 434680 251280 485780 251308
rect 434680 251268 434686 251280
rect 485774 251268 485780 251280
rect 485832 251268 485838 251320
rect 518802 251268 518808 251320
rect 518860 251308 518866 251320
rect 569954 251308 569960 251320
rect 518860 251280 569960 251308
rect 518860 251268 518866 251280
rect 569954 251268 569960 251280
rect 570012 251268 570018 251320
rect 93854 251240 93860 251252
rect 45526 251212 93860 251240
rect 93854 251200 93860 251212
rect 93912 251200 93918 251252
rect 97902 251200 97908 251252
rect 97960 251240 97966 251252
rect 149054 251240 149060 251252
rect 97960 251212 149060 251240
rect 97960 251200 97966 251212
rect 149054 251200 149060 251212
rect 149112 251200 149118 251252
rect 154482 251200 154488 251252
rect 154540 251240 154546 251252
rect 205634 251240 205640 251252
rect 154540 251212 205640 251240
rect 154540 251200 154546 251212
rect 205634 251200 205640 251212
rect 205692 251200 205698 251252
rect 209682 251200 209688 251252
rect 209740 251240 209746 251252
rect 262214 251240 262220 251252
rect 209740 251212 262220 251240
rect 209740 251200 209746 251212
rect 262214 251200 262220 251212
rect 262272 251200 262278 251252
rect 266262 251200 266268 251252
rect 266320 251240 266326 251252
rect 317414 251240 317420 251252
rect 266320 251212 317420 251240
rect 266320 251200 266326 251212
rect 317414 251200 317420 251212
rect 317472 251200 317478 251252
rect 322842 251200 322848 251252
rect 322900 251240 322906 251252
rect 373994 251240 374000 251252
rect 322900 251212 374000 251240
rect 322900 251200 322906 251212
rect 373994 251200 374000 251212
rect 374052 251200 374058 251252
rect 405642 251200 405648 251252
rect 405700 251240 405706 251252
rect 458174 251240 458180 251252
rect 405700 251212 458180 251240
rect 405700 251200 405706 251212
rect 458174 251200 458180 251212
rect 458232 251200 458238 251252
rect 489822 251200 489828 251252
rect 489880 251240 489886 251252
rect 542354 251240 542360 251252
rect 489880 251212 542360 251240
rect 489880 251200 489886 251212
rect 542354 251200 542360 251212
rect 542412 251200 542418 251252
rect 42886 249772 42892 249824
rect 42944 249812 42950 249824
rect 43622 249812 43628 249824
rect 42944 249784 43628 249812
rect 42944 249772 42950 249784
rect 43622 249772 43628 249784
rect 43680 249772 43686 249824
rect 2774 240184 2780 240236
rect 2832 240224 2838 240236
rect 5166 240224 5172 240236
rect 2832 240196 5172 240224
rect 2832 240184 2838 240196
rect 5166 240184 5172 240196
rect 5224 240184 5230 240236
rect 63586 235356 63592 235408
rect 63644 235396 63650 235408
rect 64414 235396 64420 235408
rect 63644 235368 64420 235396
rect 63644 235356 63650 235368
rect 64414 235356 64420 235368
rect 64472 235356 64478 235408
rect 147674 235356 147680 235408
rect 147732 235396 147738 235408
rect 148410 235396 148416 235408
rect 147732 235368 148416 235396
rect 147732 235356 147738 235368
rect 148410 235356 148416 235368
rect 148468 235356 148474 235408
rect 512730 234200 512736 234252
rect 512788 234240 512794 234252
rect 519630 234240 519636 234252
rect 512788 234212 519636 234240
rect 512788 234200 512794 234212
rect 519630 234200 519636 234212
rect 519688 234200 519694 234252
rect 428642 233860 428648 233912
rect 428700 233900 428706 233912
rect 435726 233900 435732 233912
rect 428700 233872 435732 233900
rect 428700 233860 428706 233872
rect 435726 233860 435732 233872
rect 435784 233860 435790 233912
rect 232682 233520 232688 233572
rect 232740 233560 232746 233572
rect 239766 233560 239772 233572
rect 232740 233532 239772 233560
rect 232740 233520 232746 233532
rect 239766 233520 239772 233532
rect 239824 233520 239830 233572
rect 287698 233520 287704 233572
rect 287756 233560 287762 233572
rect 295702 233560 295708 233572
rect 287756 233532 295708 233560
rect 287756 233520 287762 233532
rect 295702 233520 295708 233532
rect 295760 233520 295766 233572
rect 316770 233384 316776 233436
rect 316828 233424 316834 233436
rect 323670 233424 323676 233436
rect 316828 233396 323676 233424
rect 316828 233384 316834 233396
rect 323670 233384 323676 233396
rect 323728 233384 323734 233436
rect 483658 233384 483664 233436
rect 483716 233424 483722 233436
rect 491662 233424 491668 233436
rect 483716 233396 491668 233424
rect 483716 233384 483722 233396
rect 491662 233384 491668 233396
rect 491720 233384 491726 233436
rect 13538 233180 13544 233232
rect 13596 233220 13602 233232
rect 66254 233220 66260 233232
rect 13596 233192 66260 233220
rect 13596 233180 13602 233192
rect 66254 233180 66260 233192
rect 66312 233180 66318 233232
rect 70302 233180 70308 233232
rect 70360 233220 70366 233232
rect 121454 233220 121460 233232
rect 70360 233192 121460 233220
rect 70360 233180 70366 233192
rect 121454 233180 121460 233192
rect 121512 233180 121518 233232
rect 427722 233180 427728 233232
rect 427780 233220 427786 233232
rect 428550 233220 428556 233232
rect 427780 233192 428556 233220
rect 427780 233180 427786 233192
rect 428550 233180 428556 233192
rect 428608 233180 428614 233232
rect 539502 233180 539508 233232
rect 539560 233220 539566 233232
rect 541618 233220 541624 233232
rect 539560 233192 541624 233220
rect 539560 233180 539566 233192
rect 541618 233180 541624 233192
rect 541676 233180 541682 233232
rect 15102 232704 15108 232756
rect 15160 232744 15166 232756
rect 16574 232744 16580 232756
rect 15160 232716 16580 232744
rect 15160 232704 15166 232716
rect 16574 232704 16580 232716
rect 16632 232704 16638 232756
rect 343634 232704 343640 232756
rect 343692 232744 343698 232756
rect 345658 232744 345664 232756
rect 343692 232716 345664 232744
rect 343692 232704 343698 232716
rect 345658 232704 345664 232716
rect 345716 232704 345722 232756
rect 547874 232704 547880 232756
rect 547932 232744 547938 232756
rect 548150 232744 548156 232756
rect 547932 232716 548156 232744
rect 547932 232704 547938 232716
rect 548150 232704 548156 232716
rect 548208 232704 548214 232756
rect 35342 231888 35348 231940
rect 35400 231928 35406 231940
rect 36722 231928 36728 231940
rect 35400 231900 36728 231928
rect 35400 231888 35406 231900
rect 36722 231888 36728 231900
rect 36780 231888 36786 231940
rect 149698 231820 149704 231872
rect 149756 231860 149762 231872
rect 579798 231860 579804 231872
rect 149756 231832 579804 231860
rect 149756 231820 149762 231832
rect 579798 231820 579804 231832
rect 579856 231820 579862 231872
rect 71866 230392 71872 230444
rect 71924 230432 71930 230444
rect 100018 230432 100024 230444
rect 71924 230404 100024 230432
rect 71924 230392 71930 230404
rect 100018 230392 100024 230404
rect 100076 230392 100082 230444
rect 127986 230432 127992 230444
rect 103486 230404 127992 230432
rect 25682 230324 25688 230376
rect 25740 230364 25746 230376
rect 36630 230364 36636 230376
rect 25740 230336 36636 230364
rect 25740 230324 25746 230336
rect 36630 230324 36636 230336
rect 36688 230324 36694 230376
rect 42886 230324 42892 230376
rect 42944 230364 42950 230376
rect 42944 230336 45554 230364
rect 42944 230324 42950 230336
rect 15286 230256 15292 230308
rect 15344 230296 15350 230308
rect 43990 230296 43996 230308
rect 15344 230268 43996 230296
rect 15344 230256 15350 230268
rect 43990 230256 43996 230268
rect 44048 230256 44054 230308
rect 45526 230296 45554 230336
rect 53650 230324 53656 230376
rect 53708 230364 53714 230376
rect 66898 230364 66904 230376
rect 53708 230336 66904 230364
rect 53708 230324 53714 230336
rect 66898 230324 66904 230336
rect 66956 230324 66962 230376
rect 81986 230324 81992 230376
rect 82044 230364 82050 230376
rect 93118 230364 93124 230376
rect 82044 230336 93124 230364
rect 82044 230324 82050 230336
rect 93118 230324 93124 230336
rect 93176 230324 93182 230376
rect 99466 230324 99472 230376
rect 99524 230364 99530 230376
rect 103486 230364 103514 230404
rect 127986 230392 127992 230404
rect 128044 230392 128050 230444
rect 165982 230392 165988 230444
rect 166040 230432 166046 230444
rect 177298 230432 177304 230444
rect 166040 230404 177304 230432
rect 166040 230392 166046 230404
rect 177298 230392 177304 230404
rect 177356 230392 177362 230444
rect 178678 230392 178684 230444
rect 178736 230432 178742 230444
rect 184014 230432 184020 230444
rect 178736 230404 184020 230432
rect 178736 230392 178742 230404
rect 184014 230392 184020 230404
rect 184072 230392 184078 230444
rect 211706 230432 211712 230444
rect 190426 230404 211712 230432
rect 99524 230336 103514 230364
rect 99524 230324 99530 230336
rect 109678 230324 109684 230376
rect 109736 230364 109742 230376
rect 122098 230364 122104 230376
rect 109736 230336 122104 230364
rect 109736 230324 109742 230336
rect 122098 230324 122104 230336
rect 122156 230324 122162 230376
rect 137646 230324 137652 230376
rect 137704 230364 137710 230376
rect 148318 230364 148324 230376
rect 137704 230336 148324 230364
rect 137704 230324 137710 230336
rect 148318 230324 148324 230336
rect 148376 230324 148382 230376
rect 183646 230324 183652 230376
rect 183704 230364 183710 230376
rect 190426 230364 190454 230404
rect 211706 230392 211712 230404
rect 211764 230392 211770 230444
rect 277670 230392 277676 230444
rect 277728 230432 277734 230444
rect 289078 230432 289084 230444
rect 277728 230404 289084 230432
rect 277728 230392 277734 230404
rect 289078 230392 289084 230404
rect 289136 230392 289142 230444
rect 306006 230392 306012 230444
rect 306064 230432 306070 230444
rect 316678 230432 316684 230444
rect 306064 230404 316684 230432
rect 306064 230392 306070 230404
rect 316678 230392 316684 230404
rect 316736 230392 316742 230444
rect 361666 230392 361672 230444
rect 361724 230432 361730 230444
rect 373258 230432 373264 230444
rect 361724 230404 373264 230432
rect 361724 230392 361730 230404
rect 373258 230392 373264 230404
rect 373316 230392 373322 230444
rect 379606 230392 379612 230444
rect 379664 230432 379670 230444
rect 408034 230432 408040 230444
rect 379664 230404 408040 230432
rect 379664 230392 379670 230404
rect 408034 230392 408040 230404
rect 408092 230392 408098 230444
rect 473998 230392 474004 230444
rect 474056 230432 474062 230444
rect 485038 230432 485044 230444
rect 474056 230404 485044 230432
rect 474056 230392 474062 230404
rect 485038 230392 485044 230404
rect 485096 230392 485102 230444
rect 501690 230392 501696 230444
rect 501748 230432 501754 230444
rect 512638 230432 512644 230444
rect 501748 230404 512644 230432
rect 501748 230392 501754 230404
rect 512638 230392 512644 230404
rect 512696 230392 512702 230444
rect 548150 230392 548156 230444
rect 548208 230432 548214 230444
rect 557534 230432 557540 230444
rect 548208 230404 557540 230432
rect 548208 230392 548214 230404
rect 557534 230392 557540 230404
rect 557592 230392 557598 230444
rect 183704 230336 190454 230364
rect 183704 230324 183710 230336
rect 193674 230324 193680 230376
rect 193732 230364 193738 230376
rect 204990 230364 204996 230376
rect 193732 230336 204996 230364
rect 193732 230324 193738 230336
rect 204990 230324 204996 230336
rect 205048 230324 205054 230376
rect 222010 230324 222016 230376
rect 222068 230364 222074 230376
rect 232590 230364 232596 230376
rect 222068 230336 232596 230364
rect 222068 230324 222074 230336
rect 232590 230324 232596 230336
rect 232648 230324 232654 230376
rect 249702 230324 249708 230376
rect 249760 230364 249766 230376
rect 260190 230364 260196 230376
rect 249760 230336 260196 230364
rect 249760 230324 249766 230336
rect 260190 230324 260196 230336
rect 260248 230324 260254 230376
rect 333698 230324 333704 230376
rect 333756 230364 333762 230376
rect 344278 230364 344284 230376
rect 333756 230336 344284 230364
rect 333756 230324 333762 230336
rect 344278 230324 344284 230336
rect 344336 230324 344342 230376
rect 374638 230324 374644 230376
rect 374696 230364 374702 230376
rect 379698 230364 379704 230376
rect 374696 230336 379704 230364
rect 374696 230324 374702 230336
rect 379698 230324 379704 230336
rect 379756 230324 379762 230376
rect 390002 230324 390008 230376
rect 390060 230364 390066 230376
rect 400858 230364 400864 230376
rect 390060 230336 400864 230364
rect 390060 230324 390066 230336
rect 400858 230324 400864 230336
rect 400916 230324 400922 230376
rect 417694 230324 417700 230376
rect 417752 230364 417758 230376
rect 428458 230364 428464 230376
rect 417752 230336 428464 230364
rect 417752 230324 417758 230336
rect 428458 230324 428464 230336
rect 428516 230324 428522 230376
rect 445662 230324 445668 230376
rect 445720 230364 445726 230376
rect 456150 230364 456156 230376
rect 445720 230336 456156 230364
rect 445720 230324 445726 230336
rect 456150 230324 456156 230336
rect 456208 230324 456214 230376
rect 529658 230324 529664 230376
rect 529716 230364 529722 230376
rect 540238 230364 540244 230376
rect 529716 230336 540244 230364
rect 529716 230324 529722 230336
rect 540238 230324 540244 230336
rect 540296 230324 540302 230376
rect 72050 230296 72056 230308
rect 45526 230268 72056 230296
rect 72050 230256 72056 230268
rect 72108 230256 72114 230308
rect 127066 230256 127072 230308
rect 127124 230296 127130 230308
rect 156046 230296 156052 230308
rect 127124 230268 156052 230296
rect 127124 230256 127130 230268
rect 156046 230256 156052 230268
rect 156104 230256 156110 230308
rect 238846 230256 238852 230308
rect 238904 230296 238910 230308
rect 268010 230296 268016 230308
rect 238904 230268 268016 230296
rect 238904 230256 238910 230268
rect 268010 230256 268016 230268
rect 268068 230256 268074 230308
rect 323026 230256 323032 230308
rect 323084 230296 323090 230308
rect 352006 230296 352012 230308
rect 323084 230268 352012 230296
rect 323084 230256 323090 230268
rect 352006 230256 352012 230268
rect 352064 230256 352070 230308
rect 434806 230256 434812 230308
rect 434864 230296 434870 230308
rect 463694 230296 463700 230308
rect 434864 230268 463700 230296
rect 434864 230256 434870 230268
rect 463694 230256 463700 230268
rect 463752 230256 463758 230308
rect 518986 230256 518992 230308
rect 519044 230296 519050 230308
rect 547874 230296 547880 230308
rect 519044 230268 547880 230296
rect 519044 230256 519050 230268
rect 547874 230256 547880 230268
rect 547932 230256 547938 230308
rect 26234 226448 26240 226500
rect 26292 226488 26298 226500
rect 35434 226488 35440 226500
rect 26292 226460 35440 226488
rect 26292 226448 26298 226460
rect 35434 226448 35440 226460
rect 35492 226448 35498 226500
rect 71130 226448 71136 226500
rect 71188 226488 71194 226500
rect 82262 226488 82268 226500
rect 71188 226460 82268 226488
rect 71188 226448 71194 226460
rect 82262 226448 82268 226460
rect 82320 226448 82326 226500
rect 184198 226448 184204 226500
rect 184256 226488 184262 226500
rect 222286 226488 222292 226500
rect 184256 226460 222292 226488
rect 184256 226448 184262 226460
rect 222286 226448 222292 226460
rect 222344 226448 222350 226500
rect 261478 226448 261484 226500
rect 261536 226488 261542 226500
rect 268286 226488 268292 226500
rect 261536 226460 268292 226488
rect 261536 226448 261542 226460
rect 268286 226448 268292 226460
rect 268344 226448 268350 226500
rect 296162 226448 296168 226500
rect 296220 226488 296226 226500
rect 334250 226488 334256 226500
rect 296220 226460 334256 226488
rect 296220 226448 296226 226460
rect 334250 226448 334256 226460
rect 334308 226448 334314 226500
rect 352190 226448 352196 226500
rect 352248 226488 352254 226500
rect 352248 226460 364334 226488
rect 352248 226448 352254 226460
rect 36630 226380 36636 226432
rect 36688 226420 36694 226432
rect 53926 226420 53932 226432
rect 36688 226392 53932 226420
rect 36688 226380 36694 226392
rect 53926 226380 53932 226392
rect 53984 226380 53990 226432
rect 72234 226380 72240 226432
rect 72292 226420 72298 226432
rect 109954 226420 109960 226432
rect 72292 226392 109960 226420
rect 72292 226380 72298 226392
rect 109954 226380 109960 226392
rect 110012 226380 110018 226432
rect 124858 226380 124864 226432
rect 124916 226420 124922 226432
rect 128630 226420 128636 226432
rect 124916 226392 128636 226420
rect 124916 226380 124922 226392
rect 128630 226380 128636 226392
rect 128688 226380 128694 226432
rect 152458 226380 152464 226432
rect 152516 226420 152522 226432
rect 156598 226420 156604 226432
rect 152516 226392 156604 226420
rect 152516 226380 152522 226392
rect 156598 226380 156604 226392
rect 156656 226380 156662 226432
rect 182818 226380 182824 226432
rect 182876 226420 182882 226432
rect 193950 226420 193956 226432
rect 182876 226392 193956 226420
rect 182876 226380 182882 226392
rect 193950 226380 193956 226392
rect 194008 226380 194014 226432
rect 232498 226380 232504 226432
rect 232556 226420 232562 226432
rect 232556 226392 248414 226420
rect 232556 226380 232562 226392
rect 39298 226312 39304 226364
rect 39356 226352 39362 226364
rect 44266 226352 44272 226364
rect 39356 226324 44272 226352
rect 39356 226312 39362 226324
rect 44266 226312 44272 226324
rect 44324 226312 44330 226364
rect 66898 226312 66904 226364
rect 66956 226352 66962 226364
rect 72602 226352 72608 226364
rect 66956 226324 72608 226352
rect 66956 226312 66962 226324
rect 72602 226312 72608 226324
rect 72660 226312 72666 226364
rect 93118 226312 93124 226364
rect 93176 226352 93182 226364
rect 100294 226352 100300 226364
rect 93176 226324 100300 226352
rect 93176 226312 93182 226324
rect 100294 226312 100300 226324
rect 100352 226312 100358 226364
rect 138290 226352 138296 226364
rect 100404 226324 138296 226352
rect 100202 226244 100208 226296
rect 100260 226284 100266 226296
rect 100404 226284 100432 226324
rect 138290 226312 138296 226324
rect 138348 226312 138354 226364
rect 151078 226312 151084 226364
rect 151136 226352 151142 226364
rect 166258 226352 166264 226364
rect 151136 226324 166264 226352
rect 151136 226312 151142 226324
rect 166258 226312 166264 226324
rect 166316 226312 166322 226364
rect 177298 226312 177304 226364
rect 177356 226352 177362 226364
rect 184290 226352 184296 226364
rect 177356 226324 184296 226352
rect 177356 226312 177362 226324
rect 184290 226312 184296 226324
rect 184348 226312 184354 226364
rect 233970 226312 233976 226364
rect 234028 226352 234034 226364
rect 240594 226352 240600 226364
rect 234028 226324 240600 226352
rect 234028 226312 234034 226324
rect 240594 226312 240600 226324
rect 240652 226312 240658 226364
rect 248386 226352 248414 226392
rect 268194 226380 268200 226432
rect 268252 226420 268258 226432
rect 306282 226420 306288 226432
rect 268252 226392 306288 226420
rect 268252 226380 268258 226392
rect 306282 226380 306288 226392
rect 306340 226380 306346 226432
rect 347038 226380 347044 226432
rect 347096 226420 347102 226432
rect 361942 226420 361948 226432
rect 347096 226392 361948 226420
rect 347096 226380 347102 226392
rect 361942 226380 361948 226392
rect 362000 226380 362006 226432
rect 364306 226420 364334 226460
rect 380250 226448 380256 226500
rect 380308 226488 380314 226500
rect 418246 226488 418252 226500
rect 380308 226460 418252 226488
rect 380308 226448 380314 226460
rect 418246 226448 418252 226460
rect 418304 226448 418310 226500
rect 462958 226448 462964 226500
rect 463016 226488 463022 226500
rect 474274 226488 474280 226500
rect 463016 226460 474280 226488
rect 463016 226448 463022 226460
rect 474274 226448 474280 226460
rect 474332 226448 474338 226500
rect 492122 226448 492128 226500
rect 492180 226488 492186 226500
rect 529934 226488 529940 226500
rect 492180 226460 529940 226488
rect 492180 226448 492186 226460
rect 529934 226448 529940 226460
rect 529992 226448 529998 226500
rect 390278 226420 390284 226432
rect 364306 226392 390284 226420
rect 390278 226380 390284 226392
rect 390336 226380 390342 226432
rect 400950 226380 400956 226432
rect 401008 226420 401014 226432
rect 408586 226420 408592 226432
rect 401008 226392 408592 226420
rect 401008 226380 401014 226392
rect 408586 226380 408592 226392
rect 408644 226380 408650 226432
rect 429838 226380 429844 226432
rect 429896 226420 429902 226432
rect 436278 226420 436284 226432
rect 429896 226392 436284 226420
rect 429896 226380 429902 226392
rect 436278 226380 436284 226392
rect 436336 226380 436342 226432
rect 464154 226380 464160 226432
rect 464212 226420 464218 226432
rect 502242 226420 502248 226432
rect 464212 226392 502248 226420
rect 464212 226380 464218 226392
rect 502242 226380 502248 226392
rect 502300 226380 502306 226432
rect 512638 226380 512644 226432
rect 512696 226420 512702 226432
rect 520274 226420 520280 226432
rect 512696 226392 520280 226420
rect 512696 226380 512702 226392
rect 520274 226380 520280 226392
rect 520332 226380 520338 226432
rect 541618 226380 541624 226432
rect 541676 226420 541682 226432
rect 541676 226392 557534 226420
rect 541676 226380 541682 226392
rect 250254 226352 250260 226364
rect 248386 226324 250260 226352
rect 250254 226312 250260 226324
rect 250312 226312 250318 226364
rect 266998 226312 267004 226364
rect 267056 226352 267062 226364
rect 277946 226352 277952 226364
rect 267056 226324 277952 226352
rect 267056 226312 267062 226324
rect 277946 226312 277952 226324
rect 278004 226312 278010 226364
rect 289078 226312 289084 226364
rect 289136 226352 289142 226364
rect 296622 226352 296628 226364
rect 289136 226324 296628 226352
rect 289136 226312 289142 226324
rect 296622 226312 296628 226324
rect 296680 226312 296686 226364
rect 318058 226312 318064 226364
rect 318116 226352 318122 226364
rect 324590 226352 324596 226364
rect 318116 226324 324596 226352
rect 318116 226312 318122 226324
rect 324590 226312 324596 226324
rect 324648 226312 324654 226364
rect 348418 226312 348424 226364
rect 348476 226352 348482 226364
rect 352282 226352 352288 226364
rect 348476 226324 352288 226352
rect 348476 226312 348482 226324
rect 352282 226312 352288 226324
rect 352340 226312 352346 226364
rect 373258 226312 373264 226364
rect 373316 226352 373322 226364
rect 380618 226352 380624 226364
rect 373316 226324 380624 226352
rect 373316 226312 373322 226324
rect 380618 226312 380624 226324
rect 380676 226312 380682 226364
rect 428458 226312 428464 226364
rect 428516 226352 428522 226364
rect 445938 226352 445944 226364
rect 428516 226324 445944 226352
rect 428516 226312 428522 226324
rect 445938 226312 445944 226324
rect 445996 226312 446002 226364
rect 457438 226312 457444 226364
rect 457496 226352 457502 226364
rect 464614 226352 464620 226364
rect 457496 226324 464620 226352
rect 457496 226312 457502 226324
rect 464614 226312 464620 226324
rect 464672 226312 464678 226364
rect 485038 226312 485044 226364
rect 485096 226352 485102 226364
rect 492582 226352 492588 226364
rect 485096 226324 492588 226352
rect 485096 226312 485102 226324
rect 492582 226312 492588 226324
rect 492640 226312 492646 226364
rect 544378 226312 544384 226364
rect 544436 226352 544442 226364
rect 548610 226352 548616 226364
rect 544436 226324 548616 226352
rect 544436 226312 544442 226324
rect 548610 226312 548616 226324
rect 548668 226312 548674 226364
rect 557506 226352 557534 226392
rect 558270 226352 558276 226364
rect 557506 226324 558276 226352
rect 558270 226312 558276 226324
rect 558328 226312 558334 226364
rect 100260 226256 100432 226284
rect 100260 226244 100266 226256
rect 568022 224408 568028 224460
rect 568080 224408 568086 224460
rect 120166 224272 120172 224324
rect 120224 224312 120230 224324
rect 122098 224312 122104 224324
rect 120224 224284 122104 224312
rect 120224 224272 120230 224284
rect 122098 224272 122104 224284
rect 122156 224272 122162 224324
rect 210418 224272 210424 224324
rect 210476 224312 210482 224324
rect 212442 224312 212448 224324
rect 210476 224284 212448 224312
rect 210476 224272 210482 224284
rect 212442 224272 212448 224284
rect 212500 224272 212506 224324
rect 512178 224272 512184 224324
rect 512236 224312 512242 224324
rect 514018 224312 514024 224324
rect 512236 224284 514024 224312
rect 512236 224272 512242 224284
rect 514018 224272 514024 224284
rect 514076 224272 514082 224324
rect 568040 224256 568068 224408
rect 568022 224204 568028 224256
rect 568080 224204 568086 224256
rect 182082 223728 182088 223780
rect 182140 223768 182146 223780
rect 233234 223768 233240 223780
rect 182140 223740 233240 223768
rect 182140 223728 182146 223740
rect 233234 223728 233240 223740
rect 233292 223728 233298 223780
rect 350442 223728 350448 223780
rect 350500 223768 350506 223780
rect 401594 223768 401600 223780
rect 350500 223740 401600 223768
rect 350500 223728 350506 223740
rect 401594 223728 401600 223740
rect 401652 223728 401658 223780
rect 462222 223728 462228 223780
rect 462280 223768 462286 223780
rect 513374 223768 513380 223780
rect 462280 223740 513380 223768
rect 462280 223728 462286 223740
rect 513374 223728 513380 223740
rect 513432 223728 513438 223780
rect 42702 223660 42708 223712
rect 42760 223700 42766 223712
rect 93854 223700 93860 223712
rect 42760 223672 93860 223700
rect 42760 223660 42766 223672
rect 93854 223660 93860 223672
rect 93912 223660 93918 223712
rect 97902 223660 97908 223712
rect 97960 223700 97966 223712
rect 149054 223700 149060 223712
rect 97960 223672 149060 223700
rect 97960 223660 97966 223672
rect 149054 223660 149060 223672
rect 149112 223660 149118 223712
rect 154482 223660 154488 223712
rect 154540 223700 154546 223712
rect 205634 223700 205640 223712
rect 154540 223672 205640 223700
rect 154540 223660 154546 223672
rect 205634 223660 205640 223672
rect 205692 223660 205698 223712
rect 238662 223660 238668 223712
rect 238720 223700 238726 223712
rect 289814 223700 289820 223712
rect 238720 223672 289820 223700
rect 238720 223660 238726 223672
rect 289814 223660 289820 223672
rect 289872 223660 289878 223712
rect 293862 223660 293868 223712
rect 293920 223700 293926 223712
rect 345014 223700 345020 223712
rect 293920 223672 345020 223700
rect 293920 223660 293926 223672
rect 345014 223660 345020 223672
rect 345072 223660 345078 223712
rect 378042 223660 378048 223712
rect 378100 223700 378106 223712
rect 429286 223700 429292 223712
rect 378100 223672 429292 223700
rect 378100 223660 378106 223672
rect 429286 223660 429292 223672
rect 429344 223660 429350 223712
rect 434622 223660 434628 223712
rect 434680 223700 434686 223712
rect 485774 223700 485780 223712
rect 434680 223672 485780 223700
rect 434680 223660 434686 223672
rect 485774 223660 485780 223672
rect 485832 223660 485838 223712
rect 518802 223660 518808 223712
rect 518860 223700 518866 223712
rect 569954 223700 569960 223712
rect 518860 223672 569960 223700
rect 518860 223660 518866 223672
rect 569954 223660 569960 223672
rect 570012 223660 570018 223712
rect 13538 223592 13544 223644
rect 13596 223632 13602 223644
rect 66254 223632 66260 223644
rect 13596 223604 66260 223632
rect 13596 223592 13602 223604
rect 66254 223592 66260 223604
rect 66312 223592 66318 223644
rect 70302 223592 70308 223644
rect 70360 223632 70366 223644
rect 121454 223632 121460 223644
rect 70360 223604 121460 223632
rect 70360 223592 70366 223604
rect 121454 223592 121460 223604
rect 121512 223592 121518 223644
rect 126882 223592 126888 223644
rect 126940 223632 126946 223644
rect 178034 223632 178040 223644
rect 126940 223604 178040 223632
rect 126940 223592 126946 223604
rect 178034 223592 178040 223604
rect 178092 223592 178098 223644
rect 209682 223592 209688 223644
rect 209740 223632 209746 223644
rect 262214 223632 262220 223644
rect 209740 223604 262220 223632
rect 209740 223592 209746 223604
rect 262214 223592 262220 223604
rect 262272 223592 262278 223644
rect 266262 223592 266268 223644
rect 266320 223632 266326 223644
rect 317414 223632 317420 223644
rect 266320 223604 317420 223632
rect 266320 223592 266326 223604
rect 317414 223592 317420 223604
rect 317472 223592 317478 223644
rect 322842 223592 322848 223644
rect 322900 223632 322906 223644
rect 373994 223632 374000 223644
rect 322900 223604 374000 223632
rect 322900 223592 322906 223604
rect 373994 223592 374000 223604
rect 374052 223592 374058 223644
rect 405642 223592 405648 223644
rect 405700 223632 405706 223644
rect 458174 223632 458180 223644
rect 405700 223604 458180 223632
rect 405700 223592 405706 223604
rect 458174 223592 458180 223604
rect 458232 223592 458238 223644
rect 489822 223592 489828 223644
rect 489880 223632 489886 223644
rect 542354 223632 542360 223644
rect 489880 223604 542360 223632
rect 489880 223592 489886 223604
rect 542354 223592 542360 223604
rect 542412 223592 542418 223644
rect 204254 221824 204260 221876
rect 204312 221864 204318 221876
rect 204990 221864 204996 221876
rect 204312 221836 204996 221864
rect 204312 221824 204318 221836
rect 204990 221824 204996 221836
rect 205048 221824 205054 221876
rect 64046 219716 64052 219768
rect 64104 219756 64110 219768
rect 64414 219756 64420 219768
rect 64104 219728 64420 219756
rect 64104 219716 64110 219728
rect 64414 219716 64420 219728
rect 64472 219716 64478 219768
rect 231854 203940 231860 203992
rect 231912 203980 231918 203992
rect 232130 203980 232136 203992
rect 231912 203952 232136 203980
rect 231912 203940 231918 203952
rect 232130 203940 232136 203952
rect 232188 203940 232194 203992
rect 15194 202784 15200 202836
rect 15252 202824 15258 202836
rect 35894 202824 35900 202836
rect 15252 202796 35900 202824
rect 15252 202784 15258 202796
rect 35894 202784 35900 202796
rect 35952 202784 35958 202836
rect 36078 202784 36084 202836
rect 36136 202824 36142 202836
rect 63586 202824 63592 202836
rect 36136 202796 63592 202824
rect 36136 202784 36142 202796
rect 63586 202784 63592 202796
rect 63644 202784 63650 202836
rect 64414 202784 64420 202836
rect 64472 202824 64478 202836
rect 91922 202824 91928 202836
rect 64472 202796 91928 202824
rect 64472 202784 64478 202796
rect 91922 202784 91928 202796
rect 91980 202784 91986 202836
rect 92106 202784 92112 202836
rect 92164 202824 92170 202836
rect 119614 202824 119620 202836
rect 92164 202796 119620 202824
rect 92164 202784 92170 202796
rect 119614 202784 119620 202796
rect 119672 202784 119678 202836
rect 122098 202784 122104 202836
rect 122156 202824 122162 202836
rect 147674 202824 147680 202836
rect 122156 202796 147680 202824
rect 122156 202784 122162 202796
rect 147674 202784 147680 202796
rect 147732 202784 147738 202836
rect 148042 202784 148048 202836
rect 148100 202824 148106 202836
rect 175918 202824 175924 202836
rect 148100 202796 175924 202824
rect 148100 202784 148106 202796
rect 175918 202784 175924 202796
rect 175976 202784 175982 202836
rect 176102 202784 176108 202836
rect 176160 202824 176166 202836
rect 203610 202824 203616 202836
rect 176160 202796 203616 202824
rect 176160 202784 176166 202796
rect 203610 202784 203616 202796
rect 203668 202784 203674 202836
rect 204990 202784 204996 202836
rect 205048 202824 205054 202836
rect 231854 202824 231860 202836
rect 205048 202796 231860 202824
rect 205048 202784 205054 202796
rect 231854 202784 231860 202796
rect 231912 202784 231918 202836
rect 232038 202784 232044 202836
rect 232096 202824 232102 202836
rect 259914 202824 259920 202836
rect 232096 202796 259920 202824
rect 232096 202784 232102 202796
rect 259914 202784 259920 202796
rect 259972 202784 259978 202836
rect 260098 202784 260104 202836
rect 260156 202824 260162 202836
rect 287606 202824 287612 202836
rect 260156 202796 287612 202824
rect 260156 202784 260162 202796
rect 287606 202784 287612 202796
rect 287664 202784 287670 202836
rect 288066 202784 288072 202836
rect 288124 202824 288130 202836
rect 315942 202824 315948 202836
rect 288124 202796 315948 202824
rect 288124 202784 288130 202796
rect 315942 202784 315948 202796
rect 316000 202784 316006 202836
rect 316678 202784 316684 202836
rect 316736 202824 316742 202836
rect 343910 202824 343916 202836
rect 316736 202796 343916 202824
rect 316736 202784 316742 202796
rect 343910 202784 343916 202796
rect 343968 202784 343974 202836
rect 344094 202784 344100 202836
rect 344152 202824 344158 202836
rect 371602 202824 371608 202836
rect 344152 202796 371608 202824
rect 344152 202784 344158 202796
rect 371602 202784 371608 202796
rect 371660 202784 371666 202836
rect 372062 202784 372068 202836
rect 372120 202824 372126 202836
rect 399938 202824 399944 202836
rect 372120 202796 399944 202824
rect 372120 202784 372126 202796
rect 399938 202784 399944 202796
rect 399996 202784 400002 202836
rect 400858 202784 400864 202836
rect 400916 202824 400922 202836
rect 427906 202824 427912 202836
rect 400916 202796 427912 202824
rect 400916 202784 400922 202796
rect 427906 202784 427912 202796
rect 427964 202784 427970 202836
rect 428090 202784 428096 202836
rect 428148 202824 428154 202836
rect 455598 202824 455604 202836
rect 428148 202796 455604 202824
rect 428148 202784 428154 202796
rect 455598 202784 455604 202796
rect 455656 202784 455662 202836
rect 456058 202784 456064 202836
rect 456116 202824 456122 202836
rect 483934 202824 483940 202836
rect 456116 202796 483940 202824
rect 456116 202784 456122 202796
rect 483934 202784 483940 202796
rect 483992 202784 483998 202836
rect 484026 202784 484032 202836
rect 484084 202824 484090 202836
rect 511902 202824 511908 202836
rect 484084 202796 511908 202824
rect 484084 202784 484090 202796
rect 511902 202784 511908 202796
rect 511960 202784 511966 202836
rect 514018 202784 514024 202836
rect 514076 202824 514082 202836
rect 539594 202824 539600 202836
rect 514076 202796 539600 202824
rect 514076 202784 514082 202796
rect 539594 202784 539600 202796
rect 539652 202784 539658 202836
rect 540054 202784 540060 202836
rect 540112 202824 540118 202836
rect 567930 202824 567936 202836
rect 540112 202796 567936 202824
rect 540112 202784 540118 202796
rect 567930 202784 567936 202796
rect 567988 202784 567994 202836
rect 16850 202716 16856 202768
rect 16908 202756 16914 202768
rect 36630 202756 36636 202768
rect 16908 202728 36636 202756
rect 16908 202716 16914 202728
rect 36630 202716 36636 202728
rect 36688 202716 36694 202768
rect 44910 202716 44916 202768
rect 44968 202756 44974 202768
rect 71130 202756 71136 202768
rect 44968 202728 71136 202756
rect 44968 202716 44974 202728
rect 71130 202716 71136 202728
rect 71188 202716 71194 202768
rect 82262 202716 82268 202768
rect 82320 202756 82326 202768
rect 93118 202756 93124 202768
rect 82320 202728 93124 202756
rect 82320 202716 82326 202728
rect 93118 202716 93124 202728
rect 93176 202716 93182 202768
rect 110230 202716 110236 202768
rect 110288 202756 110294 202768
rect 124858 202756 124864 202768
rect 110288 202728 124864 202756
rect 110288 202716 110294 202728
rect 124858 202716 124864 202728
rect 124916 202716 124922 202768
rect 128906 202716 128912 202768
rect 128964 202756 128970 202768
rect 151078 202756 151084 202768
rect 128964 202728 151084 202756
rect 128964 202716 128970 202728
rect 151078 202716 151084 202728
rect 151136 202716 151142 202768
rect 156598 202716 156604 202768
rect 156656 202756 156662 202768
rect 182818 202756 182824 202768
rect 156656 202728 182824 202756
rect 156656 202716 156662 202728
rect 182818 202716 182824 202728
rect 182876 202716 182882 202768
rect 194502 202716 194508 202768
rect 194560 202756 194566 202768
rect 210418 202756 210424 202768
rect 194560 202728 210424 202756
rect 194560 202716 194566 202728
rect 210418 202716 210424 202728
rect 210476 202716 210482 202768
rect 212994 202716 213000 202768
rect 213052 202756 213058 202768
rect 232498 202756 232504 202768
rect 213052 202728 232504 202756
rect 213052 202716 213058 202728
rect 232498 202716 232504 202728
rect 232556 202716 232562 202768
rect 240594 202716 240600 202768
rect 240652 202756 240658 202768
rect 266998 202756 267004 202768
rect 240652 202728 267004 202756
rect 240652 202716 240658 202728
rect 266998 202716 267004 202728
rect 267056 202716 267062 202768
rect 278590 202716 278596 202768
rect 278648 202756 278654 202768
rect 289078 202756 289084 202768
rect 278648 202728 289084 202756
rect 278648 202716 278654 202728
rect 289078 202716 289084 202728
rect 289136 202716 289142 202768
rect 306282 202716 306288 202768
rect 306340 202756 306346 202768
rect 318058 202756 318064 202768
rect 306340 202728 318064 202756
rect 306340 202716 306346 202728
rect 318058 202716 318064 202728
rect 318116 202716 318122 202768
rect 324590 202716 324596 202768
rect 324648 202756 324654 202768
rect 347038 202756 347044 202768
rect 324648 202728 347044 202756
rect 324648 202716 324654 202728
rect 347038 202716 347044 202728
rect 347096 202716 347102 202768
rect 362586 202716 362592 202768
rect 362644 202756 362650 202768
rect 373258 202756 373264 202768
rect 362644 202728 373264 202756
rect 362644 202716 362650 202728
rect 373258 202716 373264 202728
rect 373316 202716 373322 202768
rect 390278 202716 390284 202768
rect 390336 202756 390342 202768
rect 400950 202756 400956 202768
rect 390336 202728 400956 202756
rect 390336 202716 390342 202728
rect 400950 202716 400956 202728
rect 401008 202716 401014 202768
rect 408586 202716 408592 202768
rect 408644 202756 408650 202768
rect 428458 202756 428464 202768
rect 408644 202728 428464 202756
rect 408644 202716 408650 202728
rect 428458 202716 428464 202728
rect 428516 202716 428522 202768
rect 436922 202716 436928 202768
rect 436980 202756 436986 202768
rect 462958 202756 462964 202768
rect 436980 202728 462964 202756
rect 436980 202716 436986 202728
rect 462958 202716 462964 202728
rect 463016 202716 463022 202768
rect 474274 202716 474280 202768
rect 474332 202756 474338 202768
rect 485038 202756 485044 202768
rect 474332 202728 485044 202756
rect 474332 202716 474338 202728
rect 485038 202716 485044 202728
rect 485096 202716 485102 202768
rect 502242 202716 502248 202768
rect 502300 202756 502306 202768
rect 512638 202756 512644 202768
rect 502300 202728 512644 202756
rect 502300 202716 502306 202728
rect 512638 202716 512644 202728
rect 512696 202716 512702 202768
rect 520918 202716 520924 202768
rect 520976 202756 520982 202768
rect 541618 202756 541624 202768
rect 520976 202728 541624 202756
rect 520976 202716 520982 202728
rect 541618 202716 541624 202728
rect 541676 202716 541682 202768
rect 26602 202648 26608 202700
rect 26660 202688 26666 202700
rect 39298 202688 39304 202700
rect 26660 202660 39304 202688
rect 26660 202648 26666 202660
rect 39298 202648 39304 202660
rect 39356 202648 39362 202700
rect 54570 202648 54576 202700
rect 54628 202688 54634 202700
rect 66898 202688 66904 202700
rect 54628 202660 66904 202688
rect 54628 202648 54634 202660
rect 66898 202648 66904 202660
rect 66956 202648 66962 202700
rect 138658 202648 138664 202700
rect 138716 202688 138722 202700
rect 152458 202688 152464 202700
rect 138716 202660 152464 202688
rect 138716 202648 138722 202660
rect 152458 202648 152464 202660
rect 152516 202648 152522 202700
rect 166258 202648 166264 202700
rect 166316 202688 166322 202700
rect 177298 202688 177304 202700
rect 166316 202660 177304 202688
rect 166316 202648 166322 202660
rect 177298 202648 177304 202660
rect 177356 202648 177362 202700
rect 222562 202648 222568 202700
rect 222620 202688 222626 202700
rect 233970 202688 233976 202700
rect 222620 202660 233976 202688
rect 222620 202648 222626 202660
rect 233970 202648 233976 202660
rect 234028 202648 234034 202700
rect 250254 202648 250260 202700
rect 250312 202688 250318 202700
rect 261478 202688 261484 202700
rect 250312 202660 261484 202688
rect 250312 202648 250318 202660
rect 261478 202648 261484 202660
rect 261536 202648 261542 202700
rect 334250 202648 334256 202700
rect 334308 202688 334314 202700
rect 348418 202688 348424 202700
rect 334308 202660 348424 202688
rect 334308 202648 334314 202660
rect 348418 202648 348424 202660
rect 348476 202648 348482 202700
rect 418246 202648 418252 202700
rect 418304 202688 418310 202700
rect 429838 202688 429844 202700
rect 418304 202660 429844 202688
rect 418304 202648 418310 202660
rect 429838 202648 429844 202660
rect 429896 202648 429902 202700
rect 446582 202648 446588 202700
rect 446640 202688 446646 202700
rect 457438 202688 457444 202700
rect 446640 202660 457444 202688
rect 446640 202648 446646 202660
rect 457438 202648 457444 202660
rect 457496 202648 457502 202700
rect 530578 202648 530584 202700
rect 530636 202688 530642 202700
rect 544378 202688 544384 202700
rect 530636 202660 544384 202688
rect 530636 202648 530642 202660
rect 544378 202648 544384 202660
rect 544436 202648 544442 202700
rect 558270 202104 558276 202156
rect 558328 202144 558334 202156
rect 567470 202144 567476 202156
rect 558328 202116 567476 202144
rect 558328 202104 558334 202116
rect 567470 202104 567476 202116
rect 567528 202104 567534 202156
rect 3050 201492 3056 201544
rect 3108 201532 3114 201544
rect 64046 201532 64052 201544
rect 3108 201504 64052 201532
rect 3108 201492 3114 201504
rect 64046 201492 64052 201504
rect 64104 201492 64110 201544
rect 548334 200744 548340 200796
rect 548392 200784 548398 200796
rect 568114 200784 568120 200796
rect 548392 200756 568120 200784
rect 548392 200744 548398 200756
rect 568114 200744 568120 200756
rect 568172 200744 568178 200796
rect 296346 200336 296352 200388
rect 296404 200376 296410 200388
rect 316770 200376 316776 200388
rect 296404 200348 316776 200376
rect 296404 200336 296410 200348
rect 316770 200336 316776 200348
rect 316828 200336 316834 200388
rect 408034 200336 408040 200388
rect 408092 200376 408098 200388
rect 428642 200376 428648 200388
rect 408092 200348 428648 200376
rect 408092 200336 408098 200348
rect 428642 200336 428648 200348
rect 428700 200336 428706 200388
rect 492030 200336 492036 200388
rect 492088 200376 492094 200388
rect 512730 200376 512736 200388
rect 492088 200348 512736 200376
rect 492088 200336 492094 200348
rect 512730 200336 512736 200348
rect 512788 200336 512794 200388
rect 148410 200268 148416 200320
rect 148468 200308 148474 200320
rect 165614 200308 165620 200320
rect 148468 200280 165620 200308
rect 148468 200268 148474 200280
rect 165614 200268 165620 200280
rect 165672 200268 165678 200320
rect 175458 200268 175464 200320
rect 175516 200308 175522 200320
rect 193674 200308 193680 200320
rect 175516 200280 193680 200308
rect 175516 200268 175522 200280
rect 193674 200268 193680 200280
rect 193732 200268 193738 200320
rect 203518 200268 203524 200320
rect 203576 200308 203582 200320
rect 221366 200308 221372 200320
rect 203576 200280 221372 200308
rect 203576 200268 203582 200280
rect 221366 200268 221372 200280
rect 221424 200268 221430 200320
rect 232498 200268 232504 200320
rect 232556 200308 232562 200320
rect 249702 200308 249708 200320
rect 232556 200280 249708 200308
rect 232556 200268 232562 200280
rect 249702 200268 249708 200280
rect 249760 200268 249766 200320
rect 260190 200268 260196 200320
rect 260248 200308 260254 200320
rect 277670 200308 277676 200320
rect 260248 200280 277676 200308
rect 260248 200268 260254 200280
rect 277670 200268 277676 200280
rect 277728 200268 277734 200320
rect 287514 200268 287520 200320
rect 287572 200308 287578 200320
rect 305362 200308 305368 200320
rect 287572 200280 305368 200308
rect 287572 200268 287578 200280
rect 305362 200268 305368 200280
rect 305420 200268 305426 200320
rect 345658 200268 345664 200320
rect 345716 200308 345722 200320
rect 361666 200308 361672 200320
rect 345716 200280 361672 200308
rect 345716 200268 345722 200280
rect 361666 200268 361672 200280
rect 361724 200268 361730 200320
rect 371510 200268 371516 200320
rect 371568 200308 371574 200320
rect 389358 200308 389364 200320
rect 371568 200280 389364 200308
rect 371568 200268 371574 200280
rect 389358 200268 389364 200280
rect 389416 200268 389422 200320
rect 399478 200268 399484 200320
rect 399536 200308 399542 200320
rect 417694 200308 417700 200320
rect 399536 200280 417700 200308
rect 399536 200268 399542 200280
rect 417694 200268 417700 200280
rect 417752 200268 417758 200320
rect 456150 200268 456156 200320
rect 456208 200308 456214 200320
rect 473538 200308 473544 200320
rect 456208 200280 473544 200308
rect 456208 200268 456214 200280
rect 473538 200268 473544 200280
rect 473596 200268 473602 200320
rect 483474 200268 483480 200320
rect 483532 200308 483538 200320
rect 501690 200308 501696 200320
rect 483532 200280 501696 200308
rect 483532 200268 483538 200280
rect 501690 200268 501696 200280
rect 501748 200268 501754 200320
rect 36722 200200 36728 200252
rect 36780 200240 36786 200252
rect 53650 200240 53656 200252
rect 36780 200212 53656 200240
rect 36780 200200 36786 200212
rect 53650 200200 53656 200212
rect 53708 200200 53714 200252
rect 64414 200200 64420 200252
rect 64472 200240 64478 200252
rect 81434 200240 81440 200252
rect 64472 200212 81440 200240
rect 64472 200200 64478 200212
rect 81434 200200 81440 200212
rect 81492 200200 81498 200252
rect 91462 200200 91468 200252
rect 91520 200240 91526 200252
rect 109678 200240 109684 200252
rect 91520 200212 109684 200240
rect 91520 200200 91526 200212
rect 109678 200200 109684 200212
rect 109736 200200 109742 200252
rect 119430 200200 119436 200252
rect 119488 200240 119494 200252
rect 137646 200240 137652 200252
rect 119488 200212 137652 200240
rect 119488 200200 119494 200212
rect 137646 200200 137652 200212
rect 137704 200200 137710 200252
rect 156322 200200 156328 200252
rect 156380 200240 156386 200252
rect 178678 200240 178684 200252
rect 156380 200212 178684 200240
rect 156380 200200 156386 200212
rect 178678 200200 178684 200212
rect 178736 200200 178742 200252
rect 212258 200200 212264 200252
rect 212316 200240 212322 200252
rect 232682 200240 232688 200252
rect 212316 200212 232688 200240
rect 212316 200200 212322 200212
rect 232682 200200 232688 200212
rect 232740 200200 232746 200252
rect 268010 200200 268016 200252
rect 268068 200240 268074 200252
rect 287698 200240 287704 200252
rect 268068 200212 287704 200240
rect 268068 200200 268074 200212
rect 287698 200200 287704 200212
rect 287756 200200 287762 200252
rect 315482 200200 315488 200252
rect 315540 200240 315546 200252
rect 333698 200240 333704 200252
rect 315540 200212 333704 200240
rect 315540 200200 315546 200212
rect 333698 200200 333704 200212
rect 333756 200200 333762 200252
rect 352006 200200 352012 200252
rect 352064 200240 352070 200252
rect 374638 200240 374644 200252
rect 352064 200212 374644 200240
rect 352064 200200 352070 200212
rect 374638 200200 374644 200212
rect 374696 200200 374702 200252
rect 428458 200200 428464 200252
rect 428516 200240 428522 200252
rect 445662 200240 445668 200252
rect 428516 200212 445668 200240
rect 428516 200200 428522 200212
rect 445662 200200 445668 200212
rect 445720 200200 445726 200252
rect 464338 200200 464344 200252
rect 464396 200240 464402 200252
rect 483658 200240 483664 200252
rect 464396 200212 483664 200240
rect 464396 200200 464402 200212
rect 483658 200200 483664 200212
rect 483716 200200 483722 200252
rect 511442 200200 511448 200252
rect 511500 200240 511506 200252
rect 529658 200240 529664 200252
rect 511500 200212 529664 200240
rect 511500 200200 511506 200212
rect 529658 200200 529664 200212
rect 529716 200200 529722 200252
rect 541618 200200 541624 200252
rect 541676 200240 541682 200252
rect 557534 200240 557540 200252
rect 541676 200212 557540 200240
rect 541676 200200 541682 200212
rect 557534 200200 557540 200212
rect 557592 200200 557598 200252
rect 15102 200132 15108 200184
rect 15160 200172 15166 200184
rect 25682 200172 25688 200184
rect 15160 200144 25688 200172
rect 15160 200132 15166 200144
rect 25682 200132 25688 200144
rect 25740 200132 25746 200184
rect 36630 200132 36636 200184
rect 36688 200172 36694 200184
rect 63310 200172 63316 200184
rect 36688 200144 63316 200172
rect 36688 200132 36694 200144
rect 63310 200132 63316 200144
rect 63368 200132 63374 200184
rect 66898 200132 66904 200184
rect 66956 200172 66962 200184
rect 91094 200172 91100 200184
rect 66956 200144 91100 200172
rect 66956 200132 66962 200144
rect 91094 200132 91100 200144
rect 91152 200132 91158 200184
rect 93118 200132 93124 200184
rect 93176 200172 93182 200184
rect 119338 200172 119344 200184
rect 93176 200144 119344 200172
rect 93176 200132 93182 200144
rect 119338 200132 119344 200144
rect 119396 200132 119402 200184
rect 124858 200132 124864 200184
rect 124916 200172 124922 200184
rect 147306 200172 147312 200184
rect 124916 200144 147312 200172
rect 124916 200132 124922 200144
rect 147306 200132 147312 200144
rect 147364 200132 147370 200184
rect 148318 200132 148324 200184
rect 148376 200172 148382 200184
rect 175274 200172 175280 200184
rect 148376 200144 175280 200172
rect 148376 200132 148382 200144
rect 175274 200132 175280 200144
rect 175332 200132 175338 200184
rect 177298 200132 177304 200184
rect 177356 200172 177362 200184
rect 203334 200172 203340 200184
rect 177356 200144 203340 200172
rect 177356 200132 177362 200144
rect 203334 200132 203340 200144
rect 203392 200132 203398 200184
rect 204990 200132 204996 200184
rect 205048 200172 205054 200184
rect 231026 200172 231032 200184
rect 205048 200144 231032 200172
rect 205048 200132 205054 200144
rect 231026 200132 231032 200144
rect 231084 200132 231090 200184
rect 232590 200132 232596 200184
rect 232648 200172 232654 200184
rect 259362 200172 259368 200184
rect 232648 200144 259368 200172
rect 232648 200132 232654 200144
rect 259362 200132 259368 200144
rect 259420 200132 259426 200184
rect 260098 200132 260104 200184
rect 260156 200172 260162 200184
rect 287330 200172 287336 200184
rect 260156 200144 287336 200172
rect 260156 200132 260162 200144
rect 287330 200132 287336 200144
rect 287388 200132 287394 200184
rect 289078 200132 289084 200184
rect 289136 200172 289142 200184
rect 315022 200172 315028 200184
rect 289136 200144 315028 200172
rect 289136 200132 289142 200144
rect 315022 200132 315028 200144
rect 315080 200132 315086 200184
rect 316678 200132 316684 200184
rect 316736 200172 316742 200184
rect 343358 200172 343364 200184
rect 316736 200144 343364 200172
rect 316736 200132 316742 200144
rect 343358 200132 343364 200144
rect 343416 200132 343422 200184
rect 344278 200132 344284 200184
rect 344336 200172 344342 200184
rect 371326 200172 371332 200184
rect 344336 200144 371332 200172
rect 344336 200132 344342 200144
rect 371326 200132 371332 200144
rect 371384 200132 371390 200184
rect 373258 200132 373264 200184
rect 373316 200172 373322 200184
rect 399018 200172 399024 200184
rect 373316 200144 399024 200172
rect 373316 200132 373322 200144
rect 399018 200132 399024 200144
rect 399076 200132 399082 200184
rect 400858 200132 400864 200184
rect 400916 200172 400922 200184
rect 427354 200172 427360 200184
rect 400916 200144 427360 200172
rect 400916 200132 400922 200144
rect 427354 200132 427360 200144
rect 427412 200132 427418 200184
rect 428550 200132 428556 200184
rect 428608 200172 428614 200184
rect 455322 200172 455328 200184
rect 428608 200144 455328 200172
rect 428608 200132 428614 200144
rect 455322 200132 455328 200144
rect 455380 200132 455386 200184
rect 456058 200132 456064 200184
rect 456116 200172 456122 200184
rect 483198 200172 483204 200184
rect 456116 200144 483204 200172
rect 456116 200132 456122 200144
rect 483198 200132 483204 200144
rect 483256 200132 483262 200184
rect 485038 200132 485044 200184
rect 485096 200172 485102 200184
rect 511350 200172 511356 200184
rect 485096 200144 511356 200172
rect 485096 200132 485102 200144
rect 511350 200132 511356 200144
rect 511408 200132 511414 200184
rect 512638 200132 512644 200184
rect 512696 200172 512702 200184
rect 539318 200172 539324 200184
rect 512696 200144 539324 200172
rect 512696 200132 512702 200144
rect 539318 200132 539324 200144
rect 539376 200132 539382 200184
rect 540238 200132 540244 200184
rect 540296 200172 540302 200184
rect 567194 200172 567200 200184
rect 540296 200144 567200 200172
rect 540296 200132 540302 200144
rect 567194 200132 567200 200144
rect 567252 200132 567258 200184
rect 42886 193808 42892 193860
rect 42944 193848 42950 193860
rect 43622 193848 43628 193860
rect 42944 193820 43628 193848
rect 42944 193808 42950 193820
rect 43622 193808 43628 193820
rect 43680 193808 43686 193860
rect 570690 191836 570696 191888
rect 570748 191876 570754 191888
rect 580166 191876 580172 191888
rect 570748 191848 580172 191876
rect 570748 191836 570754 191848
rect 580166 191836 580172 191848
rect 580224 191836 580230 191888
rect 2958 187688 2964 187740
rect 3016 187728 3022 187740
rect 11790 187728 11796 187740
rect 3016 187700 11796 187728
rect 3016 187688 3022 187700
rect 11790 187688 11796 187700
rect 11848 187688 11854 187740
rect 147674 185580 147680 185632
rect 147732 185620 147738 185632
rect 148410 185620 148416 185632
rect 147732 185592 148416 185620
rect 147732 185580 147738 185592
rect 148410 185580 148416 185592
rect 148468 185580 148474 185632
rect 259730 185580 259736 185632
rect 259788 185620 259794 185632
rect 260190 185620 260196 185632
rect 259788 185592 260196 185620
rect 259788 185580 259794 185592
rect 260190 185580 260196 185592
rect 260248 185580 260254 185632
rect 455690 185580 455696 185632
rect 455748 185620 455754 185632
rect 456150 185620 456156 185632
rect 455748 185592 456156 185620
rect 455748 185580 455754 185592
rect 456150 185580 456156 185592
rect 456208 185580 456214 185632
rect 63586 181432 63592 181484
rect 63644 181472 63650 181484
rect 64414 181472 64420 181484
rect 63644 181444 64420 181472
rect 63644 181432 63650 181444
rect 64414 181432 64420 181444
rect 64472 181432 64478 181484
rect 512730 180208 512736 180260
rect 512788 180248 512794 180260
rect 519630 180248 519636 180260
rect 512788 180220 519636 180248
rect 512788 180208 512794 180220
rect 519630 180208 519636 180220
rect 519688 180208 519694 180260
rect 428642 180072 428648 180124
rect 428700 180112 428706 180124
rect 435726 180112 435732 180124
rect 428700 180084 435732 180112
rect 428700 180072 428706 180084
rect 435726 180072 435732 180084
rect 435784 180072 435790 180124
rect 232682 179868 232688 179920
rect 232740 179908 232746 179920
rect 239766 179908 239772 179920
rect 232740 179880 239772 179908
rect 232740 179868 232746 179880
rect 239766 179868 239772 179880
rect 239824 179868 239830 179920
rect 483658 179664 483664 179716
rect 483716 179704 483722 179716
rect 491662 179704 491668 179716
rect 483716 179676 491668 179704
rect 483716 179664 483722 179676
rect 491662 179664 491668 179676
rect 491720 179664 491726 179716
rect 316770 179460 316776 179512
rect 316828 179500 316834 179512
rect 323670 179500 323676 179512
rect 316828 179472 323676 179500
rect 316828 179460 316834 179472
rect 323670 179460 323676 179472
rect 323728 179460 323734 179512
rect 287698 179392 287704 179444
rect 287756 179432 287762 179444
rect 295702 179432 295708 179444
rect 287756 179404 295708 179432
rect 287756 179392 287762 179404
rect 295702 179392 295708 179404
rect 295760 179392 295766 179444
rect 13538 179324 13544 179376
rect 13596 179364 13602 179376
rect 66254 179364 66260 179376
rect 13596 179336 66260 179364
rect 13596 179324 13602 179336
rect 66254 179324 66260 179336
rect 66312 179324 66318 179376
rect 70302 179324 70308 179376
rect 70360 179364 70366 179376
rect 121454 179364 121460 179376
rect 70360 179336 121460 179364
rect 70360 179324 70366 179336
rect 121454 179324 121460 179336
rect 121512 179324 121518 179376
rect 126882 179324 126888 179376
rect 126940 179364 126946 179376
rect 178034 179364 178040 179376
rect 126940 179336 178040 179364
rect 126940 179324 126946 179336
rect 178034 179324 178040 179336
rect 178092 179324 178098 179376
rect 209682 179324 209688 179376
rect 209740 179364 209746 179376
rect 262214 179364 262220 179376
rect 209740 179336 262220 179364
rect 209740 179324 209746 179336
rect 262214 179324 262220 179336
rect 262272 179324 262278 179376
rect 266262 179324 266268 179376
rect 266320 179364 266326 179376
rect 317414 179364 317420 179376
rect 266320 179336 317420 179364
rect 266320 179324 266326 179336
rect 317414 179324 317420 179336
rect 317472 179324 317478 179376
rect 322842 179324 322848 179376
rect 322900 179364 322906 179376
rect 373994 179364 374000 179376
rect 322900 179336 374000 179364
rect 322900 179324 322906 179336
rect 373994 179324 374000 179336
rect 374052 179324 374058 179376
rect 405642 179324 405648 179376
rect 405700 179364 405706 179376
rect 458174 179364 458180 179376
rect 405700 179336 458180 179364
rect 405700 179324 405706 179336
rect 458174 179324 458180 179336
rect 458232 179324 458238 179376
rect 489822 179324 489828 179376
rect 489880 179364 489886 179376
rect 489880 179336 539364 179364
rect 489880 179324 489886 179336
rect 42702 179256 42708 179308
rect 42760 179296 42766 179308
rect 93854 179296 93860 179308
rect 42760 179268 93860 179296
rect 42760 179256 42766 179268
rect 93854 179256 93860 179268
rect 93912 179256 93918 179308
rect 97902 179256 97908 179308
rect 97960 179296 97966 179308
rect 149054 179296 149060 179308
rect 97960 179268 149060 179296
rect 97960 179256 97966 179268
rect 149054 179256 149060 179268
rect 149112 179256 149118 179308
rect 154482 179256 154488 179308
rect 154540 179296 154546 179308
rect 205634 179296 205640 179308
rect 154540 179268 205640 179296
rect 154540 179256 154546 179268
rect 205634 179256 205640 179268
rect 205692 179256 205698 179308
rect 238662 179256 238668 179308
rect 238720 179296 238726 179308
rect 289814 179296 289820 179308
rect 238720 179268 289820 179296
rect 238720 179256 238726 179268
rect 289814 179256 289820 179268
rect 289872 179256 289878 179308
rect 293862 179256 293868 179308
rect 293920 179296 293926 179308
rect 293920 179268 335354 179296
rect 293920 179256 293926 179268
rect 182082 179188 182088 179240
rect 182140 179228 182146 179240
rect 233234 179228 233240 179240
rect 182140 179200 233240 179228
rect 182140 179188 182146 179200
rect 233234 179188 233240 179200
rect 233292 179188 233298 179240
rect 335326 179228 335354 179268
rect 343542 179256 343548 179308
rect 343600 179296 343606 179308
rect 345658 179296 345664 179308
rect 343600 179268 345664 179296
rect 343600 179256 343606 179268
rect 345658 179256 345664 179268
rect 345716 179256 345722 179308
rect 378042 179256 378048 179308
rect 378100 179296 378106 179308
rect 429286 179296 429292 179308
rect 378100 179268 429292 179296
rect 378100 179256 378106 179268
rect 429286 179256 429292 179268
rect 429344 179256 429350 179308
rect 434622 179256 434628 179308
rect 434680 179296 434686 179308
rect 485774 179296 485780 179308
rect 434680 179268 485780 179296
rect 434680 179256 434686 179268
rect 485774 179256 485780 179268
rect 485832 179256 485838 179308
rect 518802 179256 518808 179308
rect 518860 179296 518866 179308
rect 518860 179268 528554 179296
rect 518860 179256 518866 179268
rect 345014 179228 345020 179240
rect 335326 179200 345020 179228
rect 345014 179188 345020 179200
rect 345072 179188 345078 179240
rect 350442 179188 350448 179240
rect 350500 179228 350506 179240
rect 401594 179228 401600 179240
rect 350500 179200 401600 179228
rect 350500 179188 350506 179200
rect 401594 179188 401600 179200
rect 401652 179188 401658 179240
rect 462222 179188 462228 179240
rect 462280 179228 462286 179240
rect 513374 179228 513380 179240
rect 462280 179200 513380 179228
rect 462280 179188 462286 179200
rect 513374 179188 513380 179200
rect 513432 179188 513438 179240
rect 528526 179160 528554 179268
rect 539336 179228 539364 179336
rect 539502 179324 539508 179376
rect 539560 179364 539566 179376
rect 541618 179364 541624 179376
rect 539560 179336 541624 179364
rect 539560 179324 539566 179336
rect 541618 179324 541624 179336
rect 541676 179324 541682 179376
rect 569954 179296 569960 179308
rect 547846 179268 569960 179296
rect 542354 179228 542360 179240
rect 539336 179200 542360 179228
rect 542354 179188 542360 179200
rect 542412 179188 542418 179240
rect 547846 179160 547874 179268
rect 569954 179256 569960 179268
rect 570012 179256 570018 179308
rect 528526 179132 547874 179160
rect 15102 178712 15108 178764
rect 15160 178752 15166 178764
rect 16574 178752 16580 178764
rect 15160 178724 16580 178752
rect 15160 178712 15166 178724
rect 16574 178712 16580 178724
rect 16632 178712 16638 178764
rect 35250 178712 35256 178764
rect 35308 178752 35314 178764
rect 36722 178752 36728 178764
rect 35308 178724 36728 178752
rect 35308 178712 35314 178724
rect 36722 178712 36728 178724
rect 36780 178712 36786 178764
rect 547874 178712 547880 178764
rect 547932 178752 547938 178764
rect 548150 178752 548156 178764
rect 547932 178724 548156 178752
rect 547932 178712 547938 178724
rect 548150 178712 548156 178724
rect 548208 178712 548214 178764
rect 71866 176604 71872 176656
rect 71924 176644 71930 176656
rect 100018 176644 100024 176656
rect 71924 176616 100024 176644
rect 71924 176604 71930 176616
rect 100018 176604 100024 176616
rect 100076 176604 100082 176656
rect 127986 176644 127992 176656
rect 103486 176616 127992 176644
rect 25682 176536 25688 176588
rect 25740 176576 25746 176588
rect 36630 176576 36636 176588
rect 25740 176548 36636 176576
rect 25740 176536 25746 176548
rect 36630 176536 36636 176548
rect 36688 176536 36694 176588
rect 42886 176536 42892 176588
rect 42944 176576 42950 176588
rect 42944 176548 45554 176576
rect 42944 176536 42950 176548
rect 15286 176468 15292 176520
rect 15344 176508 15350 176520
rect 43990 176508 43996 176520
rect 15344 176480 43996 176508
rect 15344 176468 15350 176480
rect 43990 176468 43996 176480
rect 44048 176468 44054 176520
rect 45526 176508 45554 176548
rect 53650 176536 53656 176588
rect 53708 176576 53714 176588
rect 66898 176576 66904 176588
rect 53708 176548 66904 176576
rect 53708 176536 53714 176548
rect 66898 176536 66904 176548
rect 66956 176536 66962 176588
rect 81986 176536 81992 176588
rect 82044 176576 82050 176588
rect 93118 176576 93124 176588
rect 82044 176548 93124 176576
rect 82044 176536 82050 176548
rect 93118 176536 93124 176548
rect 93176 176536 93182 176588
rect 99466 176536 99472 176588
rect 99524 176576 99530 176588
rect 103486 176576 103514 176616
rect 127986 176604 127992 176616
rect 128044 176604 128050 176656
rect 165982 176604 165988 176656
rect 166040 176644 166046 176656
rect 177298 176644 177304 176656
rect 166040 176616 177304 176644
rect 166040 176604 166046 176616
rect 177298 176604 177304 176616
rect 177356 176604 177362 176656
rect 178678 176604 178684 176656
rect 178736 176644 178742 176656
rect 184014 176644 184020 176656
rect 178736 176616 184020 176644
rect 178736 176604 178742 176616
rect 184014 176604 184020 176616
rect 184072 176604 184078 176656
rect 211706 176644 211712 176656
rect 190426 176616 211712 176644
rect 99524 176548 103514 176576
rect 99524 176536 99530 176548
rect 109678 176536 109684 176588
rect 109736 176576 109742 176588
rect 124858 176576 124864 176588
rect 109736 176548 124864 176576
rect 109736 176536 109742 176548
rect 124858 176536 124864 176548
rect 124916 176536 124922 176588
rect 137646 176536 137652 176588
rect 137704 176576 137710 176588
rect 148318 176576 148324 176588
rect 137704 176548 148324 176576
rect 137704 176536 137710 176548
rect 148318 176536 148324 176548
rect 148376 176536 148382 176588
rect 183646 176536 183652 176588
rect 183704 176576 183710 176588
rect 190426 176576 190454 176616
rect 211706 176604 211712 176616
rect 211764 176604 211770 176656
rect 277670 176604 277676 176656
rect 277728 176644 277734 176656
rect 289078 176644 289084 176656
rect 277728 176616 289084 176644
rect 277728 176604 277734 176616
rect 289078 176604 289084 176616
rect 289136 176604 289142 176656
rect 306006 176604 306012 176656
rect 306064 176644 306070 176656
rect 316678 176644 316684 176656
rect 306064 176616 316684 176644
rect 306064 176604 306070 176616
rect 316678 176604 316684 176616
rect 316736 176604 316742 176656
rect 361666 176604 361672 176656
rect 361724 176644 361730 176656
rect 373258 176644 373264 176656
rect 361724 176616 373264 176644
rect 361724 176604 361730 176616
rect 373258 176604 373264 176616
rect 373316 176604 373322 176656
rect 374638 176604 374644 176656
rect 374696 176644 374702 176656
rect 379698 176644 379704 176656
rect 374696 176616 379704 176644
rect 374696 176604 374702 176616
rect 379698 176604 379704 176616
rect 379756 176604 379762 176656
rect 408034 176644 408040 176656
rect 383626 176616 408040 176644
rect 183704 176548 190454 176576
rect 183704 176536 183710 176548
rect 193674 176536 193680 176588
rect 193732 176576 193738 176588
rect 204990 176576 204996 176588
rect 193732 176548 204996 176576
rect 193732 176536 193738 176548
rect 204990 176536 204996 176548
rect 205048 176536 205054 176588
rect 222010 176536 222016 176588
rect 222068 176576 222074 176588
rect 232590 176576 232596 176588
rect 222068 176548 232596 176576
rect 222068 176536 222074 176548
rect 232590 176536 232596 176548
rect 232648 176536 232654 176588
rect 249702 176536 249708 176588
rect 249760 176576 249766 176588
rect 260098 176576 260104 176588
rect 249760 176548 260104 176576
rect 249760 176536 249766 176548
rect 260098 176536 260104 176548
rect 260156 176536 260162 176588
rect 333698 176536 333704 176588
rect 333756 176576 333762 176588
rect 344278 176576 344284 176588
rect 333756 176548 344284 176576
rect 333756 176536 333762 176548
rect 344278 176536 344284 176548
rect 344336 176536 344342 176588
rect 379606 176536 379612 176588
rect 379664 176576 379670 176588
rect 383626 176576 383654 176616
rect 408034 176604 408040 176616
rect 408092 176604 408098 176656
rect 473998 176604 474004 176656
rect 474056 176644 474062 176656
rect 485038 176644 485044 176656
rect 474056 176616 485044 176644
rect 474056 176604 474062 176616
rect 485038 176604 485044 176616
rect 485096 176604 485102 176656
rect 501690 176604 501696 176656
rect 501748 176644 501754 176656
rect 512638 176644 512644 176656
rect 501748 176616 512644 176644
rect 501748 176604 501754 176616
rect 512638 176604 512644 176616
rect 512696 176604 512702 176656
rect 548150 176604 548156 176656
rect 548208 176644 548214 176656
rect 557534 176644 557540 176656
rect 548208 176616 557540 176644
rect 548208 176604 548214 176616
rect 557534 176604 557540 176616
rect 557592 176604 557598 176656
rect 379664 176548 383654 176576
rect 379664 176536 379670 176548
rect 390002 176536 390008 176588
rect 390060 176576 390066 176588
rect 400858 176576 400864 176588
rect 390060 176548 400864 176576
rect 390060 176536 390066 176548
rect 400858 176536 400864 176548
rect 400916 176536 400922 176588
rect 417694 176536 417700 176588
rect 417752 176576 417758 176588
rect 428550 176576 428556 176588
rect 417752 176548 428556 176576
rect 417752 176536 417758 176548
rect 428550 176536 428556 176548
rect 428608 176536 428614 176588
rect 445662 176536 445668 176588
rect 445720 176576 445726 176588
rect 456058 176576 456064 176588
rect 445720 176548 456064 176576
rect 445720 176536 445726 176548
rect 456058 176536 456064 176548
rect 456116 176536 456122 176588
rect 529658 176536 529664 176588
rect 529716 176576 529722 176588
rect 540238 176576 540244 176588
rect 529716 176548 540244 176576
rect 529716 176536 529722 176548
rect 540238 176536 540244 176548
rect 540296 176536 540302 176588
rect 72050 176508 72056 176520
rect 45526 176480 72056 176508
rect 72050 176468 72056 176480
rect 72108 176468 72114 176520
rect 127066 176468 127072 176520
rect 127124 176508 127130 176520
rect 156046 176508 156052 176520
rect 127124 176480 156052 176508
rect 127124 176468 127130 176480
rect 156046 176468 156052 176480
rect 156104 176468 156110 176520
rect 238846 176468 238852 176520
rect 238904 176508 238910 176520
rect 268010 176508 268016 176520
rect 238904 176480 268016 176508
rect 238904 176468 238910 176480
rect 268010 176468 268016 176480
rect 268068 176468 268074 176520
rect 323026 176468 323032 176520
rect 323084 176508 323090 176520
rect 352006 176508 352012 176520
rect 323084 176480 352012 176508
rect 323084 176468 323090 176480
rect 352006 176468 352012 176480
rect 352064 176468 352070 176520
rect 434806 176468 434812 176520
rect 434864 176508 434870 176520
rect 463694 176508 463700 176520
rect 434864 176480 463700 176508
rect 434864 176468 434870 176480
rect 463694 176468 463700 176480
rect 463752 176468 463758 176520
rect 518986 176468 518992 176520
rect 519044 176508 519050 176520
rect 547874 176508 547880 176520
rect 519044 176480 547880 176508
rect 519044 176468 519050 176480
rect 547874 176468 547880 176480
rect 547932 176468 547938 176520
rect 26234 172796 26240 172848
rect 26292 172836 26298 172848
rect 35434 172836 35440 172848
rect 26292 172808 35440 172836
rect 26292 172796 26298 172808
rect 35434 172796 35440 172808
rect 35492 172796 35498 172848
rect 71130 172660 71136 172712
rect 71188 172700 71194 172712
rect 82262 172700 82268 172712
rect 71188 172672 82268 172700
rect 71188 172660 71194 172672
rect 82262 172660 82268 172672
rect 82320 172660 82326 172712
rect 99374 172660 99380 172712
rect 99432 172700 99438 172712
rect 100294 172700 100300 172712
rect 99432 172672 100300 172700
rect 99432 172660 99438 172672
rect 100294 172660 100300 172672
rect 100352 172660 100358 172712
rect 183646 172660 183652 172712
rect 183704 172700 183710 172712
rect 222286 172700 222292 172712
rect 183704 172672 222292 172700
rect 183704 172660 183710 172672
rect 222286 172660 222292 172672
rect 222344 172660 222350 172712
rect 261478 172660 261484 172712
rect 261536 172700 261542 172712
rect 268286 172700 268292 172712
rect 261536 172672 268292 172700
rect 261536 172660 261542 172672
rect 268286 172660 268292 172672
rect 268344 172660 268350 172712
rect 295426 172660 295432 172712
rect 295484 172700 295490 172712
rect 334250 172700 334256 172712
rect 295484 172672 334256 172700
rect 295484 172660 295490 172672
rect 334250 172660 334256 172672
rect 334308 172660 334314 172712
rect 352006 172660 352012 172712
rect 352064 172700 352070 172712
rect 352064 172672 364334 172700
rect 352064 172660 352070 172672
rect 36630 172592 36636 172644
rect 36688 172632 36694 172644
rect 53926 172632 53932 172644
rect 36688 172604 53932 172632
rect 36688 172592 36694 172604
rect 53926 172592 53932 172604
rect 53984 172592 53990 172644
rect 71866 172592 71872 172644
rect 71924 172632 71930 172644
rect 109954 172632 109960 172644
rect 71924 172604 109960 172632
rect 71924 172592 71930 172604
rect 109954 172592 109960 172604
rect 110012 172592 110018 172644
rect 124858 172592 124864 172644
rect 124916 172632 124922 172644
rect 128630 172632 128636 172644
rect 124916 172604 128636 172632
rect 124916 172592 124922 172604
rect 128630 172592 128636 172604
rect 128688 172592 128694 172644
rect 152458 172592 152464 172644
rect 152516 172632 152522 172644
rect 156598 172632 156604 172644
rect 152516 172604 156604 172632
rect 152516 172592 152522 172604
rect 156598 172592 156604 172604
rect 156656 172592 156662 172644
rect 182818 172592 182824 172644
rect 182876 172632 182882 172644
rect 193950 172632 193956 172644
rect 182876 172604 193956 172632
rect 182876 172592 182882 172604
rect 193950 172592 193956 172604
rect 194008 172592 194014 172644
rect 232498 172592 232504 172644
rect 232556 172632 232562 172644
rect 232556 172604 248414 172632
rect 232556 172592 232562 172604
rect 39298 172524 39304 172576
rect 39356 172564 39362 172576
rect 44266 172564 44272 172576
rect 39356 172536 44272 172564
rect 39356 172524 39362 172536
rect 44266 172524 44272 172536
rect 44324 172524 44330 172576
rect 66898 172524 66904 172576
rect 66956 172564 66962 172576
rect 72602 172564 72608 172576
rect 66956 172536 72608 172564
rect 66956 172524 66962 172536
rect 72602 172524 72608 172536
rect 72660 172524 72666 172576
rect 93118 172524 93124 172576
rect 93176 172564 93182 172576
rect 99374 172564 99380 172576
rect 93176 172536 99380 172564
rect 93176 172524 93182 172536
rect 99374 172524 99380 172536
rect 99432 172524 99438 172576
rect 99466 172524 99472 172576
rect 99524 172564 99530 172576
rect 138290 172564 138296 172576
rect 99524 172536 138296 172564
rect 99524 172524 99530 172536
rect 138290 172524 138296 172536
rect 138348 172524 138354 172576
rect 151078 172524 151084 172576
rect 151136 172564 151142 172576
rect 166258 172564 166264 172576
rect 151136 172536 166264 172564
rect 151136 172524 151142 172536
rect 166258 172524 166264 172536
rect 166316 172524 166322 172576
rect 177298 172524 177304 172576
rect 177356 172564 177362 172576
rect 184290 172564 184296 172576
rect 177356 172536 184296 172564
rect 177356 172524 177362 172536
rect 184290 172524 184296 172536
rect 184348 172524 184354 172576
rect 233970 172524 233976 172576
rect 234028 172564 234034 172576
rect 240594 172564 240600 172576
rect 234028 172536 240600 172564
rect 234028 172524 234034 172536
rect 240594 172524 240600 172536
rect 240652 172524 240658 172576
rect 248386 172564 248414 172604
rect 267826 172592 267832 172644
rect 267884 172632 267890 172644
rect 306282 172632 306288 172644
rect 267884 172604 306288 172632
rect 267884 172592 267890 172604
rect 306282 172592 306288 172604
rect 306340 172592 306346 172644
rect 345658 172592 345664 172644
rect 345716 172632 345722 172644
rect 361942 172632 361948 172644
rect 345716 172604 361948 172632
rect 345716 172592 345722 172604
rect 361942 172592 361948 172604
rect 362000 172592 362006 172644
rect 364306 172632 364334 172672
rect 379606 172660 379612 172712
rect 379664 172700 379670 172712
rect 418246 172700 418252 172712
rect 379664 172672 418252 172700
rect 379664 172660 379670 172672
rect 418246 172660 418252 172672
rect 418304 172660 418310 172712
rect 463786 172660 463792 172712
rect 463844 172700 463850 172712
rect 463844 172672 470594 172700
rect 463844 172660 463850 172672
rect 390278 172632 390284 172644
rect 364306 172604 390284 172632
rect 390278 172592 390284 172604
rect 390336 172592 390342 172644
rect 400950 172592 400956 172644
rect 401008 172632 401014 172644
rect 408586 172632 408592 172644
rect 401008 172604 408592 172632
rect 401008 172592 401014 172604
rect 408586 172592 408592 172604
rect 408644 172592 408650 172644
rect 429838 172592 429844 172644
rect 429896 172632 429902 172644
rect 436278 172632 436284 172644
rect 429896 172604 436284 172632
rect 429896 172592 429902 172604
rect 436278 172592 436284 172604
rect 436336 172592 436342 172644
rect 457438 172592 457444 172644
rect 457496 172632 457502 172644
rect 464614 172632 464620 172644
rect 457496 172604 464620 172632
rect 457496 172592 457502 172604
rect 464614 172592 464620 172604
rect 464672 172592 464678 172644
rect 470566 172632 470594 172672
rect 485038 172660 485044 172712
rect 485096 172700 485102 172712
rect 492582 172700 492588 172712
rect 485096 172672 492588 172700
rect 485096 172660 485102 172672
rect 492582 172660 492588 172672
rect 492640 172660 492646 172712
rect 502242 172632 502248 172644
rect 470566 172604 502248 172632
rect 502242 172592 502248 172604
rect 502300 172592 502306 172644
rect 514018 172592 514024 172644
rect 514076 172632 514082 172644
rect 520274 172632 520280 172644
rect 514076 172604 520280 172632
rect 514076 172592 514082 172604
rect 520274 172592 520280 172604
rect 520332 172592 520338 172644
rect 541618 172592 541624 172644
rect 541676 172632 541682 172644
rect 541676 172604 557534 172632
rect 541676 172592 541682 172604
rect 250254 172564 250260 172576
rect 248386 172536 250260 172564
rect 250254 172524 250260 172536
rect 250312 172524 250318 172576
rect 266998 172524 267004 172576
rect 267056 172564 267062 172576
rect 277946 172564 277952 172576
rect 267056 172536 277952 172564
rect 267056 172524 267062 172536
rect 277946 172524 277952 172536
rect 278004 172524 278010 172576
rect 289078 172524 289084 172576
rect 289136 172564 289142 172576
rect 296622 172564 296628 172576
rect 289136 172536 296628 172564
rect 289136 172524 289142 172536
rect 296622 172524 296628 172536
rect 296680 172524 296686 172576
rect 318058 172524 318064 172576
rect 318116 172564 318122 172576
rect 324590 172564 324596 172576
rect 318116 172536 324596 172564
rect 318116 172524 318122 172536
rect 324590 172524 324596 172536
rect 324648 172524 324654 172576
rect 347038 172524 347044 172576
rect 347096 172564 347102 172576
rect 352282 172564 352288 172576
rect 347096 172536 352288 172564
rect 347096 172524 347102 172536
rect 352282 172524 352288 172536
rect 352340 172524 352346 172576
rect 373258 172524 373264 172576
rect 373316 172564 373322 172576
rect 380618 172564 380624 172576
rect 373316 172536 380624 172564
rect 373316 172524 373322 172536
rect 380618 172524 380624 172536
rect 380676 172524 380682 172576
rect 428458 172524 428464 172576
rect 428516 172564 428522 172576
rect 445938 172564 445944 172576
rect 428516 172536 445944 172564
rect 428516 172524 428522 172536
rect 445938 172524 445944 172536
rect 445996 172524 446002 172576
rect 462958 172524 462964 172576
rect 463016 172564 463022 172576
rect 474274 172564 474280 172576
rect 463016 172536 474280 172564
rect 463016 172524 463022 172536
rect 474274 172524 474280 172536
rect 474332 172524 474338 172576
rect 491386 172524 491392 172576
rect 491444 172564 491450 172576
rect 529934 172564 529940 172576
rect 491444 172536 529940 172564
rect 491444 172524 491450 172536
rect 529934 172524 529940 172536
rect 529992 172524 529998 172576
rect 544378 172524 544384 172576
rect 544436 172564 544442 172576
rect 548610 172564 548616 172576
rect 544436 172536 548616 172564
rect 544436 172524 544442 172536
rect 548610 172524 548616 172536
rect 548668 172524 548674 172576
rect 557506 172564 557534 172604
rect 558270 172564 558276 172576
rect 557506 172536 558276 172564
rect 558270 172524 558276 172536
rect 558328 172524 558334 172576
rect 210418 171096 210424 171148
rect 210476 171136 210482 171148
rect 212626 171136 212632 171148
rect 210476 171108 212632 171136
rect 210476 171096 210482 171108
rect 212626 171096 212632 171108
rect 212684 171096 212690 171148
rect 568022 170416 568028 170468
rect 568080 170416 568086 170468
rect 63770 170280 63776 170332
rect 63828 170320 63834 170332
rect 65794 170320 65800 170332
rect 63828 170292 65800 170320
rect 63828 170280 63834 170292
rect 65794 170280 65800 170292
rect 65852 170280 65858 170332
rect 120166 170280 120172 170332
rect 120224 170320 120230 170332
rect 122098 170320 122104 170332
rect 120224 170292 122104 170320
rect 120224 170280 120230 170292
rect 122098 170280 122104 170292
rect 122156 170280 122162 170332
rect 568040 170264 568068 170416
rect 568022 170212 568028 170264
rect 568080 170212 568086 170264
rect 204254 165860 204260 165912
rect 204312 165900 204318 165912
rect 204990 165900 204996 165912
rect 204312 165872 204996 165900
rect 204312 165860 204318 165872
rect 204990 165860 204996 165872
rect 205048 165860 205054 165912
rect 13538 151716 13544 151768
rect 13596 151756 13602 151768
rect 66254 151756 66260 151768
rect 13596 151728 66260 151756
rect 13596 151716 13602 151728
rect 66254 151716 66260 151728
rect 66312 151716 66318 151768
rect 70302 151716 70308 151768
rect 70360 151756 70366 151768
rect 121454 151756 121460 151768
rect 70360 151728 121460 151756
rect 70360 151716 70366 151728
rect 121454 151716 121460 151728
rect 121512 151716 121518 151768
rect 126882 151716 126888 151768
rect 126940 151756 126946 151768
rect 178034 151756 178040 151768
rect 126940 151728 178040 151756
rect 126940 151716 126946 151728
rect 178034 151716 178040 151728
rect 178092 151716 178098 151768
rect 209682 151716 209688 151768
rect 209740 151756 209746 151768
rect 262214 151756 262220 151768
rect 209740 151728 262220 151756
rect 209740 151716 209746 151728
rect 262214 151716 262220 151728
rect 262272 151716 262278 151768
rect 266262 151716 266268 151768
rect 266320 151756 266326 151768
rect 317414 151756 317420 151768
rect 266320 151728 317420 151756
rect 266320 151716 266326 151728
rect 317414 151716 317420 151728
rect 317472 151716 317478 151768
rect 322842 151716 322848 151768
rect 322900 151756 322906 151768
rect 373994 151756 374000 151768
rect 322900 151728 374000 151756
rect 322900 151716 322906 151728
rect 373994 151716 374000 151728
rect 374052 151716 374058 151768
rect 405642 151716 405648 151768
rect 405700 151756 405706 151768
rect 458174 151756 458180 151768
rect 405700 151728 458180 151756
rect 405700 151716 405706 151728
rect 458174 151716 458180 151728
rect 458232 151716 458238 151768
rect 489822 151716 489828 151768
rect 489880 151756 489886 151768
rect 542354 151756 542360 151768
rect 489880 151728 542360 151756
rect 489880 151716 489886 151728
rect 542354 151716 542360 151728
rect 542412 151716 542418 151768
rect 42702 151648 42708 151700
rect 42760 151688 42766 151700
rect 93854 151688 93860 151700
rect 42760 151660 93860 151688
rect 42760 151648 42766 151660
rect 93854 151648 93860 151660
rect 93912 151648 93918 151700
rect 97902 151648 97908 151700
rect 97960 151688 97966 151700
rect 149054 151688 149060 151700
rect 97960 151660 149060 151688
rect 97960 151648 97966 151660
rect 149054 151648 149060 151660
rect 149112 151648 149118 151700
rect 154482 151648 154488 151700
rect 154540 151688 154546 151700
rect 205634 151688 205640 151700
rect 154540 151660 205640 151688
rect 154540 151648 154546 151660
rect 205634 151648 205640 151660
rect 205692 151648 205698 151700
rect 238662 151648 238668 151700
rect 238720 151688 238726 151700
rect 289814 151688 289820 151700
rect 238720 151660 289820 151688
rect 238720 151648 238726 151660
rect 289814 151648 289820 151660
rect 289872 151648 289878 151700
rect 293862 151648 293868 151700
rect 293920 151688 293926 151700
rect 345014 151688 345020 151700
rect 293920 151660 345020 151688
rect 293920 151648 293926 151660
rect 345014 151648 345020 151660
rect 345072 151648 345078 151700
rect 378042 151648 378048 151700
rect 378100 151688 378106 151700
rect 429286 151688 429292 151700
rect 378100 151660 429292 151688
rect 378100 151648 378106 151660
rect 429286 151648 429292 151660
rect 429344 151648 429350 151700
rect 434622 151648 434628 151700
rect 434680 151688 434686 151700
rect 485774 151688 485780 151700
rect 434680 151660 485780 151688
rect 434680 151648 434686 151660
rect 485774 151648 485780 151660
rect 485832 151648 485838 151700
rect 518802 151648 518808 151700
rect 518860 151688 518866 151700
rect 569954 151688 569960 151700
rect 518860 151660 569960 151688
rect 518860 151648 518866 151660
rect 569954 151648 569960 151660
rect 570012 151648 570018 151700
rect 182082 151580 182088 151632
rect 182140 151620 182146 151632
rect 233234 151620 233240 151632
rect 182140 151592 233240 151620
rect 182140 151580 182146 151592
rect 233234 151580 233240 151592
rect 233292 151580 233298 151632
rect 350442 151580 350448 151632
rect 350500 151620 350506 151632
rect 401594 151620 401600 151632
rect 350500 151592 401600 151620
rect 350500 151580 350506 151592
rect 401594 151580 401600 151592
rect 401652 151580 401658 151632
rect 462222 151580 462228 151632
rect 462280 151620 462286 151632
rect 513374 151620 513380 151632
rect 462280 151592 513380 151620
rect 462280 151580 462286 151592
rect 513374 151580 513380 151592
rect 513432 151580 513438 151632
rect 15194 148996 15200 149048
rect 15252 149036 15258 149048
rect 35894 149036 35900 149048
rect 15252 149008 35900 149036
rect 15252 148996 15258 149008
rect 35894 148996 35900 149008
rect 35952 148996 35958 149048
rect 36078 148996 36084 149048
rect 36136 149036 36142 149048
rect 63586 149036 63592 149048
rect 36136 149008 63592 149036
rect 36136 148996 36142 149008
rect 63586 148996 63592 149008
rect 63644 148996 63650 149048
rect 65794 148996 65800 149048
rect 65852 149036 65858 149048
rect 91922 149036 91928 149048
rect 65852 149008 91928 149036
rect 65852 148996 65858 149008
rect 91922 148996 91928 149008
rect 91980 148996 91986 149048
rect 92106 148996 92112 149048
rect 92164 149036 92170 149048
rect 119614 149036 119620 149048
rect 92164 149008 119620 149036
rect 92164 148996 92170 149008
rect 119614 148996 119620 149008
rect 119672 148996 119678 149048
rect 122098 148996 122104 149048
rect 122156 149036 122162 149048
rect 147950 149036 147956 149048
rect 122156 149008 147956 149036
rect 122156 148996 122162 149008
rect 147950 148996 147956 149008
rect 148008 148996 148014 149048
rect 148042 148996 148048 149048
rect 148100 149036 148106 149048
rect 175918 149036 175924 149048
rect 148100 149008 175924 149036
rect 148100 148996 148106 149008
rect 175918 148996 175924 149008
rect 175976 148996 175982 149048
rect 176102 148996 176108 149048
rect 176160 149036 176166 149048
rect 203610 149036 203616 149048
rect 176160 149008 203616 149036
rect 176160 148996 176166 149008
rect 203610 148996 203616 149008
rect 203668 148996 203674 149048
rect 204990 148996 204996 149048
rect 205048 149036 205054 149048
rect 231946 149036 231952 149048
rect 205048 149008 231952 149036
rect 205048 148996 205054 149008
rect 231946 148996 231952 149008
rect 232004 148996 232010 149048
rect 232038 148996 232044 149048
rect 232096 149036 232102 149048
rect 259914 149036 259920 149048
rect 232096 149008 259920 149036
rect 232096 148996 232102 149008
rect 259914 148996 259920 149008
rect 259972 148996 259978 149048
rect 260098 148996 260104 149048
rect 260156 149036 260162 149048
rect 287606 149036 287612 149048
rect 260156 149008 287612 149036
rect 260156 148996 260162 149008
rect 287606 148996 287612 149008
rect 287664 148996 287670 149048
rect 288066 148996 288072 149048
rect 288124 149036 288130 149048
rect 315942 149036 315948 149048
rect 288124 149008 315948 149036
rect 288124 148996 288130 149008
rect 315942 148996 315948 149008
rect 316000 148996 316006 149048
rect 316678 148996 316684 149048
rect 316736 149036 316742 149048
rect 343910 149036 343916 149048
rect 316736 149008 343916 149036
rect 316736 148996 316742 149008
rect 343910 148996 343916 149008
rect 343968 148996 343974 149048
rect 344094 148996 344100 149048
rect 344152 149036 344158 149048
rect 371602 149036 371608 149048
rect 344152 149008 371608 149036
rect 344152 148996 344158 149008
rect 371602 148996 371608 149008
rect 371660 148996 371666 149048
rect 372062 148996 372068 149048
rect 372120 149036 372126 149048
rect 399938 149036 399944 149048
rect 372120 149008 399944 149036
rect 372120 148996 372126 149008
rect 399938 148996 399944 149008
rect 399996 148996 400002 149048
rect 400858 148996 400864 149048
rect 400916 149036 400922 149048
rect 427906 149036 427912 149048
rect 400916 149008 427912 149036
rect 400916 148996 400922 149008
rect 427906 148996 427912 149008
rect 427964 148996 427970 149048
rect 428090 148996 428096 149048
rect 428148 149036 428154 149048
rect 455598 149036 455604 149048
rect 428148 149008 455604 149036
rect 428148 148996 428154 149008
rect 455598 148996 455604 149008
rect 455656 148996 455662 149048
rect 456058 148996 456064 149048
rect 456116 149036 456122 149048
rect 483934 149036 483940 149048
rect 456116 149008 483940 149036
rect 456116 148996 456122 149008
rect 483934 148996 483940 149008
rect 483992 148996 483998 149048
rect 484026 148996 484032 149048
rect 484084 149036 484090 149048
rect 511902 149036 511908 149048
rect 484084 149008 511908 149036
rect 484084 148996 484090 149008
rect 511902 148996 511908 149008
rect 511960 148996 511966 149048
rect 512086 148996 512092 149048
rect 512144 149036 512150 149048
rect 539594 149036 539600 149048
rect 512144 149008 539600 149036
rect 512144 148996 512150 149008
rect 539594 148996 539600 149008
rect 539652 148996 539658 149048
rect 540054 148996 540060 149048
rect 540112 149036 540118 149048
rect 567930 149036 567936 149048
rect 540112 149008 567936 149036
rect 540112 148996 540118 149008
rect 567930 148996 567936 149008
rect 567988 148996 567994 149048
rect 16574 148928 16580 148980
rect 16632 148968 16638 148980
rect 36630 148968 36636 148980
rect 16632 148940 36636 148968
rect 16632 148928 16638 148940
rect 36630 148928 36636 148940
rect 36688 148928 36694 148980
rect 44910 148928 44916 148980
rect 44968 148968 44974 148980
rect 71130 148968 71136 148980
rect 44968 148940 71136 148968
rect 44968 148928 44974 148940
rect 71130 148928 71136 148940
rect 71188 148928 71194 148980
rect 82262 148928 82268 148980
rect 82320 148968 82326 148980
rect 93118 148968 93124 148980
rect 82320 148940 93124 148968
rect 82320 148928 82326 148940
rect 93118 148928 93124 148940
rect 93176 148928 93182 148980
rect 110230 148928 110236 148980
rect 110288 148968 110294 148980
rect 124858 148968 124864 148980
rect 110288 148940 124864 148968
rect 110288 148928 110294 148940
rect 124858 148928 124864 148940
rect 124916 148928 124922 148980
rect 128630 148928 128636 148980
rect 128688 148968 128694 148980
rect 151078 148968 151084 148980
rect 128688 148940 151084 148968
rect 128688 148928 128694 148940
rect 151078 148928 151084 148940
rect 151136 148928 151142 148980
rect 156598 148928 156604 148980
rect 156656 148968 156662 148980
rect 182818 148968 182824 148980
rect 156656 148940 182824 148968
rect 156656 148928 156662 148940
rect 182818 148928 182824 148940
rect 182876 148928 182882 148980
rect 194502 148928 194508 148980
rect 194560 148968 194566 148980
rect 210418 148968 210424 148980
rect 194560 148940 210424 148968
rect 194560 148928 194566 148940
rect 210418 148928 210424 148940
rect 210476 148928 210482 148980
rect 212626 148928 212632 148980
rect 212684 148968 212690 148980
rect 232498 148968 232504 148980
rect 212684 148940 232504 148968
rect 212684 148928 212690 148940
rect 232498 148928 232504 148940
rect 232556 148928 232562 148980
rect 240594 148928 240600 148980
rect 240652 148968 240658 148980
rect 266998 148968 267004 148980
rect 240652 148940 267004 148968
rect 240652 148928 240658 148940
rect 266998 148928 267004 148940
rect 267056 148928 267062 148980
rect 278590 148928 278596 148980
rect 278648 148968 278654 148980
rect 289078 148968 289084 148980
rect 278648 148940 289084 148968
rect 278648 148928 278654 148940
rect 289078 148928 289084 148940
rect 289136 148928 289142 148980
rect 306282 148928 306288 148980
rect 306340 148968 306346 148980
rect 318058 148968 318064 148980
rect 306340 148940 318064 148968
rect 306340 148928 306346 148940
rect 318058 148928 318064 148940
rect 318116 148928 318122 148980
rect 324590 148928 324596 148980
rect 324648 148968 324654 148980
rect 345658 148968 345664 148980
rect 324648 148940 345664 148968
rect 324648 148928 324654 148940
rect 345658 148928 345664 148940
rect 345716 148928 345722 148980
rect 362586 148928 362592 148980
rect 362644 148968 362650 148980
rect 373258 148968 373264 148980
rect 362644 148940 373264 148968
rect 362644 148928 362650 148940
rect 373258 148928 373264 148940
rect 373316 148928 373322 148980
rect 390278 148928 390284 148980
rect 390336 148968 390342 148980
rect 400950 148968 400956 148980
rect 390336 148940 400956 148968
rect 390336 148928 390342 148940
rect 400950 148928 400956 148940
rect 401008 148928 401014 148980
rect 408586 148928 408592 148980
rect 408644 148968 408650 148980
rect 428458 148968 428464 148980
rect 408644 148940 428464 148968
rect 408644 148928 408650 148940
rect 428458 148928 428464 148940
rect 428516 148928 428522 148980
rect 436922 148928 436928 148980
rect 436980 148968 436986 148980
rect 462958 148968 462964 148980
rect 436980 148940 462964 148968
rect 436980 148928 436986 148940
rect 462958 148928 462964 148940
rect 463016 148928 463022 148980
rect 474274 148928 474280 148980
rect 474332 148968 474338 148980
rect 485038 148968 485044 148980
rect 474332 148940 485044 148968
rect 474332 148928 474338 148940
rect 485038 148928 485044 148940
rect 485096 148928 485102 148980
rect 502242 148928 502248 148980
rect 502300 148968 502306 148980
rect 514018 148968 514024 148980
rect 502300 148940 514024 148968
rect 502300 148928 502306 148940
rect 514018 148928 514024 148940
rect 514076 148928 514082 148980
rect 520918 148928 520924 148980
rect 520976 148968 520982 148980
rect 541618 148968 541624 148980
rect 520976 148940 541624 148968
rect 520976 148928 520982 148940
rect 541618 148928 541624 148940
rect 541676 148928 541682 148980
rect 26234 148860 26240 148912
rect 26292 148900 26298 148912
rect 39298 148900 39304 148912
rect 26292 148872 39304 148900
rect 26292 148860 26298 148872
rect 39298 148860 39304 148872
rect 39356 148860 39362 148912
rect 54570 148860 54576 148912
rect 54628 148900 54634 148912
rect 66898 148900 66904 148912
rect 54628 148872 66904 148900
rect 54628 148860 54634 148872
rect 66898 148860 66904 148872
rect 66956 148860 66962 148912
rect 138290 148860 138296 148912
rect 138348 148900 138354 148912
rect 152458 148900 152464 148912
rect 138348 148872 152464 148900
rect 138348 148860 138354 148872
rect 152458 148860 152464 148872
rect 152516 148860 152522 148912
rect 166258 148860 166264 148912
rect 166316 148900 166322 148912
rect 177298 148900 177304 148912
rect 166316 148872 177304 148900
rect 166316 148860 166322 148872
rect 177298 148860 177304 148872
rect 177356 148860 177362 148912
rect 222286 148860 222292 148912
rect 222344 148900 222350 148912
rect 233970 148900 233976 148912
rect 222344 148872 233976 148900
rect 222344 148860 222350 148872
rect 233970 148860 233976 148872
rect 234028 148860 234034 148912
rect 250254 148860 250260 148912
rect 250312 148900 250318 148912
rect 261478 148900 261484 148912
rect 250312 148872 261484 148900
rect 250312 148860 250318 148872
rect 261478 148860 261484 148872
rect 261536 148860 261542 148912
rect 334250 148860 334256 148912
rect 334308 148900 334314 148912
rect 347038 148900 347044 148912
rect 334308 148872 347044 148900
rect 334308 148860 334314 148872
rect 347038 148860 347044 148872
rect 347096 148860 347102 148912
rect 418246 148860 418252 148912
rect 418304 148900 418310 148912
rect 429838 148900 429844 148912
rect 418304 148872 429844 148900
rect 418304 148860 418310 148872
rect 429838 148860 429844 148872
rect 429896 148860 429902 148912
rect 446582 148860 446588 148912
rect 446640 148900 446646 148912
rect 457438 148900 457444 148912
rect 446640 148872 457444 148900
rect 446640 148860 446646 148872
rect 457438 148860 457444 148872
rect 457496 148860 457502 148912
rect 530578 148860 530584 148912
rect 530636 148900 530642 148912
rect 544378 148900 544384 148912
rect 530636 148872 544384 148900
rect 530636 148860 530642 148872
rect 544378 148860 544384 148872
rect 544436 148860 544442 148912
rect 558270 148316 558276 148368
rect 558328 148356 558334 148368
rect 567470 148356 567476 148368
rect 558328 148328 567476 148356
rect 558328 148316 558334 148328
rect 567470 148316 567476 148328
rect 567528 148316 567534 148368
rect 548334 146888 548340 146940
rect 548392 146928 548398 146940
rect 568114 146928 568120 146940
rect 548392 146900 568120 146928
rect 548392 146888 548398 146900
rect 568114 146888 568120 146900
rect 568172 146888 568178 146940
rect 212350 146480 212356 146532
rect 212408 146520 212414 146532
rect 232682 146520 232688 146532
rect 212408 146492 232688 146520
rect 212408 146480 212414 146492
rect 232682 146480 232688 146492
rect 232740 146480 232746 146532
rect 296346 146480 296352 146532
rect 296404 146520 296410 146532
rect 316770 146520 316776 146532
rect 296404 146492 316776 146520
rect 296404 146480 296410 146492
rect 316770 146480 316776 146492
rect 316828 146480 316834 146532
rect 408034 146480 408040 146532
rect 408092 146520 408098 146532
rect 428642 146520 428648 146532
rect 408092 146492 428648 146520
rect 408092 146480 408098 146492
rect 428642 146480 428648 146492
rect 428700 146480 428706 146532
rect 492030 146480 492036 146532
rect 492088 146520 492094 146532
rect 512730 146520 512736 146532
rect 492088 146492 512736 146520
rect 492088 146480 492094 146492
rect 512730 146480 512736 146492
rect 512788 146480 512794 146532
rect 148318 146412 148324 146464
rect 148376 146452 148382 146464
rect 165706 146452 165712 146464
rect 148376 146424 165712 146452
rect 148376 146412 148382 146424
rect 165706 146412 165712 146424
rect 165764 146412 165770 146464
rect 175458 146412 175464 146464
rect 175516 146452 175522 146464
rect 193674 146452 193680 146464
rect 175516 146424 193680 146452
rect 175516 146412 175522 146424
rect 193674 146412 193680 146424
rect 193732 146412 193738 146464
rect 203518 146412 203524 146464
rect 203576 146452 203582 146464
rect 221366 146452 221372 146464
rect 203576 146424 221372 146452
rect 203576 146412 203582 146424
rect 221366 146412 221372 146424
rect 221424 146412 221430 146464
rect 260190 146412 260196 146464
rect 260248 146452 260254 146464
rect 277670 146452 277676 146464
rect 260248 146424 277676 146452
rect 260248 146412 260254 146424
rect 277670 146412 277676 146424
rect 277728 146412 277734 146464
rect 287514 146412 287520 146464
rect 287572 146452 287578 146464
rect 305362 146452 305368 146464
rect 287572 146424 305368 146452
rect 287572 146412 287578 146424
rect 305362 146412 305368 146424
rect 305420 146412 305426 146464
rect 345658 146412 345664 146464
rect 345716 146452 345722 146464
rect 361666 146452 361672 146464
rect 345716 146424 361672 146452
rect 345716 146412 345722 146424
rect 361666 146412 361672 146424
rect 361724 146412 361730 146464
rect 371510 146412 371516 146464
rect 371568 146452 371574 146464
rect 389358 146452 389364 146464
rect 371568 146424 389364 146452
rect 371568 146412 371574 146424
rect 389358 146412 389364 146424
rect 389416 146412 389422 146464
rect 399478 146412 399484 146464
rect 399536 146452 399542 146464
rect 417694 146452 417700 146464
rect 399536 146424 417700 146452
rect 399536 146412 399542 146424
rect 417694 146412 417700 146424
rect 417752 146412 417758 146464
rect 456150 146412 456156 146464
rect 456208 146452 456214 146464
rect 473354 146452 473360 146464
rect 456208 146424 473360 146452
rect 456208 146412 456214 146424
rect 473354 146412 473360 146424
rect 473412 146412 473418 146464
rect 483474 146412 483480 146464
rect 483532 146452 483538 146464
rect 501690 146452 501696 146464
rect 483532 146424 501696 146452
rect 483532 146412 483538 146424
rect 501690 146412 501696 146424
rect 501748 146412 501754 146464
rect 36630 146344 36636 146396
rect 36688 146384 36694 146396
rect 53650 146384 53656 146396
rect 36688 146356 53656 146384
rect 36688 146344 36694 146356
rect 53650 146344 53656 146356
rect 53708 146344 53714 146396
rect 64414 146344 64420 146396
rect 64472 146384 64478 146396
rect 81434 146384 81440 146396
rect 64472 146356 81440 146384
rect 64472 146344 64478 146356
rect 81434 146344 81440 146356
rect 81492 146344 81498 146396
rect 91462 146344 91468 146396
rect 91520 146384 91526 146396
rect 109678 146384 109684 146396
rect 91520 146356 109684 146384
rect 91520 146344 91526 146356
rect 109678 146344 109684 146356
rect 109736 146344 109742 146396
rect 119430 146344 119436 146396
rect 119488 146384 119494 146396
rect 137646 146384 137652 146396
rect 119488 146356 137652 146384
rect 119488 146344 119494 146356
rect 137646 146344 137652 146356
rect 137704 146344 137710 146396
rect 156322 146344 156328 146396
rect 156380 146384 156386 146396
rect 178678 146384 178684 146396
rect 156380 146356 178684 146384
rect 156380 146344 156386 146356
rect 178678 146344 178684 146356
rect 178736 146344 178742 146396
rect 232498 146344 232504 146396
rect 232556 146384 232562 146396
rect 249702 146384 249708 146396
rect 232556 146356 249708 146384
rect 232556 146344 232562 146356
rect 249702 146344 249708 146356
rect 249760 146344 249766 146396
rect 268010 146344 268016 146396
rect 268068 146384 268074 146396
rect 287698 146384 287704 146396
rect 268068 146356 287704 146384
rect 268068 146344 268074 146356
rect 287698 146344 287704 146356
rect 287756 146344 287762 146396
rect 315482 146344 315488 146396
rect 315540 146384 315546 146396
rect 333698 146384 333704 146396
rect 315540 146356 333704 146384
rect 315540 146344 315546 146356
rect 333698 146344 333704 146356
rect 333756 146344 333762 146396
rect 352006 146344 352012 146396
rect 352064 146384 352070 146396
rect 374638 146384 374644 146396
rect 352064 146356 374644 146384
rect 352064 146344 352070 146356
rect 374638 146344 374644 146356
rect 374696 146344 374702 146396
rect 428458 146344 428464 146396
rect 428516 146384 428522 146396
rect 445662 146384 445668 146396
rect 428516 146356 445668 146384
rect 428516 146344 428522 146356
rect 445662 146344 445668 146356
rect 445720 146344 445726 146396
rect 464338 146344 464344 146396
rect 464396 146384 464402 146396
rect 483658 146384 483664 146396
rect 464396 146356 483664 146384
rect 464396 146344 464402 146356
rect 483658 146344 483664 146356
rect 483716 146344 483722 146396
rect 511442 146344 511448 146396
rect 511500 146384 511506 146396
rect 529658 146384 529664 146396
rect 511500 146356 529664 146384
rect 511500 146344 511506 146356
rect 529658 146344 529664 146356
rect 529716 146344 529722 146396
rect 541618 146344 541624 146396
rect 541676 146384 541682 146396
rect 557534 146384 557540 146396
rect 541676 146356 557540 146384
rect 541676 146344 541682 146356
rect 557534 146344 557540 146356
rect 557592 146344 557598 146396
rect 15102 146276 15108 146328
rect 15160 146316 15166 146328
rect 25682 146316 25688 146328
rect 15160 146288 25688 146316
rect 15160 146276 15166 146288
rect 25682 146276 25688 146288
rect 25740 146276 25746 146328
rect 36722 146276 36728 146328
rect 36780 146316 36786 146328
rect 63310 146316 63316 146328
rect 36780 146288 63316 146316
rect 36780 146276 36786 146288
rect 63310 146276 63316 146288
rect 63368 146276 63374 146328
rect 66898 146276 66904 146328
rect 66956 146316 66962 146328
rect 91094 146316 91100 146328
rect 66956 146288 91100 146316
rect 66956 146276 66962 146288
rect 91094 146276 91100 146288
rect 91152 146276 91158 146328
rect 93118 146276 93124 146328
rect 93176 146316 93182 146328
rect 119338 146316 119344 146328
rect 93176 146288 119344 146316
rect 93176 146276 93182 146288
rect 119338 146276 119344 146288
rect 119396 146276 119402 146328
rect 124858 146276 124864 146328
rect 124916 146316 124922 146328
rect 147306 146316 147312 146328
rect 124916 146288 147312 146316
rect 124916 146276 124922 146288
rect 147306 146276 147312 146288
rect 147364 146276 147370 146328
rect 148410 146276 148416 146328
rect 148468 146316 148474 146328
rect 175366 146316 175372 146328
rect 148468 146288 175372 146316
rect 148468 146276 148474 146288
rect 175366 146276 175372 146288
rect 175424 146276 175430 146328
rect 177298 146276 177304 146328
rect 177356 146316 177362 146328
rect 203334 146316 203340 146328
rect 177356 146288 203340 146316
rect 177356 146276 177362 146288
rect 203334 146276 203340 146288
rect 203392 146276 203398 146328
rect 204990 146276 204996 146328
rect 205048 146316 205054 146328
rect 231026 146316 231032 146328
rect 205048 146288 231032 146316
rect 205048 146276 205054 146288
rect 231026 146276 231032 146288
rect 231084 146276 231090 146328
rect 232590 146276 232596 146328
rect 232648 146316 232654 146328
rect 259362 146316 259368 146328
rect 232648 146288 259368 146316
rect 232648 146276 232654 146288
rect 259362 146276 259368 146288
rect 259420 146276 259426 146328
rect 260098 146276 260104 146328
rect 260156 146316 260162 146328
rect 287330 146316 287336 146328
rect 260156 146288 287336 146316
rect 260156 146276 260162 146288
rect 287330 146276 287336 146288
rect 287388 146276 287394 146328
rect 289078 146276 289084 146328
rect 289136 146316 289142 146328
rect 315022 146316 315028 146328
rect 289136 146288 315028 146316
rect 289136 146276 289142 146288
rect 315022 146276 315028 146288
rect 315080 146276 315086 146328
rect 316678 146276 316684 146328
rect 316736 146316 316742 146328
rect 343358 146316 343364 146328
rect 316736 146288 343364 146316
rect 316736 146276 316742 146288
rect 343358 146276 343364 146288
rect 343416 146276 343422 146328
rect 344278 146276 344284 146328
rect 344336 146316 344342 146328
rect 371326 146316 371332 146328
rect 344336 146288 371332 146316
rect 344336 146276 344342 146288
rect 371326 146276 371332 146288
rect 371384 146276 371390 146328
rect 373258 146276 373264 146328
rect 373316 146316 373322 146328
rect 399018 146316 399024 146328
rect 373316 146288 399024 146316
rect 373316 146276 373322 146288
rect 399018 146276 399024 146288
rect 399076 146276 399082 146328
rect 400858 146276 400864 146328
rect 400916 146316 400922 146328
rect 427354 146316 427360 146328
rect 400916 146288 427360 146316
rect 400916 146276 400922 146288
rect 427354 146276 427360 146288
rect 427412 146276 427418 146328
rect 428550 146276 428556 146328
rect 428608 146316 428614 146328
rect 455322 146316 455328 146328
rect 428608 146288 455328 146316
rect 428608 146276 428614 146288
rect 455322 146276 455328 146288
rect 455380 146276 455386 146328
rect 456058 146276 456064 146328
rect 456116 146316 456122 146328
rect 483014 146316 483020 146328
rect 456116 146288 483020 146316
rect 456116 146276 456122 146288
rect 483014 146276 483020 146288
rect 483072 146276 483078 146328
rect 485038 146276 485044 146328
rect 485096 146316 485102 146328
rect 511350 146316 511356 146328
rect 485096 146288 511356 146316
rect 485096 146276 485102 146288
rect 511350 146276 511356 146288
rect 511408 146276 511414 146328
rect 512638 146276 512644 146328
rect 512696 146316 512702 146328
rect 539318 146316 539324 146328
rect 512696 146288 539324 146316
rect 512696 146276 512702 146288
rect 539318 146276 539324 146288
rect 539376 146276 539382 146328
rect 540238 146276 540244 146328
rect 540296 146316 540302 146328
rect 567194 146316 567200 146328
rect 540296 146288 567200 146316
rect 540296 146276 540302 146288
rect 567194 146276 567200 146288
rect 567252 146276 567258 146328
rect 3326 136688 3332 136740
rect 3384 136728 3390 136740
rect 9030 136728 9036 136740
rect 3384 136700 9036 136728
rect 3384 136688 3390 136700
rect 9030 136688 9036 136700
rect 9088 136688 9094 136740
rect 42886 135464 42892 135516
rect 42944 135504 42950 135516
rect 43622 135504 43628 135516
rect 42944 135476 43628 135504
rect 42944 135464 42950 135476
rect 43622 135464 43628 135476
rect 43680 135464 43686 135516
rect 63586 128256 63592 128308
rect 63644 128296 63650 128308
rect 64414 128296 64420 128308
rect 63644 128268 64420 128296
rect 63644 128256 63650 128268
rect 64414 128256 64420 128268
rect 64472 128256 64478 128308
rect 259730 128256 259736 128308
rect 259788 128296 259794 128308
rect 260190 128296 260196 128308
rect 259788 128268 260196 128296
rect 259788 128256 259794 128268
rect 260190 128256 260196 128268
rect 260248 128256 260254 128308
rect 455690 128256 455696 128308
rect 455748 128296 455754 128308
rect 456150 128296 456156 128308
rect 455748 128268 456156 128296
rect 455748 128256 455754 128268
rect 456150 128256 456156 128268
rect 456208 128256 456214 128308
rect 232682 126896 232688 126948
rect 232740 126936 232746 126948
rect 239766 126936 239772 126948
rect 232740 126908 239772 126936
rect 232740 126896 232746 126908
rect 239766 126896 239772 126908
rect 239824 126896 239830 126948
rect 483658 126896 483664 126948
rect 483716 126936 483722 126948
rect 491662 126936 491668 126948
rect 483716 126908 491668 126936
rect 483716 126896 483722 126908
rect 491662 126896 491668 126908
rect 491720 126896 491726 126948
rect 512730 126896 512736 126948
rect 512788 126936 512794 126948
rect 519630 126936 519636 126948
rect 512788 126908 519636 126936
rect 512788 126896 512794 126908
rect 519630 126896 519636 126908
rect 519688 126896 519694 126948
rect 428642 126216 428648 126268
rect 428700 126256 428706 126268
rect 435726 126256 435732 126268
rect 428700 126228 435732 126256
rect 428700 126216 428706 126228
rect 435726 126216 435732 126228
rect 435784 126216 435790 126268
rect 287698 126080 287704 126132
rect 287756 126120 287762 126132
rect 295702 126120 295708 126132
rect 287756 126092 295708 126120
rect 287756 126080 287762 126092
rect 295702 126080 295708 126092
rect 295760 126080 295766 126132
rect 316770 126080 316776 126132
rect 316828 126120 316834 126132
rect 323670 126120 323676 126132
rect 316828 126092 323676 126120
rect 316828 126080 316834 126092
rect 323670 126080 323676 126092
rect 323728 126080 323734 126132
rect 13538 125536 13544 125588
rect 13596 125576 13602 125588
rect 66254 125576 66260 125588
rect 13596 125548 66260 125576
rect 13596 125536 13602 125548
rect 66254 125536 66260 125548
rect 66312 125536 66318 125588
rect 70302 125536 70308 125588
rect 70360 125576 70366 125588
rect 121454 125576 121460 125588
rect 70360 125548 121460 125576
rect 70360 125536 70366 125548
rect 121454 125536 121460 125548
rect 121512 125536 121518 125588
rect 126882 125536 126888 125588
rect 126940 125576 126946 125588
rect 178034 125576 178040 125588
rect 126940 125548 178040 125576
rect 126940 125536 126946 125548
rect 178034 125536 178040 125548
rect 178092 125536 178098 125588
rect 209682 125536 209688 125588
rect 209740 125576 209746 125588
rect 262214 125576 262220 125588
rect 209740 125548 262220 125576
rect 209740 125536 209746 125548
rect 262214 125536 262220 125548
rect 262272 125536 262278 125588
rect 266262 125536 266268 125588
rect 266320 125576 266326 125588
rect 317414 125576 317420 125588
rect 266320 125548 317420 125576
rect 266320 125536 266326 125548
rect 317414 125536 317420 125548
rect 317472 125536 317478 125588
rect 322842 125536 322848 125588
rect 322900 125576 322906 125588
rect 373994 125576 374000 125588
rect 322900 125548 374000 125576
rect 322900 125536 322906 125548
rect 373994 125536 374000 125548
rect 374052 125536 374058 125588
rect 405642 125536 405648 125588
rect 405700 125576 405706 125588
rect 458174 125576 458180 125588
rect 405700 125548 458180 125576
rect 405700 125536 405706 125548
rect 458174 125536 458180 125548
rect 458232 125536 458238 125588
rect 489822 125536 489828 125588
rect 489880 125576 489886 125588
rect 542354 125576 542360 125588
rect 489880 125548 542360 125576
rect 489880 125536 489886 125548
rect 542354 125536 542360 125548
rect 542412 125536 542418 125588
rect 42702 125468 42708 125520
rect 42760 125508 42766 125520
rect 93854 125508 93860 125520
rect 42760 125480 93860 125508
rect 42760 125468 42766 125480
rect 93854 125468 93860 125480
rect 93912 125468 93918 125520
rect 97902 125468 97908 125520
rect 97960 125508 97966 125520
rect 149054 125508 149060 125520
rect 97960 125480 149060 125508
rect 97960 125468 97966 125480
rect 149054 125468 149060 125480
rect 149112 125468 149118 125520
rect 154482 125468 154488 125520
rect 154540 125508 154546 125520
rect 205634 125508 205640 125520
rect 154540 125480 205640 125508
rect 154540 125468 154546 125480
rect 205634 125468 205640 125480
rect 205692 125468 205698 125520
rect 238662 125468 238668 125520
rect 238720 125508 238726 125520
rect 289814 125508 289820 125520
rect 238720 125480 289820 125508
rect 238720 125468 238726 125480
rect 289814 125468 289820 125480
rect 289872 125468 289878 125520
rect 293862 125468 293868 125520
rect 293920 125508 293926 125520
rect 345014 125508 345020 125520
rect 293920 125480 345020 125508
rect 293920 125468 293926 125480
rect 345014 125468 345020 125480
rect 345072 125468 345078 125520
rect 378042 125468 378048 125520
rect 378100 125508 378106 125520
rect 429286 125508 429292 125520
rect 378100 125480 429292 125508
rect 378100 125468 378106 125480
rect 429286 125468 429292 125480
rect 429344 125468 429350 125520
rect 434622 125468 434628 125520
rect 434680 125508 434686 125520
rect 485774 125508 485780 125520
rect 434680 125480 485780 125508
rect 434680 125468 434686 125480
rect 485774 125468 485780 125480
rect 485832 125468 485838 125520
rect 518802 125468 518808 125520
rect 518860 125508 518866 125520
rect 569954 125508 569960 125520
rect 518860 125480 569960 125508
rect 518860 125468 518866 125480
rect 569954 125468 569960 125480
rect 570012 125468 570018 125520
rect 182082 125400 182088 125452
rect 182140 125440 182146 125452
rect 233234 125440 233240 125452
rect 182140 125412 233240 125440
rect 182140 125400 182146 125412
rect 233234 125400 233240 125412
rect 233292 125400 233298 125452
rect 350442 125400 350448 125452
rect 350500 125440 350506 125452
rect 401594 125440 401600 125452
rect 350500 125412 401600 125440
rect 350500 125400 350506 125412
rect 401594 125400 401600 125412
rect 401652 125400 401658 125452
rect 462222 125400 462228 125452
rect 462280 125440 462286 125452
rect 513374 125440 513380 125452
rect 462280 125412 513380 125440
rect 462280 125400 462286 125412
rect 513374 125400 513380 125412
rect 513432 125400 513438 125452
rect 343542 124788 343548 124840
rect 343600 124828 343606 124840
rect 345658 124828 345664 124840
rect 343600 124800 345664 124828
rect 343600 124788 343606 124800
rect 345658 124788 345664 124800
rect 345716 124788 345722 124840
rect 35250 124652 35256 124704
rect 35308 124692 35314 124704
rect 36630 124692 36636 124704
rect 35308 124664 36636 124692
rect 35308 124652 35314 124664
rect 36630 124652 36636 124664
rect 36688 124652 36694 124704
rect 547874 124652 547880 124704
rect 547932 124692 547938 124704
rect 548150 124692 548156 124704
rect 547932 124664 548156 124692
rect 547932 124652 547938 124664
rect 548150 124652 548156 124664
rect 548208 124652 548214 124704
rect 15102 124176 15108 124228
rect 15160 124216 15166 124228
rect 16574 124216 16580 124228
rect 15160 124188 16580 124216
rect 15160 124176 15166 124188
rect 16574 124176 16580 124188
rect 16632 124176 16638 124228
rect 71866 122748 71872 122800
rect 71924 122788 71930 122800
rect 100018 122788 100024 122800
rect 71924 122760 100024 122788
rect 71924 122748 71930 122760
rect 100018 122748 100024 122760
rect 100076 122748 100082 122800
rect 127986 122788 127992 122800
rect 103486 122760 127992 122788
rect 25682 122680 25688 122732
rect 25740 122720 25746 122732
rect 36722 122720 36728 122732
rect 25740 122692 36728 122720
rect 25740 122680 25746 122692
rect 36722 122680 36728 122692
rect 36780 122680 36786 122732
rect 42886 122680 42892 122732
rect 42944 122720 42950 122732
rect 42944 122692 45554 122720
rect 42944 122680 42950 122692
rect 15286 122612 15292 122664
rect 15344 122652 15350 122664
rect 43990 122652 43996 122664
rect 15344 122624 43996 122652
rect 15344 122612 15350 122624
rect 43990 122612 43996 122624
rect 44048 122612 44054 122664
rect 45526 122652 45554 122692
rect 53650 122680 53656 122732
rect 53708 122720 53714 122732
rect 66898 122720 66904 122732
rect 53708 122692 66904 122720
rect 53708 122680 53714 122692
rect 66898 122680 66904 122692
rect 66956 122680 66962 122732
rect 81986 122680 81992 122732
rect 82044 122720 82050 122732
rect 93118 122720 93124 122732
rect 82044 122692 93124 122720
rect 82044 122680 82050 122692
rect 93118 122680 93124 122692
rect 93176 122680 93182 122732
rect 99466 122680 99472 122732
rect 99524 122720 99530 122732
rect 103486 122720 103514 122760
rect 127986 122748 127992 122760
rect 128044 122748 128050 122800
rect 165982 122748 165988 122800
rect 166040 122788 166046 122800
rect 177298 122788 177304 122800
rect 166040 122760 177304 122788
rect 166040 122748 166046 122760
rect 177298 122748 177304 122760
rect 177356 122748 177362 122800
rect 178678 122748 178684 122800
rect 178736 122788 178742 122800
rect 184014 122788 184020 122800
rect 178736 122760 184020 122788
rect 178736 122748 178742 122760
rect 184014 122748 184020 122760
rect 184072 122748 184078 122800
rect 211706 122788 211712 122800
rect 190426 122760 211712 122788
rect 99524 122692 103514 122720
rect 99524 122680 99530 122692
rect 109678 122680 109684 122732
rect 109736 122720 109742 122732
rect 124858 122720 124864 122732
rect 109736 122692 124864 122720
rect 109736 122680 109742 122692
rect 124858 122680 124864 122692
rect 124916 122680 124922 122732
rect 137646 122680 137652 122732
rect 137704 122720 137710 122732
rect 148410 122720 148416 122732
rect 137704 122692 148416 122720
rect 137704 122680 137710 122692
rect 148410 122680 148416 122692
rect 148468 122680 148474 122732
rect 183646 122680 183652 122732
rect 183704 122720 183710 122732
rect 190426 122720 190454 122760
rect 211706 122748 211712 122760
rect 211764 122748 211770 122800
rect 231578 122748 231584 122800
rect 231636 122788 231642 122800
rect 232498 122788 232504 122800
rect 231636 122760 232504 122788
rect 231636 122748 231642 122760
rect 232498 122748 232504 122760
rect 232556 122748 232562 122800
rect 277670 122748 277676 122800
rect 277728 122788 277734 122800
rect 289078 122788 289084 122800
rect 277728 122760 289084 122788
rect 277728 122748 277734 122760
rect 289078 122748 289084 122760
rect 289136 122748 289142 122800
rect 306006 122748 306012 122800
rect 306064 122788 306070 122800
rect 316678 122788 316684 122800
rect 306064 122760 316684 122788
rect 306064 122748 306070 122760
rect 316678 122748 316684 122760
rect 316736 122748 316742 122800
rect 361666 122748 361672 122800
rect 361724 122788 361730 122800
rect 373258 122788 373264 122800
rect 361724 122760 373264 122788
rect 361724 122748 361730 122760
rect 373258 122748 373264 122760
rect 373316 122748 373322 122800
rect 379606 122748 379612 122800
rect 379664 122788 379670 122800
rect 408034 122788 408040 122800
rect 379664 122760 408040 122788
rect 379664 122748 379670 122760
rect 408034 122748 408040 122760
rect 408092 122748 408098 122800
rect 473998 122748 474004 122800
rect 474056 122788 474062 122800
rect 485038 122788 485044 122800
rect 474056 122760 485044 122788
rect 474056 122748 474062 122760
rect 485038 122748 485044 122760
rect 485096 122748 485102 122800
rect 501690 122748 501696 122800
rect 501748 122788 501754 122800
rect 512638 122788 512644 122800
rect 501748 122760 512644 122788
rect 501748 122748 501754 122760
rect 512638 122748 512644 122760
rect 512696 122748 512702 122800
rect 539318 122748 539324 122800
rect 539376 122788 539382 122800
rect 541618 122788 541624 122800
rect 539376 122760 541624 122788
rect 539376 122748 539382 122760
rect 541618 122748 541624 122760
rect 541676 122748 541682 122800
rect 548150 122748 548156 122800
rect 548208 122788 548214 122800
rect 557534 122788 557540 122800
rect 548208 122760 557540 122788
rect 548208 122748 548214 122760
rect 557534 122748 557540 122760
rect 557592 122748 557598 122800
rect 183704 122692 190454 122720
rect 183704 122680 183710 122692
rect 193674 122680 193680 122732
rect 193732 122720 193738 122732
rect 204990 122720 204996 122732
rect 193732 122692 204996 122720
rect 193732 122680 193738 122692
rect 204990 122680 204996 122692
rect 205048 122680 205054 122732
rect 221918 122680 221924 122732
rect 221976 122720 221982 122732
rect 232590 122720 232596 122732
rect 221976 122692 232596 122720
rect 221976 122680 221982 122692
rect 232590 122680 232596 122692
rect 232648 122680 232654 122732
rect 249702 122680 249708 122732
rect 249760 122720 249766 122732
rect 260098 122720 260104 122732
rect 249760 122692 260104 122720
rect 249760 122680 249766 122692
rect 260098 122680 260104 122692
rect 260156 122680 260162 122732
rect 333698 122680 333704 122732
rect 333756 122720 333762 122732
rect 344278 122720 344284 122732
rect 333756 122692 344284 122720
rect 333756 122680 333762 122692
rect 344278 122680 344284 122692
rect 344336 122680 344342 122732
rect 374638 122680 374644 122732
rect 374696 122720 374702 122732
rect 379698 122720 379704 122732
rect 374696 122692 379704 122720
rect 374696 122680 374702 122692
rect 379698 122680 379704 122692
rect 379756 122680 379762 122732
rect 390002 122680 390008 122732
rect 390060 122720 390066 122732
rect 400858 122720 400864 122732
rect 390060 122692 400864 122720
rect 390060 122680 390066 122692
rect 400858 122680 400864 122692
rect 400916 122680 400922 122732
rect 417694 122680 417700 122732
rect 417752 122720 417758 122732
rect 428550 122720 428556 122732
rect 417752 122692 428556 122720
rect 417752 122680 417758 122692
rect 428550 122680 428556 122692
rect 428608 122680 428614 122732
rect 445662 122680 445668 122732
rect 445720 122720 445726 122732
rect 456058 122720 456064 122732
rect 445720 122692 456064 122720
rect 445720 122680 445726 122692
rect 456058 122680 456064 122692
rect 456116 122680 456122 122732
rect 529658 122680 529664 122732
rect 529716 122720 529722 122732
rect 540238 122720 540244 122732
rect 529716 122692 540244 122720
rect 529716 122680 529722 122692
rect 540238 122680 540244 122692
rect 540296 122680 540302 122732
rect 71958 122652 71964 122664
rect 45526 122624 71964 122652
rect 71958 122612 71964 122624
rect 72016 122612 72022 122664
rect 127066 122612 127072 122664
rect 127124 122652 127130 122664
rect 155954 122652 155960 122664
rect 127124 122624 155960 122652
rect 127124 122612 127130 122624
rect 155954 122612 155960 122624
rect 156012 122612 156018 122664
rect 238846 122612 238852 122664
rect 238904 122652 238910 122664
rect 268010 122652 268016 122664
rect 238904 122624 268016 122652
rect 238904 122612 238910 122624
rect 268010 122612 268016 122624
rect 268068 122612 268074 122664
rect 323026 122612 323032 122664
rect 323084 122652 323090 122664
rect 352006 122652 352012 122664
rect 323084 122624 352012 122652
rect 323084 122612 323090 122624
rect 352006 122612 352012 122624
rect 352064 122612 352070 122664
rect 434806 122612 434812 122664
rect 434864 122652 434870 122664
rect 463786 122652 463792 122664
rect 434864 122624 463792 122652
rect 434864 122612 434870 122624
rect 463786 122612 463792 122624
rect 463844 122612 463850 122664
rect 518986 122612 518992 122664
rect 519044 122652 519050 122664
rect 547874 122652 547880 122664
rect 519044 122624 547880 122652
rect 519044 122612 519050 122624
rect 547874 122612 547880 122624
rect 547932 122612 547938 122664
rect 489886 118884 499574 118912
rect 71130 118804 71136 118856
rect 71188 118844 71194 118856
rect 82262 118844 82268 118856
rect 71188 118816 82268 118844
rect 71188 118804 71194 118816
rect 82262 118804 82268 118816
rect 82320 118804 82326 118856
rect 99466 118804 99472 118856
rect 99524 118844 99530 118856
rect 138290 118844 138296 118856
rect 99524 118816 138296 118844
rect 99524 118804 99530 118816
rect 138290 118804 138296 118816
rect 138348 118804 138354 118856
rect 183646 118804 183652 118856
rect 183704 118844 183710 118856
rect 222286 118844 222292 118856
rect 183704 118816 222292 118844
rect 183704 118804 183710 118816
rect 222286 118804 222292 118816
rect 222344 118804 222350 118856
rect 266998 118804 267004 118856
rect 267056 118844 267062 118856
rect 277946 118844 277952 118856
rect 267056 118816 277952 118844
rect 267056 118804 267062 118816
rect 277946 118804 277952 118816
rect 278004 118804 278010 118856
rect 295426 118804 295432 118856
rect 295484 118844 295490 118856
rect 334250 118844 334256 118856
rect 295484 118816 334256 118844
rect 295484 118804 295490 118816
rect 334250 118804 334256 118816
rect 334308 118804 334314 118856
rect 352006 118804 352012 118856
rect 352064 118844 352070 118856
rect 352064 118816 364334 118844
rect 352064 118804 352070 118816
rect 26234 118736 26240 118788
rect 26292 118776 26298 118788
rect 35434 118776 35440 118788
rect 26292 118748 35440 118776
rect 26292 118736 26298 118748
rect 35434 118736 35440 118748
rect 35492 118736 35498 118788
rect 36630 118736 36636 118788
rect 36688 118776 36694 118788
rect 53926 118776 53932 118788
rect 36688 118748 53932 118776
rect 36688 118736 36694 118748
rect 53926 118736 53932 118748
rect 53984 118736 53990 118788
rect 71866 118736 71872 118788
rect 71924 118776 71930 118788
rect 109954 118776 109960 118788
rect 71924 118748 109960 118776
rect 71924 118736 71930 118748
rect 109954 118736 109960 118748
rect 110012 118736 110018 118788
rect 120718 118736 120724 118788
rect 120776 118776 120782 118788
rect 128630 118776 128636 118788
rect 120776 118748 128636 118776
rect 120776 118736 120782 118748
rect 128630 118736 128636 118748
rect 128688 118736 128694 118788
rect 151078 118736 151084 118788
rect 151136 118776 151142 118788
rect 156598 118776 156604 118788
rect 151136 118748 156604 118776
rect 151136 118736 151142 118748
rect 156598 118736 156604 118748
rect 156656 118736 156662 118788
rect 182818 118736 182824 118788
rect 182876 118776 182882 118788
rect 193950 118776 193956 118788
rect 182876 118748 193956 118776
rect 182876 118736 182882 118748
rect 193950 118736 193956 118748
rect 194008 118736 194014 118788
rect 232498 118736 232504 118788
rect 232556 118776 232562 118788
rect 232556 118748 248414 118776
rect 232556 118736 232562 118748
rect 39298 118668 39304 118720
rect 39356 118708 39362 118720
rect 44266 118708 44272 118720
rect 39356 118680 44272 118708
rect 39356 118668 39362 118680
rect 44266 118668 44272 118680
rect 44324 118668 44330 118720
rect 66898 118668 66904 118720
rect 66956 118708 66962 118720
rect 72602 118708 72608 118720
rect 66956 118680 72608 118708
rect 66956 118668 66962 118680
rect 72602 118668 72608 118680
rect 72660 118668 72666 118720
rect 93118 118668 93124 118720
rect 93176 118708 93182 118720
rect 100294 118708 100300 118720
rect 93176 118680 100300 118708
rect 93176 118668 93182 118680
rect 100294 118668 100300 118680
rect 100352 118668 100358 118720
rect 148318 118668 148324 118720
rect 148376 118708 148382 118720
rect 166258 118708 166264 118720
rect 148376 118680 166264 118708
rect 148376 118668 148382 118680
rect 166258 118668 166264 118680
rect 166316 118668 166322 118720
rect 177298 118668 177304 118720
rect 177356 118708 177362 118720
rect 184290 118708 184296 118720
rect 177356 118680 184296 118708
rect 177356 118668 177362 118680
rect 184290 118668 184296 118680
rect 184348 118668 184354 118720
rect 233970 118668 233976 118720
rect 234028 118708 234034 118720
rect 240594 118708 240600 118720
rect 234028 118680 240600 118708
rect 234028 118668 234034 118680
rect 240594 118668 240600 118680
rect 240652 118668 240658 118720
rect 248386 118708 248414 118748
rect 267826 118736 267832 118788
rect 267884 118776 267890 118788
rect 306282 118776 306288 118788
rect 267884 118748 306288 118776
rect 267884 118736 267890 118748
rect 306282 118736 306288 118748
rect 306340 118736 306346 118788
rect 345658 118736 345664 118788
rect 345716 118776 345722 118788
rect 361942 118776 361948 118788
rect 345716 118748 361948 118776
rect 345716 118736 345722 118748
rect 361942 118736 361948 118748
rect 362000 118736 362006 118788
rect 364306 118776 364334 118816
rect 379606 118804 379612 118856
rect 379664 118844 379670 118856
rect 418246 118844 418252 118856
rect 379664 118816 418252 118844
rect 379664 118804 379670 118816
rect 418246 118804 418252 118816
rect 418304 118804 418310 118856
rect 463786 118804 463792 118856
rect 463844 118844 463850 118856
rect 463844 118816 470594 118844
rect 463844 118804 463850 118816
rect 390278 118776 390284 118788
rect 364306 118748 390284 118776
rect 390278 118736 390284 118748
rect 390336 118736 390342 118788
rect 400950 118736 400956 118788
rect 401008 118776 401014 118788
rect 408586 118776 408592 118788
rect 401008 118748 408592 118776
rect 401008 118736 401014 118748
rect 408586 118736 408592 118748
rect 408644 118736 408650 118788
rect 429838 118736 429844 118788
rect 429896 118776 429902 118788
rect 436278 118776 436284 118788
rect 429896 118748 436284 118776
rect 429896 118736 429902 118748
rect 436278 118736 436284 118748
rect 436336 118736 436342 118788
rect 457438 118736 457444 118788
rect 457496 118776 457502 118788
rect 464614 118776 464620 118788
rect 457496 118748 464620 118776
rect 457496 118736 457502 118748
rect 464614 118736 464620 118748
rect 464672 118736 464678 118788
rect 470566 118776 470594 118816
rect 489886 118776 489914 118884
rect 491386 118804 491392 118856
rect 491444 118844 491450 118856
rect 491444 118816 492812 118844
rect 491444 118804 491450 118816
rect 470566 118748 489914 118776
rect 250254 118708 250260 118720
rect 248386 118680 250260 118708
rect 250254 118668 250260 118680
rect 250312 118668 250318 118720
rect 261478 118668 261484 118720
rect 261536 118708 261542 118720
rect 268286 118708 268292 118720
rect 261536 118680 268292 118708
rect 261536 118668 261542 118680
rect 268286 118668 268292 118680
rect 268344 118668 268350 118720
rect 289078 118668 289084 118720
rect 289136 118708 289142 118720
rect 296622 118708 296628 118720
rect 289136 118680 296628 118708
rect 289136 118668 289142 118680
rect 296622 118668 296628 118680
rect 296680 118668 296686 118720
rect 318058 118668 318064 118720
rect 318116 118708 318122 118720
rect 324590 118708 324596 118720
rect 318116 118680 324596 118708
rect 318116 118668 318122 118680
rect 324590 118668 324596 118680
rect 324648 118668 324654 118720
rect 347038 118668 347044 118720
rect 347096 118708 347102 118720
rect 352282 118708 352288 118720
rect 347096 118680 352288 118708
rect 347096 118668 347102 118680
rect 352282 118668 352288 118680
rect 352340 118668 352346 118720
rect 373258 118668 373264 118720
rect 373316 118708 373322 118720
rect 380618 118708 380624 118720
rect 373316 118680 380624 118708
rect 373316 118668 373322 118680
rect 380618 118668 380624 118680
rect 380676 118668 380682 118720
rect 428458 118668 428464 118720
rect 428516 118708 428522 118720
rect 445938 118708 445944 118720
rect 428516 118680 445944 118708
rect 428516 118668 428522 118680
rect 445938 118668 445944 118680
rect 445996 118668 446002 118720
rect 462958 118668 462964 118720
rect 463016 118708 463022 118720
rect 474274 118708 474280 118720
rect 463016 118680 474280 118708
rect 463016 118668 463022 118680
rect 474274 118668 474280 118680
rect 474332 118668 474338 118720
rect 485038 118668 485044 118720
rect 485096 118708 485102 118720
rect 492582 118708 492588 118720
rect 485096 118680 492588 118708
rect 485096 118668 485102 118680
rect 492582 118668 492588 118680
rect 492640 118668 492646 118720
rect 492784 118708 492812 118816
rect 499546 118776 499574 118884
rect 541618 118804 541624 118856
rect 541676 118844 541682 118856
rect 541676 118816 547874 118844
rect 541676 118804 541682 118816
rect 502242 118776 502248 118788
rect 499546 118748 502248 118776
rect 502242 118736 502248 118748
rect 502300 118736 502306 118788
rect 514018 118736 514024 118788
rect 514076 118776 514082 118788
rect 520274 118776 520280 118788
rect 514076 118748 520280 118776
rect 514076 118736 514082 118748
rect 520274 118736 520280 118748
rect 520332 118736 520338 118788
rect 547846 118776 547874 118816
rect 558270 118776 558276 118788
rect 547846 118748 558276 118776
rect 558270 118736 558276 118748
rect 558328 118736 558334 118788
rect 529934 118708 529940 118720
rect 492784 118680 529940 118708
rect 529934 118668 529940 118680
rect 529992 118668 529998 118720
rect 544378 118668 544384 118720
rect 544436 118708 544442 118720
rect 548610 118708 548616 118720
rect 544436 118680 548616 118708
rect 544436 118668 544442 118680
rect 548610 118668 548616 118680
rect 548668 118668 548674 118720
rect 567930 118708 567936 118720
rect 548720 118680 567936 118708
rect 547966 118600 547972 118652
rect 548024 118640 548030 118652
rect 548720 118640 548748 118680
rect 567930 118668 567936 118680
rect 567988 118668 567994 118720
rect 548024 118612 548748 118640
rect 548024 118600 548030 118612
rect 63770 116288 63776 116340
rect 63828 116328 63834 116340
rect 65794 116328 65800 116340
rect 63828 116300 65800 116328
rect 63828 116288 63834 116300
rect 65794 116288 65800 116300
rect 65852 116288 65858 116340
rect 120074 116288 120080 116340
rect 120132 116328 120138 116340
rect 122098 116328 122104 116340
rect 120132 116300 122104 116328
rect 120132 116288 120138 116300
rect 122098 116288 122104 116300
rect 122156 116288 122162 116340
rect 210418 116288 210424 116340
rect 210476 116328 210482 116340
rect 212350 116328 212356 116340
rect 210476 116300 212356 116328
rect 210476 116288 210482 116300
rect 212350 116288 212356 116300
rect 212408 116288 212414 116340
rect 204254 114724 204260 114776
rect 204312 114764 204318 114776
rect 204990 114764 204996 114776
rect 204312 114736 204996 114764
rect 204312 114724 204318 114736
rect 204990 114724 204996 114736
rect 205048 114724 205054 114776
rect 13538 97928 13544 97980
rect 13596 97968 13602 97980
rect 66254 97968 66260 97980
rect 13596 97940 66260 97968
rect 13596 97928 13602 97940
rect 66254 97928 66260 97940
rect 66312 97928 66318 97980
rect 97902 97928 97908 97980
rect 97960 97968 97966 97980
rect 149054 97968 149060 97980
rect 97960 97940 149060 97968
rect 97960 97928 97966 97940
rect 149054 97928 149060 97940
rect 149112 97928 149118 97980
rect 154482 97928 154488 97980
rect 154540 97968 154546 97980
rect 205634 97968 205640 97980
rect 154540 97940 205640 97968
rect 154540 97928 154546 97940
rect 205634 97928 205640 97940
rect 205692 97928 205698 97980
rect 209682 97928 209688 97980
rect 209740 97968 209746 97980
rect 262214 97968 262220 97980
rect 209740 97940 262220 97968
rect 209740 97928 209746 97940
rect 262214 97928 262220 97940
rect 262272 97928 262278 97980
rect 266262 97928 266268 97980
rect 266320 97968 266326 97980
rect 317414 97968 317420 97980
rect 266320 97940 317420 97968
rect 266320 97928 266326 97940
rect 317414 97928 317420 97940
rect 317472 97928 317478 97980
rect 322842 97928 322848 97980
rect 322900 97968 322906 97980
rect 373994 97968 374000 97980
rect 322900 97940 374000 97968
rect 322900 97928 322906 97940
rect 373994 97928 374000 97940
rect 374052 97928 374058 97980
rect 405642 97928 405648 97980
rect 405700 97968 405706 97980
rect 458174 97968 458180 97980
rect 405700 97940 458180 97968
rect 405700 97928 405706 97940
rect 458174 97928 458180 97940
rect 458232 97928 458238 97980
rect 489822 97928 489828 97980
rect 489880 97968 489886 97980
rect 542354 97968 542360 97980
rect 489880 97940 542360 97968
rect 489880 97928 489886 97940
rect 542354 97928 542360 97940
rect 542412 97928 542418 97980
rect 70302 97860 70308 97912
rect 70360 97900 70366 97912
rect 121454 97900 121460 97912
rect 70360 97872 121460 97900
rect 70360 97860 70366 97872
rect 121454 97860 121460 97872
rect 121512 97860 121518 97912
rect 126882 97860 126888 97912
rect 126940 97900 126946 97912
rect 178034 97900 178040 97912
rect 126940 97872 178040 97900
rect 126940 97860 126946 97872
rect 178034 97860 178040 97872
rect 178092 97860 178098 97912
rect 182082 97860 182088 97912
rect 182140 97900 182146 97912
rect 233234 97900 233240 97912
rect 182140 97872 233240 97900
rect 182140 97860 182146 97872
rect 233234 97860 233240 97872
rect 233292 97860 233298 97912
rect 238662 97860 238668 97912
rect 238720 97900 238726 97912
rect 289814 97900 289820 97912
rect 238720 97872 289820 97900
rect 238720 97860 238726 97872
rect 289814 97860 289820 97872
rect 289872 97860 289878 97912
rect 293862 97860 293868 97912
rect 293920 97900 293926 97912
rect 345014 97900 345020 97912
rect 293920 97872 345020 97900
rect 293920 97860 293926 97872
rect 345014 97860 345020 97872
rect 345072 97860 345078 97912
rect 378042 97860 378048 97912
rect 378100 97900 378106 97912
rect 429286 97900 429292 97912
rect 378100 97872 429292 97900
rect 378100 97860 378106 97872
rect 429286 97860 429292 97872
rect 429344 97860 429350 97912
rect 434622 97860 434628 97912
rect 434680 97900 434686 97912
rect 485774 97900 485780 97912
rect 434680 97872 485780 97900
rect 434680 97860 434686 97872
rect 485774 97860 485780 97872
rect 485832 97860 485838 97912
rect 518802 97860 518808 97912
rect 518860 97900 518866 97912
rect 569954 97900 569960 97912
rect 518860 97872 569960 97900
rect 518860 97860 518866 97872
rect 569954 97860 569960 97872
rect 570012 97860 570018 97912
rect 42702 97792 42708 97844
rect 42760 97832 42766 97844
rect 93854 97832 93860 97844
rect 42760 97804 93860 97832
rect 42760 97792 42766 97804
rect 93854 97792 93860 97804
rect 93912 97792 93918 97844
rect 350442 97792 350448 97844
rect 350500 97832 350506 97844
rect 401594 97832 401600 97844
rect 350500 97804 401600 97832
rect 350500 97792 350506 97804
rect 401594 97792 401600 97804
rect 401652 97792 401658 97844
rect 462222 97792 462228 97844
rect 462280 97832 462286 97844
rect 513374 97832 513380 97844
rect 462280 97804 513380 97832
rect 462280 97792 462286 97804
rect 513374 97792 513380 97804
rect 513432 97792 513438 97844
rect 547874 95412 547880 95464
rect 547932 95452 547938 95464
rect 548334 95452 548340 95464
rect 547932 95424 548340 95452
rect 547932 95412 547938 95424
rect 548334 95412 548340 95424
rect 548392 95412 548398 95464
rect 15194 95140 15200 95192
rect 15252 95180 15258 95192
rect 35894 95180 35900 95192
rect 15252 95152 35900 95180
rect 15252 95140 15258 95152
rect 35894 95140 35900 95152
rect 35952 95140 35958 95192
rect 36078 95140 36084 95192
rect 36136 95180 36142 95192
rect 63586 95180 63592 95192
rect 36136 95152 63592 95180
rect 36136 95140 36142 95152
rect 63586 95140 63592 95152
rect 63644 95140 63650 95192
rect 65794 95140 65800 95192
rect 65852 95180 65858 95192
rect 91922 95180 91928 95192
rect 65852 95152 91928 95180
rect 65852 95140 65858 95152
rect 91922 95140 91928 95152
rect 91980 95140 91986 95192
rect 92106 95140 92112 95192
rect 92164 95180 92170 95192
rect 119614 95180 119620 95192
rect 92164 95152 119620 95180
rect 92164 95140 92170 95152
rect 119614 95140 119620 95152
rect 119672 95140 119678 95192
rect 122098 95140 122104 95192
rect 122156 95180 122162 95192
rect 147950 95180 147956 95192
rect 122156 95152 147956 95180
rect 122156 95140 122162 95152
rect 147950 95140 147956 95152
rect 148008 95140 148014 95192
rect 148042 95140 148048 95192
rect 148100 95180 148106 95192
rect 175918 95180 175924 95192
rect 148100 95152 175924 95180
rect 148100 95140 148106 95152
rect 175918 95140 175924 95152
rect 175976 95140 175982 95192
rect 176102 95140 176108 95192
rect 176160 95180 176166 95192
rect 203610 95180 203616 95192
rect 176160 95152 203616 95180
rect 176160 95140 176166 95152
rect 203610 95140 203616 95152
rect 203668 95140 203674 95192
rect 204990 95140 204996 95192
rect 205048 95180 205054 95192
rect 231946 95180 231952 95192
rect 205048 95152 231952 95180
rect 205048 95140 205054 95152
rect 231946 95140 231952 95152
rect 232004 95140 232010 95192
rect 232038 95140 232044 95192
rect 232096 95180 232102 95192
rect 259914 95180 259920 95192
rect 232096 95152 259920 95180
rect 232096 95140 232102 95152
rect 259914 95140 259920 95152
rect 259972 95140 259978 95192
rect 260098 95140 260104 95192
rect 260156 95180 260162 95192
rect 287606 95180 287612 95192
rect 260156 95152 287612 95180
rect 260156 95140 260162 95152
rect 287606 95140 287612 95152
rect 287664 95140 287670 95192
rect 288066 95140 288072 95192
rect 288124 95180 288130 95192
rect 315942 95180 315948 95192
rect 288124 95152 315948 95180
rect 288124 95140 288130 95152
rect 315942 95140 315948 95152
rect 316000 95140 316006 95192
rect 316678 95140 316684 95192
rect 316736 95180 316742 95192
rect 343910 95180 343916 95192
rect 316736 95152 343916 95180
rect 316736 95140 316742 95152
rect 343910 95140 343916 95152
rect 343968 95140 343974 95192
rect 344094 95140 344100 95192
rect 344152 95180 344158 95192
rect 371602 95180 371608 95192
rect 344152 95152 371608 95180
rect 344152 95140 344158 95152
rect 371602 95140 371608 95152
rect 371660 95140 371666 95192
rect 372062 95140 372068 95192
rect 372120 95180 372126 95192
rect 399938 95180 399944 95192
rect 372120 95152 399944 95180
rect 372120 95140 372126 95152
rect 399938 95140 399944 95152
rect 399996 95140 400002 95192
rect 400858 95140 400864 95192
rect 400916 95180 400922 95192
rect 427906 95180 427912 95192
rect 400916 95152 427912 95180
rect 400916 95140 400922 95152
rect 427906 95140 427912 95152
rect 427964 95140 427970 95192
rect 428090 95140 428096 95192
rect 428148 95180 428154 95192
rect 455598 95180 455604 95192
rect 428148 95152 455604 95180
rect 428148 95140 428154 95152
rect 455598 95140 455604 95152
rect 455656 95140 455662 95192
rect 456058 95140 456064 95192
rect 456116 95180 456122 95192
rect 483934 95180 483940 95192
rect 456116 95152 483940 95180
rect 456116 95140 456122 95152
rect 483934 95140 483940 95152
rect 483992 95140 483998 95192
rect 484026 95140 484032 95192
rect 484084 95180 484090 95192
rect 511902 95180 511908 95192
rect 484084 95152 511908 95180
rect 484084 95140 484090 95152
rect 511902 95140 511908 95152
rect 511960 95140 511966 95192
rect 512086 95140 512092 95192
rect 512144 95180 512150 95192
rect 539594 95180 539600 95192
rect 512144 95152 539600 95180
rect 512144 95140 512150 95152
rect 539594 95140 539600 95152
rect 539652 95140 539658 95192
rect 540054 95140 540060 95192
rect 540112 95180 540118 95192
rect 567930 95180 567936 95192
rect 540112 95152 567936 95180
rect 540112 95140 540118 95152
rect 567930 95140 567936 95152
rect 567988 95140 567994 95192
rect 16574 95072 16580 95124
rect 16632 95112 16638 95124
rect 36630 95112 36636 95124
rect 16632 95084 36636 95112
rect 16632 95072 16638 95084
rect 36630 95072 36636 95084
rect 36688 95072 36694 95124
rect 44910 95072 44916 95124
rect 44968 95112 44974 95124
rect 71130 95112 71136 95124
rect 44968 95084 71136 95112
rect 44968 95072 44974 95084
rect 71130 95072 71136 95084
rect 71188 95072 71194 95124
rect 82262 95072 82268 95124
rect 82320 95112 82326 95124
rect 93118 95112 93124 95124
rect 82320 95084 93124 95112
rect 82320 95072 82326 95084
rect 93118 95072 93124 95084
rect 93176 95072 93182 95124
rect 110230 95072 110236 95124
rect 110288 95112 110294 95124
rect 120718 95112 120724 95124
rect 110288 95084 120724 95112
rect 110288 95072 110294 95084
rect 120718 95072 120724 95084
rect 120776 95072 120782 95124
rect 128630 95072 128636 95124
rect 128688 95112 128694 95124
rect 148318 95112 148324 95124
rect 128688 95084 148324 95112
rect 128688 95072 128694 95084
rect 148318 95072 148324 95084
rect 148376 95072 148382 95124
rect 156598 95072 156604 95124
rect 156656 95112 156662 95124
rect 182818 95112 182824 95124
rect 156656 95084 182824 95112
rect 156656 95072 156662 95084
rect 182818 95072 182824 95084
rect 182876 95072 182882 95124
rect 194502 95072 194508 95124
rect 194560 95112 194566 95124
rect 210418 95112 210424 95124
rect 194560 95084 210424 95112
rect 194560 95072 194566 95084
rect 210418 95072 210424 95084
rect 210476 95072 210482 95124
rect 212626 95072 212632 95124
rect 212684 95112 212690 95124
rect 232498 95112 232504 95124
rect 212684 95084 232504 95112
rect 212684 95072 212690 95084
rect 232498 95072 232504 95084
rect 232556 95072 232562 95124
rect 240594 95072 240600 95124
rect 240652 95112 240658 95124
rect 266998 95112 267004 95124
rect 240652 95084 267004 95112
rect 240652 95072 240658 95084
rect 266998 95072 267004 95084
rect 267056 95072 267062 95124
rect 278590 95072 278596 95124
rect 278648 95112 278654 95124
rect 289078 95112 289084 95124
rect 278648 95084 289084 95112
rect 278648 95072 278654 95084
rect 289078 95072 289084 95084
rect 289136 95072 289142 95124
rect 306282 95072 306288 95124
rect 306340 95112 306346 95124
rect 318058 95112 318064 95124
rect 306340 95084 318064 95112
rect 306340 95072 306346 95084
rect 318058 95072 318064 95084
rect 318116 95072 318122 95124
rect 324590 95072 324596 95124
rect 324648 95112 324654 95124
rect 345658 95112 345664 95124
rect 324648 95084 345664 95112
rect 324648 95072 324654 95084
rect 345658 95072 345664 95084
rect 345716 95072 345722 95124
rect 362586 95072 362592 95124
rect 362644 95112 362650 95124
rect 373258 95112 373264 95124
rect 362644 95084 373264 95112
rect 362644 95072 362650 95084
rect 373258 95072 373264 95084
rect 373316 95072 373322 95124
rect 390278 95072 390284 95124
rect 390336 95112 390342 95124
rect 400950 95112 400956 95124
rect 390336 95084 400956 95112
rect 390336 95072 390342 95084
rect 400950 95072 400956 95084
rect 401008 95072 401014 95124
rect 408586 95072 408592 95124
rect 408644 95112 408650 95124
rect 428458 95112 428464 95124
rect 408644 95084 428464 95112
rect 408644 95072 408650 95084
rect 428458 95072 428464 95084
rect 428516 95072 428522 95124
rect 436922 95072 436928 95124
rect 436980 95112 436986 95124
rect 462958 95112 462964 95124
rect 436980 95084 462964 95112
rect 436980 95072 436986 95084
rect 462958 95072 462964 95084
rect 463016 95072 463022 95124
rect 474274 95072 474280 95124
rect 474332 95112 474338 95124
rect 485038 95112 485044 95124
rect 474332 95084 485044 95112
rect 474332 95072 474338 95084
rect 485038 95072 485044 95084
rect 485096 95072 485102 95124
rect 502242 95072 502248 95124
rect 502300 95112 502306 95124
rect 514018 95112 514024 95124
rect 502300 95084 514024 95112
rect 502300 95072 502306 95084
rect 514018 95072 514024 95084
rect 514076 95072 514082 95124
rect 520918 95072 520924 95124
rect 520976 95112 520982 95124
rect 541618 95112 541624 95124
rect 520976 95084 541624 95112
rect 520976 95072 520982 95084
rect 541618 95072 541624 95084
rect 541676 95072 541682 95124
rect 26234 95004 26240 95056
rect 26292 95044 26298 95056
rect 39298 95044 39304 95056
rect 26292 95016 39304 95044
rect 26292 95004 26298 95016
rect 39298 95004 39304 95016
rect 39356 95004 39362 95056
rect 54570 95004 54576 95056
rect 54628 95044 54634 95056
rect 66898 95044 66904 95056
rect 54628 95016 66904 95044
rect 54628 95004 54634 95016
rect 66898 95004 66904 95016
rect 66956 95004 66962 95056
rect 138290 95004 138296 95056
rect 138348 95044 138354 95056
rect 151078 95044 151084 95056
rect 138348 95016 151084 95044
rect 138348 95004 138354 95016
rect 151078 95004 151084 95016
rect 151136 95004 151142 95056
rect 166258 95004 166264 95056
rect 166316 95044 166322 95056
rect 177298 95044 177304 95056
rect 166316 95016 177304 95044
rect 166316 95004 166322 95016
rect 177298 95004 177304 95016
rect 177356 95004 177362 95056
rect 222286 95004 222292 95056
rect 222344 95044 222350 95056
rect 233970 95044 233976 95056
rect 222344 95016 233976 95044
rect 222344 95004 222350 95016
rect 233970 95004 233976 95016
rect 234028 95004 234034 95056
rect 250254 95004 250260 95056
rect 250312 95044 250318 95056
rect 261478 95044 261484 95056
rect 250312 95016 261484 95044
rect 250312 95004 250318 95016
rect 261478 95004 261484 95016
rect 261536 95004 261542 95056
rect 334250 95004 334256 95056
rect 334308 95044 334314 95056
rect 347038 95044 347044 95056
rect 334308 95016 347044 95044
rect 334308 95004 334314 95016
rect 347038 95004 347044 95016
rect 347096 95004 347102 95056
rect 418246 95004 418252 95056
rect 418304 95044 418310 95056
rect 429838 95044 429844 95056
rect 418304 95016 429844 95044
rect 418304 95004 418310 95016
rect 429838 95004 429844 95016
rect 429896 95004 429902 95056
rect 446582 95004 446588 95056
rect 446640 95044 446646 95056
rect 457438 95044 457444 95056
rect 446640 95016 457444 95044
rect 446640 95004 446646 95016
rect 457438 95004 457444 95016
rect 457496 95004 457502 95056
rect 530578 95004 530584 95056
rect 530636 95044 530642 95056
rect 544378 95044 544384 95056
rect 530636 95016 544384 95044
rect 530636 95004 530642 95016
rect 544378 95004 544384 95016
rect 544436 95004 544442 95056
rect 558270 94460 558276 94512
rect 558328 94500 558334 94512
rect 567470 94500 567476 94512
rect 558328 94472 567476 94500
rect 558328 94460 558334 94472
rect 567470 94460 567476 94472
rect 567528 94460 567534 94512
rect 408034 91264 408040 91316
rect 408092 91304 408098 91316
rect 428642 91304 428648 91316
rect 408092 91276 428648 91304
rect 408092 91264 408098 91276
rect 428642 91264 428648 91276
rect 428700 91264 428706 91316
rect 148410 91196 148416 91248
rect 148468 91236 148474 91248
rect 165706 91236 165712 91248
rect 148468 91208 165712 91236
rect 148468 91196 148474 91208
rect 165706 91196 165712 91208
rect 165764 91196 165770 91248
rect 175458 91196 175464 91248
rect 175516 91236 175522 91248
rect 193674 91236 193680 91248
rect 175516 91208 193680 91236
rect 175516 91196 175522 91208
rect 193674 91196 193680 91208
rect 193732 91196 193738 91248
rect 203518 91196 203524 91248
rect 203576 91236 203582 91248
rect 221366 91236 221372 91248
rect 203576 91208 221372 91236
rect 203576 91196 203582 91208
rect 221366 91196 221372 91208
rect 221424 91196 221430 91248
rect 232590 91196 232596 91248
rect 232648 91236 232654 91248
rect 249702 91236 249708 91248
rect 232648 91208 249708 91236
rect 232648 91196 232654 91208
rect 249702 91196 249708 91208
rect 249760 91196 249766 91248
rect 260190 91196 260196 91248
rect 260248 91236 260254 91248
rect 277670 91236 277676 91248
rect 260248 91208 277676 91236
rect 260248 91196 260254 91208
rect 277670 91196 277676 91208
rect 277728 91196 277734 91248
rect 287514 91196 287520 91248
rect 287572 91236 287578 91248
rect 305362 91236 305368 91248
rect 287572 91208 305368 91236
rect 287572 91196 287578 91208
rect 305362 91196 305368 91208
rect 305420 91196 305426 91248
rect 315482 91196 315488 91248
rect 315540 91236 315546 91248
rect 333698 91236 333704 91248
rect 315540 91208 333704 91236
rect 315540 91196 315546 91208
rect 333698 91196 333704 91208
rect 333756 91196 333762 91248
rect 345658 91196 345664 91248
rect 345716 91236 345722 91248
rect 361666 91236 361672 91248
rect 345716 91208 361672 91236
rect 345716 91196 345722 91208
rect 361666 91196 361672 91208
rect 361724 91196 361730 91248
rect 371510 91196 371516 91248
rect 371568 91236 371574 91248
rect 389358 91236 389364 91248
rect 371568 91208 389364 91236
rect 371568 91196 371574 91208
rect 389358 91196 389364 91208
rect 389416 91196 389422 91248
rect 399478 91196 399484 91248
rect 399536 91236 399542 91248
rect 417694 91236 417700 91248
rect 399536 91208 417700 91236
rect 399536 91196 399542 91208
rect 417694 91196 417700 91208
rect 417752 91196 417758 91248
rect 456150 91196 456156 91248
rect 456208 91236 456214 91248
rect 473354 91236 473360 91248
rect 456208 91208 473360 91236
rect 456208 91196 456214 91208
rect 473354 91196 473360 91208
rect 473412 91196 473418 91248
rect 483474 91196 483480 91248
rect 483532 91236 483538 91248
rect 501690 91236 501696 91248
rect 483532 91208 501696 91236
rect 483532 91196 483538 91208
rect 501690 91196 501696 91208
rect 501748 91196 501754 91248
rect 511442 91196 511448 91248
rect 511500 91236 511506 91248
rect 529658 91236 529664 91248
rect 511500 91208 529664 91236
rect 511500 91196 511506 91208
rect 529658 91196 529664 91208
rect 529716 91196 529722 91248
rect 36722 91128 36728 91180
rect 36780 91168 36786 91180
rect 53650 91168 53656 91180
rect 36780 91140 53656 91168
rect 36780 91128 36786 91140
rect 53650 91128 53656 91140
rect 53708 91128 53714 91180
rect 64414 91128 64420 91180
rect 64472 91168 64478 91180
rect 81434 91168 81440 91180
rect 64472 91140 81440 91168
rect 64472 91128 64478 91140
rect 81434 91128 81440 91140
rect 81492 91128 81498 91180
rect 91462 91128 91468 91180
rect 91520 91168 91526 91180
rect 109678 91168 109684 91180
rect 91520 91140 109684 91168
rect 91520 91128 91526 91140
rect 109678 91128 109684 91140
rect 109736 91128 109742 91180
rect 119430 91128 119436 91180
rect 119488 91168 119494 91180
rect 137646 91168 137652 91180
rect 119488 91140 137652 91168
rect 119488 91128 119494 91140
rect 137646 91128 137652 91140
rect 137704 91128 137710 91180
rect 156322 91128 156328 91180
rect 156380 91168 156386 91180
rect 178678 91168 178684 91180
rect 156380 91140 178684 91168
rect 156380 91128 156386 91140
rect 178678 91128 178684 91140
rect 178736 91128 178742 91180
rect 212350 91128 212356 91180
rect 212408 91168 212414 91180
rect 232682 91168 232688 91180
rect 212408 91140 232688 91168
rect 212408 91128 212414 91140
rect 232682 91128 232688 91140
rect 232740 91128 232746 91180
rect 268010 91128 268016 91180
rect 268068 91168 268074 91180
rect 287698 91168 287704 91180
rect 268068 91140 287704 91168
rect 268068 91128 268074 91140
rect 287698 91128 287704 91140
rect 287756 91128 287762 91180
rect 296346 91128 296352 91180
rect 296404 91168 296410 91180
rect 316770 91168 316776 91180
rect 296404 91140 316776 91168
rect 296404 91128 296410 91140
rect 316770 91128 316776 91140
rect 316828 91128 316834 91180
rect 352006 91128 352012 91180
rect 352064 91168 352070 91180
rect 374638 91168 374644 91180
rect 352064 91140 374644 91168
rect 352064 91128 352070 91140
rect 374638 91128 374644 91140
rect 374696 91128 374702 91180
rect 428458 91128 428464 91180
rect 428516 91168 428522 91180
rect 445662 91168 445668 91180
rect 428516 91140 445668 91168
rect 428516 91128 428522 91140
rect 445662 91128 445668 91140
rect 445720 91128 445726 91180
rect 464338 91128 464344 91180
rect 464396 91168 464402 91180
rect 483658 91168 483664 91180
rect 464396 91140 483664 91168
rect 464396 91128 464402 91140
rect 483658 91128 483664 91140
rect 483716 91128 483722 91180
rect 492030 91128 492036 91180
rect 492088 91168 492094 91180
rect 512730 91168 512736 91180
rect 492088 91140 512736 91168
rect 492088 91128 492094 91140
rect 512730 91128 512736 91140
rect 512788 91128 512794 91180
rect 541618 91128 541624 91180
rect 541676 91168 541682 91180
rect 557534 91168 557540 91180
rect 541676 91140 557540 91168
rect 541676 91128 541682 91140
rect 557534 91128 557540 91140
rect 557592 91128 557598 91180
rect 15102 91060 15108 91112
rect 15160 91100 15166 91112
rect 25682 91100 25688 91112
rect 15160 91072 25688 91100
rect 15160 91060 15166 91072
rect 25682 91060 25688 91072
rect 25740 91060 25746 91112
rect 36630 91060 36636 91112
rect 36688 91100 36694 91112
rect 63310 91100 63316 91112
rect 36688 91072 63316 91100
rect 36688 91060 36694 91072
rect 63310 91060 63316 91072
rect 63368 91060 63374 91112
rect 66898 91060 66904 91112
rect 66956 91100 66962 91112
rect 91094 91100 91100 91112
rect 66956 91072 91100 91100
rect 66956 91060 66962 91072
rect 91094 91060 91100 91072
rect 91152 91060 91158 91112
rect 93118 91060 93124 91112
rect 93176 91100 93182 91112
rect 119338 91100 119344 91112
rect 93176 91072 119344 91100
rect 93176 91060 93182 91072
rect 119338 91060 119344 91072
rect 119396 91060 119402 91112
rect 124858 91060 124864 91112
rect 124916 91100 124922 91112
rect 147306 91100 147312 91112
rect 124916 91072 147312 91100
rect 124916 91060 124922 91072
rect 147306 91060 147312 91072
rect 147364 91060 147370 91112
rect 148318 91060 148324 91112
rect 148376 91100 148382 91112
rect 175366 91100 175372 91112
rect 148376 91072 175372 91100
rect 148376 91060 148382 91072
rect 175366 91060 175372 91072
rect 175424 91060 175430 91112
rect 177298 91060 177304 91112
rect 177356 91100 177362 91112
rect 203334 91100 203340 91112
rect 177356 91072 203340 91100
rect 177356 91060 177362 91072
rect 203334 91060 203340 91072
rect 203392 91060 203398 91112
rect 204990 91060 204996 91112
rect 205048 91100 205054 91112
rect 231026 91100 231032 91112
rect 205048 91072 231032 91100
rect 205048 91060 205054 91072
rect 231026 91060 231032 91072
rect 231084 91060 231090 91112
rect 232498 91060 232504 91112
rect 232556 91100 232562 91112
rect 259362 91100 259368 91112
rect 232556 91072 259368 91100
rect 232556 91060 232562 91072
rect 259362 91060 259368 91072
rect 259420 91060 259426 91112
rect 260098 91060 260104 91112
rect 260156 91100 260162 91112
rect 287330 91100 287336 91112
rect 260156 91072 287336 91100
rect 260156 91060 260162 91072
rect 287330 91060 287336 91072
rect 287388 91060 287394 91112
rect 289078 91060 289084 91112
rect 289136 91100 289142 91112
rect 315022 91100 315028 91112
rect 289136 91072 315028 91100
rect 289136 91060 289142 91072
rect 315022 91060 315028 91072
rect 315080 91060 315086 91112
rect 316678 91060 316684 91112
rect 316736 91100 316742 91112
rect 343358 91100 343364 91112
rect 316736 91072 343364 91100
rect 316736 91060 316742 91072
rect 343358 91060 343364 91072
rect 343416 91060 343422 91112
rect 344278 91060 344284 91112
rect 344336 91100 344342 91112
rect 371326 91100 371332 91112
rect 344336 91072 371332 91100
rect 344336 91060 344342 91072
rect 371326 91060 371332 91072
rect 371384 91060 371390 91112
rect 373258 91060 373264 91112
rect 373316 91100 373322 91112
rect 399018 91100 399024 91112
rect 373316 91072 399024 91100
rect 373316 91060 373322 91072
rect 399018 91060 399024 91072
rect 399076 91060 399082 91112
rect 400858 91060 400864 91112
rect 400916 91100 400922 91112
rect 427354 91100 427360 91112
rect 400916 91072 427360 91100
rect 400916 91060 400922 91072
rect 427354 91060 427360 91072
rect 427412 91060 427418 91112
rect 428550 91060 428556 91112
rect 428608 91100 428614 91112
rect 455322 91100 455328 91112
rect 428608 91072 455328 91100
rect 428608 91060 428614 91072
rect 455322 91060 455328 91072
rect 455380 91060 455386 91112
rect 456058 91060 456064 91112
rect 456116 91100 456122 91112
rect 483014 91100 483020 91112
rect 456116 91072 483020 91100
rect 456116 91060 456122 91072
rect 483014 91060 483020 91072
rect 483072 91060 483078 91112
rect 485038 91060 485044 91112
rect 485096 91100 485102 91112
rect 511350 91100 511356 91112
rect 485096 91072 511356 91100
rect 485096 91060 485102 91072
rect 511350 91060 511356 91072
rect 511408 91060 511414 91112
rect 512638 91060 512644 91112
rect 512696 91100 512702 91112
rect 539318 91100 539324 91112
rect 512696 91072 539324 91100
rect 512696 91060 512702 91072
rect 539318 91060 539324 91072
rect 539376 91060 539382 91112
rect 540238 91060 540244 91112
rect 540296 91100 540302 91112
rect 567194 91100 567200 91112
rect 540296 91072 567200 91100
rect 540296 91060 540302 91072
rect 567194 91060 567200 91072
rect 567252 91060 567258 91112
rect 434622 88816 434628 88868
rect 434680 88856 434686 88868
rect 485774 88856 485780 88868
rect 434680 88828 485780 88856
rect 434680 88816 434686 88828
rect 485774 88816 485780 88828
rect 485832 88816 485838 88868
rect 405642 88748 405648 88800
rect 405700 88788 405706 88800
rect 458174 88788 458180 88800
rect 405700 88760 458180 88788
rect 405700 88748 405706 88760
rect 458174 88748 458180 88760
rect 458232 88748 458238 88800
rect 42702 88340 42708 88392
rect 42760 88380 42766 88392
rect 93854 88380 93860 88392
rect 42760 88352 93860 88380
rect 42760 88340 42766 88352
rect 93854 88340 93860 88352
rect 93912 88340 93918 88392
rect 97902 88340 97908 88392
rect 97960 88380 97966 88392
rect 149054 88380 149060 88392
rect 97960 88352 149060 88380
rect 97960 88340 97966 88352
rect 149054 88340 149060 88352
rect 149112 88340 149118 88392
rect 154482 88340 154488 88392
rect 154540 88380 154546 88392
rect 205634 88380 205640 88392
rect 154540 88352 205640 88380
rect 154540 88340 154546 88352
rect 205634 88340 205640 88352
rect 205692 88340 205698 88392
rect 209682 88340 209688 88392
rect 209740 88380 209746 88392
rect 262214 88380 262220 88392
rect 209740 88352 262220 88380
rect 209740 88340 209746 88352
rect 262214 88340 262220 88352
rect 262272 88340 262278 88392
rect 266262 88340 266268 88392
rect 266320 88380 266326 88392
rect 317414 88380 317420 88392
rect 266320 88352 317420 88380
rect 266320 88340 266326 88352
rect 317414 88340 317420 88352
rect 317472 88340 317478 88392
rect 322842 88340 322848 88392
rect 322900 88380 322906 88392
rect 373994 88380 374000 88392
rect 322900 88352 374000 88380
rect 322900 88340 322906 88352
rect 373994 88340 374000 88352
rect 374052 88340 374058 88392
rect 378042 88340 378048 88392
rect 378100 88380 378106 88392
rect 429286 88380 429292 88392
rect 378100 88352 429292 88380
rect 378100 88340 378106 88352
rect 429286 88340 429292 88352
rect 429344 88340 429350 88392
rect 489822 88340 489828 88392
rect 489880 88380 489886 88392
rect 542354 88380 542360 88392
rect 489880 88352 542360 88380
rect 489880 88340 489886 88352
rect 542354 88340 542360 88352
rect 542412 88340 542418 88392
rect 42886 85892 42892 85944
rect 42944 85932 42950 85944
rect 43622 85932 43628 85944
rect 42944 85904 43628 85932
rect 42944 85892 42950 85904
rect 43622 85892 43628 85904
rect 43680 85892 43686 85944
rect 3142 84192 3148 84244
rect 3200 84232 3206 84244
rect 14550 84232 14556 84244
rect 3200 84204 14556 84232
rect 3200 84192 3206 84204
rect 14550 84192 14556 84204
rect 14608 84192 14614 84244
rect 428642 72428 428648 72480
rect 428700 72468 428706 72480
rect 435726 72468 435732 72480
rect 428700 72440 435732 72468
rect 428700 72428 428706 72440
rect 435726 72428 435732 72440
rect 435784 72428 435790 72480
rect 63586 72292 63592 72344
rect 63644 72332 63650 72344
rect 64414 72332 64420 72344
rect 63644 72304 64420 72332
rect 63644 72292 63650 72304
rect 64414 72292 64420 72304
rect 64472 72292 64478 72344
rect 147674 72292 147680 72344
rect 147732 72332 147738 72344
rect 148410 72332 148416 72344
rect 147732 72304 148416 72332
rect 147732 72292 147738 72304
rect 148410 72292 148416 72304
rect 148468 72292 148474 72344
rect 232682 72292 232688 72344
rect 232740 72332 232746 72344
rect 239766 72332 239772 72344
rect 232740 72304 239772 72332
rect 232740 72292 232746 72304
rect 239766 72292 239772 72304
rect 239824 72292 239830 72344
rect 259730 72292 259736 72344
rect 259788 72332 259794 72344
rect 260190 72332 260196 72344
rect 259788 72304 260196 72332
rect 259788 72292 259794 72304
rect 260190 72292 260196 72304
rect 260248 72292 260254 72344
rect 316770 72292 316776 72344
rect 316828 72332 316834 72344
rect 323670 72332 323676 72344
rect 316828 72304 323676 72332
rect 316828 72292 316834 72304
rect 323670 72292 323676 72304
rect 323728 72292 323734 72344
rect 455690 72292 455696 72344
rect 455748 72332 455754 72344
rect 456150 72332 456156 72344
rect 455748 72304 456156 72332
rect 455748 72292 455754 72304
rect 456150 72292 456156 72304
rect 456208 72292 456214 72344
rect 483658 72224 483664 72276
rect 483716 72264 483722 72276
rect 491662 72264 491668 72276
rect 483716 72236 491668 72264
rect 483716 72224 483722 72236
rect 491662 72224 491668 72236
rect 491720 72224 491726 72276
rect 287698 72088 287704 72140
rect 287756 72128 287762 72140
rect 295702 72128 295708 72140
rect 287756 72100 295708 72128
rect 287756 72088 287762 72100
rect 295702 72088 295708 72100
rect 295760 72088 295766 72140
rect 512730 72088 512736 72140
rect 512788 72128 512794 72140
rect 519630 72128 519636 72140
rect 512788 72100 519636 72128
rect 512788 72088 512794 72100
rect 519630 72088 519636 72100
rect 519688 72088 519694 72140
rect 13538 71680 13544 71732
rect 13596 71720 13602 71732
rect 66254 71720 66260 71732
rect 13596 71692 66260 71720
rect 13596 71680 13602 71692
rect 66254 71680 66260 71692
rect 66312 71680 66318 71732
rect 70302 71680 70308 71732
rect 70360 71720 70366 71732
rect 121454 71720 121460 71732
rect 70360 71692 121460 71720
rect 70360 71680 70366 71692
rect 121454 71680 121460 71692
rect 121512 71680 121518 71732
rect 126882 71680 126888 71732
rect 126940 71720 126946 71732
rect 178034 71720 178040 71732
rect 126940 71692 178040 71720
rect 126940 71680 126946 71692
rect 178034 71680 178040 71692
rect 178092 71680 178098 71732
rect 182082 71680 182088 71732
rect 182140 71720 182146 71732
rect 233234 71720 233240 71732
rect 182140 71692 233240 71720
rect 182140 71680 182146 71692
rect 233234 71680 233240 71692
rect 233292 71680 233298 71732
rect 238662 71680 238668 71732
rect 238720 71720 238726 71732
rect 289814 71720 289820 71732
rect 238720 71692 289820 71720
rect 238720 71680 238726 71692
rect 289814 71680 289820 71692
rect 289872 71680 289878 71732
rect 293862 71680 293868 71732
rect 293920 71720 293926 71732
rect 345014 71720 345020 71732
rect 293920 71692 345020 71720
rect 293920 71680 293926 71692
rect 345014 71680 345020 71692
rect 345072 71680 345078 71732
rect 350442 71680 350448 71732
rect 350500 71720 350506 71732
rect 401594 71720 401600 71732
rect 350500 71692 401600 71720
rect 350500 71680 350506 71692
rect 401594 71680 401600 71692
rect 401652 71680 401658 71732
rect 462222 71680 462228 71732
rect 462280 71720 462286 71732
rect 513374 71720 513380 71732
rect 462280 71692 513380 71720
rect 462280 71680 462286 71692
rect 513374 71680 513380 71692
rect 513432 71680 513438 71732
rect 518802 71680 518808 71732
rect 518860 71720 518866 71732
rect 569954 71720 569960 71732
rect 518860 71692 569960 71720
rect 518860 71680 518866 71692
rect 569954 71680 569960 71692
rect 570012 71680 570018 71732
rect 231670 71612 231676 71664
rect 231728 71652 231734 71664
rect 232590 71652 232596 71664
rect 231728 71624 232596 71652
rect 231728 71612 231734 71624
rect 232590 71612 232596 71624
rect 232648 71612 232654 71664
rect 343542 71612 343548 71664
rect 343600 71652 343606 71664
rect 345658 71652 345664 71664
rect 343600 71624 345664 71652
rect 343600 71612 343606 71624
rect 345658 71612 345664 71624
rect 345716 71612 345722 71664
rect 539502 71612 539508 71664
rect 539560 71652 539566 71664
rect 541618 71652 541624 71664
rect 539560 71624 541624 71652
rect 539560 71612 539566 71624
rect 541618 71612 541624 71624
rect 541676 71612 541682 71664
rect 15102 70660 15108 70712
rect 15160 70700 15166 70712
rect 16574 70700 16580 70712
rect 15160 70672 16580 70700
rect 15160 70660 15166 70672
rect 16574 70660 16580 70672
rect 16632 70660 16638 70712
rect 35250 70660 35256 70712
rect 35308 70700 35314 70712
rect 36722 70700 36728 70712
rect 35308 70672 36728 70700
rect 35308 70660 35314 70672
rect 36722 70660 36728 70672
rect 36780 70660 36786 70712
rect 547874 70660 547880 70712
rect 547932 70700 547938 70712
rect 548150 70700 548156 70712
rect 547932 70672 548156 70700
rect 547932 70660 547938 70672
rect 548150 70660 548156 70672
rect 548208 70660 548214 70712
rect 71866 68960 71872 69012
rect 71924 69000 71930 69012
rect 100018 69000 100024 69012
rect 71924 68972 100024 69000
rect 71924 68960 71930 68972
rect 100018 68960 100024 68972
rect 100076 68960 100082 69012
rect 127986 69000 127992 69012
rect 103486 68972 127992 69000
rect 25682 68892 25688 68944
rect 25740 68932 25746 68944
rect 36630 68932 36636 68944
rect 25740 68904 36636 68932
rect 25740 68892 25746 68904
rect 36630 68892 36636 68904
rect 36688 68892 36694 68944
rect 42886 68892 42892 68944
rect 42944 68932 42950 68944
rect 42944 68904 45554 68932
rect 42944 68892 42950 68904
rect 15286 68824 15292 68876
rect 15344 68864 15350 68876
rect 43990 68864 43996 68876
rect 15344 68836 43996 68864
rect 15344 68824 15350 68836
rect 43990 68824 43996 68836
rect 44048 68824 44054 68876
rect 45526 68864 45554 68904
rect 53650 68892 53656 68944
rect 53708 68932 53714 68944
rect 66898 68932 66904 68944
rect 53708 68904 66904 68932
rect 53708 68892 53714 68904
rect 66898 68892 66904 68904
rect 66956 68892 66962 68944
rect 81986 68892 81992 68944
rect 82044 68932 82050 68944
rect 93118 68932 93124 68944
rect 82044 68904 93124 68932
rect 82044 68892 82050 68904
rect 93118 68892 93124 68904
rect 93176 68892 93182 68944
rect 99466 68892 99472 68944
rect 99524 68932 99530 68944
rect 103486 68932 103514 68972
rect 127986 68960 127992 68972
rect 128044 68960 128050 69012
rect 165982 68960 165988 69012
rect 166040 69000 166046 69012
rect 177298 69000 177304 69012
rect 166040 68972 177304 69000
rect 166040 68960 166046 68972
rect 177298 68960 177304 68972
rect 177356 68960 177362 69012
rect 178678 68960 178684 69012
rect 178736 69000 178742 69012
rect 184014 69000 184020 69012
rect 178736 68972 184020 69000
rect 178736 68960 178742 68972
rect 184014 68960 184020 68972
rect 184072 68960 184078 69012
rect 211706 69000 211712 69012
rect 190426 68972 211712 69000
rect 99524 68904 103514 68932
rect 99524 68892 99530 68904
rect 109678 68892 109684 68944
rect 109736 68932 109742 68944
rect 124858 68932 124864 68944
rect 109736 68904 124864 68932
rect 109736 68892 109742 68904
rect 124858 68892 124864 68904
rect 124916 68892 124922 68944
rect 137646 68892 137652 68944
rect 137704 68932 137710 68944
rect 148318 68932 148324 68944
rect 137704 68904 148324 68932
rect 137704 68892 137710 68904
rect 148318 68892 148324 68904
rect 148376 68892 148382 68944
rect 183646 68892 183652 68944
rect 183704 68932 183710 68944
rect 190426 68932 190454 68972
rect 211706 68960 211712 68972
rect 211764 68960 211770 69012
rect 222010 68960 222016 69012
rect 222068 69000 222074 69012
rect 232498 69000 232504 69012
rect 222068 68972 232504 69000
rect 222068 68960 222074 68972
rect 232498 68960 232504 68972
rect 232556 68960 232562 69012
rect 277670 68960 277676 69012
rect 277728 69000 277734 69012
rect 289078 69000 289084 69012
rect 277728 68972 289084 69000
rect 277728 68960 277734 68972
rect 289078 68960 289084 68972
rect 289136 68960 289142 69012
rect 306006 68960 306012 69012
rect 306064 69000 306070 69012
rect 316678 69000 316684 69012
rect 306064 68972 316684 69000
rect 306064 68960 306070 68972
rect 316678 68960 316684 68972
rect 316736 68960 316742 69012
rect 361666 68960 361672 69012
rect 361724 69000 361730 69012
rect 373258 69000 373264 69012
rect 361724 68972 373264 69000
rect 361724 68960 361730 68972
rect 373258 68960 373264 68972
rect 373316 68960 373322 69012
rect 379606 68960 379612 69012
rect 379664 69000 379670 69012
rect 408034 69000 408040 69012
rect 379664 68972 408040 69000
rect 379664 68960 379670 68972
rect 408034 68960 408040 68972
rect 408092 68960 408098 69012
rect 473998 68960 474004 69012
rect 474056 69000 474062 69012
rect 485038 69000 485044 69012
rect 474056 68972 485044 69000
rect 474056 68960 474062 68972
rect 485038 68960 485044 68972
rect 485096 68960 485102 69012
rect 501690 68960 501696 69012
rect 501748 69000 501754 69012
rect 512638 69000 512644 69012
rect 501748 68972 512644 69000
rect 501748 68960 501754 68972
rect 512638 68960 512644 68972
rect 512696 68960 512702 69012
rect 548150 68960 548156 69012
rect 548208 69000 548214 69012
rect 557534 69000 557540 69012
rect 548208 68972 557540 69000
rect 548208 68960 548214 68972
rect 557534 68960 557540 68972
rect 557592 68960 557598 69012
rect 183704 68904 190454 68932
rect 183704 68892 183710 68904
rect 193674 68892 193680 68944
rect 193732 68932 193738 68944
rect 204990 68932 204996 68944
rect 193732 68904 204996 68932
rect 193732 68892 193738 68904
rect 204990 68892 204996 68904
rect 205048 68892 205054 68944
rect 249702 68892 249708 68944
rect 249760 68932 249766 68944
rect 260098 68932 260104 68944
rect 249760 68904 260104 68932
rect 249760 68892 249766 68904
rect 260098 68892 260104 68904
rect 260156 68892 260162 68944
rect 333698 68892 333704 68944
rect 333756 68932 333762 68944
rect 344278 68932 344284 68944
rect 333756 68904 344284 68932
rect 333756 68892 333762 68904
rect 344278 68892 344284 68904
rect 344336 68892 344342 68944
rect 374638 68892 374644 68944
rect 374696 68932 374702 68944
rect 379698 68932 379704 68944
rect 374696 68904 379704 68932
rect 374696 68892 374702 68904
rect 379698 68892 379704 68904
rect 379756 68892 379762 68944
rect 390002 68892 390008 68944
rect 390060 68932 390066 68944
rect 400858 68932 400864 68944
rect 390060 68904 400864 68932
rect 390060 68892 390066 68904
rect 400858 68892 400864 68904
rect 400916 68892 400922 68944
rect 417694 68892 417700 68944
rect 417752 68932 417758 68944
rect 428550 68932 428556 68944
rect 417752 68904 428556 68932
rect 417752 68892 417758 68904
rect 428550 68892 428556 68904
rect 428608 68892 428614 68944
rect 445662 68892 445668 68944
rect 445720 68932 445726 68944
rect 456058 68932 456064 68944
rect 445720 68904 456064 68932
rect 445720 68892 445726 68904
rect 456058 68892 456064 68904
rect 456116 68892 456122 68944
rect 529658 68892 529664 68944
rect 529716 68932 529722 68944
rect 540238 68932 540244 68944
rect 529716 68904 540244 68932
rect 529716 68892 529722 68904
rect 540238 68892 540244 68904
rect 540296 68892 540302 68944
rect 72050 68864 72056 68876
rect 45526 68836 72056 68864
rect 72050 68824 72056 68836
rect 72108 68824 72114 68876
rect 127066 68824 127072 68876
rect 127124 68864 127130 68876
rect 156046 68864 156052 68876
rect 127124 68836 156052 68864
rect 127124 68824 127130 68836
rect 156046 68824 156052 68836
rect 156104 68824 156110 68876
rect 238846 68824 238852 68876
rect 238904 68864 238910 68876
rect 268010 68864 268016 68876
rect 238904 68836 268016 68864
rect 238904 68824 238910 68836
rect 268010 68824 268016 68836
rect 268068 68824 268074 68876
rect 323026 68824 323032 68876
rect 323084 68864 323090 68876
rect 352006 68864 352012 68876
rect 323084 68836 352012 68864
rect 323084 68824 323090 68836
rect 352006 68824 352012 68836
rect 352064 68824 352070 68876
rect 434806 68824 434812 68876
rect 434864 68864 434870 68876
rect 463694 68864 463700 68876
rect 434864 68836 463700 68864
rect 434864 68824 434870 68836
rect 463694 68824 463700 68836
rect 463752 68824 463758 68876
rect 518986 68824 518992 68876
rect 519044 68864 519050 68876
rect 547874 68864 547880 68876
rect 519044 68836 547880 68864
rect 519044 68824 519050 68836
rect 547874 68824 547880 68836
rect 547932 68824 547938 68876
rect 26234 65288 26240 65340
rect 26292 65328 26298 65340
rect 35434 65328 35440 65340
rect 26292 65300 35440 65328
rect 26292 65288 26298 65300
rect 35434 65288 35440 65300
rect 35492 65288 35498 65340
rect 71130 65016 71136 65068
rect 71188 65056 71194 65068
rect 82262 65056 82268 65068
rect 71188 65028 82268 65056
rect 71188 65016 71194 65028
rect 82262 65016 82268 65028
rect 82320 65016 82326 65068
rect 99374 65016 99380 65068
rect 99432 65056 99438 65068
rect 100294 65056 100300 65068
rect 99432 65028 100300 65056
rect 99432 65016 99438 65028
rect 100294 65016 100300 65028
rect 100352 65016 100358 65068
rect 183646 65016 183652 65068
rect 183704 65056 183710 65068
rect 222286 65056 222292 65068
rect 183704 65028 222292 65056
rect 183704 65016 183710 65028
rect 222286 65016 222292 65028
rect 222344 65016 222350 65068
rect 261478 65016 261484 65068
rect 261536 65056 261542 65068
rect 268286 65056 268292 65068
rect 261536 65028 268292 65056
rect 261536 65016 261542 65028
rect 268286 65016 268292 65028
rect 268344 65016 268350 65068
rect 295426 65016 295432 65068
rect 295484 65056 295490 65068
rect 334250 65056 334256 65068
rect 295484 65028 334256 65056
rect 295484 65016 295490 65028
rect 334250 65016 334256 65028
rect 334308 65016 334314 65068
rect 352006 65016 352012 65068
rect 352064 65056 352070 65068
rect 352064 65028 364334 65056
rect 352064 65016 352070 65028
rect 36630 64948 36636 65000
rect 36688 64988 36694 65000
rect 53926 64988 53932 65000
rect 36688 64960 53932 64988
rect 36688 64948 36694 64960
rect 53926 64948 53932 64960
rect 53984 64948 53990 65000
rect 71866 64948 71872 65000
rect 71924 64988 71930 65000
rect 109954 64988 109960 65000
rect 71924 64960 109960 64988
rect 71924 64948 71930 64960
rect 109954 64948 109960 64960
rect 110012 64948 110018 65000
rect 124858 64948 124864 65000
rect 124916 64988 124922 65000
rect 128630 64988 128636 65000
rect 124916 64960 128636 64988
rect 124916 64948 124922 64960
rect 128630 64948 128636 64960
rect 128688 64948 128694 65000
rect 152458 64948 152464 65000
rect 152516 64988 152522 65000
rect 156598 64988 156604 65000
rect 152516 64960 156604 64988
rect 152516 64948 152522 64960
rect 156598 64948 156604 64960
rect 156656 64948 156662 65000
rect 182818 64948 182824 65000
rect 182876 64988 182882 65000
rect 193950 64988 193956 65000
rect 182876 64960 193956 64988
rect 182876 64948 182882 64960
rect 193950 64948 193956 64960
rect 194008 64948 194014 65000
rect 232498 64948 232504 65000
rect 232556 64988 232562 65000
rect 232556 64960 248414 64988
rect 232556 64948 232562 64960
rect 39298 64880 39304 64932
rect 39356 64920 39362 64932
rect 44266 64920 44272 64932
rect 39356 64892 44272 64920
rect 39356 64880 39362 64892
rect 44266 64880 44272 64892
rect 44324 64880 44330 64932
rect 66898 64880 66904 64932
rect 66956 64920 66962 64932
rect 72602 64920 72608 64932
rect 66956 64892 72608 64920
rect 66956 64880 66962 64892
rect 72602 64880 72608 64892
rect 72660 64880 72666 64932
rect 93118 64880 93124 64932
rect 93176 64920 93182 64932
rect 99374 64920 99380 64932
rect 93176 64892 99380 64920
rect 93176 64880 93182 64892
rect 99374 64880 99380 64892
rect 99432 64880 99438 64932
rect 99466 64880 99472 64932
rect 99524 64920 99530 64932
rect 138290 64920 138296 64932
rect 99524 64892 138296 64920
rect 99524 64880 99530 64892
rect 138290 64880 138296 64892
rect 138348 64880 138354 64932
rect 151078 64880 151084 64932
rect 151136 64920 151142 64932
rect 166258 64920 166264 64932
rect 151136 64892 166264 64920
rect 151136 64880 151142 64892
rect 166258 64880 166264 64892
rect 166316 64880 166322 64932
rect 177298 64880 177304 64932
rect 177356 64920 177362 64932
rect 184290 64920 184296 64932
rect 177356 64892 184296 64920
rect 177356 64880 177362 64892
rect 184290 64880 184296 64892
rect 184348 64880 184354 64932
rect 210418 64880 210424 64932
rect 210476 64920 210482 64932
rect 212626 64920 212632 64932
rect 210476 64892 212632 64920
rect 210476 64880 210482 64892
rect 212626 64880 212632 64892
rect 212684 64880 212690 64932
rect 233970 64880 233976 64932
rect 234028 64920 234034 64932
rect 240594 64920 240600 64932
rect 234028 64892 240600 64920
rect 234028 64880 234034 64892
rect 240594 64880 240600 64892
rect 240652 64880 240658 64932
rect 248386 64920 248414 64960
rect 267826 64948 267832 65000
rect 267884 64988 267890 65000
rect 306282 64988 306288 65000
rect 267884 64960 306288 64988
rect 267884 64948 267890 64960
rect 306282 64948 306288 64960
rect 306340 64948 306346 65000
rect 345658 64948 345664 65000
rect 345716 64988 345722 65000
rect 361942 64988 361948 65000
rect 345716 64960 361948 64988
rect 345716 64948 345722 64960
rect 361942 64948 361948 64960
rect 362000 64948 362006 65000
rect 364306 64988 364334 65028
rect 379606 65016 379612 65068
rect 379664 65056 379670 65068
rect 418246 65056 418252 65068
rect 379664 65028 418252 65056
rect 379664 65016 379670 65028
rect 418246 65016 418252 65028
rect 418304 65016 418310 65068
rect 463786 65016 463792 65068
rect 463844 65056 463850 65068
rect 463844 65028 470594 65056
rect 463844 65016 463850 65028
rect 390278 64988 390284 65000
rect 364306 64960 390284 64988
rect 390278 64948 390284 64960
rect 390336 64948 390342 65000
rect 400858 64948 400864 65000
rect 400916 64988 400922 65000
rect 408586 64988 408592 65000
rect 400916 64960 408592 64988
rect 400916 64948 400922 64960
rect 408586 64948 408592 64960
rect 408644 64948 408650 65000
rect 429838 64948 429844 65000
rect 429896 64988 429902 65000
rect 436278 64988 436284 65000
rect 429896 64960 436284 64988
rect 429896 64948 429902 64960
rect 436278 64948 436284 64960
rect 436336 64948 436342 65000
rect 457438 64948 457444 65000
rect 457496 64988 457502 65000
rect 464614 64988 464620 65000
rect 457496 64960 464620 64988
rect 457496 64948 457502 64960
rect 464614 64948 464620 64960
rect 464672 64948 464678 65000
rect 470566 64988 470594 65028
rect 485038 65016 485044 65068
rect 485096 65056 485102 65068
rect 492582 65056 492588 65068
rect 485096 65028 492588 65056
rect 485096 65016 485102 65028
rect 492582 65016 492588 65028
rect 492640 65016 492646 65068
rect 502242 64988 502248 65000
rect 470566 64960 502248 64988
rect 502242 64948 502248 64960
rect 502300 64948 502306 65000
rect 514018 64948 514024 65000
rect 514076 64988 514082 65000
rect 520274 64988 520280 65000
rect 514076 64960 520280 64988
rect 514076 64948 514082 64960
rect 520274 64948 520280 64960
rect 520332 64948 520338 65000
rect 541618 64948 541624 65000
rect 541676 64988 541682 65000
rect 558270 64988 558276 65000
rect 541676 64960 558276 64988
rect 541676 64948 541682 64960
rect 558270 64948 558276 64960
rect 558328 64948 558334 65000
rect 250254 64920 250260 64932
rect 248386 64892 250260 64920
rect 250254 64880 250260 64892
rect 250312 64880 250318 64932
rect 266998 64880 267004 64932
rect 267056 64920 267062 64932
rect 277946 64920 277952 64932
rect 267056 64892 277952 64920
rect 267056 64880 267062 64892
rect 277946 64880 277952 64892
rect 278004 64880 278010 64932
rect 289078 64880 289084 64932
rect 289136 64920 289142 64932
rect 296622 64920 296628 64932
rect 289136 64892 296628 64920
rect 289136 64880 289142 64892
rect 296622 64880 296628 64892
rect 296680 64880 296686 64932
rect 318058 64880 318064 64932
rect 318116 64920 318122 64932
rect 324590 64920 324596 64932
rect 318116 64892 324596 64920
rect 318116 64880 318122 64892
rect 324590 64880 324596 64892
rect 324648 64880 324654 64932
rect 347038 64880 347044 64932
rect 347096 64920 347102 64932
rect 352282 64920 352288 64932
rect 347096 64892 352288 64920
rect 347096 64880 347102 64892
rect 352282 64880 352288 64892
rect 352340 64880 352346 64932
rect 373258 64880 373264 64932
rect 373316 64920 373322 64932
rect 380618 64920 380624 64932
rect 373316 64892 380624 64920
rect 373316 64880 373322 64892
rect 380618 64880 380624 64892
rect 380676 64880 380682 64932
rect 428458 64880 428464 64932
rect 428516 64920 428522 64932
rect 445938 64920 445944 64932
rect 428516 64892 445944 64920
rect 428516 64880 428522 64892
rect 445938 64880 445944 64892
rect 445996 64880 446002 64932
rect 462958 64880 462964 64932
rect 463016 64920 463022 64932
rect 474274 64920 474280 64932
rect 463016 64892 474280 64920
rect 463016 64880 463022 64892
rect 474274 64880 474280 64892
rect 474332 64880 474338 64932
rect 491386 64880 491392 64932
rect 491444 64920 491450 64932
rect 529934 64920 529940 64932
rect 491444 64892 529940 64920
rect 491444 64880 491450 64892
rect 529934 64880 529940 64892
rect 529992 64880 529998 64932
rect 547966 64880 547972 64932
rect 548024 64920 548030 64932
rect 567930 64920 567936 64932
rect 548024 64892 567936 64920
rect 548024 64880 548030 64892
rect 567930 64880 567936 64892
rect 567988 64880 567994 64932
rect 63770 62296 63776 62348
rect 63828 62336 63834 62348
rect 65794 62336 65800 62348
rect 63828 62308 65800 62336
rect 63828 62296 63834 62308
rect 65794 62296 65800 62308
rect 65852 62296 65858 62348
rect 120258 62160 120264 62212
rect 120316 62200 120322 62212
rect 122098 62200 122104 62212
rect 120316 62172 122104 62200
rect 120316 62160 120322 62172
rect 122098 62160 122104 62172
rect 122156 62160 122162 62212
rect 42702 62092 42708 62144
rect 42760 62132 42766 62144
rect 93854 62132 93860 62144
rect 42760 62104 93860 62132
rect 42760 62092 42766 62104
rect 93854 62092 93860 62104
rect 93912 62092 93918 62144
rect 97902 62092 97908 62144
rect 97960 62132 97966 62144
rect 149054 62132 149060 62144
rect 97960 62104 149060 62132
rect 97960 62092 97966 62104
rect 149054 62092 149060 62104
rect 149112 62092 149118 62144
rect 154482 62092 154488 62144
rect 154540 62132 154546 62144
rect 205634 62132 205640 62144
rect 154540 62104 205640 62132
rect 154540 62092 154546 62104
rect 205634 62092 205640 62104
rect 205692 62092 205698 62144
rect 209682 62092 209688 62144
rect 209740 62132 209746 62144
rect 262214 62132 262220 62144
rect 209740 62104 262220 62132
rect 209740 62092 209746 62104
rect 262214 62092 262220 62104
rect 262272 62092 262278 62144
rect 266262 62092 266268 62144
rect 266320 62132 266326 62144
rect 317414 62132 317420 62144
rect 266320 62104 317420 62132
rect 266320 62092 266326 62104
rect 317414 62092 317420 62104
rect 317472 62092 317478 62144
rect 322842 62092 322848 62144
rect 322900 62132 322906 62144
rect 373994 62132 374000 62144
rect 322900 62104 374000 62132
rect 322900 62092 322906 62104
rect 373994 62092 374000 62104
rect 374052 62092 374058 62144
rect 378042 62092 378048 62144
rect 378100 62132 378106 62144
rect 429286 62132 429292 62144
rect 378100 62104 429292 62132
rect 378100 62092 378106 62104
rect 429286 62092 429292 62104
rect 429344 62092 429350 62144
rect 434622 62092 434628 62144
rect 434680 62132 434686 62144
rect 485774 62132 485780 62144
rect 434680 62104 485780 62132
rect 434680 62092 434686 62104
rect 485774 62092 485780 62104
rect 485832 62092 485838 62144
rect 489822 62092 489828 62144
rect 489880 62132 489886 62144
rect 542354 62132 542360 62144
rect 489880 62104 542360 62132
rect 489880 62092 489886 62104
rect 542354 62092 542360 62104
rect 542412 62092 542418 62144
rect 544378 62092 544384 62144
rect 544436 62132 544442 62144
rect 548334 62132 548340 62144
rect 544436 62104 548340 62132
rect 544436 62092 544442 62104
rect 548334 62092 548340 62104
rect 548392 62092 548398 62144
rect 400306 58692 400312 58744
rect 400364 58732 400370 58744
rect 400950 58732 400956 58744
rect 400364 58704 400956 58732
rect 400364 58692 400370 58704
rect 400950 58692 400956 58704
rect 401008 58692 401014 58744
rect 204254 57876 204260 57928
rect 204312 57916 204318 57928
rect 204990 57916 204996 57928
rect 204312 57888 204996 57916
rect 204312 57876 204318 57888
rect 204990 57876 204996 57888
rect 205048 57876 205054 57928
rect 2958 44140 2964 44192
rect 3016 44180 3022 44192
rect 11882 44180 11888 44192
rect 3016 44152 11888 44180
rect 3016 44140 3022 44152
rect 11882 44140 11888 44152
rect 11940 44140 11946 44192
rect 13538 44072 13544 44124
rect 13596 44112 13602 44124
rect 66254 44112 66260 44124
rect 13596 44084 66260 44112
rect 13596 44072 13602 44084
rect 66254 44072 66260 44084
rect 66312 44072 66318 44124
rect 70302 44072 70308 44124
rect 70360 44112 70366 44124
rect 121454 44112 121460 44124
rect 70360 44084 121460 44112
rect 70360 44072 70366 44084
rect 121454 44072 121460 44084
rect 121512 44072 121518 44124
rect 126882 44072 126888 44124
rect 126940 44112 126946 44124
rect 178034 44112 178040 44124
rect 126940 44084 178040 44112
rect 126940 44072 126946 44084
rect 178034 44072 178040 44084
rect 178092 44072 178098 44124
rect 182082 44072 182088 44124
rect 182140 44112 182146 44124
rect 233234 44112 233240 44124
rect 182140 44084 233240 44112
rect 182140 44072 182146 44084
rect 233234 44072 233240 44084
rect 233292 44072 233298 44124
rect 238662 44072 238668 44124
rect 238720 44112 238726 44124
rect 289814 44112 289820 44124
rect 238720 44084 289820 44112
rect 238720 44072 238726 44084
rect 289814 44072 289820 44084
rect 289872 44072 289878 44124
rect 293862 44072 293868 44124
rect 293920 44112 293926 44124
rect 345014 44112 345020 44124
rect 293920 44084 345020 44112
rect 293920 44072 293926 44084
rect 345014 44072 345020 44084
rect 345072 44072 345078 44124
rect 350442 44072 350448 44124
rect 350500 44112 350506 44124
rect 401594 44112 401600 44124
rect 350500 44084 401600 44112
rect 350500 44072 350506 44084
rect 401594 44072 401600 44084
rect 401652 44072 401658 44124
rect 405642 44072 405648 44124
rect 405700 44112 405706 44124
rect 458174 44112 458180 44124
rect 405700 44084 458180 44112
rect 405700 44072 405706 44084
rect 458174 44072 458180 44084
rect 458232 44072 458238 44124
rect 462222 44072 462228 44124
rect 462280 44112 462286 44124
rect 513374 44112 513380 44124
rect 462280 44084 513380 44112
rect 462280 44072 462286 44084
rect 513374 44072 513380 44084
rect 513432 44072 513438 44124
rect 518802 44072 518808 44124
rect 518860 44112 518866 44124
rect 569954 44112 569960 44124
rect 518860 44084 569960 44112
rect 518860 44072 518866 44084
rect 569954 44072 569960 44084
rect 570012 44072 570018 44124
rect 15194 41352 15200 41404
rect 15252 41392 15258 41404
rect 35894 41392 35900 41404
rect 15252 41364 35900 41392
rect 15252 41352 15258 41364
rect 35894 41352 35900 41364
rect 35952 41352 35958 41404
rect 36078 41352 36084 41404
rect 36136 41392 36142 41404
rect 63586 41392 63592 41404
rect 36136 41364 63592 41392
rect 36136 41352 36142 41364
rect 63586 41352 63592 41364
rect 63644 41352 63650 41404
rect 65794 41352 65800 41404
rect 65852 41392 65858 41404
rect 91922 41392 91928 41404
rect 65852 41364 91928 41392
rect 65852 41352 65858 41364
rect 91922 41352 91928 41364
rect 91980 41352 91986 41404
rect 92106 41352 92112 41404
rect 92164 41392 92170 41404
rect 119614 41392 119620 41404
rect 92164 41364 119620 41392
rect 92164 41352 92170 41364
rect 119614 41352 119620 41364
rect 119672 41352 119678 41404
rect 122098 41352 122104 41404
rect 122156 41392 122162 41404
rect 147950 41392 147956 41404
rect 122156 41364 147956 41392
rect 122156 41352 122162 41364
rect 147950 41352 147956 41364
rect 148008 41352 148014 41404
rect 148042 41352 148048 41404
rect 148100 41392 148106 41404
rect 175918 41392 175924 41404
rect 148100 41364 175924 41392
rect 148100 41352 148106 41364
rect 175918 41352 175924 41364
rect 175976 41352 175982 41404
rect 176102 41352 176108 41404
rect 176160 41392 176166 41404
rect 203610 41392 203616 41404
rect 176160 41364 203616 41392
rect 176160 41352 176166 41364
rect 203610 41352 203616 41364
rect 203668 41352 203674 41404
rect 204990 41352 204996 41404
rect 205048 41392 205054 41404
rect 231946 41392 231952 41404
rect 205048 41364 231952 41392
rect 205048 41352 205054 41364
rect 231946 41352 231952 41364
rect 232004 41352 232010 41404
rect 232038 41352 232044 41404
rect 232096 41392 232102 41404
rect 259914 41392 259920 41404
rect 232096 41364 259920 41392
rect 232096 41352 232102 41364
rect 259914 41352 259920 41364
rect 259972 41352 259978 41404
rect 260098 41352 260104 41404
rect 260156 41392 260162 41404
rect 287606 41392 287612 41404
rect 260156 41364 287612 41392
rect 260156 41352 260162 41364
rect 287606 41352 287612 41364
rect 287664 41352 287670 41404
rect 288066 41352 288072 41404
rect 288124 41392 288130 41404
rect 315942 41392 315948 41404
rect 288124 41364 315948 41392
rect 288124 41352 288130 41364
rect 315942 41352 315948 41364
rect 316000 41352 316006 41404
rect 316678 41352 316684 41404
rect 316736 41392 316742 41404
rect 343910 41392 343916 41404
rect 316736 41364 343916 41392
rect 316736 41352 316742 41364
rect 343910 41352 343916 41364
rect 343968 41352 343974 41404
rect 344094 41352 344100 41404
rect 344152 41392 344158 41404
rect 371602 41392 371608 41404
rect 344152 41364 371608 41392
rect 344152 41352 344158 41364
rect 371602 41352 371608 41364
rect 371660 41352 371666 41404
rect 372062 41352 372068 41404
rect 372120 41392 372126 41404
rect 399938 41392 399944 41404
rect 372120 41364 399944 41392
rect 372120 41352 372126 41364
rect 399938 41352 399944 41364
rect 399996 41352 400002 41404
rect 400950 41352 400956 41404
rect 401008 41392 401014 41404
rect 427906 41392 427912 41404
rect 401008 41364 427912 41392
rect 401008 41352 401014 41364
rect 427906 41352 427912 41364
rect 427964 41352 427970 41404
rect 428090 41352 428096 41404
rect 428148 41392 428154 41404
rect 455598 41392 455604 41404
rect 428148 41364 455604 41392
rect 428148 41352 428154 41364
rect 455598 41352 455604 41364
rect 455656 41352 455662 41404
rect 456058 41352 456064 41404
rect 456116 41392 456122 41404
rect 483934 41392 483940 41404
rect 456116 41364 483940 41392
rect 456116 41352 456122 41364
rect 483934 41352 483940 41364
rect 483992 41352 483998 41404
rect 484026 41352 484032 41404
rect 484084 41392 484090 41404
rect 511902 41392 511908 41404
rect 484084 41364 511908 41392
rect 484084 41352 484090 41364
rect 511902 41352 511908 41364
rect 511960 41352 511966 41404
rect 512086 41352 512092 41404
rect 512144 41392 512150 41404
rect 539594 41392 539600 41404
rect 512144 41364 539600 41392
rect 512144 41352 512150 41364
rect 539594 41352 539600 41364
rect 539652 41352 539658 41404
rect 540054 41352 540060 41404
rect 540112 41392 540118 41404
rect 567930 41392 567936 41404
rect 540112 41364 567936 41392
rect 540112 41352 540118 41364
rect 567930 41352 567936 41364
rect 567988 41352 567994 41404
rect 16574 41284 16580 41336
rect 16632 41324 16638 41336
rect 36630 41324 36636 41336
rect 16632 41296 36636 41324
rect 16632 41284 16638 41296
rect 36630 41284 36636 41296
rect 36688 41284 36694 41336
rect 44910 41284 44916 41336
rect 44968 41324 44974 41336
rect 71130 41324 71136 41336
rect 44968 41296 71136 41324
rect 44968 41284 44974 41296
rect 71130 41284 71136 41296
rect 71188 41284 71194 41336
rect 82262 41284 82268 41336
rect 82320 41324 82326 41336
rect 93118 41324 93124 41336
rect 82320 41296 93124 41324
rect 82320 41284 82326 41296
rect 93118 41284 93124 41296
rect 93176 41284 93182 41336
rect 110230 41284 110236 41336
rect 110288 41324 110294 41336
rect 124858 41324 124864 41336
rect 110288 41296 124864 41324
rect 110288 41284 110294 41296
rect 124858 41284 124864 41296
rect 124916 41284 124922 41336
rect 128630 41284 128636 41336
rect 128688 41324 128694 41336
rect 151078 41324 151084 41336
rect 128688 41296 151084 41324
rect 128688 41284 128694 41296
rect 151078 41284 151084 41296
rect 151136 41284 151142 41336
rect 156598 41284 156604 41336
rect 156656 41324 156662 41336
rect 182818 41324 182824 41336
rect 156656 41296 182824 41324
rect 156656 41284 156662 41296
rect 182818 41284 182824 41296
rect 182876 41284 182882 41336
rect 194502 41284 194508 41336
rect 194560 41324 194566 41336
rect 210418 41324 210424 41336
rect 194560 41296 210424 41324
rect 194560 41284 194566 41296
rect 210418 41284 210424 41296
rect 210476 41284 210482 41336
rect 212626 41284 212632 41336
rect 212684 41324 212690 41336
rect 232498 41324 232504 41336
rect 212684 41296 232504 41324
rect 212684 41284 212690 41296
rect 232498 41284 232504 41296
rect 232556 41284 232562 41336
rect 240594 41284 240600 41336
rect 240652 41324 240658 41336
rect 266998 41324 267004 41336
rect 240652 41296 267004 41324
rect 240652 41284 240658 41296
rect 266998 41284 267004 41296
rect 267056 41284 267062 41336
rect 278590 41284 278596 41336
rect 278648 41324 278654 41336
rect 289078 41324 289084 41336
rect 278648 41296 289084 41324
rect 278648 41284 278654 41296
rect 289078 41284 289084 41296
rect 289136 41284 289142 41336
rect 306282 41284 306288 41336
rect 306340 41324 306346 41336
rect 318058 41324 318064 41336
rect 306340 41296 318064 41324
rect 306340 41284 306346 41296
rect 318058 41284 318064 41296
rect 318116 41284 318122 41336
rect 324590 41284 324596 41336
rect 324648 41324 324654 41336
rect 345658 41324 345664 41336
rect 324648 41296 345664 41324
rect 324648 41284 324654 41296
rect 345658 41284 345664 41296
rect 345716 41284 345722 41336
rect 362586 41284 362592 41336
rect 362644 41324 362650 41336
rect 373258 41324 373264 41336
rect 362644 41296 373264 41324
rect 362644 41284 362650 41296
rect 373258 41284 373264 41296
rect 373316 41284 373322 41336
rect 390278 41284 390284 41336
rect 390336 41324 390342 41336
rect 400858 41324 400864 41336
rect 390336 41296 400864 41324
rect 390336 41284 390342 41296
rect 400858 41284 400864 41296
rect 400916 41284 400922 41336
rect 408586 41284 408592 41336
rect 408644 41324 408650 41336
rect 428458 41324 428464 41336
rect 408644 41296 428464 41324
rect 408644 41284 408650 41296
rect 428458 41284 428464 41296
rect 428516 41284 428522 41336
rect 436922 41284 436928 41336
rect 436980 41324 436986 41336
rect 462958 41324 462964 41336
rect 436980 41296 462964 41324
rect 436980 41284 436986 41296
rect 462958 41284 462964 41296
rect 463016 41284 463022 41336
rect 474274 41284 474280 41336
rect 474332 41324 474338 41336
rect 485038 41324 485044 41336
rect 474332 41296 485044 41324
rect 474332 41284 474338 41296
rect 485038 41284 485044 41296
rect 485096 41284 485102 41336
rect 502242 41284 502248 41336
rect 502300 41324 502306 41336
rect 514018 41324 514024 41336
rect 502300 41296 514024 41324
rect 502300 41284 502306 41296
rect 514018 41284 514024 41296
rect 514076 41284 514082 41336
rect 520918 41284 520924 41336
rect 520976 41324 520982 41336
rect 541618 41324 541624 41336
rect 520976 41296 541624 41324
rect 520976 41284 520982 41296
rect 541618 41284 541624 41296
rect 541676 41284 541682 41336
rect 26234 41216 26240 41268
rect 26292 41256 26298 41268
rect 39298 41256 39304 41268
rect 26292 41228 39304 41256
rect 26292 41216 26298 41228
rect 39298 41216 39304 41228
rect 39356 41216 39362 41268
rect 54570 41216 54576 41268
rect 54628 41256 54634 41268
rect 66898 41256 66904 41268
rect 54628 41228 66904 41256
rect 54628 41216 54634 41228
rect 66898 41216 66904 41228
rect 66956 41216 66962 41268
rect 138290 41216 138296 41268
rect 138348 41256 138354 41268
rect 152458 41256 152464 41268
rect 138348 41228 152464 41256
rect 138348 41216 138354 41228
rect 152458 41216 152464 41228
rect 152516 41216 152522 41268
rect 166258 41216 166264 41268
rect 166316 41256 166322 41268
rect 177298 41256 177304 41268
rect 166316 41228 177304 41256
rect 166316 41216 166322 41228
rect 177298 41216 177304 41228
rect 177356 41216 177362 41268
rect 222286 41216 222292 41268
rect 222344 41256 222350 41268
rect 233970 41256 233976 41268
rect 222344 41228 233976 41256
rect 222344 41216 222350 41228
rect 233970 41216 233976 41228
rect 234028 41216 234034 41268
rect 250254 41216 250260 41268
rect 250312 41256 250318 41268
rect 261478 41256 261484 41268
rect 250312 41228 261484 41256
rect 250312 41216 250318 41228
rect 261478 41216 261484 41228
rect 261536 41216 261542 41268
rect 334250 41216 334256 41268
rect 334308 41256 334314 41268
rect 347038 41256 347044 41268
rect 334308 41228 347044 41256
rect 334308 41216 334314 41228
rect 347038 41216 347044 41228
rect 347096 41216 347102 41268
rect 418246 41216 418252 41268
rect 418304 41256 418310 41268
rect 429838 41256 429844 41268
rect 418304 41228 429844 41256
rect 418304 41216 418310 41228
rect 429838 41216 429844 41228
rect 429896 41216 429902 41268
rect 446582 41216 446588 41268
rect 446640 41256 446646 41268
rect 457438 41256 457444 41268
rect 446640 41228 457444 41256
rect 446640 41216 446646 41228
rect 457438 41216 457444 41228
rect 457496 41216 457502 41268
rect 530578 41216 530584 41268
rect 530636 41256 530642 41268
rect 544378 41256 544384 41268
rect 530636 41228 544384 41256
rect 530636 41216 530642 41228
rect 544378 41216 544384 41228
rect 544436 41216 544442 41268
rect 558270 40672 558276 40724
rect 558328 40712 558334 40724
rect 567470 40712 567476 40724
rect 558328 40684 567476 40712
rect 558328 40672 558334 40684
rect 567470 40672 567476 40684
rect 567528 40672 567534 40724
rect 46934 39380 46940 39432
rect 46992 39420 46998 39432
rect 204898 39420 204904 39432
rect 46992 39392 204904 39420
rect 46992 39380 46998 39392
rect 204898 39380 204904 39392
rect 204956 39380 204962 39432
rect 19242 39312 19248 39364
rect 19300 39352 19306 39364
rect 234614 39352 234620 39364
rect 19300 39324 234620 39352
rect 19300 39312 19306 39324
rect 234614 39312 234620 39324
rect 234672 39312 234678 39364
rect 547874 38496 547880 38548
rect 547932 38536 547938 38548
rect 548334 38536 548340 38548
rect 547932 38508 548340 38536
rect 547932 38496 547938 38508
rect 548334 38496 548340 38508
rect 548392 38496 548398 38548
rect 26970 38428 26976 38480
rect 27028 38468 27034 38480
rect 36538 38468 36544 38480
rect 27028 38440 36544 38468
rect 27028 38428 27034 38440
rect 36538 38428 36544 38440
rect 36596 38428 36602 38480
rect 53374 38428 53380 38480
rect 53432 38468 53438 38480
rect 65702 38468 65708 38480
rect 53432 38440 65708 38468
rect 53432 38428 53438 38440
rect 65702 38428 65708 38440
rect 65760 38428 65766 38480
rect 5074 38360 5080 38412
rect 5132 38400 5138 38412
rect 33410 38400 33416 38412
rect 5132 38372 33416 38400
rect 5132 38360 5138 38372
rect 33410 38360 33416 38372
rect 33468 38360 33474 38412
rect 35342 38360 35348 38412
rect 35400 38400 35406 38412
rect 149698 38400 149704 38412
rect 35400 38372 149704 38400
rect 35400 38360 35406 38372
rect 149698 38360 149704 38372
rect 149756 38360 149762 38412
rect 5166 38292 5172 38344
rect 5224 38332 5230 38344
rect 38562 38332 38568 38344
rect 5224 38304 38568 38332
rect 5224 38292 5230 38304
rect 38562 38292 38568 38304
rect 38620 38292 38626 38344
rect 43438 38292 43444 38344
rect 43496 38332 43502 38344
rect 54662 38332 54668 38344
rect 43496 38304 54668 38332
rect 43496 38292 43502 38304
rect 54662 38292 54668 38304
rect 54720 38292 54726 38344
rect 59814 38292 59820 38344
rect 59872 38332 59878 38344
rect 322198 38332 322204 38344
rect 59872 38304 322204 38332
rect 59872 38292 59878 38304
rect 322198 38292 322204 38304
rect 322256 38292 322262 38344
rect 14458 38224 14464 38276
rect 14516 38264 14522 38276
rect 20530 38264 20536 38276
rect 14516 38236 20536 38264
rect 14516 38224 14522 38236
rect 20530 38224 20536 38236
rect 20588 38224 20594 38276
rect 23750 38224 23756 38276
rect 23808 38264 23814 38276
rect 462314 38264 462320 38276
rect 23808 38236 462320 38264
rect 23808 38224 23814 38236
rect 462314 38224 462320 38236
rect 462372 38224 462378 38276
rect 11790 38156 11796 38208
rect 11848 38196 11854 38208
rect 45002 38196 45008 38208
rect 11848 38168 45008 38196
rect 11848 38156 11854 38168
rect 45002 38156 45008 38168
rect 45060 38156 45066 38208
rect 61102 38156 61108 38208
rect 61160 38196 61166 38208
rect 570690 38196 570696 38208
rect 61160 38168 570696 38196
rect 61160 38156 61166 38168
rect 570690 38156 570696 38168
rect 570748 38156 570754 38208
rect 10318 38088 10324 38140
rect 10376 38128 10382 38140
rect 30190 38128 30196 38140
rect 10376 38100 30196 38128
rect 10376 38088 10382 38100
rect 30190 38088 30196 38100
rect 30248 38088 30254 38140
rect 32122 38088 32128 38140
rect 32180 38128 32186 38140
rect 542998 38128 543004 38140
rect 32180 38100 543004 38128
rect 32180 38088 32186 38100
rect 542998 38088 543004 38100
rect 543056 38088 543062 38140
rect 4890 38020 4896 38072
rect 4948 38060 4954 38072
rect 41782 38060 41788 38072
rect 4948 38032 41788 38060
rect 4948 38020 4954 38032
rect 41782 38020 41788 38032
rect 41840 38020 41846 38072
rect 51442 38020 51448 38072
rect 51500 38060 51506 38072
rect 580902 38060 580908 38072
rect 51500 38032 580908 38060
rect 51500 38020 51506 38032
rect 580902 38020 580908 38032
rect 580960 38020 580966 38072
rect 6178 37952 6184 38004
rect 6236 37992 6242 38004
rect 22462 37992 22468 38004
rect 6236 37964 22468 37992
rect 6236 37952 6242 37964
rect 22462 37952 22468 37964
rect 22520 37952 22526 38004
rect 25682 37952 25688 38004
rect 25740 37992 25746 38004
rect 580442 37992 580448 38004
rect 25740 37964 580448 37992
rect 25740 37952 25746 37964
rect 580442 37952 580448 37964
rect 580500 37952 580506 38004
rect 16022 37884 16028 37936
rect 16080 37924 16086 37936
rect 580718 37924 580724 37936
rect 16080 37896 580724 37924
rect 16080 37884 16086 37896
rect 580718 37884 580724 37896
rect 580776 37884 580782 37936
rect 57882 37816 57888 37868
rect 57940 37856 57946 37868
rect 64230 37856 64236 37868
rect 57940 37828 64236 37856
rect 57940 37816 57946 37828
rect 64230 37816 64236 37828
rect 64288 37816 64294 37868
rect 50154 37408 50160 37460
rect 50212 37448 50218 37460
rect 61378 37448 61384 37460
rect 50212 37420 61384 37448
rect 50212 37408 50218 37420
rect 61378 37408 61384 37420
rect 61436 37408 61442 37460
rect 149790 37408 149796 37460
rect 149848 37448 149854 37460
rect 165706 37448 165712 37460
rect 149848 37420 165712 37448
rect 149848 37408 149854 37420
rect 165706 37408 165712 37420
rect 165764 37408 165770 37460
rect 175458 37408 175464 37460
rect 175516 37448 175522 37460
rect 193674 37448 193680 37460
rect 175516 37420 193680 37448
rect 175516 37408 175522 37420
rect 193674 37408 193680 37420
rect 193732 37408 193738 37460
rect 203518 37408 203524 37460
rect 203576 37448 203582 37460
rect 221366 37448 221372 37460
rect 203576 37420 221372 37448
rect 203576 37408 203582 37420
rect 221366 37408 221372 37420
rect 221424 37408 221430 37460
rect 232498 37408 232504 37460
rect 232556 37448 232562 37460
rect 249702 37448 249708 37460
rect 232556 37420 249708 37448
rect 232556 37408 232562 37420
rect 249702 37408 249708 37420
rect 249760 37408 249766 37460
rect 260190 37408 260196 37460
rect 260248 37448 260254 37460
rect 277670 37448 277676 37460
rect 260248 37420 277676 37448
rect 260248 37408 260254 37420
rect 277670 37408 277676 37420
rect 277728 37408 277734 37460
rect 287514 37408 287520 37460
rect 287572 37448 287578 37460
rect 305362 37448 305368 37460
rect 287572 37420 305368 37448
rect 287572 37408 287578 37420
rect 305362 37408 305368 37420
rect 305420 37408 305426 37460
rect 345658 37408 345664 37460
rect 345716 37448 345722 37460
rect 361666 37448 361672 37460
rect 345716 37420 361672 37448
rect 345716 37408 345722 37420
rect 361666 37408 361672 37420
rect 361724 37408 361730 37460
rect 371510 37408 371516 37460
rect 371568 37448 371574 37460
rect 389358 37448 389364 37460
rect 371568 37420 389364 37448
rect 371568 37408 371574 37420
rect 389358 37408 389364 37420
rect 389416 37408 389422 37460
rect 399478 37408 399484 37460
rect 399536 37448 399542 37460
rect 417694 37448 417700 37460
rect 399536 37420 417700 37448
rect 399536 37408 399542 37420
rect 417694 37408 417700 37420
rect 417752 37408 417758 37460
rect 456058 37408 456064 37460
rect 456116 37448 456122 37460
rect 473354 37448 473360 37460
rect 456116 37420 473360 37448
rect 456116 37408 456122 37420
rect 473354 37408 473360 37420
rect 473412 37408 473418 37460
rect 483474 37408 483480 37460
rect 483532 37448 483538 37460
rect 501690 37448 501696 37460
rect 483532 37420 501696 37448
rect 483532 37408 483538 37420
rect 501690 37408 501696 37420
rect 501748 37408 501754 37460
rect 42058 37340 42064 37392
rect 42116 37380 42122 37392
rect 48222 37380 48228 37392
rect 42116 37352 48228 37380
rect 42116 37340 42122 37352
rect 48222 37340 48228 37352
rect 48280 37340 48286 37392
rect 56594 37340 56600 37392
rect 56652 37380 56658 37392
rect 91094 37380 91100 37392
rect 56652 37352 91100 37380
rect 56652 37340 56658 37352
rect 91094 37340 91100 37352
rect 91152 37340 91158 37392
rect 91462 37340 91468 37392
rect 91520 37380 91526 37392
rect 109678 37380 109684 37392
rect 91520 37352 109684 37380
rect 91520 37340 91526 37352
rect 109678 37340 109684 37352
rect 109736 37340 109742 37392
rect 122098 37340 122104 37392
rect 122156 37380 122162 37392
rect 137646 37380 137652 37392
rect 122156 37352 137652 37380
rect 122156 37340 122162 37352
rect 137646 37340 137652 37352
rect 137704 37340 137710 37392
rect 156322 37340 156328 37392
rect 156380 37380 156386 37392
rect 178678 37380 178684 37392
rect 156380 37352 178684 37380
rect 156380 37340 156386 37352
rect 178678 37340 178684 37352
rect 178736 37340 178742 37392
rect 212350 37340 212356 37392
rect 212408 37380 212414 37392
rect 232590 37380 232596 37392
rect 212408 37352 232596 37380
rect 212408 37340 212414 37352
rect 232590 37340 232596 37352
rect 232648 37340 232654 37392
rect 268010 37340 268016 37392
rect 268068 37380 268074 37392
rect 287698 37380 287704 37392
rect 268068 37352 287704 37380
rect 268068 37340 268074 37352
rect 287698 37340 287704 37352
rect 287756 37340 287762 37392
rect 296162 37340 296168 37392
rect 296220 37380 296226 37392
rect 316770 37380 316776 37392
rect 296220 37352 316776 37380
rect 296220 37340 296226 37352
rect 316770 37340 316776 37352
rect 316828 37340 316834 37392
rect 322290 37340 322296 37392
rect 322348 37380 322354 37392
rect 333698 37380 333704 37392
rect 322348 37352 333704 37380
rect 322348 37340 322354 37352
rect 333698 37340 333704 37352
rect 333756 37340 333762 37392
rect 352006 37340 352012 37392
rect 352064 37380 352070 37392
rect 374638 37380 374644 37392
rect 352064 37352 374644 37380
rect 352064 37340 352070 37352
rect 374638 37340 374644 37352
rect 374696 37340 374702 37392
rect 408034 37340 408040 37392
rect 408092 37380 408098 37392
rect 428550 37380 428556 37392
rect 408092 37352 428556 37380
rect 408092 37340 408098 37352
rect 428550 37340 428556 37352
rect 428608 37340 428614 37392
rect 429838 37340 429844 37392
rect 429896 37380 429902 37392
rect 445662 37380 445668 37392
rect 429896 37352 445668 37380
rect 429896 37340 429902 37352
rect 445662 37340 445668 37352
rect 445720 37340 445726 37392
rect 464338 37340 464344 37392
rect 464396 37380 464402 37392
rect 483658 37380 483664 37392
rect 464396 37352 483664 37380
rect 464396 37340 464402 37352
rect 483658 37340 483664 37352
rect 483716 37340 483722 37392
rect 492030 37340 492036 37392
rect 492088 37380 492094 37392
rect 512730 37380 512736 37392
rect 492088 37352 512736 37380
rect 492088 37340 492094 37352
rect 512730 37340 512736 37352
rect 512788 37340 512794 37392
rect 518250 37340 518256 37392
rect 518308 37380 518314 37392
rect 529658 37380 529664 37392
rect 518308 37352 529664 37380
rect 518308 37340 518314 37352
rect 529658 37340 529664 37352
rect 529716 37340 529722 37392
rect 541618 37340 541624 37392
rect 541676 37380 541682 37392
rect 557534 37380 557540 37392
rect 541676 37352 557540 37380
rect 541676 37340 541682 37352
rect 557534 37340 557540 37352
rect 557592 37340 557598 37392
rect 13538 37272 13544 37324
rect 13596 37312 13602 37324
rect 81434 37312 81440 37324
rect 13596 37284 81440 37312
rect 13596 37272 13602 37284
rect 81434 37272 81440 37284
rect 81492 37272 81498 37324
rect 93118 37272 93124 37324
rect 93176 37312 93182 37324
rect 119338 37312 119344 37324
rect 93176 37284 119344 37312
rect 93176 37272 93182 37284
rect 119338 37272 119344 37284
rect 119396 37272 119402 37324
rect 120718 37272 120724 37324
rect 120776 37312 120782 37324
rect 147306 37312 147312 37324
rect 120776 37284 147312 37312
rect 120776 37272 120782 37284
rect 147306 37272 147312 37284
rect 147364 37272 147370 37324
rect 148318 37272 148324 37324
rect 148376 37312 148382 37324
rect 175366 37312 175372 37324
rect 148376 37284 175372 37312
rect 148376 37272 148382 37284
rect 175366 37272 175372 37284
rect 175424 37272 175430 37324
rect 177298 37272 177304 37324
rect 177356 37312 177362 37324
rect 203334 37312 203340 37324
rect 177356 37284 203340 37312
rect 177356 37272 177362 37284
rect 203334 37272 203340 37284
rect 203392 37272 203398 37324
rect 204898 37272 204904 37324
rect 204956 37312 204962 37324
rect 231026 37312 231032 37324
rect 204956 37284 231032 37312
rect 204956 37272 204962 37284
rect 231026 37272 231032 37284
rect 231084 37272 231090 37324
rect 239398 37272 239404 37324
rect 239456 37312 239462 37324
rect 259362 37312 259368 37324
rect 239456 37284 259368 37312
rect 239456 37272 239462 37284
rect 259362 37272 259368 37284
rect 259420 37272 259426 37324
rect 260098 37272 260104 37324
rect 260156 37312 260162 37324
rect 287330 37312 287336 37324
rect 260156 37284 287336 37312
rect 260156 37272 260162 37284
rect 287330 37272 287336 37284
rect 287388 37272 287394 37324
rect 289078 37272 289084 37324
rect 289136 37312 289142 37324
rect 315022 37312 315028 37324
rect 289136 37284 315028 37312
rect 289136 37272 289142 37284
rect 315022 37272 315028 37284
rect 315080 37272 315086 37324
rect 316678 37272 316684 37324
rect 316736 37312 316742 37324
rect 343358 37312 343364 37324
rect 316736 37284 343364 37312
rect 316736 37272 316742 37284
rect 343358 37272 343364 37284
rect 343416 37272 343422 37324
rect 344278 37272 344284 37324
rect 344336 37312 344342 37324
rect 371326 37312 371332 37324
rect 344336 37284 371332 37312
rect 344336 37272 344342 37284
rect 371326 37272 371332 37284
rect 371384 37272 371390 37324
rect 373258 37272 373264 37324
rect 373316 37312 373322 37324
rect 399018 37312 399024 37324
rect 373316 37284 399024 37312
rect 373316 37272 373322 37284
rect 399018 37272 399024 37284
rect 399076 37272 399082 37324
rect 400858 37272 400864 37324
rect 400916 37312 400922 37324
rect 427354 37312 427360 37324
rect 400916 37284 427360 37312
rect 400916 37272 400922 37284
rect 427354 37272 427360 37284
rect 427412 37272 427418 37324
rect 428458 37272 428464 37324
rect 428516 37312 428522 37324
rect 455322 37312 455328 37324
rect 428516 37284 455328 37312
rect 428516 37272 428522 37284
rect 455322 37272 455328 37284
rect 455380 37272 455386 37324
rect 456150 37272 456156 37324
rect 456208 37312 456214 37324
rect 483014 37312 483020 37324
rect 456208 37284 483020 37312
rect 456208 37272 456214 37284
rect 483014 37272 483020 37284
rect 483072 37272 483078 37324
rect 485038 37272 485044 37324
rect 485096 37312 485102 37324
rect 511350 37312 511356 37324
rect 485096 37284 511356 37312
rect 485096 37272 485102 37284
rect 511350 37272 511356 37284
rect 511408 37272 511414 37324
rect 512638 37272 512644 37324
rect 512696 37312 512702 37324
rect 539318 37312 539324 37324
rect 512696 37284 539324 37312
rect 512696 37272 512702 37284
rect 539318 37272 539324 37284
rect 539376 37272 539382 37324
rect 540238 37272 540244 37324
rect 540296 37312 540302 37324
rect 567194 37312 567200 37324
rect 540296 37284 567200 37312
rect 540296 37272 540302 37284
rect 567194 37272 567200 37284
rect 567252 37272 567258 37324
rect 64230 36728 64236 36780
rect 64288 36768 64294 36780
rect 568022 36768 568028 36780
rect 64288 36740 568028 36768
rect 64288 36728 64294 36740
rect 568022 36728 568028 36740
rect 568080 36728 568086 36780
rect 64598 36660 64604 36712
rect 64656 36700 64662 36712
rect 580166 36700 580172 36712
rect 64656 36672 580172 36700
rect 64656 36660 64662 36672
rect 580166 36660 580172 36672
rect 580224 36660 580230 36712
rect 64506 36592 64512 36644
rect 64564 36632 64570 36644
rect 580258 36632 580264 36644
rect 64564 36604 580264 36632
rect 64564 36592 64570 36604
rect 580258 36592 580264 36604
rect 580316 36592 580322 36644
rect 13722 36524 13728 36576
rect 13780 36564 13786 36576
rect 580626 36564 580632 36576
rect 13780 36536 580632 36564
rect 13780 36524 13786 36536
rect 580626 36524 580632 36536
rect 580684 36524 580690 36576
rect 39850 36048 39856 36100
rect 39908 36088 39914 36100
rect 61470 36088 61476 36100
rect 39908 36060 61476 36088
rect 39908 36048 39914 36060
rect 61470 36048 61476 36060
rect 61528 36048 61534 36100
rect 36906 35980 36912 36032
rect 36964 36020 36970 36032
rect 93854 36020 93860 36032
rect 36964 35992 93860 36020
rect 36964 35980 36970 35992
rect 93854 35980 93860 35992
rect 93912 35980 93918 36032
rect 28718 35912 28724 35964
rect 28776 35952 28782 35964
rect 579982 35952 579988 35964
rect 28776 35924 579988 35952
rect 28776 35912 28782 35924
rect 579982 35912 579988 35924
rect 580040 35912 580046 35964
rect 3786 35164 3792 35216
rect 3844 35204 3850 35216
rect 61286 35204 61292 35216
rect 3844 35176 61292 35204
rect 3844 35164 3850 35176
rect 61286 35164 61292 35176
rect 61344 35164 61350 35216
rect 63494 35164 63500 35216
rect 63552 35204 63558 35216
rect 580350 35204 580356 35216
rect 63552 35176 580356 35204
rect 63552 35164 63558 35176
rect 580350 35164 580356 35176
rect 580408 35164 580414 35216
rect 266262 34620 266268 34672
rect 266320 34660 266326 34672
rect 317414 34660 317420 34672
rect 266320 34632 317420 34660
rect 266320 34620 266326 34632
rect 317414 34620 317420 34632
rect 317472 34620 317478 34672
rect 434622 34620 434628 34672
rect 434680 34660 434686 34672
rect 485774 34660 485780 34672
rect 434680 34632 485780 34660
rect 434680 34620 434686 34632
rect 485774 34620 485780 34632
rect 485832 34620 485838 34672
rect 70302 34552 70308 34604
rect 70360 34592 70366 34604
rect 121454 34592 121460 34604
rect 70360 34564 121460 34592
rect 70360 34552 70366 34564
rect 121454 34552 121460 34564
rect 121512 34552 121518 34604
rect 126882 34552 126888 34604
rect 126940 34592 126946 34604
rect 178034 34592 178040 34604
rect 126940 34564 178040 34592
rect 126940 34552 126946 34564
rect 178034 34552 178040 34564
rect 178092 34552 178098 34604
rect 182082 34552 182088 34604
rect 182140 34592 182146 34604
rect 233234 34592 233240 34604
rect 182140 34564 233240 34592
rect 182140 34552 182146 34564
rect 233234 34552 233240 34564
rect 233292 34552 233298 34604
rect 238662 34552 238668 34604
rect 238720 34592 238726 34604
rect 289814 34592 289820 34604
rect 238720 34564 289820 34592
rect 238720 34552 238726 34564
rect 289814 34552 289820 34564
rect 289872 34552 289878 34604
rect 322842 34552 322848 34604
rect 322900 34592 322906 34604
rect 373994 34592 374000 34604
rect 322900 34564 374000 34592
rect 322900 34552 322906 34564
rect 373994 34552 374000 34564
rect 374052 34552 374058 34604
rect 378042 34552 378048 34604
rect 378100 34592 378106 34604
rect 429286 34592 429292 34604
rect 378100 34564 429292 34592
rect 378100 34552 378106 34564
rect 429286 34552 429292 34564
rect 429344 34552 429350 34604
rect 462222 34552 462228 34604
rect 462280 34592 462286 34604
rect 513374 34592 513380 34604
rect 462280 34564 513380 34592
rect 462280 34552 462286 34564
rect 513374 34552 513380 34564
rect 513432 34552 513438 34604
rect 518802 34552 518808 34604
rect 518860 34592 518866 34604
rect 569954 34592 569960 34604
rect 518860 34564 569960 34592
rect 518860 34552 518866 34564
rect 569954 34552 569960 34564
rect 570012 34552 570018 34604
rect 97902 34484 97908 34536
rect 97960 34524 97966 34536
rect 149054 34524 149060 34536
rect 97960 34496 149060 34524
rect 97960 34484 97966 34496
rect 149054 34484 149060 34496
rect 149112 34484 149118 34536
rect 154482 34484 154488 34536
rect 154540 34524 154546 34536
rect 205634 34524 205640 34536
rect 154540 34496 205640 34524
rect 154540 34484 154546 34496
rect 205634 34484 205640 34496
rect 205692 34484 205698 34536
rect 209682 34484 209688 34536
rect 209740 34524 209746 34536
rect 262214 34524 262220 34536
rect 209740 34496 262220 34524
rect 209740 34484 209746 34496
rect 262214 34484 262220 34496
rect 262272 34484 262278 34536
rect 293862 34484 293868 34536
rect 293920 34524 293926 34536
rect 345014 34524 345020 34536
rect 293920 34496 345020 34524
rect 293920 34484 293926 34496
rect 345014 34484 345020 34496
rect 345072 34484 345078 34536
rect 350442 34484 350448 34536
rect 350500 34524 350506 34536
rect 401594 34524 401600 34536
rect 350500 34496 401600 34524
rect 350500 34484 350506 34496
rect 401594 34484 401600 34496
rect 401652 34484 401658 34536
rect 405642 34484 405648 34536
rect 405700 34524 405706 34536
rect 458174 34524 458180 34536
rect 405700 34496 458180 34524
rect 405700 34484 405706 34496
rect 458174 34484 458180 34496
rect 458232 34484 458238 34536
rect 489822 34484 489828 34536
rect 489880 34524 489886 34536
rect 542354 34524 542360 34536
rect 489880 34496 542360 34524
rect 489880 34484 489886 34496
rect 542354 34484 542360 34496
rect 542412 34484 542418 34536
rect 3326 31696 3332 31748
rect 3384 31736 3390 31748
rect 12434 31736 12440 31748
rect 3384 31708 12440 31736
rect 3384 31696 3390 31708
rect 12434 31696 12440 31708
rect 12492 31696 12498 31748
rect 238846 30744 238852 30796
rect 238904 30784 238910 30796
rect 239766 30784 239772 30796
rect 238904 30756 239772 30784
rect 238904 30744 238910 30756
rect 239766 30744 239772 30756
rect 239824 30744 239830 30796
rect 63494 27548 63500 27600
rect 63552 27588 63558 27600
rect 71038 27588 71044 27600
rect 63552 27560 71044 27588
rect 63552 27548 63558 27560
rect 71038 27548 71044 27560
rect 71096 27548 71102 27600
rect 4982 23400 4988 23452
rect 5040 23440 5046 23452
rect 12434 23440 12440 23452
rect 5040 23412 12440 23440
rect 5040 23400 5046 23412
rect 12434 23400 12440 23412
rect 12492 23400 12498 23452
rect 4798 22040 4804 22092
rect 4856 22080 4862 22092
rect 12434 22080 12440 22092
rect 4856 22052 12440 22080
rect 4856 22040 4862 22052
rect 12434 22040 12440 22052
rect 12492 22040 12498 22092
rect 259730 21428 259736 21480
rect 259788 21468 259794 21480
rect 260190 21468 260196 21480
rect 259788 21440 260196 21468
rect 259788 21428 259794 21440
rect 260190 21428 260196 21440
rect 260248 21428 260254 21480
rect 9030 20612 9036 20664
rect 9088 20652 9094 20664
rect 12618 20652 12624 20664
rect 9088 20624 12624 20652
rect 9088 20612 9094 20624
rect 12618 20612 12624 20624
rect 12676 20612 12682 20664
rect 428550 18572 428556 18624
rect 428608 18612 428614 18624
rect 435726 18612 435732 18624
rect 428608 18584 435732 18612
rect 428608 18572 428614 18584
rect 435726 18572 435732 18584
rect 435784 18572 435790 18624
rect 287698 18232 287704 18284
rect 287756 18272 287762 18284
rect 295702 18272 295708 18284
rect 287756 18244 295708 18272
rect 287756 18232 287762 18244
rect 295702 18232 295708 18244
rect 295760 18232 295766 18284
rect 316770 18096 316776 18148
rect 316828 18136 316834 18148
rect 323670 18136 323676 18148
rect 316828 18108 323676 18136
rect 316828 18096 316834 18108
rect 323670 18096 323676 18108
rect 323728 18096 323734 18148
rect 232590 17960 232596 18012
rect 232648 18000 232654 18012
rect 239766 18000 239772 18012
rect 232648 17972 239772 18000
rect 232648 17960 232654 17972
rect 239766 17960 239772 17972
rect 239824 17960 239830 18012
rect 483658 17960 483664 18012
rect 483716 18000 483722 18012
rect 491662 18000 491668 18012
rect 483716 17972 491668 18000
rect 483716 17960 483722 17972
rect 491662 17960 491668 17972
rect 491720 17960 491726 18012
rect 512730 17960 512736 18012
rect 512788 18000 512794 18012
rect 519630 18000 519636 18012
rect 512788 17972 519636 18000
rect 512788 17960 512794 17972
rect 519630 17960 519636 17972
rect 519688 17960 519694 18012
rect 7558 17892 7564 17944
rect 7616 17932 7622 17944
rect 12434 17932 12440 17944
rect 7616 17904 12440 17932
rect 7616 17892 7622 17904
rect 12434 17892 12440 17904
rect 12492 17892 12498 17944
rect 3786 16532 3792 16584
rect 3844 16572 3850 16584
rect 63494 16572 63500 16584
rect 3844 16544 63500 16572
rect 3844 16532 3850 16544
rect 63494 16532 63500 16544
rect 63552 16532 63558 16584
rect 119706 16532 119712 16584
rect 119764 16572 119770 16584
rect 122098 16572 122104 16584
rect 119764 16544 122104 16572
rect 119764 16532 119770 16544
rect 122098 16532 122104 16544
rect 122156 16532 122162 16584
rect 147582 16532 147588 16584
rect 147640 16572 147646 16584
rect 149790 16572 149796 16584
rect 147640 16544 149796 16572
rect 147640 16532 147646 16544
rect 149790 16532 149796 16544
rect 149848 16532 149854 16584
rect 343542 16532 343548 16584
rect 343600 16572 343606 16584
rect 345658 16572 345664 16584
rect 343600 16544 345664 16572
rect 343600 16532 343606 16544
rect 345658 16532 345664 16544
rect 345716 16532 345722 16584
rect 427722 16532 427728 16584
rect 427780 16572 427786 16584
rect 429838 16572 429844 16584
rect 427780 16544 429844 16572
rect 427780 16532 427786 16544
rect 429838 16532 429844 16544
rect 429896 16532 429902 16584
rect 539502 16532 539508 16584
rect 539560 16572 539566 16584
rect 541618 16572 541624 16584
rect 539560 16544 541624 16572
rect 539560 16532 539566 16544
rect 541618 16532 541624 16544
rect 541676 16532 541682 16584
rect 41782 15104 41788 15156
rect 41840 15144 41846 15156
rect 429194 15144 429200 15156
rect 41840 15116 429200 15144
rect 41840 15104 41846 15116
rect 429194 15104 429200 15116
rect 429252 15104 429258 15156
rect 52730 15036 52736 15088
rect 52788 15076 52794 15088
rect 233878 15076 233884 15088
rect 52788 15048 233884 15076
rect 52788 15036 52794 15048
rect 233878 15036 233884 15048
rect 233936 15036 233942 15088
rect 39850 13744 39856 13796
rect 39908 13784 39914 13796
rect 65610 13784 65616 13796
rect 39908 13756 65616 13784
rect 39908 13744 39914 13756
rect 65610 13744 65616 13756
rect 65668 13744 65674 13796
rect 81986 13744 81992 13796
rect 82044 13784 82050 13796
rect 93118 13784 93124 13796
rect 82044 13756 93124 13784
rect 82044 13744 82050 13756
rect 93118 13744 93124 13756
rect 93176 13744 93182 13796
rect 165982 13744 165988 13796
rect 166040 13784 166046 13796
rect 177298 13784 177304 13796
rect 166040 13756 177304 13784
rect 166040 13744 166046 13756
rect 177298 13744 177304 13756
rect 177356 13744 177362 13796
rect 178678 13744 178684 13796
rect 178736 13784 178742 13796
rect 184014 13784 184020 13796
rect 178736 13756 184020 13784
rect 178736 13744 178742 13756
rect 184014 13744 184020 13756
rect 184072 13744 184078 13796
rect 193674 13744 193680 13796
rect 193732 13784 193738 13796
rect 204898 13784 204904 13796
rect 193732 13756 204904 13784
rect 193732 13744 193738 13756
rect 204898 13744 204904 13756
rect 204956 13744 204962 13796
rect 249702 13744 249708 13796
rect 249760 13784 249766 13796
rect 260098 13784 260104 13796
rect 249760 13756 260104 13784
rect 249760 13744 249766 13756
rect 260098 13744 260104 13756
rect 260156 13744 260162 13796
rect 277670 13744 277676 13796
rect 277728 13784 277734 13796
rect 289078 13784 289084 13796
rect 277728 13756 289084 13784
rect 277728 13744 277734 13756
rect 289078 13744 289084 13756
rect 289136 13744 289142 13796
rect 306006 13744 306012 13796
rect 306064 13784 306070 13796
rect 316678 13784 316684 13796
rect 306064 13756 316684 13784
rect 306064 13744 306070 13756
rect 316678 13744 316684 13756
rect 316736 13744 316742 13796
rect 361666 13744 361672 13796
rect 361724 13784 361730 13796
rect 373258 13784 373264 13796
rect 361724 13756 373264 13784
rect 361724 13744 361730 13756
rect 373258 13744 373264 13756
rect 373316 13744 373322 13796
rect 374638 13744 374644 13796
rect 374696 13784 374702 13796
rect 379698 13784 379704 13796
rect 374696 13756 379704 13784
rect 374696 13744 374702 13756
rect 379698 13744 379704 13756
rect 379756 13744 379762 13796
rect 390002 13744 390008 13796
rect 390060 13784 390066 13796
rect 400858 13784 400864 13796
rect 390060 13756 400864 13784
rect 390060 13744 390066 13756
rect 400858 13744 400864 13756
rect 400916 13744 400922 13796
rect 473998 13744 474004 13796
rect 474056 13784 474062 13796
rect 485038 13784 485044 13796
rect 474056 13756 485044 13784
rect 474056 13744 474062 13756
rect 485038 13744 485044 13756
rect 485096 13744 485102 13796
rect 501690 13744 501696 13796
rect 501748 13784 501754 13796
rect 512638 13784 512644 13796
rect 501748 13756 512644 13784
rect 501748 13744 501754 13756
rect 512638 13744 512644 13756
rect 512696 13744 512702 13796
rect 529658 13744 529664 13796
rect 529716 13784 529722 13796
rect 540238 13784 540244 13796
rect 529716 13756 540244 13784
rect 529716 13744 529722 13756
rect 540238 13744 540244 13756
rect 540296 13744 540302 13796
rect 547874 13744 547880 13796
rect 547932 13784 547938 13796
rect 557534 13784 557540 13796
rect 547932 13756 557540 13784
rect 547932 13744 547938 13756
rect 557534 13744 557540 13756
rect 557592 13744 557598 13796
rect 17310 13676 17316 13728
rect 17368 13716 17374 13728
rect 570598 13716 570604 13728
rect 17368 13688 570604 13716
rect 17368 13676 17374 13688
rect 570598 13676 570604 13688
rect 570656 13676 570662 13728
rect 3418 13608 3424 13660
rect 3476 13648 3482 13660
rect 28902 13648 28908 13660
rect 3476 13620 28908 13648
rect 3476 13608 3482 13620
rect 28902 13608 28908 13620
rect 28960 13608 28966 13660
rect 32122 13608 32128 13660
rect 32180 13648 32186 13660
rect 580074 13648 580080 13660
rect 32180 13620 580080 13648
rect 32180 13608 32186 13620
rect 580074 13608 580080 13620
rect 580132 13608 580138 13660
rect 4062 13540 4068 13592
rect 4120 13580 4126 13592
rect 25682 13580 25688 13592
rect 4120 13552 25688 13580
rect 4120 13540 4126 13552
rect 25682 13540 25688 13552
rect 25740 13540 25746 13592
rect 36630 13540 36636 13592
rect 36688 13580 36694 13592
rect 580534 13580 580540 13592
rect 36688 13552 580540 13580
rect 36688 13540 36694 13552
rect 580534 13540 580540 13552
rect 580592 13540 580598 13592
rect 8938 13472 8944 13524
rect 8996 13512 9002 13524
rect 30190 13512 30196 13524
rect 8996 13484 30196 13512
rect 8996 13472 9002 13484
rect 30190 13472 30196 13484
rect 30248 13472 30254 13524
rect 43070 13472 43076 13524
rect 43128 13512 43134 13524
rect 580810 13512 580816 13524
rect 43128 13484 580816 13512
rect 43128 13472 43134 13484
rect 580810 13472 580816 13484
rect 580868 13472 580874 13524
rect 26970 13404 26976 13456
rect 27028 13444 27034 13456
rect 378778 13444 378784 13456
rect 27028 13416 378784 13444
rect 27028 13404 27034 13416
rect 378778 13404 378784 13416
rect 378836 13404 378842 13456
rect 379606 13404 379612 13456
rect 379664 13444 379670 13456
rect 408034 13444 408040 13456
rect 379664 13416 408040 13444
rect 379664 13404 379670 13416
rect 408034 13404 408040 13416
rect 408092 13404 408098 13456
rect 417694 13404 417700 13456
rect 417752 13444 417758 13456
rect 428458 13444 428464 13456
rect 417752 13416 428464 13444
rect 417752 13404 417758 13416
rect 428458 13404 428464 13416
rect 428516 13404 428522 13456
rect 434806 13404 434812 13456
rect 434864 13444 434870 13456
rect 463694 13444 463700 13456
rect 434864 13416 463700 13444
rect 434864 13404 434870 13416
rect 463694 13404 463700 13416
rect 463752 13404 463758 13456
rect 511350 13404 511356 13456
rect 511408 13444 511414 13456
rect 518250 13444 518256 13456
rect 511408 13416 518256 13444
rect 511408 13404 511414 13416
rect 518250 13404 518256 13416
rect 518308 13404 518314 13456
rect 518986 13404 518992 13456
rect 519044 13444 519050 13456
rect 547966 13444 547972 13456
rect 519044 13416 547972 13444
rect 519044 13404 519050 13416
rect 547966 13404 547972 13416
rect 548024 13404 548030 13456
rect 3602 13336 3608 13388
rect 3660 13376 3666 13388
rect 57882 13376 57888 13388
rect 3660 13348 57888 13376
rect 3660 13336 3666 13348
rect 57882 13336 57888 13348
rect 57940 13336 57946 13388
rect 71866 13336 71872 13388
rect 71924 13376 71930 13388
rect 100018 13376 100024 13388
rect 71924 13348 100024 13376
rect 71924 13336 71930 13348
rect 100018 13336 100024 13348
rect 100076 13336 100082 13388
rect 127986 13376 127992 13388
rect 103486 13348 127992 13376
rect 3694 13268 3700 13320
rect 3752 13308 3758 13320
rect 54662 13308 54668 13320
rect 3752 13280 54668 13308
rect 3752 13268 3758 13280
rect 54662 13268 54668 13280
rect 54720 13268 54726 13320
rect 99466 13268 99472 13320
rect 99524 13308 99530 13320
rect 103486 13308 103514 13348
rect 127986 13336 127992 13348
rect 128044 13336 128050 13388
rect 156046 13376 156052 13388
rect 132466 13348 156052 13376
rect 99524 13280 103514 13308
rect 99524 13268 99530 13280
rect 109678 13268 109684 13320
rect 109736 13308 109742 13320
rect 120718 13308 120724 13320
rect 109736 13280 120724 13308
rect 109736 13268 109742 13280
rect 120718 13268 120724 13280
rect 120776 13268 120782 13320
rect 127066 13268 127072 13320
rect 127124 13308 127130 13320
rect 132466 13308 132494 13348
rect 156046 13336 156052 13348
rect 156104 13336 156110 13388
rect 183646 13336 183652 13388
rect 183704 13376 183710 13388
rect 211706 13376 211712 13388
rect 183704 13348 211712 13376
rect 183704 13336 183710 13348
rect 211706 13336 211712 13348
rect 211764 13336 211770 13388
rect 222010 13336 222016 13388
rect 222068 13376 222074 13388
rect 239398 13376 239404 13388
rect 222068 13348 239404 13376
rect 222068 13336 222074 13348
rect 239398 13336 239404 13348
rect 239456 13336 239462 13388
rect 315666 13336 315672 13388
rect 315724 13376 315730 13388
rect 322290 13376 322296 13388
rect 315724 13348 322296 13376
rect 315724 13336 315730 13348
rect 322290 13336 322296 13348
rect 322348 13336 322354 13388
rect 323026 13336 323032 13388
rect 323084 13376 323090 13388
rect 352006 13376 352012 13388
rect 323084 13348 352012 13376
rect 323084 13336 323090 13348
rect 352006 13336 352012 13348
rect 352064 13336 352070 13388
rect 445662 13336 445668 13388
rect 445720 13376 445726 13388
rect 456150 13376 456156 13388
rect 445720 13348 456156 13376
rect 445720 13336 445726 13348
rect 456150 13336 456156 13348
rect 456208 13336 456214 13388
rect 127124 13280 132494 13308
rect 127124 13268 127130 13280
rect 137646 13268 137652 13320
rect 137704 13308 137710 13320
rect 148318 13308 148324 13320
rect 137704 13280 148324 13308
rect 137704 13268 137710 13280
rect 148318 13268 148324 13280
rect 148376 13268 148382 13320
rect 333698 13268 333704 13320
rect 333756 13308 333762 13320
rect 344278 13308 344284 13320
rect 333756 13280 344284 13308
rect 333756 13268 333762 13280
rect 344278 13268 344284 13280
rect 344336 13268 344342 13320
rect 6914 13200 6920 13252
rect 6972 13240 6978 13252
rect 55950 13240 55956 13252
rect 6972 13212 55956 13240
rect 6972 13200 6978 13212
rect 55950 13200 55956 13212
rect 56008 13200 56014 13252
rect 238846 13200 238852 13252
rect 238904 13240 238910 13252
rect 268010 13240 268016 13252
rect 238904 13212 268016 13240
rect 238904 13200 238910 13212
rect 268010 13200 268016 13212
rect 268068 13200 268074 13252
rect 3970 13132 3976 13184
rect 4028 13172 4034 13184
rect 22462 13172 22468 13184
rect 4028 13144 22468 13172
rect 4028 13132 4034 13144
rect 22462 13132 22468 13144
rect 22520 13132 22526 13184
rect 23750 13132 23756 13184
rect 23808 13172 23814 13184
rect 65518 13172 65524 13184
rect 23808 13144 65524 13172
rect 23808 13132 23814 13144
rect 65518 13132 65524 13144
rect 65576 13132 65582 13184
rect 1394 13064 1400 13116
rect 1452 13104 1458 13116
rect 33410 13104 33416 13116
rect 1452 13076 33416 13104
rect 1452 13064 1458 13076
rect 33410 13064 33416 13076
rect 33468 13064 33474 13116
rect 38562 13064 38568 13116
rect 38620 13104 38626 13116
rect 72050 13104 72056 13116
rect 38620 13076 72056 13104
rect 38620 13064 38626 13076
rect 72050 13064 72056 13076
rect 72108 13064 72114 13116
rect 20530 12996 20536 13048
rect 20588 13036 20594 13048
rect 578878 13036 578884 13048
rect 20588 13008 578884 13036
rect 20588 12996 20594 13008
rect 578878 12996 578884 13008
rect 578936 12996 578942 13048
rect 3510 12928 3516 12980
rect 3568 12968 3574 12980
rect 46290 12968 46296 12980
rect 3568 12940 46296 12968
rect 3568 12928 3574 12940
rect 46290 12928 46296 12940
rect 46348 12928 46354 12980
rect 3878 12860 3884 12912
rect 3936 12900 3942 12912
rect 51442 12900 51448 12912
rect 3936 12872 51448 12900
rect 3936 12860 3942 12872
rect 51442 12860 51448 12872
rect 51500 12860 51506 12912
rect 11698 12792 11704 12844
rect 11756 12832 11762 12844
rect 35342 12832 35348 12844
rect 11756 12804 35348 12832
rect 11756 12792 11762 12804
rect 35342 12792 35348 12804
rect 35400 12792 35406 12844
rect 64414 3680 64420 3732
rect 64472 3720 64478 3732
rect 125870 3720 125876 3732
rect 64472 3692 125876 3720
rect 64472 3680 64478 3692
rect 125870 3680 125876 3692
rect 125928 3680 125934 3732
rect 64230 3612 64236 3664
rect 64288 3652 64294 3664
rect 126974 3652 126980 3664
rect 64288 3624 126980 3652
rect 64288 3612 64294 3624
rect 126974 3612 126980 3624
rect 127032 3612 127038 3664
rect 61378 3544 61384 3596
rect 61436 3584 61442 3596
rect 132954 3584 132960 3596
rect 61436 3556 132960 3584
rect 61436 3544 61442 3556
rect 132954 3544 132960 3556
rect 133012 3544 133018 3596
rect 13722 3476 13728 3528
rect 13780 3516 13786 3528
rect 129366 3516 129372 3528
rect 13780 3488 129372 3516
rect 13780 3476 13786 3488
rect 129366 3476 129372 3488
rect 129424 3476 129430 3528
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 48314 3448 48320 3460
rect 624 3420 48320 3448
rect 624 3408 630 3420
rect 48314 3408 48320 3420
rect 48372 3408 48378 3460
rect 61470 3408 61476 3460
rect 61528 3448 61534 3460
rect 136450 3448 136456 3460
rect 61528 3420 136456 3448
rect 61528 3408 61534 3420
rect 136450 3408 136456 3420
rect 136508 3408 136514 3460
<< via1 >>
rect 36544 700612 36596 700664
rect 105452 700612 105504 700664
rect 71044 700544 71096 700596
rect 267648 700544 267700 700596
rect 13452 700476 13504 700528
rect 300124 700476 300176 700528
rect 322204 700476 322256 700528
rect 332508 700476 332560 700528
rect 65524 700408 65576 700460
rect 137836 700408 137888 700460
rect 153844 700408 153896 700460
rect 170312 700408 170364 700460
rect 204904 700408 204956 700460
rect 494796 700408 494848 700460
rect 64144 700340 64196 700392
rect 364984 700340 365036 700392
rect 378784 700340 378836 700392
rect 397460 700340 397512 700392
rect 518164 700340 518216 700392
rect 527180 700340 527232 700392
rect 64236 700272 64288 700324
rect 202788 700272 202840 700324
rect 233884 700272 233936 700324
rect 559656 700272 559708 700324
rect 40500 699932 40552 699984
rect 42064 699932 42116 699984
rect 65616 699660 65668 699712
rect 72976 699660 73028 699712
rect 65708 696940 65760 696992
rect 580172 696940 580224 696992
rect 212356 686060 212408 686112
rect 232688 686060 232740 686112
rect 296352 686060 296404 686112
rect 316776 686060 316828 686112
rect 408040 686060 408092 686112
rect 428648 686060 428700 686112
rect 492036 686060 492088 686112
rect 512736 686060 512788 686112
rect 148324 685992 148376 686044
rect 165712 685992 165764 686044
rect 175464 685992 175516 686044
rect 193680 685992 193732 686044
rect 203524 685992 203576 686044
rect 221372 685992 221424 686044
rect 260104 685992 260156 686044
rect 277676 685992 277728 686044
rect 287520 685992 287572 686044
rect 305368 685992 305420 686044
rect 345664 685992 345716 686044
rect 361672 685992 361724 686044
rect 371516 685992 371568 686044
rect 389364 685992 389416 686044
rect 399484 685992 399536 686044
rect 417700 685992 417752 686044
rect 456064 685992 456116 686044
rect 473360 685992 473412 686044
rect 483480 685992 483532 686044
rect 501696 685992 501748 686044
rect 36728 685924 36780 685976
rect 53656 685924 53708 685976
rect 64328 685924 64380 685976
rect 81440 685924 81492 685976
rect 91468 685924 91520 685976
rect 109684 685924 109736 685976
rect 119436 685924 119488 685976
rect 137652 685924 137704 685976
rect 156328 685924 156380 685976
rect 178684 685924 178736 685976
rect 232596 685924 232648 685976
rect 249708 685924 249760 685976
rect 268016 685924 268068 685976
rect 287704 685924 287756 685976
rect 315488 685924 315540 685976
rect 333704 685924 333756 685976
rect 352012 685924 352064 685976
rect 374644 685924 374696 685976
rect 428556 685924 428608 685976
rect 445668 685924 445720 685976
rect 464344 685924 464396 685976
rect 483664 685924 483716 685976
rect 511448 685924 511500 685976
rect 529664 685924 529716 685976
rect 541624 685924 541676 685976
rect 557540 685924 557592 685976
rect 16120 685856 16172 685908
rect 25688 685856 25740 685908
rect 36636 685856 36688 685908
rect 63316 685856 63368 685908
rect 66904 685856 66956 685908
rect 91100 685856 91152 685908
rect 93124 685856 93176 685908
rect 119344 685856 119396 685908
rect 122104 685856 122156 685908
rect 147312 685856 147364 685908
rect 148416 685856 148468 685908
rect 175372 685856 175424 685908
rect 177304 685856 177356 685908
rect 203340 685856 203392 685908
rect 204996 685856 205048 685908
rect 231032 685856 231084 685908
rect 232504 685856 232556 685908
rect 259368 685856 259420 685908
rect 260196 685856 260248 685908
rect 287336 685856 287388 685908
rect 289084 685856 289136 685908
rect 315028 685856 315080 685908
rect 316684 685856 316736 685908
rect 343364 685856 343416 685908
rect 344284 685856 344336 685908
rect 371332 685856 371384 685908
rect 373264 685856 373316 685908
rect 399024 685856 399076 685908
rect 400864 685856 400916 685908
rect 427360 685856 427412 685908
rect 428464 685856 428516 685908
rect 455328 685856 455380 685908
rect 456156 685856 456208 685908
rect 483020 685856 483072 685908
rect 485044 685856 485096 685908
rect 511356 685856 511408 685908
rect 512644 685856 512696 685908
rect 539324 685856 539376 685908
rect 540244 685856 540296 685908
rect 567200 685856 567252 685908
rect 15844 683272 15896 683324
rect 16120 683272 16172 683324
rect 3424 683204 3476 683256
rect 43444 683204 43496 683256
rect 182088 683204 182140 683256
rect 233240 683204 233292 683256
rect 350448 683204 350500 683256
rect 401600 683204 401652 683256
rect 42708 683136 42760 683188
rect 93860 683136 93912 683188
rect 97908 683136 97960 683188
rect 149060 683136 149112 683188
rect 154488 683136 154540 683188
rect 205640 683136 205692 683188
rect 238668 683136 238720 683188
rect 289820 683136 289872 683188
rect 293868 683136 293920 683188
rect 345020 683136 345072 683188
rect 378048 683136 378100 683188
rect 429292 683136 429344 683188
rect 434628 683136 434680 683188
rect 485780 683136 485832 683188
rect 489828 683136 489880 683188
rect 542360 683136 542412 683188
rect 543004 673752 543056 673804
rect 545120 673752 545172 673804
rect 63592 668720 63644 668772
rect 64328 668720 64380 668772
rect 428648 665796 428700 665848
rect 435732 665796 435784 665848
rect 287704 665456 287756 665508
rect 295708 665456 295760 665508
rect 316776 665456 316828 665508
rect 323676 665456 323728 665508
rect 232688 665252 232740 665304
rect 239772 665252 239824 665304
rect 483664 665252 483716 665304
rect 491668 665252 491720 665304
rect 512736 665252 512788 665304
rect 519636 665252 519688 665304
rect 13636 665116 13688 665168
rect 66260 665116 66312 665168
rect 70308 665116 70360 665168
rect 121460 665116 121512 665168
rect 126888 665116 126940 665168
rect 178040 665116 178092 665168
rect 209688 665116 209740 665168
rect 262220 665116 262272 665168
rect 266268 665116 266320 665168
rect 317420 665116 317472 665168
rect 322848 665116 322900 665168
rect 374000 665116 374052 665168
rect 405648 665116 405700 665168
rect 458180 665116 458232 665168
rect 462228 665116 462280 665168
rect 513380 665116 513432 665168
rect 518808 665116 518860 665168
rect 569960 665116 570012 665168
rect 343548 665048 343600 665100
rect 345664 665048 345716 665100
rect 427728 665048 427780 665100
rect 428556 665048 428608 665100
rect 35256 664708 35308 664760
rect 36728 664708 36780 664760
rect 15844 664096 15896 664148
rect 16580 664096 16632 664148
rect 231584 663688 231636 663740
rect 232596 663688 232648 663740
rect 539324 663688 539376 663740
rect 541624 663688 541676 663740
rect 71872 662328 71924 662380
rect 100024 662328 100076 662380
rect 25688 662260 25740 662312
rect 36636 662260 36688 662312
rect 42892 662260 42944 662312
rect 15292 662192 15344 662244
rect 43628 662192 43680 662244
rect 53748 662260 53800 662312
rect 66904 662260 66956 662312
rect 81992 662260 82044 662312
rect 93124 662260 93176 662312
rect 99472 662260 99524 662312
rect 127716 662328 127768 662380
rect 165988 662328 166040 662380
rect 177304 662328 177356 662380
rect 178684 662328 178736 662380
rect 184020 662328 184072 662380
rect 109684 662260 109736 662312
rect 122104 662260 122156 662312
rect 137928 662260 137980 662312
rect 148416 662260 148468 662312
rect 183652 662260 183704 662312
rect 211712 662328 211764 662380
rect 277676 662328 277728 662380
rect 289084 662328 289136 662380
rect 306012 662328 306064 662380
rect 316684 662328 316736 662380
rect 361672 662328 361724 662380
rect 373264 662328 373316 662380
rect 379612 662328 379664 662380
rect 408040 662328 408092 662380
rect 474004 662328 474056 662380
rect 485044 662328 485096 662380
rect 501696 662328 501748 662380
rect 512644 662328 512696 662380
rect 193680 662260 193732 662312
rect 204996 662260 205048 662312
rect 222016 662260 222068 662312
rect 232504 662260 232556 662312
rect 249616 662260 249668 662312
rect 260196 662260 260248 662312
rect 333888 662260 333940 662312
rect 344284 662260 344336 662312
rect 374644 662260 374696 662312
rect 379704 662260 379756 662312
rect 390008 662260 390060 662312
rect 400864 662260 400916 662312
rect 417700 662260 417752 662312
rect 428464 662260 428516 662312
rect 445668 662260 445720 662312
rect 456156 662260 456208 662312
rect 529664 662260 529716 662312
rect 540244 662260 540296 662312
rect 71964 662192 72016 662244
rect 127072 662192 127124 662244
rect 155960 662192 156012 662244
rect 238852 662192 238904 662244
rect 268016 662192 268068 662244
rect 323032 662192 323084 662244
rect 352012 662192 352064 662244
rect 434812 662192 434864 662244
rect 463792 662192 463844 662244
rect 518992 662192 519044 662244
rect 547880 662192 547932 662244
rect 13636 661648 13688 661700
rect 557540 661648 557592 661700
rect 267832 658452 267884 658504
rect 71136 658384 71188 658436
rect 82268 658384 82320 658436
rect 99472 658384 99524 658436
rect 100392 658384 100444 658436
rect 183652 658384 183704 658436
rect 222292 658384 222344 658436
rect 267004 658384 267056 658436
rect 26240 658316 26292 658368
rect 35440 658316 35492 658368
rect 36636 658316 36688 658368
rect 53932 658316 53984 658368
rect 71872 658316 71924 658368
rect 109960 658316 110012 658368
rect 124864 658316 124916 658368
rect 128636 658316 128688 658368
rect 151084 658316 151136 658368
rect 156604 658316 156656 658368
rect 182824 658316 182876 658368
rect 193956 658316 194008 658368
rect 232504 658316 232556 658368
rect 66904 658248 66956 658300
rect 72608 658248 72660 658300
rect 93124 658248 93176 658300
rect 100300 658248 100352 658300
rect 100392 658248 100444 658300
rect 138296 658248 138348 658300
rect 149704 658248 149756 658300
rect 166264 658248 166316 658300
rect 177304 658248 177356 658300
rect 184296 658248 184348 658300
rect 233976 658248 234028 658300
rect 240600 658248 240652 658300
rect 250260 658248 250312 658300
rect 261484 658248 261536 658300
rect 268292 658248 268344 658300
rect 295432 658384 295484 658436
rect 334256 658384 334308 658436
rect 352012 658384 352064 658436
rect 306288 658316 306340 658368
rect 347044 658316 347096 658368
rect 361948 658316 362000 658368
rect 379612 658384 379664 658436
rect 418252 658384 418304 658436
rect 463792 658384 463844 658436
rect 390284 658316 390336 658368
rect 400864 658316 400916 658368
rect 408592 658316 408644 658368
rect 429844 658316 429896 658368
rect 436284 658316 436336 658368
rect 457444 658316 457496 658368
rect 464620 658316 464672 658368
rect 491392 658384 491444 658436
rect 529940 658384 529992 658436
rect 502248 658316 502300 658368
rect 512644 658316 512696 658368
rect 520280 658316 520332 658368
rect 541624 658316 541676 658368
rect 277952 658248 278004 658300
rect 289084 658248 289136 658300
rect 296628 658248 296680 658300
rect 318064 658248 318116 658300
rect 324596 658248 324648 658300
rect 348424 658248 348476 658300
rect 352288 658248 352340 658300
rect 373264 658248 373316 658300
rect 380624 658248 380676 658300
rect 428464 658248 428516 658300
rect 445944 658248 445996 658300
rect 462964 658248 463016 658300
rect 474280 658248 474332 658300
rect 485044 658248 485096 658300
rect 492588 658248 492640 658300
rect 544384 658248 544436 658300
rect 548616 658248 548668 658300
rect 558276 658248 558328 658300
rect 2780 657500 2832 657552
rect 6184 657500 6236 657552
rect 120172 656208 120224 656260
rect 122104 656208 122156 656260
rect 210424 656208 210476 656260
rect 212356 656208 212408 656260
rect 512092 656208 512144 656260
rect 514024 656208 514076 656260
rect 184388 655664 184440 655716
rect 233240 655664 233292 655716
rect 350448 655664 350500 655716
rect 401600 655664 401652 655716
rect 464436 655664 464488 655716
rect 513380 655664 513432 655716
rect 42708 655596 42760 655648
rect 93860 655596 93912 655648
rect 97908 655596 97960 655648
rect 149060 655596 149112 655648
rect 156420 655596 156472 655648
rect 205640 655596 205692 655648
rect 238668 655596 238720 655648
rect 289820 655596 289872 655648
rect 293868 655596 293920 655648
rect 345020 655596 345072 655648
rect 378048 655596 378100 655648
rect 429292 655596 429344 655648
rect 436468 655596 436520 655648
rect 485780 655596 485832 655648
rect 518808 655596 518860 655648
rect 569960 655596 570012 655648
rect 13728 655528 13780 655580
rect 66260 655528 66312 655580
rect 70308 655528 70360 655580
rect 121460 655528 121512 655580
rect 126888 655528 126940 655580
rect 178040 655528 178092 655580
rect 209688 655528 209740 655580
rect 262220 655528 262272 655580
rect 266268 655528 266320 655580
rect 317420 655528 317472 655580
rect 322848 655528 322900 655580
rect 374000 655528 374052 655580
rect 408408 655528 408460 655580
rect 458180 655528 458232 655580
rect 489828 655528 489880 655580
rect 542360 655528 542412 655580
rect 400312 655188 400364 655240
rect 400956 655188 401008 655240
rect 204260 654304 204312 654356
rect 204996 654304 205048 654356
rect 434628 654032 434680 654084
rect 436468 654032 436520 654084
rect 15200 634720 15252 634772
rect 35900 634720 35952 634772
rect 36084 634720 36136 634772
rect 63592 634720 63644 634772
rect 64052 634720 64104 634772
rect 91928 634720 91980 634772
rect 92112 634720 92164 634772
rect 119620 634720 119672 634772
rect 122104 634720 122156 634772
rect 147956 634720 148008 634772
rect 148048 634720 148100 634772
rect 175924 634720 175976 634772
rect 176108 634720 176160 634772
rect 203616 634720 203668 634772
rect 204996 634720 205048 634772
rect 231952 634720 232004 634772
rect 232044 634720 232096 634772
rect 259920 634720 259972 634772
rect 260104 634720 260156 634772
rect 287612 634720 287664 634772
rect 288072 634720 288124 634772
rect 315948 634720 316000 634772
rect 316684 634720 316736 634772
rect 343916 634720 343968 634772
rect 344100 634720 344152 634772
rect 371608 634720 371660 634772
rect 372068 634720 372120 634772
rect 399944 634720 399996 634772
rect 400956 634720 401008 634772
rect 427912 634720 427964 634772
rect 428096 634720 428148 634772
rect 455604 634720 455656 634772
rect 456064 634720 456116 634772
rect 483940 634720 483992 634772
rect 484032 634720 484084 634772
rect 511908 634720 511960 634772
rect 514024 634720 514076 634772
rect 539600 634720 539652 634772
rect 540060 634720 540112 634772
rect 567936 634720 567988 634772
rect 16580 634652 16632 634704
rect 36636 634652 36688 634704
rect 44916 634652 44968 634704
rect 71136 634652 71188 634704
rect 82268 634652 82320 634704
rect 93124 634652 93176 634704
rect 110328 634652 110380 634704
rect 124864 634652 124916 634704
rect 128636 634652 128688 634704
rect 149704 634652 149756 634704
rect 156604 634652 156656 634704
rect 182824 634652 182876 634704
rect 194508 634652 194560 634704
rect 210424 634652 210476 634704
rect 212632 634652 212684 634704
rect 232504 634652 232556 634704
rect 240600 634652 240652 634704
rect 267004 634652 267056 634704
rect 278596 634652 278648 634704
rect 289084 634652 289136 634704
rect 306288 634652 306340 634704
rect 318064 634652 318116 634704
rect 324596 634652 324648 634704
rect 347044 634652 347096 634704
rect 362592 634652 362644 634704
rect 373264 634652 373316 634704
rect 390284 634652 390336 634704
rect 400864 634652 400916 634704
rect 408592 634652 408644 634704
rect 428464 634652 428516 634704
rect 436928 634652 436980 634704
rect 462964 634652 463016 634704
rect 474280 634652 474332 634704
rect 485044 634652 485096 634704
rect 502248 634652 502300 634704
rect 512644 634652 512696 634704
rect 520924 634652 520976 634704
rect 541624 634652 541676 634704
rect 26240 634584 26292 634636
rect 43536 634584 43588 634636
rect 54576 634584 54628 634636
rect 66904 634584 66956 634636
rect 138296 634584 138348 634636
rect 151084 634584 151136 634636
rect 166264 634584 166316 634636
rect 177304 634584 177356 634636
rect 222292 634584 222344 634636
rect 233976 634584 234028 634636
rect 250260 634584 250312 634636
rect 261484 634584 261536 634636
rect 334256 634584 334308 634636
rect 348424 634584 348476 634636
rect 418252 634584 418304 634636
rect 429844 634584 429896 634636
rect 446588 634584 446640 634636
rect 457444 634584 457496 634636
rect 530584 634584 530636 634636
rect 544384 634584 544436 634636
rect 558276 634040 558328 634092
rect 567476 634040 567528 634092
rect 548340 632680 548392 632732
rect 568028 632680 568080 632732
rect 212356 632272 212408 632324
rect 232688 632272 232740 632324
rect 296352 632272 296404 632324
rect 316776 632272 316828 632324
rect 408040 632272 408092 632324
rect 428648 632272 428700 632324
rect 492036 632272 492088 632324
rect 512736 632272 512788 632324
rect 148324 632204 148376 632256
rect 165712 632204 165764 632256
rect 175464 632204 175516 632256
rect 193680 632204 193732 632256
rect 203524 632204 203576 632256
rect 221372 632204 221424 632256
rect 260104 632204 260156 632256
rect 277676 632204 277728 632256
rect 287520 632204 287572 632256
rect 305368 632204 305420 632256
rect 345664 632204 345716 632256
rect 361672 632204 361724 632256
rect 371516 632204 371568 632256
rect 389364 632204 389416 632256
rect 399484 632204 399536 632256
rect 417700 632204 417752 632256
rect 456156 632204 456208 632256
rect 473360 632204 473412 632256
rect 483480 632204 483532 632256
rect 501696 632204 501748 632256
rect 36728 632136 36780 632188
rect 53656 632136 53708 632188
rect 64328 632136 64380 632188
rect 81440 632136 81492 632188
rect 91468 632136 91520 632188
rect 109684 632136 109736 632188
rect 119436 632136 119488 632188
rect 137652 632136 137704 632188
rect 156328 632136 156380 632188
rect 178684 632136 178736 632188
rect 232504 632136 232556 632188
rect 249708 632136 249760 632188
rect 268016 632136 268068 632188
rect 287704 632136 287756 632188
rect 315488 632136 315540 632188
rect 333704 632136 333756 632188
rect 352012 632136 352064 632188
rect 374644 632136 374696 632188
rect 428464 632136 428516 632188
rect 445668 632136 445720 632188
rect 464344 632136 464396 632188
rect 483664 632136 483716 632188
rect 511448 632136 511500 632188
rect 529664 632136 529716 632188
rect 541624 632136 541676 632188
rect 557540 632136 557592 632188
rect 3424 632068 3476 632120
rect 14464 632068 14516 632120
rect 16120 632068 16172 632120
rect 25688 632068 25740 632120
rect 36636 632068 36688 632120
rect 63316 632068 63368 632120
rect 66904 632068 66956 632120
rect 91100 632068 91152 632120
rect 93124 632068 93176 632120
rect 119344 632068 119396 632120
rect 124864 632068 124916 632120
rect 147312 632068 147364 632120
rect 148416 632068 148468 632120
rect 175372 632068 175424 632120
rect 177304 632068 177356 632120
rect 203340 632068 203392 632120
rect 204996 632068 205048 632120
rect 231032 632068 231084 632120
rect 232596 632068 232648 632120
rect 259368 632068 259420 632120
rect 260196 632068 260248 632120
rect 287336 632068 287388 632120
rect 289084 632068 289136 632120
rect 315028 632068 315080 632120
rect 316684 632068 316736 632120
rect 343364 632068 343416 632120
rect 344284 632068 344336 632120
rect 371332 632068 371384 632120
rect 373264 632068 373316 632120
rect 399024 632068 399076 632120
rect 400864 632068 400916 632120
rect 427360 632068 427412 632120
rect 428556 632068 428608 632120
rect 455328 632068 455380 632120
rect 456064 632068 456116 632120
rect 483020 632068 483072 632120
rect 485044 632068 485096 632120
rect 511356 632068 511408 632120
rect 512644 632068 512696 632120
rect 539324 632068 539376 632120
rect 540244 632068 540296 632120
rect 567200 632068 567252 632120
rect 15844 629280 15896 629332
rect 16120 629280 16172 629332
rect 42892 627240 42944 627292
rect 43628 627240 43680 627292
rect 63592 612756 63644 612808
rect 64328 612756 64380 612808
rect 455696 612756 455748 612808
rect 456156 612756 456208 612808
rect 428648 612008 428700 612060
rect 435732 612008 435784 612060
rect 232688 611940 232740 611992
rect 239772 611940 239824 611992
rect 287704 611872 287756 611924
rect 295708 611872 295760 611924
rect 316776 611872 316828 611924
rect 323676 611872 323728 611924
rect 483664 611736 483716 611788
rect 491668 611736 491720 611788
rect 512736 611736 512788 611788
rect 519636 611736 519688 611788
rect 13544 611260 13596 611312
rect 66260 611260 66312 611312
rect 70308 611260 70360 611312
rect 121460 611260 121512 611312
rect 126888 611260 126940 611312
rect 178040 611260 178092 611312
rect 209688 611260 209740 611312
rect 262220 611260 262272 611312
rect 266268 611260 266320 611312
rect 317420 611260 317472 611312
rect 322848 611260 322900 611312
rect 374000 611260 374052 611312
rect 405648 611260 405700 611312
rect 458180 611260 458232 611312
rect 489828 611260 489880 611312
rect 42708 611192 42760 611244
rect 93860 611192 93912 611244
rect 97908 611192 97960 611244
rect 149060 611192 149112 611244
rect 154488 611192 154540 611244
rect 205640 611192 205692 611244
rect 238668 611192 238720 611244
rect 289820 611192 289872 611244
rect 293868 611192 293920 611244
rect 345020 611192 345072 611244
rect 378048 611192 378100 611244
rect 429292 611192 429344 611244
rect 434628 611192 434680 611244
rect 485780 611192 485832 611244
rect 518808 611192 518860 611244
rect 182088 611124 182140 611176
rect 233240 611124 233292 611176
rect 350448 611124 350500 611176
rect 401600 611124 401652 611176
rect 462228 611124 462280 611176
rect 513380 611124 513432 611176
rect 539508 611260 539560 611312
rect 541624 611260 541676 611312
rect 542360 611124 542412 611176
rect 569960 611192 570012 611244
rect 15844 610648 15896 610700
rect 16580 610648 16632 610700
rect 35256 610648 35308 610700
rect 36728 610648 36780 610700
rect 547880 610648 547932 610700
rect 548156 610648 548208 610700
rect 71872 608540 71924 608592
rect 100024 608540 100076 608592
rect 25688 608472 25740 608524
rect 36636 608472 36688 608524
rect 42892 608472 42944 608524
rect 15292 608404 15344 608456
rect 43996 608404 44048 608456
rect 53656 608472 53708 608524
rect 66904 608472 66956 608524
rect 81992 608472 82044 608524
rect 93124 608472 93176 608524
rect 99472 608472 99524 608524
rect 127992 608540 128044 608592
rect 165988 608540 166040 608592
rect 177304 608540 177356 608592
rect 178684 608540 178736 608592
rect 184020 608540 184072 608592
rect 109684 608472 109736 608524
rect 124864 608472 124916 608524
rect 137652 608472 137704 608524
rect 148416 608472 148468 608524
rect 183652 608472 183704 608524
rect 211712 608540 211764 608592
rect 277676 608540 277728 608592
rect 289084 608540 289136 608592
rect 306012 608540 306064 608592
rect 316684 608540 316736 608592
rect 343364 608540 343416 608592
rect 345664 608540 345716 608592
rect 361672 608540 361724 608592
rect 373264 608540 373316 608592
rect 379612 608540 379664 608592
rect 408040 608540 408092 608592
rect 474004 608540 474056 608592
rect 485044 608540 485096 608592
rect 501696 608540 501748 608592
rect 512644 608540 512696 608592
rect 548156 608540 548208 608592
rect 557540 608540 557592 608592
rect 193680 608472 193732 608524
rect 204996 608472 205048 608524
rect 222016 608472 222068 608524
rect 232596 608472 232648 608524
rect 249708 608472 249760 608524
rect 260196 608472 260248 608524
rect 333704 608472 333756 608524
rect 344284 608472 344336 608524
rect 374644 608472 374696 608524
rect 379704 608472 379756 608524
rect 390008 608472 390060 608524
rect 400864 608472 400916 608524
rect 417700 608472 417752 608524
rect 428556 608472 428608 608524
rect 445668 608472 445720 608524
rect 456064 608472 456116 608524
rect 529664 608472 529716 608524
rect 540244 608472 540296 608524
rect 72056 608404 72108 608456
rect 127072 608404 127124 608456
rect 156052 608404 156104 608456
rect 238852 608404 238904 608456
rect 268016 608404 268068 608456
rect 323032 608404 323084 608456
rect 352012 608404 352064 608456
rect 434812 608404 434864 608456
rect 463700 608404 463752 608456
rect 518992 608404 519044 608456
rect 547880 608404 547932 608456
rect 3240 605820 3292 605872
rect 11704 605820 11756 605872
rect 71136 604596 71188 604648
rect 82268 604596 82320 604648
rect 99472 604596 99524 604648
rect 100392 604596 100444 604648
rect 183652 604596 183704 604648
rect 222292 604596 222344 604648
rect 267004 604596 267056 604648
rect 277952 604596 278004 604648
rect 295432 604596 295484 604648
rect 334256 604596 334308 604648
rect 352012 604596 352064 604648
rect 36636 604528 36688 604580
rect 53932 604528 53984 604580
rect 71872 604528 71924 604580
rect 109960 604528 110012 604580
rect 151084 604528 151136 604580
rect 156604 604528 156656 604580
rect 182824 604528 182876 604580
rect 193956 604528 194008 604580
rect 232504 604528 232556 604580
rect 26240 604460 26292 604512
rect 35440 604460 35492 604512
rect 66904 604460 66956 604512
rect 72608 604460 72660 604512
rect 93124 604460 93176 604512
rect 100300 604460 100352 604512
rect 100392 604460 100444 604512
rect 138296 604460 138348 604512
rect 149704 604460 149756 604512
rect 166264 604460 166316 604512
rect 177304 604460 177356 604512
rect 184296 604460 184348 604512
rect 233976 604460 234028 604512
rect 240600 604460 240652 604512
rect 267832 604528 267884 604580
rect 306288 604528 306340 604580
rect 347044 604528 347096 604580
rect 361948 604528 362000 604580
rect 379612 604596 379664 604648
rect 418252 604596 418304 604648
rect 462964 604596 463016 604648
rect 474280 604596 474332 604648
rect 491392 604596 491444 604648
rect 529940 604596 529992 604648
rect 390284 604528 390336 604580
rect 400956 604528 401008 604580
rect 408592 604528 408644 604580
rect 429844 604528 429896 604580
rect 436284 604528 436336 604580
rect 463792 604528 463844 604580
rect 502248 604528 502300 604580
rect 512644 604528 512696 604580
rect 520280 604528 520332 604580
rect 541624 604528 541676 604580
rect 250260 604460 250312 604512
rect 261484 604460 261536 604512
rect 268292 604460 268344 604512
rect 289084 604460 289136 604512
rect 296628 604460 296680 604512
rect 318064 604460 318116 604512
rect 324596 604460 324648 604512
rect 348424 604460 348476 604512
rect 352288 604460 352340 604512
rect 373264 604460 373316 604512
rect 380624 604460 380676 604512
rect 428464 604460 428516 604512
rect 445944 604460 445996 604512
rect 457444 604460 457496 604512
rect 464620 604460 464672 604512
rect 485044 604460 485096 604512
rect 492588 604460 492640 604512
rect 544384 604460 544436 604512
rect 548616 604460 548668 604512
rect 558276 604460 558328 604512
rect 120172 602216 120224 602268
rect 122104 602216 122156 602268
rect 124864 602216 124916 602268
rect 128268 602216 128320 602268
rect 210424 602216 210476 602268
rect 212356 602216 212408 602268
rect 512092 602216 512144 602268
rect 514024 602216 514076 602268
rect 182088 601808 182140 601860
rect 233240 601808 233292 601860
rect 350448 601808 350500 601860
rect 401600 601808 401652 601860
rect 462228 601808 462280 601860
rect 513380 601808 513432 601860
rect 42708 601740 42760 601792
rect 93860 601740 93912 601792
rect 97908 601740 97960 601792
rect 149060 601740 149112 601792
rect 154488 601740 154540 601792
rect 205640 601740 205692 601792
rect 238668 601740 238720 601792
rect 289820 601740 289872 601792
rect 293868 601740 293920 601792
rect 345020 601740 345072 601792
rect 378048 601740 378100 601792
rect 429292 601740 429344 601792
rect 434628 601740 434680 601792
rect 485780 601740 485832 601792
rect 518808 601740 518860 601792
rect 569960 601740 570012 601792
rect 13544 601672 13596 601724
rect 66260 601672 66312 601724
rect 70308 601672 70360 601724
rect 121460 601672 121512 601724
rect 126888 601672 126940 601724
rect 178040 601672 178092 601724
rect 209688 601672 209740 601724
rect 262220 601672 262272 601724
rect 266268 601672 266320 601724
rect 317420 601672 317472 601724
rect 322848 601672 322900 601724
rect 374000 601672 374052 601724
rect 405648 601672 405700 601724
rect 458180 601672 458232 601724
rect 489828 601672 489880 601724
rect 542360 601672 542412 601724
rect 204260 599224 204312 599276
rect 204996 599224 205048 599276
rect 15200 580932 15252 580984
rect 35900 580932 35952 580984
rect 36084 580932 36136 580984
rect 63592 580932 63644 580984
rect 64052 580932 64104 580984
rect 91928 580932 91980 580984
rect 92112 580932 92164 580984
rect 119620 580932 119672 580984
rect 122104 580932 122156 580984
rect 147956 580932 148008 580984
rect 148048 580932 148100 580984
rect 175924 580932 175976 580984
rect 176108 580932 176160 580984
rect 203616 580932 203668 580984
rect 204996 580932 205048 580984
rect 231952 580932 232004 580984
rect 232044 580932 232096 580984
rect 259920 580932 259972 580984
rect 260104 580932 260156 580984
rect 287612 580932 287664 580984
rect 288072 580932 288124 580984
rect 315948 580932 316000 580984
rect 316684 580932 316736 580984
rect 343916 580932 343968 580984
rect 344100 580932 344152 580984
rect 371608 580932 371660 580984
rect 372068 580932 372120 580984
rect 399944 580932 399996 580984
rect 400864 580932 400916 580984
rect 427912 580932 427964 580984
rect 428096 580932 428148 580984
rect 455604 580932 455656 580984
rect 456064 580932 456116 580984
rect 483940 580932 483992 580984
rect 484032 580932 484084 580984
rect 511908 580932 511960 580984
rect 514024 580932 514076 580984
rect 539600 580932 539652 580984
rect 540060 580932 540112 580984
rect 567936 580932 567988 580984
rect 16580 580864 16632 580916
rect 36636 580864 36688 580916
rect 44916 580864 44968 580916
rect 71136 580864 71188 580916
rect 82268 580864 82320 580916
rect 93124 580864 93176 580916
rect 110236 580864 110288 580916
rect 124864 580864 124916 580916
rect 128636 580864 128688 580916
rect 149704 580864 149756 580916
rect 156604 580864 156656 580916
rect 182824 580864 182876 580916
rect 194508 580864 194560 580916
rect 210424 580864 210476 580916
rect 212632 580864 212684 580916
rect 232504 580864 232556 580916
rect 240600 580864 240652 580916
rect 267004 580864 267056 580916
rect 278596 580864 278648 580916
rect 289084 580864 289136 580916
rect 306288 580864 306340 580916
rect 318064 580864 318116 580916
rect 324596 580864 324648 580916
rect 347044 580864 347096 580916
rect 362592 580864 362644 580916
rect 373264 580864 373316 580916
rect 390284 580864 390336 580916
rect 400956 580864 401008 580916
rect 408592 580864 408644 580916
rect 428464 580864 428516 580916
rect 436928 580864 436980 580916
rect 462964 580864 463016 580916
rect 474280 580864 474332 580916
rect 485044 580864 485096 580916
rect 502248 580864 502300 580916
rect 512644 580864 512696 580916
rect 520924 580864 520976 580916
rect 541624 580864 541676 580916
rect 26240 580796 26292 580848
rect 43536 580796 43588 580848
rect 54576 580796 54628 580848
rect 66904 580796 66956 580848
rect 138296 580796 138348 580848
rect 151084 580796 151136 580848
rect 166264 580796 166316 580848
rect 177304 580796 177356 580848
rect 222292 580796 222344 580848
rect 233976 580796 234028 580848
rect 250260 580796 250312 580848
rect 261484 580796 261536 580848
rect 334256 580796 334308 580848
rect 348424 580796 348476 580848
rect 418252 580796 418304 580848
rect 429844 580796 429896 580848
rect 446588 580796 446640 580848
rect 457444 580796 457496 580848
rect 530584 580796 530636 580848
rect 544384 580796 544436 580848
rect 558276 580252 558328 580304
rect 567476 580252 567528 580304
rect 548340 578892 548392 578944
rect 568028 578892 568080 578944
rect 212264 578416 212316 578468
rect 232688 578416 232740 578468
rect 296352 578416 296404 578468
rect 316776 578416 316828 578468
rect 408040 578416 408092 578468
rect 428648 578416 428700 578468
rect 492036 578416 492088 578468
rect 512736 578416 512788 578468
rect 148416 578348 148468 578400
rect 165620 578348 165672 578400
rect 175464 578348 175516 578400
rect 193680 578348 193732 578400
rect 203524 578348 203576 578400
rect 221372 578348 221424 578400
rect 260196 578348 260248 578400
rect 277676 578348 277728 578400
rect 287520 578348 287572 578400
rect 305368 578348 305420 578400
rect 345664 578348 345716 578400
rect 361672 578348 361724 578400
rect 371516 578348 371568 578400
rect 389364 578348 389416 578400
rect 399484 578348 399536 578400
rect 417700 578348 417752 578400
rect 456156 578348 456208 578400
rect 473544 578348 473596 578400
rect 483480 578348 483532 578400
rect 501696 578348 501748 578400
rect 36728 578280 36780 578332
rect 53656 578280 53708 578332
rect 64328 578280 64380 578332
rect 81440 578280 81492 578332
rect 91468 578280 91520 578332
rect 109684 578280 109736 578332
rect 119436 578280 119488 578332
rect 137652 578280 137704 578332
rect 156328 578280 156380 578332
rect 178684 578280 178736 578332
rect 232504 578280 232556 578332
rect 249708 578280 249760 578332
rect 268016 578280 268068 578332
rect 287704 578280 287756 578332
rect 315488 578280 315540 578332
rect 333704 578280 333756 578332
rect 352012 578280 352064 578332
rect 374644 578280 374696 578332
rect 428464 578280 428516 578332
rect 445668 578280 445720 578332
rect 464344 578280 464396 578332
rect 483664 578280 483716 578332
rect 511448 578280 511500 578332
rect 529664 578280 529716 578332
rect 541624 578280 541676 578332
rect 557540 578280 557592 578332
rect 15844 578212 15896 578264
rect 25688 578212 25740 578264
rect 36636 578212 36688 578264
rect 63316 578212 63368 578264
rect 66904 578212 66956 578264
rect 91100 578212 91152 578264
rect 93124 578212 93176 578264
rect 119344 578212 119396 578264
rect 124864 578212 124916 578264
rect 147312 578212 147364 578264
rect 148324 578212 148376 578264
rect 175280 578212 175332 578264
rect 177304 578212 177356 578264
rect 203340 578212 203392 578264
rect 204996 578212 205048 578264
rect 231032 578212 231084 578264
rect 232596 578212 232648 578264
rect 259368 578212 259420 578264
rect 260104 578212 260156 578264
rect 287336 578212 287388 578264
rect 289084 578212 289136 578264
rect 315028 578212 315080 578264
rect 316684 578212 316736 578264
rect 343364 578212 343416 578264
rect 344284 578212 344336 578264
rect 371332 578212 371384 578264
rect 373264 578212 373316 578264
rect 399024 578212 399076 578264
rect 400864 578212 400916 578264
rect 427360 578212 427412 578264
rect 428556 578212 428608 578264
rect 455328 578212 455380 578264
rect 456064 578212 456116 578264
rect 483204 578212 483256 578264
rect 485044 578212 485096 578264
rect 511356 578212 511408 578264
rect 512644 578212 512696 578264
rect 539324 578212 539376 578264
rect 540244 578212 540296 578264
rect 567200 578212 567252 578264
rect 15292 575220 15344 575272
rect 15936 575220 15988 575272
rect 42892 571208 42944 571260
rect 43628 571208 43680 571260
rect 147680 562300 147732 562352
rect 148416 562300 148468 562352
rect 259736 562300 259788 562352
rect 260196 562300 260248 562352
rect 455696 562300 455748 562352
rect 456156 562300 456208 562352
rect 287704 558832 287756 558884
rect 295708 558832 295760 558884
rect 316776 558832 316828 558884
rect 323676 558832 323728 558884
rect 63592 558288 63644 558340
rect 64328 558288 64380 558340
rect 232688 558152 232740 558204
rect 239772 558152 239824 558204
rect 428648 558152 428700 558204
rect 435732 558152 435784 558204
rect 483664 558152 483716 558204
rect 491668 558152 491720 558204
rect 512736 558152 512788 558204
rect 519636 558152 519688 558204
rect 13544 557472 13596 557524
rect 66260 557472 66312 557524
rect 70308 557472 70360 557524
rect 121460 557472 121512 557524
rect 126888 557472 126940 557524
rect 178040 557472 178092 557524
rect 209688 557472 209740 557524
rect 262220 557472 262272 557524
rect 266268 557472 266320 557524
rect 317420 557472 317472 557524
rect 322848 557472 322900 557524
rect 374000 557472 374052 557524
rect 405648 557472 405700 557524
rect 458180 557472 458232 557524
rect 489828 557472 489880 557524
rect 542360 557472 542412 557524
rect 42708 557404 42760 557456
rect 93860 557404 93912 557456
rect 97908 557404 97960 557456
rect 149060 557404 149112 557456
rect 154488 557404 154540 557456
rect 205640 557404 205692 557456
rect 238668 557404 238720 557456
rect 289820 557404 289872 557456
rect 293868 557404 293920 557456
rect 182088 557336 182140 557388
rect 233240 557336 233292 557388
rect 343548 557404 343600 557456
rect 345664 557404 345716 557456
rect 378048 557404 378100 557456
rect 429292 557404 429344 557456
rect 434628 557404 434680 557456
rect 485780 557404 485832 557456
rect 518808 557404 518860 557456
rect 569960 557404 570012 557456
rect 345020 557336 345072 557388
rect 350448 557336 350500 557388
rect 401600 557336 401652 557388
rect 462228 557336 462280 557388
rect 513380 557336 513432 557388
rect 539508 556724 539560 556776
rect 541624 556724 541676 556776
rect 35256 556656 35308 556708
rect 36728 556656 36780 556708
rect 15844 556180 15896 556232
rect 16580 556180 16632 556232
rect 547880 556112 547932 556164
rect 548156 556112 548208 556164
rect 71872 554684 71924 554736
rect 100024 554684 100076 554736
rect 25688 554616 25740 554668
rect 36636 554616 36688 554668
rect 42892 554616 42944 554668
rect 15292 554548 15344 554600
rect 43996 554548 44048 554600
rect 53656 554616 53708 554668
rect 66904 554616 66956 554668
rect 81992 554616 82044 554668
rect 93124 554616 93176 554668
rect 99472 554616 99524 554668
rect 127992 554684 128044 554736
rect 165988 554684 166040 554736
rect 177304 554684 177356 554736
rect 178684 554684 178736 554736
rect 184020 554684 184072 554736
rect 109684 554616 109736 554668
rect 124864 554616 124916 554668
rect 137652 554616 137704 554668
rect 148324 554616 148376 554668
rect 183652 554616 183704 554668
rect 211712 554684 211764 554736
rect 277676 554684 277728 554736
rect 289084 554684 289136 554736
rect 306012 554684 306064 554736
rect 316684 554684 316736 554736
rect 361672 554684 361724 554736
rect 373264 554684 373316 554736
rect 374644 554684 374696 554736
rect 379704 554684 379756 554736
rect 193680 554616 193732 554668
rect 204996 554616 205048 554668
rect 222016 554616 222068 554668
rect 232596 554616 232648 554668
rect 249708 554616 249760 554668
rect 260104 554616 260156 554668
rect 333704 554616 333756 554668
rect 344284 554616 344336 554668
rect 379612 554616 379664 554668
rect 408040 554684 408092 554736
rect 474004 554684 474056 554736
rect 485044 554684 485096 554736
rect 501696 554684 501748 554736
rect 512644 554684 512696 554736
rect 548156 554684 548208 554736
rect 557540 554684 557592 554736
rect 390008 554616 390060 554668
rect 400864 554616 400916 554668
rect 417700 554616 417752 554668
rect 428556 554616 428608 554668
rect 445668 554616 445720 554668
rect 456064 554616 456116 554668
rect 529664 554616 529716 554668
rect 540244 554616 540296 554668
rect 72056 554548 72108 554600
rect 127072 554548 127124 554600
rect 156052 554548 156104 554600
rect 238852 554548 238904 554600
rect 268016 554548 268068 554600
rect 323032 554548 323084 554600
rect 352012 554548 352064 554600
rect 434812 554548 434864 554600
rect 463700 554548 463752 554600
rect 518992 554548 519044 554600
rect 547880 554548 547932 554600
rect 3332 553392 3384 553444
rect 10324 553392 10376 553444
rect 26240 550876 26292 550928
rect 35440 550876 35492 550928
rect 352012 550808 352064 550860
rect 71136 550740 71188 550792
rect 82268 550740 82320 550792
rect 99472 550740 99524 550792
rect 100392 550740 100444 550792
rect 183652 550740 183704 550792
rect 222292 550740 222344 550792
rect 267832 550740 267884 550792
rect 36636 550672 36688 550724
rect 53932 550672 53984 550724
rect 71872 550672 71924 550724
rect 109960 550672 110012 550724
rect 151084 550672 151136 550724
rect 156604 550672 156656 550724
rect 182824 550672 182876 550724
rect 193956 550672 194008 550724
rect 232504 550672 232556 550724
rect 66904 550604 66956 550656
rect 72608 550604 72660 550656
rect 93124 550604 93176 550656
rect 100300 550604 100352 550656
rect 100392 550604 100444 550656
rect 138296 550604 138348 550656
rect 149704 550604 149756 550656
rect 166264 550604 166316 550656
rect 177304 550604 177356 550656
rect 184296 550604 184348 550656
rect 233976 550604 234028 550656
rect 240600 550604 240652 550656
rect 267004 550672 267056 550724
rect 295432 550740 295484 550792
rect 334256 550740 334308 550792
rect 345664 550740 345716 550792
rect 250260 550604 250312 550656
rect 261484 550604 261536 550656
rect 268292 550604 268344 550656
rect 306288 550672 306340 550724
rect 277952 550604 278004 550656
rect 289084 550604 289136 550656
rect 296628 550604 296680 550656
rect 318064 550604 318116 550656
rect 324596 550604 324648 550656
rect 347044 550604 347096 550656
rect 352288 550604 352340 550656
rect 463792 550808 463844 550860
rect 379612 550740 379664 550792
rect 418252 550740 418304 550792
rect 390284 550672 390336 550724
rect 400956 550672 401008 550724
rect 408592 550672 408644 550724
rect 429844 550672 429896 550724
rect 436284 550672 436336 550724
rect 457444 550672 457496 550724
rect 464620 550672 464672 550724
rect 491392 550740 491444 550792
rect 361948 550604 362000 550656
rect 373264 550604 373316 550656
rect 380624 550604 380676 550656
rect 428464 550604 428516 550656
rect 445944 550604 445996 550656
rect 462964 550604 463016 550656
rect 474280 550604 474332 550656
rect 485044 550604 485096 550656
rect 492588 550604 492640 550656
rect 502248 550672 502300 550724
rect 529940 550740 529992 550792
rect 541624 550672 541676 550724
rect 514024 550604 514076 550656
rect 520280 550604 520332 550656
rect 544384 550604 544436 550656
rect 548616 550604 548668 550656
rect 558276 550604 558328 550656
rect 120080 548224 120132 548276
rect 122104 548224 122156 548276
rect 124864 548224 124916 548276
rect 128268 548224 128320 548276
rect 210424 548224 210476 548276
rect 212356 548224 212408 548276
rect 204260 547068 204312 547120
rect 204996 547068 205048 547120
rect 13544 529864 13596 529916
rect 66260 529864 66312 529916
rect 70308 529864 70360 529916
rect 121460 529864 121512 529916
rect 126888 529864 126940 529916
rect 178040 529864 178092 529916
rect 209688 529864 209740 529916
rect 262220 529864 262272 529916
rect 266268 529864 266320 529916
rect 317420 529864 317472 529916
rect 322848 529864 322900 529916
rect 374000 529864 374052 529916
rect 405648 529864 405700 529916
rect 458180 529864 458232 529916
rect 489828 529864 489880 529916
rect 542360 529864 542412 529916
rect 42708 529796 42760 529848
rect 93860 529796 93912 529848
rect 97908 529796 97960 529848
rect 149060 529796 149112 529848
rect 154488 529796 154540 529848
rect 205640 529796 205692 529848
rect 238668 529796 238720 529848
rect 289820 529796 289872 529848
rect 293868 529796 293920 529848
rect 345020 529796 345072 529848
rect 378048 529796 378100 529848
rect 429292 529796 429344 529848
rect 434628 529796 434680 529848
rect 485780 529796 485832 529848
rect 518808 529796 518860 529848
rect 569960 529796 570012 529848
rect 182088 529728 182140 529780
rect 233240 529728 233292 529780
rect 350448 529728 350500 529780
rect 401600 529728 401652 529780
rect 462228 529728 462280 529780
rect 513380 529728 513432 529780
rect 2780 527144 2832 527196
rect 4804 527144 4856 527196
rect 15200 527076 15252 527128
rect 35900 527076 35952 527128
rect 36084 527076 36136 527128
rect 63592 527076 63644 527128
rect 64052 527076 64104 527128
rect 91928 527076 91980 527128
rect 92112 527076 92164 527128
rect 119620 527076 119672 527128
rect 122104 527076 122156 527128
rect 147956 527076 148008 527128
rect 148048 527076 148100 527128
rect 175924 527076 175976 527128
rect 176108 527076 176160 527128
rect 203616 527076 203668 527128
rect 204996 527076 205048 527128
rect 231952 527076 232004 527128
rect 232044 527076 232096 527128
rect 259920 527076 259972 527128
rect 260104 527076 260156 527128
rect 287612 527076 287664 527128
rect 288072 527076 288124 527128
rect 315948 527076 316000 527128
rect 316684 527076 316736 527128
rect 343916 527076 343968 527128
rect 344100 527076 344152 527128
rect 371608 527076 371660 527128
rect 372068 527076 372120 527128
rect 399944 527076 399996 527128
rect 400864 527076 400916 527128
rect 427912 527076 427964 527128
rect 428096 527076 428148 527128
rect 455604 527076 455656 527128
rect 456064 527076 456116 527128
rect 483940 527076 483992 527128
rect 484032 527076 484084 527128
rect 511908 527076 511960 527128
rect 512092 527076 512144 527128
rect 539600 527076 539652 527128
rect 540060 527076 540112 527128
rect 567936 527076 567988 527128
rect 16580 527008 16632 527060
rect 36636 527008 36688 527060
rect 44916 527008 44968 527060
rect 71136 527008 71188 527060
rect 82268 527008 82320 527060
rect 93124 527008 93176 527060
rect 110328 527008 110380 527060
rect 124864 527008 124916 527060
rect 128636 527008 128688 527060
rect 149704 527008 149756 527060
rect 156604 527008 156656 527060
rect 182824 527008 182876 527060
rect 194508 527008 194560 527060
rect 210424 527008 210476 527060
rect 212632 527008 212684 527060
rect 232504 527008 232556 527060
rect 240600 527008 240652 527060
rect 267004 527008 267056 527060
rect 278596 527008 278648 527060
rect 289084 527008 289136 527060
rect 306288 527008 306340 527060
rect 318064 527008 318116 527060
rect 324596 527008 324648 527060
rect 345664 527008 345716 527060
rect 362592 527008 362644 527060
rect 373264 527008 373316 527060
rect 390284 527008 390336 527060
rect 400956 527008 401008 527060
rect 408592 527008 408644 527060
rect 428464 527008 428516 527060
rect 436928 527008 436980 527060
rect 462964 527008 463016 527060
rect 474280 527008 474332 527060
rect 485044 527008 485096 527060
rect 502248 527008 502300 527060
rect 514024 527008 514076 527060
rect 520924 527008 520976 527060
rect 541624 527008 541676 527060
rect 26240 526940 26292 526992
rect 43536 526940 43588 526992
rect 54576 526940 54628 526992
rect 66904 526940 66956 526992
rect 138296 526940 138348 526992
rect 151084 526940 151136 526992
rect 166264 526940 166316 526992
rect 177304 526940 177356 526992
rect 222292 526940 222344 526992
rect 233976 526940 234028 526992
rect 250260 526940 250312 526992
rect 261484 526940 261536 526992
rect 334256 526940 334308 526992
rect 347044 526940 347096 526992
rect 418252 526940 418304 526992
rect 429844 526940 429896 526992
rect 446588 526940 446640 526992
rect 457444 526940 457496 526992
rect 530584 526940 530636 526992
rect 544384 526940 544436 526992
rect 558276 526396 558328 526448
rect 567476 526396 567528 526448
rect 548340 523676 548392 523728
rect 568028 523676 568080 523728
rect 212356 523200 212408 523252
rect 232688 523200 232740 523252
rect 296352 523200 296404 523252
rect 316776 523200 316828 523252
rect 408040 523200 408092 523252
rect 428648 523200 428700 523252
rect 492036 523200 492088 523252
rect 512736 523200 512788 523252
rect 148416 523132 148468 523184
rect 165712 523132 165764 523184
rect 175464 523132 175516 523184
rect 193680 523132 193732 523184
rect 203524 523132 203576 523184
rect 221372 523132 221424 523184
rect 260196 523132 260248 523184
rect 277676 523132 277728 523184
rect 287520 523132 287572 523184
rect 305368 523132 305420 523184
rect 345664 523132 345716 523184
rect 361672 523132 361724 523184
rect 371516 523132 371568 523184
rect 389364 523132 389416 523184
rect 399484 523132 399536 523184
rect 417700 523132 417752 523184
rect 456156 523132 456208 523184
rect 473360 523132 473412 523184
rect 483480 523132 483532 523184
rect 501696 523132 501748 523184
rect 36636 523064 36688 523116
rect 53656 523064 53708 523116
rect 64328 523064 64380 523116
rect 81440 523064 81492 523116
rect 91468 523064 91520 523116
rect 109684 523064 109736 523116
rect 119436 523064 119488 523116
rect 137652 523064 137704 523116
rect 156328 523064 156380 523116
rect 178684 523064 178736 523116
rect 232504 523064 232556 523116
rect 249708 523064 249760 523116
rect 268016 523064 268068 523116
rect 287704 523064 287756 523116
rect 315488 523064 315540 523116
rect 333704 523064 333756 523116
rect 352012 523064 352064 523116
rect 374644 523064 374696 523116
rect 428464 523064 428516 523116
rect 445668 523064 445720 523116
rect 464344 523064 464396 523116
rect 483664 523064 483716 523116
rect 511448 523064 511500 523116
rect 529664 523064 529716 523116
rect 541624 523064 541676 523116
rect 557540 523064 557592 523116
rect 15108 522996 15160 523048
rect 25688 522996 25740 523048
rect 36728 522996 36780 523048
rect 63316 522996 63368 523048
rect 66904 522996 66956 523048
rect 91100 522996 91152 523048
rect 93124 522996 93176 523048
rect 119344 522996 119396 523048
rect 124864 522996 124916 523048
rect 147312 522996 147364 523048
rect 148324 522996 148376 523048
rect 175372 522996 175424 523048
rect 177304 522996 177356 523048
rect 203340 522996 203392 523048
rect 204996 522996 205048 523048
rect 231032 522996 231084 523048
rect 232596 522996 232648 523048
rect 259368 522996 259420 523048
rect 260104 522996 260156 523048
rect 287336 522996 287388 523048
rect 289084 522996 289136 523048
rect 315028 522996 315080 523048
rect 316684 522996 316736 523048
rect 343364 522996 343416 523048
rect 344284 522996 344336 523048
rect 371332 522996 371384 523048
rect 373264 522996 373316 523048
rect 399024 522996 399076 523048
rect 400864 522996 400916 523048
rect 427360 522996 427412 523048
rect 428556 522996 428608 523048
rect 455328 522996 455380 523048
rect 456064 522996 456116 523048
rect 483020 522996 483072 523048
rect 485044 522996 485096 523048
rect 511356 522996 511408 523048
rect 512644 522996 512696 523048
rect 539324 522996 539376 523048
rect 540244 522996 540296 523048
rect 567200 522996 567252 523048
rect 42708 520276 42760 520328
rect 93860 520276 93912 520328
rect 97908 520276 97960 520328
rect 149060 520276 149112 520328
rect 155868 520276 155920 520328
rect 205640 520276 205692 520328
rect 209688 520276 209740 520328
rect 262220 520276 262272 520328
rect 266268 520276 266320 520328
rect 317420 520276 317472 520328
rect 322848 520276 322900 520328
rect 374000 520276 374052 520328
rect 378048 520276 378100 520328
rect 429292 520276 429344 520328
rect 434628 520276 434680 520328
rect 485780 520276 485832 520328
rect 489828 520276 489880 520328
rect 542360 520276 542412 520328
rect 154488 518848 154540 518900
rect 155868 518848 155920 518900
rect 42892 514020 42944 514072
rect 43628 514020 43680 514072
rect 63592 505588 63644 505640
rect 64328 505588 64380 505640
rect 147680 505588 147732 505640
rect 148416 505588 148468 505640
rect 259736 505588 259788 505640
rect 260196 505588 260248 505640
rect 455696 505588 455748 505640
rect 456156 505588 456208 505640
rect 287704 504568 287756 504620
rect 295708 504568 295760 504620
rect 428648 504364 428700 504416
rect 435732 504364 435784 504416
rect 483664 504296 483716 504348
rect 491668 504296 491720 504348
rect 512736 504296 512788 504348
rect 519636 504296 519688 504348
rect 232688 504228 232740 504280
rect 239772 504228 239824 504280
rect 316776 503752 316828 503804
rect 323676 503752 323728 503804
rect 13544 503616 13596 503668
rect 66260 503616 66312 503668
rect 70308 503616 70360 503668
rect 121460 503616 121512 503668
rect 126888 503616 126940 503668
rect 178040 503616 178092 503668
rect 182088 503616 182140 503668
rect 233240 503616 233292 503668
rect 238668 503616 238720 503668
rect 289820 503616 289872 503668
rect 293868 503616 293920 503668
rect 345020 503616 345072 503668
rect 350448 503616 350500 503668
rect 401600 503616 401652 503668
rect 405648 503616 405700 503668
rect 458180 503616 458232 503668
rect 462228 503616 462280 503668
rect 513380 503616 513432 503668
rect 518808 503616 518860 503668
rect 569960 503616 570012 503668
rect 539508 503548 539560 503600
rect 541624 503548 541676 503600
rect 15108 502664 15160 502716
rect 16580 502664 16632 502716
rect 547880 502664 547932 502716
rect 548156 502664 548208 502716
rect 35256 502256 35308 502308
rect 36636 502256 36688 502308
rect 71872 500896 71924 500948
rect 100024 500896 100076 500948
rect 25688 500828 25740 500880
rect 36728 500828 36780 500880
rect 42892 500828 42944 500880
rect 15292 500760 15344 500812
rect 43996 500760 44048 500812
rect 53656 500828 53708 500880
rect 66904 500828 66956 500880
rect 81992 500828 82044 500880
rect 93124 500828 93176 500880
rect 99472 500828 99524 500880
rect 127992 500896 128044 500948
rect 165988 500896 166040 500948
rect 177304 500896 177356 500948
rect 178684 500896 178736 500948
rect 184020 500896 184072 500948
rect 109684 500828 109736 500880
rect 124864 500828 124916 500880
rect 137652 500828 137704 500880
rect 148324 500828 148376 500880
rect 183652 500828 183704 500880
rect 211712 500896 211764 500948
rect 277676 500896 277728 500948
rect 289084 500896 289136 500948
rect 306012 500896 306064 500948
rect 316684 500896 316736 500948
rect 343364 500896 343416 500948
rect 345664 500896 345716 500948
rect 361672 500896 361724 500948
rect 373264 500896 373316 500948
rect 379612 500896 379664 500948
rect 408040 500896 408092 500948
rect 474004 500896 474056 500948
rect 485044 500896 485096 500948
rect 501696 500896 501748 500948
rect 512644 500896 512696 500948
rect 548156 500896 548208 500948
rect 557540 500896 557592 500948
rect 193680 500828 193732 500880
rect 204996 500828 205048 500880
rect 222016 500828 222068 500880
rect 232596 500828 232648 500880
rect 249708 500828 249760 500880
rect 260104 500828 260156 500880
rect 333704 500828 333756 500880
rect 344284 500828 344336 500880
rect 374644 500828 374696 500880
rect 379704 500828 379756 500880
rect 390008 500828 390060 500880
rect 400864 500828 400916 500880
rect 417700 500828 417752 500880
rect 428556 500828 428608 500880
rect 445668 500828 445720 500880
rect 456064 500828 456116 500880
rect 529664 500828 529716 500880
rect 540244 500828 540296 500880
rect 72056 500760 72108 500812
rect 127072 500760 127124 500812
rect 156052 500760 156104 500812
rect 238852 500760 238904 500812
rect 268016 500760 268068 500812
rect 323032 500760 323084 500812
rect 352012 500760 352064 500812
rect 434812 500760 434864 500812
rect 463700 500760 463752 500812
rect 518992 500760 519044 500812
rect 547880 500760 547932 500812
rect 71136 496952 71188 497004
rect 82268 496952 82320 497004
rect 184204 496952 184256 497004
rect 222292 496952 222344 497004
rect 267004 496952 267056 497004
rect 277952 496952 278004 497004
rect 296168 496952 296220 497004
rect 334256 496952 334308 497004
rect 352196 496952 352248 497004
rect 26240 496884 26292 496936
rect 35440 496884 35492 496936
rect 36636 496884 36688 496936
rect 53932 496884 53984 496936
rect 72240 496884 72292 496936
rect 109960 496884 110012 496936
rect 151084 496884 151136 496936
rect 156604 496884 156656 496936
rect 182824 496884 182876 496936
rect 193956 496884 194008 496936
rect 232504 496884 232556 496936
rect 66904 496816 66956 496868
rect 72608 496816 72660 496868
rect 93124 496816 93176 496868
rect 100300 496816 100352 496868
rect 100208 496748 100260 496800
rect 138296 496816 138348 496868
rect 149704 496816 149756 496868
rect 166264 496816 166316 496868
rect 177304 496816 177356 496868
rect 184296 496816 184348 496868
rect 233976 496816 234028 496868
rect 240600 496816 240652 496868
rect 268200 496884 268252 496936
rect 306288 496884 306340 496936
rect 345664 496884 345716 496936
rect 361948 496884 362000 496936
rect 380256 496952 380308 497004
rect 418252 496952 418304 497004
rect 464160 496952 464212 497004
rect 390284 496884 390336 496936
rect 400956 496884 401008 496936
rect 408592 496884 408644 496936
rect 429844 496884 429896 496936
rect 436284 496884 436336 496936
rect 457444 496884 457496 496936
rect 464620 496884 464672 496936
rect 485044 496952 485096 497004
rect 492588 496952 492640 497004
rect 502248 496884 502300 496936
rect 514024 496884 514076 496936
rect 520280 496884 520332 496936
rect 250260 496816 250312 496868
rect 261484 496816 261536 496868
rect 268292 496816 268344 496868
rect 289084 496816 289136 496868
rect 296628 496816 296680 496868
rect 318064 496816 318116 496868
rect 324596 496816 324648 496868
rect 347044 496816 347096 496868
rect 352288 496816 352340 496868
rect 373264 496816 373316 496868
rect 380624 496816 380676 496868
rect 428464 496816 428516 496868
rect 445944 496816 445996 496868
rect 462964 496816 463016 496868
rect 474280 496816 474332 496868
rect 492128 496816 492180 496868
rect 529940 496816 529992 496868
rect 541624 496816 541676 496868
rect 558276 496816 558328 496868
rect 120172 494232 120224 494284
rect 122104 494232 122156 494284
rect 124864 494232 124916 494284
rect 128268 494232 128320 494284
rect 210424 494232 210476 494284
rect 212356 494232 212408 494284
rect 544384 494028 544436 494080
rect 548340 494028 548392 494080
rect 204260 492056 204312 492108
rect 204996 492056 205048 492108
rect 13544 476008 13596 476060
rect 66260 476008 66312 476060
rect 70308 476008 70360 476060
rect 121460 476008 121512 476060
rect 126888 476008 126940 476060
rect 178040 476008 178092 476060
rect 209688 476008 209740 476060
rect 262220 476008 262272 476060
rect 266268 476008 266320 476060
rect 317420 476008 317472 476060
rect 322848 476008 322900 476060
rect 374000 476008 374052 476060
rect 405648 476008 405700 476060
rect 458180 476008 458232 476060
rect 489828 476008 489880 476060
rect 542360 476008 542412 476060
rect 42708 475940 42760 475992
rect 93860 475940 93912 475992
rect 97908 475940 97960 475992
rect 149060 475940 149112 475992
rect 154488 475940 154540 475992
rect 205640 475940 205692 475992
rect 238668 475940 238720 475992
rect 289820 475940 289872 475992
rect 293868 475940 293920 475992
rect 345020 475940 345072 475992
rect 378048 475940 378100 475992
rect 429292 475940 429344 475992
rect 462228 475940 462280 475992
rect 513380 475940 513432 475992
rect 518808 475940 518860 475992
rect 569960 475940 570012 475992
rect 182088 475872 182140 475924
rect 233240 475872 233292 475924
rect 350448 475872 350500 475924
rect 401600 475872 401652 475924
rect 434628 475872 434680 475924
rect 485780 475872 485832 475924
rect 15200 473288 15252 473340
rect 35900 473288 35952 473340
rect 36084 473288 36136 473340
rect 63592 473288 63644 473340
rect 64052 473288 64104 473340
rect 91928 473288 91980 473340
rect 92112 473288 92164 473340
rect 119620 473288 119672 473340
rect 122104 473288 122156 473340
rect 147956 473288 148008 473340
rect 148048 473288 148100 473340
rect 175924 473288 175976 473340
rect 176108 473288 176160 473340
rect 203616 473288 203668 473340
rect 204996 473288 205048 473340
rect 231952 473288 232004 473340
rect 232044 473288 232096 473340
rect 259920 473288 259972 473340
rect 260104 473288 260156 473340
rect 287612 473288 287664 473340
rect 288072 473288 288124 473340
rect 315948 473288 316000 473340
rect 316684 473288 316736 473340
rect 343916 473288 343968 473340
rect 344100 473288 344152 473340
rect 371608 473288 371660 473340
rect 372068 473288 372120 473340
rect 399944 473288 399996 473340
rect 400864 473288 400916 473340
rect 427912 473288 427964 473340
rect 428096 473288 428148 473340
rect 455604 473288 455656 473340
rect 456064 473288 456116 473340
rect 483940 473288 483992 473340
rect 484032 473288 484084 473340
rect 511908 473288 511960 473340
rect 512092 473288 512144 473340
rect 539600 473288 539652 473340
rect 540060 473288 540112 473340
rect 567936 473288 567988 473340
rect 16580 473220 16632 473272
rect 36636 473220 36688 473272
rect 44916 473220 44968 473272
rect 71136 473220 71188 473272
rect 82268 473220 82320 473272
rect 93124 473220 93176 473272
rect 110236 473220 110288 473272
rect 124864 473220 124916 473272
rect 128636 473220 128688 473272
rect 149704 473220 149756 473272
rect 156604 473220 156656 473272
rect 182824 473220 182876 473272
rect 194508 473220 194560 473272
rect 210424 473220 210476 473272
rect 212632 473220 212684 473272
rect 232504 473220 232556 473272
rect 240600 473220 240652 473272
rect 267004 473220 267056 473272
rect 278596 473220 278648 473272
rect 289084 473220 289136 473272
rect 306288 473220 306340 473272
rect 318064 473220 318116 473272
rect 324596 473220 324648 473272
rect 345664 473220 345716 473272
rect 362592 473220 362644 473272
rect 373264 473220 373316 473272
rect 390284 473220 390336 473272
rect 400956 473220 401008 473272
rect 408592 473220 408644 473272
rect 428464 473220 428516 473272
rect 436928 473220 436980 473272
rect 462964 473220 463016 473272
rect 474280 473220 474332 473272
rect 485044 473220 485096 473272
rect 502248 473220 502300 473272
rect 514024 473220 514076 473272
rect 520924 473220 520976 473272
rect 541624 473220 541676 473272
rect 26240 473152 26292 473204
rect 43536 473152 43588 473204
rect 54576 473152 54628 473204
rect 66904 473152 66956 473204
rect 138296 473152 138348 473204
rect 151084 473152 151136 473204
rect 166264 473152 166316 473204
rect 177304 473152 177356 473204
rect 222292 473152 222344 473204
rect 233976 473152 234028 473204
rect 250260 473152 250312 473204
rect 261484 473152 261536 473204
rect 334256 473152 334308 473204
rect 347044 473152 347096 473204
rect 418252 473152 418304 473204
rect 429844 473152 429896 473204
rect 446588 473152 446640 473204
rect 457444 473152 457496 473204
rect 530584 473152 530636 473204
rect 544384 473152 544436 473204
rect 558276 472608 558328 472660
rect 567476 472608 567528 472660
rect 64328 470568 64380 470620
rect 579988 470568 580040 470620
rect 548340 469820 548392 469872
rect 568028 469820 568080 469872
rect 212356 469412 212408 469464
rect 232688 469412 232740 469464
rect 296352 469412 296404 469464
rect 316776 469412 316828 469464
rect 408040 469412 408092 469464
rect 428648 469412 428700 469464
rect 148324 469344 148376 469396
rect 165712 469344 165764 469396
rect 175464 469344 175516 469396
rect 193680 469344 193732 469396
rect 203524 469344 203576 469396
rect 221372 469344 221424 469396
rect 260104 469344 260156 469396
rect 277676 469344 277728 469396
rect 287520 469344 287572 469396
rect 305368 469344 305420 469396
rect 345664 469344 345716 469396
rect 361672 469344 361724 469396
rect 371516 469344 371568 469396
rect 389364 469344 389416 469396
rect 399484 469344 399536 469396
rect 417700 469344 417752 469396
rect 456156 469344 456208 469396
rect 473360 469344 473412 469396
rect 483480 469344 483532 469396
rect 501696 469344 501748 469396
rect 511448 469344 511500 469396
rect 529664 469344 529716 469396
rect 36728 469276 36780 469328
rect 53656 469276 53708 469328
rect 64420 469276 64472 469328
rect 81440 469276 81492 469328
rect 91468 469276 91520 469328
rect 109684 469276 109736 469328
rect 119436 469276 119488 469328
rect 137652 469276 137704 469328
rect 156328 469276 156380 469328
rect 178684 469276 178736 469328
rect 232596 469276 232648 469328
rect 249708 469276 249760 469328
rect 268016 469276 268068 469328
rect 287704 469276 287756 469328
rect 315488 469276 315540 469328
rect 333704 469276 333756 469328
rect 352012 469276 352064 469328
rect 374644 469276 374696 469328
rect 428464 469276 428516 469328
rect 445668 469276 445720 469328
rect 464344 469276 464396 469328
rect 483664 469276 483716 469328
rect 492036 469276 492088 469328
rect 512736 469276 512788 469328
rect 541624 469276 541676 469328
rect 557540 469276 557592 469328
rect 15660 469208 15712 469260
rect 25688 469208 25740 469260
rect 36636 469208 36688 469260
rect 63316 469208 63368 469260
rect 66904 469208 66956 469260
rect 91100 469208 91152 469260
rect 93124 469208 93176 469260
rect 119344 469208 119396 469260
rect 124864 469208 124916 469260
rect 147312 469208 147364 469260
rect 148416 469208 148468 469260
rect 175372 469208 175424 469260
rect 177304 469208 177356 469260
rect 203340 469208 203392 469260
rect 204996 469208 205048 469260
rect 231032 469208 231084 469260
rect 232504 469208 232556 469260
rect 259368 469208 259420 469260
rect 260196 469208 260248 469260
rect 287336 469208 287388 469260
rect 289084 469208 289136 469260
rect 315028 469208 315080 469260
rect 316684 469208 316736 469260
rect 343364 469208 343416 469260
rect 344284 469208 344336 469260
rect 371332 469208 371384 469260
rect 373264 469208 373316 469260
rect 399024 469208 399076 469260
rect 400864 469208 400916 469260
rect 427360 469208 427412 469260
rect 428556 469208 428608 469260
rect 455328 469208 455380 469260
rect 456064 469208 456116 469260
rect 483020 469208 483072 469260
rect 485044 469208 485096 469260
rect 511356 469208 511408 469260
rect 512644 469208 512696 469260
rect 539324 469208 539376 469260
rect 540244 469208 540296 469260
rect 567200 469208 567252 469260
rect 15292 467236 15344 467288
rect 15936 467236 15988 467288
rect 182088 466556 182140 466608
rect 233240 466556 233292 466608
rect 350448 466556 350500 466608
rect 401600 466556 401652 466608
rect 462228 466556 462280 466608
rect 513380 466556 513432 466608
rect 42708 466488 42760 466540
rect 93860 466488 93912 466540
rect 97908 466488 97960 466540
rect 149060 466488 149112 466540
rect 154488 466488 154540 466540
rect 205640 466488 205692 466540
rect 238668 466488 238720 466540
rect 289820 466488 289872 466540
rect 293868 466488 293920 466540
rect 345020 466488 345072 466540
rect 378048 466488 378100 466540
rect 429292 466488 429344 466540
rect 434628 466488 434680 466540
rect 485780 466488 485832 466540
rect 518808 466488 518860 466540
rect 569960 466488 570012 466540
rect 13544 466420 13596 466472
rect 66260 466420 66312 466472
rect 70308 466420 70360 466472
rect 121460 466420 121512 466472
rect 126888 466420 126940 466472
rect 178040 466420 178092 466472
rect 209688 466420 209740 466472
rect 262220 466420 262272 466472
rect 266268 466420 266320 466472
rect 317420 466420 317472 466472
rect 322848 466420 322900 466472
rect 374000 466420 374052 466472
rect 405648 466420 405700 466472
rect 458180 466420 458232 466472
rect 489828 466420 489880 466472
rect 542360 466420 542412 466472
rect 42892 464040 42944 464092
rect 43628 464040 43680 464092
rect 428648 450508 428700 450560
rect 435732 450508 435784 450560
rect 512736 450440 512788 450492
rect 519636 450440 519688 450492
rect 483664 450304 483716 450356
rect 491668 450304 491720 450356
rect 232688 449896 232740 449948
rect 239772 449896 239824 449948
rect 287704 449896 287756 449948
rect 295708 449896 295760 449948
rect 316776 449896 316828 449948
rect 323676 449896 323728 449948
rect 63592 449624 63644 449676
rect 64420 449624 64472 449676
rect 455696 449624 455748 449676
rect 456156 449624 456208 449676
rect 15844 448672 15896 448724
rect 16672 448672 16724 448724
rect 2780 448604 2832 448656
rect 4896 448604 4948 448656
rect 35256 448468 35308 448520
rect 36728 448468 36780 448520
rect 231676 448468 231728 448520
rect 232596 448468 232648 448520
rect 343640 448468 343692 448520
rect 345664 448468 345716 448520
rect 539508 448468 539560 448520
rect 541624 448468 541676 448520
rect 547880 448468 547932 448520
rect 548156 448468 548208 448520
rect 71872 445680 71924 445732
rect 100024 445680 100076 445732
rect 25688 445612 25740 445664
rect 36636 445612 36688 445664
rect 42892 445612 42944 445664
rect 15292 445544 15344 445596
rect 43996 445544 44048 445596
rect 53656 445612 53708 445664
rect 66904 445612 66956 445664
rect 81992 445612 82044 445664
rect 93124 445612 93176 445664
rect 99472 445612 99524 445664
rect 127992 445680 128044 445732
rect 165988 445680 166040 445732
rect 177304 445680 177356 445732
rect 178684 445680 178736 445732
rect 184020 445680 184072 445732
rect 109684 445612 109736 445664
rect 124864 445612 124916 445664
rect 137652 445612 137704 445664
rect 148416 445612 148468 445664
rect 183652 445612 183704 445664
rect 211712 445680 211764 445732
rect 222016 445680 222068 445732
rect 232504 445680 232556 445732
rect 277676 445680 277728 445732
rect 289084 445680 289136 445732
rect 306012 445680 306064 445732
rect 316684 445680 316736 445732
rect 361672 445680 361724 445732
rect 373264 445680 373316 445732
rect 379612 445680 379664 445732
rect 408040 445680 408092 445732
rect 474004 445680 474056 445732
rect 485044 445680 485096 445732
rect 501696 445680 501748 445732
rect 512644 445680 512696 445732
rect 548156 445680 548208 445732
rect 557540 445680 557592 445732
rect 193680 445612 193732 445664
rect 204996 445612 205048 445664
rect 249708 445612 249760 445664
rect 260196 445612 260248 445664
rect 333704 445612 333756 445664
rect 344284 445612 344336 445664
rect 374644 445612 374696 445664
rect 379704 445612 379756 445664
rect 390008 445612 390060 445664
rect 400864 445612 400916 445664
rect 417700 445612 417752 445664
rect 428556 445612 428608 445664
rect 445668 445612 445720 445664
rect 456064 445612 456116 445664
rect 529664 445612 529716 445664
rect 540244 445612 540296 445664
rect 72056 445544 72108 445596
rect 127072 445544 127124 445596
rect 156052 445544 156104 445596
rect 238852 445544 238904 445596
rect 268016 445544 268068 445596
rect 323032 445544 323084 445596
rect 352012 445544 352064 445596
rect 434812 445544 434864 445596
rect 463700 445544 463752 445596
rect 518992 445544 519044 445596
rect 547880 445544 547932 445596
rect 26608 443368 26660 443420
rect 35440 443368 35492 443420
rect 71136 443096 71188 443148
rect 82268 443096 82320 443148
rect 99380 443096 99432 443148
rect 100300 443096 100352 443148
rect 183652 443096 183704 443148
rect 222200 443096 222252 443148
rect 267004 443096 267056 443148
rect 277952 443096 278004 443148
rect 295432 443096 295484 443148
rect 334256 443096 334308 443148
rect 352012 443096 352064 443148
rect 36636 443028 36688 443080
rect 53932 443028 53984 443080
rect 71872 443028 71924 443080
rect 109960 443028 110012 443080
rect 124864 443028 124916 443080
rect 128360 443028 128412 443080
rect 151084 443028 151136 443080
rect 156604 443028 156656 443080
rect 182824 443028 182876 443080
rect 193956 443028 194008 443080
rect 232504 443028 232556 443080
rect 66904 442960 66956 443012
rect 72608 442960 72660 443012
rect 93124 442960 93176 443012
rect 99380 442960 99432 443012
rect 99472 442960 99524 443012
rect 138020 442960 138072 443012
rect 149704 442960 149756 443012
rect 166264 442960 166316 443012
rect 177304 442960 177356 443012
rect 184296 442960 184348 443012
rect 233976 442960 234028 443012
rect 240600 442960 240652 443012
rect 267832 443028 267884 443080
rect 306288 443028 306340 443080
rect 345664 443028 345716 443080
rect 361948 443028 362000 443080
rect 379612 443096 379664 443148
rect 418252 443096 418304 443148
rect 462964 443096 463016 443148
rect 474280 443096 474332 443148
rect 485044 443096 485096 443148
rect 492588 443096 492640 443148
rect 390284 443028 390336 443080
rect 400864 443028 400916 443080
rect 408592 443028 408644 443080
rect 429844 443028 429896 443080
rect 436284 443028 436336 443080
rect 463792 443028 463844 443080
rect 502248 443028 502300 443080
rect 514024 443028 514076 443080
rect 520280 443028 520332 443080
rect 250260 442960 250312 443012
rect 261484 442960 261536 443012
rect 268292 442960 268344 443012
rect 289084 442960 289136 443012
rect 296628 442960 296680 443012
rect 318064 442960 318116 443012
rect 324596 442960 324648 443012
rect 347044 442960 347096 443012
rect 352288 442960 352340 443012
rect 373264 442960 373316 443012
rect 380624 442960 380676 443012
rect 428464 442960 428516 443012
rect 445944 442960 445996 443012
rect 457444 442960 457496 443012
rect 464620 442960 464672 443012
rect 491392 442960 491444 443012
rect 529940 442960 529992 443012
rect 541624 442960 541676 443012
rect 558276 442960 558328 443012
rect 210424 441600 210476 441652
rect 212540 441600 212592 441652
rect 42708 440240 42760 440292
rect 93860 440240 93912 440292
rect 97908 440240 97960 440292
rect 149060 440240 149112 440292
rect 154488 440240 154540 440292
rect 205640 440240 205692 440292
rect 209688 440240 209740 440292
rect 262220 440240 262272 440292
rect 266268 440240 266320 440292
rect 317420 440240 317472 440292
rect 322848 440240 322900 440292
rect 374000 440240 374052 440292
rect 378048 440240 378100 440292
rect 429292 440240 429344 440292
rect 434628 440240 434680 440292
rect 485780 440240 485832 440292
rect 489828 440240 489880 440292
rect 542360 440240 542412 440292
rect 544384 440240 544436 440292
rect 548340 440240 548392 440292
rect 120264 440172 120316 440224
rect 122104 440172 122156 440224
rect 204260 436092 204312 436144
rect 204996 436092 205048 436144
rect 400312 436092 400364 436144
rect 400956 436092 401008 436144
rect 13544 422220 13596 422272
rect 66260 422220 66312 422272
rect 70308 422220 70360 422272
rect 121460 422220 121512 422272
rect 126888 422220 126940 422272
rect 178040 422220 178092 422272
rect 182088 422220 182140 422272
rect 233240 422220 233292 422272
rect 238668 422220 238720 422272
rect 289820 422220 289872 422272
rect 293868 422220 293920 422272
rect 345020 422220 345072 422272
rect 350448 422220 350500 422272
rect 401600 422220 401652 422272
rect 405648 422220 405700 422272
rect 458180 422220 458232 422272
rect 462228 422220 462280 422272
rect 513380 422220 513432 422272
rect 518808 422220 518860 422272
rect 569960 422220 570012 422272
rect 15200 419432 15252 419484
rect 35900 419432 35952 419484
rect 36084 419432 36136 419484
rect 63592 419432 63644 419484
rect 64052 419432 64104 419484
rect 91928 419432 91980 419484
rect 92112 419432 92164 419484
rect 119620 419432 119672 419484
rect 122104 419432 122156 419484
rect 147956 419432 148008 419484
rect 148048 419432 148100 419484
rect 175924 419432 175976 419484
rect 176108 419432 176160 419484
rect 203616 419432 203668 419484
rect 204996 419432 205048 419484
rect 231952 419432 232004 419484
rect 232044 419432 232096 419484
rect 259920 419432 259972 419484
rect 260104 419432 260156 419484
rect 287612 419432 287664 419484
rect 288072 419432 288124 419484
rect 315948 419432 316000 419484
rect 316684 419432 316736 419484
rect 343916 419432 343968 419484
rect 344100 419432 344152 419484
rect 371608 419432 371660 419484
rect 372068 419432 372120 419484
rect 399944 419432 399996 419484
rect 400956 419432 401008 419484
rect 427912 419432 427964 419484
rect 428096 419432 428148 419484
rect 455604 419432 455656 419484
rect 456064 419432 456116 419484
rect 483940 419432 483992 419484
rect 484032 419432 484084 419484
rect 511908 419432 511960 419484
rect 512092 419432 512144 419484
rect 539600 419432 539652 419484
rect 540060 419432 540112 419484
rect 567936 419432 567988 419484
rect 16580 419364 16632 419416
rect 36636 419364 36688 419416
rect 44916 419364 44968 419416
rect 71136 419364 71188 419416
rect 82268 419364 82320 419416
rect 93124 419364 93176 419416
rect 110236 419364 110288 419416
rect 124864 419364 124916 419416
rect 128636 419364 128688 419416
rect 149704 419364 149756 419416
rect 156604 419364 156656 419416
rect 182824 419364 182876 419416
rect 194508 419364 194560 419416
rect 210424 419364 210476 419416
rect 212632 419364 212684 419416
rect 232504 419364 232556 419416
rect 240600 419364 240652 419416
rect 267004 419364 267056 419416
rect 278596 419364 278648 419416
rect 289084 419364 289136 419416
rect 306288 419364 306340 419416
rect 318064 419364 318116 419416
rect 324596 419364 324648 419416
rect 345664 419364 345716 419416
rect 362592 419364 362644 419416
rect 373264 419364 373316 419416
rect 390284 419364 390336 419416
rect 400864 419364 400916 419416
rect 408592 419364 408644 419416
rect 428464 419364 428516 419416
rect 436928 419364 436980 419416
rect 462964 419364 463016 419416
rect 474280 419364 474332 419416
rect 485044 419364 485096 419416
rect 502248 419364 502300 419416
rect 514024 419364 514076 419416
rect 520924 419364 520976 419416
rect 541624 419364 541676 419416
rect 26240 419296 26292 419348
rect 43536 419296 43588 419348
rect 54576 419296 54628 419348
rect 66904 419296 66956 419348
rect 138296 419296 138348 419348
rect 151084 419296 151136 419348
rect 166264 419296 166316 419348
rect 177304 419296 177356 419348
rect 222292 419296 222344 419348
rect 233976 419296 234028 419348
rect 250260 419296 250312 419348
rect 261484 419296 261536 419348
rect 334256 419296 334308 419348
rect 347044 419296 347096 419348
rect 418252 419296 418304 419348
rect 429844 419296 429896 419348
rect 446588 419296 446640 419348
rect 457444 419296 457496 419348
rect 530584 419296 530636 419348
rect 544384 419296 544436 419348
rect 558276 418752 558328 418804
rect 567476 418752 567528 418804
rect 548340 416032 548392 416084
rect 568028 416032 568080 416084
rect 212356 415624 212408 415676
rect 232688 415624 232740 415676
rect 296352 415624 296404 415676
rect 316776 415624 316828 415676
rect 408040 415624 408092 415676
rect 428648 415624 428700 415676
rect 119436 415556 119488 415608
rect 137652 415556 137704 415608
rect 148324 415556 148376 415608
rect 165712 415556 165764 415608
rect 175464 415556 175516 415608
rect 193680 415556 193732 415608
rect 203524 415556 203576 415608
rect 221372 415556 221424 415608
rect 260104 415556 260156 415608
rect 277676 415556 277728 415608
rect 287520 415556 287572 415608
rect 305368 415556 305420 415608
rect 345664 415556 345716 415608
rect 361672 415556 361724 415608
rect 371516 415556 371568 415608
rect 389364 415556 389416 415608
rect 399484 415556 399536 415608
rect 417700 415556 417752 415608
rect 456064 415556 456116 415608
rect 473360 415556 473412 415608
rect 483480 415556 483532 415608
rect 501696 415556 501748 415608
rect 511448 415556 511500 415608
rect 529664 415556 529716 415608
rect 36728 415488 36780 415540
rect 53656 415488 53708 415540
rect 64420 415488 64472 415540
rect 81440 415488 81492 415540
rect 91468 415488 91520 415540
rect 109684 415488 109736 415540
rect 127992 415488 128044 415540
rect 148508 415488 148560 415540
rect 156328 415488 156380 415540
rect 178684 415488 178736 415540
rect 232596 415488 232648 415540
rect 249708 415488 249760 415540
rect 268016 415488 268068 415540
rect 287704 415488 287756 415540
rect 315488 415488 315540 415540
rect 333704 415488 333756 415540
rect 352012 415488 352064 415540
rect 374644 415488 374696 415540
rect 428464 415488 428516 415540
rect 445668 415488 445720 415540
rect 464344 415488 464396 415540
rect 483664 415488 483716 415540
rect 492036 415488 492088 415540
rect 512736 415488 512788 415540
rect 541624 415488 541676 415540
rect 557540 415488 557592 415540
rect 15108 415420 15160 415472
rect 25688 415420 25740 415472
rect 36636 415420 36688 415472
rect 63316 415420 63368 415472
rect 66904 415420 66956 415472
rect 91100 415420 91152 415472
rect 93124 415420 93176 415472
rect 119344 415420 119396 415472
rect 122104 415420 122156 415472
rect 147312 415420 147364 415472
rect 148416 415420 148468 415472
rect 175372 415420 175424 415472
rect 177304 415420 177356 415472
rect 203340 415420 203392 415472
rect 204996 415420 205048 415472
rect 231032 415420 231084 415472
rect 232504 415420 232556 415472
rect 259368 415420 259420 415472
rect 260196 415420 260248 415472
rect 287336 415420 287388 415472
rect 289084 415420 289136 415472
rect 315028 415420 315080 415472
rect 316684 415420 316736 415472
rect 343364 415420 343416 415472
rect 344284 415420 344336 415472
rect 371332 415420 371384 415472
rect 373264 415420 373316 415472
rect 399024 415420 399076 415472
rect 400864 415420 400916 415472
rect 427360 415420 427412 415472
rect 428556 415420 428608 415472
rect 455328 415420 455380 415472
rect 456156 415420 456208 415472
rect 483020 415420 483072 415472
rect 485044 415420 485096 415472
rect 511356 415420 511408 415472
rect 512644 415420 512696 415472
rect 539324 415420 539376 415472
rect 540244 415420 540296 415472
rect 567200 415420 567252 415472
rect 3148 410320 3200 410372
rect 8944 410320 8996 410372
rect 42892 405900 42944 405952
rect 43628 405900 43680 405952
rect 148508 395292 148560 395344
rect 155868 395292 155920 395344
rect 428648 395292 428700 395344
rect 435732 395292 435784 395344
rect 287704 395088 287756 395140
rect 295800 395088 295852 395140
rect 316776 395088 316828 395140
rect 323676 395088 323728 395140
rect 232688 395020 232740 395072
rect 239772 395020 239824 395072
rect 483664 395020 483716 395072
rect 491668 395020 491720 395072
rect 512736 395020 512788 395072
rect 519636 395020 519688 395072
rect 547880 394680 547932 394732
rect 548156 394680 548208 394732
rect 13544 394612 13596 394664
rect 35256 394544 35308 394596
rect 36728 394544 36780 394596
rect 42708 394544 42760 394596
rect 63592 394612 63644 394664
rect 64420 394612 64472 394664
rect 70308 394612 70360 394664
rect 121460 394612 121512 394664
rect 126888 394612 126940 394664
rect 178040 394612 178092 394664
rect 209688 394612 209740 394664
rect 262220 394612 262272 394664
rect 266268 394612 266320 394664
rect 317420 394612 317472 394664
rect 322848 394612 322900 394664
rect 374000 394612 374052 394664
rect 405648 394612 405700 394664
rect 458180 394612 458232 394664
rect 489828 394612 489880 394664
rect 542360 394612 542412 394664
rect 66260 394476 66312 394528
rect 93860 394544 93912 394596
rect 97908 394544 97960 394596
rect 149060 394544 149112 394596
rect 182088 394544 182140 394596
rect 233240 394544 233292 394596
rect 238668 394544 238720 394596
rect 289820 394544 289872 394596
rect 293868 394544 293920 394596
rect 154488 394476 154540 394528
rect 205640 394476 205692 394528
rect 343640 394544 343692 394596
rect 345664 394544 345716 394596
rect 378048 394544 378100 394596
rect 429292 394544 429344 394596
rect 462228 394544 462280 394596
rect 513380 394544 513432 394596
rect 518808 394544 518860 394596
rect 569960 394544 570012 394596
rect 345020 394476 345072 394528
rect 350448 394476 350500 394528
rect 401600 394476 401652 394528
rect 434628 394476 434680 394528
rect 485780 394476 485832 394528
rect 231584 393252 231636 393304
rect 232596 393252 232648 393304
rect 539324 393252 539376 393304
rect 541624 393252 541676 393304
rect 71872 391892 71924 391944
rect 100024 391892 100076 391944
rect 25688 391824 25740 391876
rect 36636 391824 36688 391876
rect 42892 391824 42944 391876
rect 15292 391756 15344 391808
rect 43996 391756 44048 391808
rect 53656 391824 53708 391876
rect 66904 391824 66956 391876
rect 81992 391824 82044 391876
rect 93124 391824 93176 391876
rect 99472 391824 99524 391876
rect 127992 391892 128044 391944
rect 165988 391892 166040 391944
rect 177304 391892 177356 391944
rect 178684 391892 178736 391944
rect 184020 391892 184072 391944
rect 109684 391824 109736 391876
rect 122104 391824 122156 391876
rect 137652 391824 137704 391876
rect 148416 391824 148468 391876
rect 183652 391824 183704 391876
rect 211712 391892 211764 391944
rect 221924 391892 221976 391944
rect 232504 391892 232556 391944
rect 277676 391892 277728 391944
rect 289084 391892 289136 391944
rect 306012 391892 306064 391944
rect 316684 391892 316736 391944
rect 361672 391892 361724 391944
rect 373264 391892 373316 391944
rect 379612 391892 379664 391944
rect 408040 391892 408092 391944
rect 474004 391892 474056 391944
rect 485044 391892 485096 391944
rect 501696 391892 501748 391944
rect 512644 391892 512696 391944
rect 548156 391892 548208 391944
rect 557540 391892 557592 391944
rect 193680 391824 193732 391876
rect 204996 391824 205048 391876
rect 249708 391824 249760 391876
rect 260196 391824 260248 391876
rect 333704 391824 333756 391876
rect 344284 391824 344336 391876
rect 374644 391824 374696 391876
rect 379704 391824 379756 391876
rect 390008 391824 390060 391876
rect 400864 391824 400916 391876
rect 417700 391824 417752 391876
rect 428556 391824 428608 391876
rect 445668 391824 445720 391876
rect 456156 391824 456208 391876
rect 529664 391824 529716 391876
rect 540244 391824 540296 391876
rect 71964 391756 72016 391808
rect 238852 391756 238904 391808
rect 268016 391756 268068 391808
rect 323032 391756 323084 391808
rect 352012 391756 352064 391808
rect 434812 391756 434864 391808
rect 463792 391756 463844 391808
rect 518992 391756 519044 391808
rect 547880 391756 547932 391808
rect 15108 390396 15160 390448
rect 16580 390396 16632 390448
rect 26240 389784 26292 389836
rect 35440 389784 35492 389836
rect 71136 389308 71188 389360
rect 82268 389308 82320 389360
rect 99472 389308 99524 389360
rect 100392 389308 100444 389360
rect 183652 389308 183704 389360
rect 222292 389308 222344 389360
rect 267004 389308 267056 389360
rect 277952 389308 278004 389360
rect 295432 389308 295484 389360
rect 334256 389308 334308 389360
rect 352012 389308 352064 389360
rect 36636 389240 36688 389292
rect 53932 389240 53984 389292
rect 71872 389240 71924 389292
rect 109960 389240 110012 389292
rect 151084 389240 151136 389292
rect 156604 389240 156656 389292
rect 182824 389240 182876 389292
rect 193956 389240 194008 389292
rect 232504 389240 232556 389292
rect 66904 389172 66956 389224
rect 72608 389172 72660 389224
rect 93124 389172 93176 389224
rect 100300 389172 100352 389224
rect 100392 389172 100444 389224
rect 138296 389172 138348 389224
rect 149704 389172 149756 389224
rect 166264 389172 166316 389224
rect 177304 389172 177356 389224
rect 184296 389172 184348 389224
rect 233976 389172 234028 389224
rect 240600 389172 240652 389224
rect 267832 389240 267884 389292
rect 306288 389240 306340 389292
rect 345664 389240 345716 389292
rect 361948 389240 362000 389292
rect 379612 389308 379664 389360
rect 418252 389308 418304 389360
rect 463792 389308 463844 389360
rect 390284 389240 390336 389292
rect 400956 389240 401008 389292
rect 408592 389240 408644 389292
rect 429844 389240 429896 389292
rect 436284 389240 436336 389292
rect 457444 389240 457496 389292
rect 464620 389240 464672 389292
rect 491392 389308 491444 389360
rect 250260 389172 250312 389224
rect 261484 389172 261536 389224
rect 268292 389172 268344 389224
rect 289084 389172 289136 389224
rect 296628 389172 296680 389224
rect 318064 389172 318116 389224
rect 324596 389172 324648 389224
rect 347044 389172 347096 389224
rect 352288 389172 352340 389224
rect 373264 389172 373316 389224
rect 380624 389172 380676 389224
rect 428464 389172 428516 389224
rect 445944 389172 445996 389224
rect 462964 389172 463016 389224
rect 474280 389172 474332 389224
rect 485044 389172 485096 389224
rect 492588 389172 492640 389224
rect 502248 389240 502300 389292
rect 514024 389240 514076 389292
rect 520280 389240 520332 389292
rect 529940 389172 529992 389224
rect 541624 389172 541676 389224
rect 558276 389172 558328 389224
rect 42708 386452 42760 386504
rect 93860 386452 93912 386504
rect 97908 386452 97960 386504
rect 126888 386520 126940 386572
rect 13544 386384 13596 386436
rect 66260 386384 66312 386436
rect 70308 386384 70360 386436
rect 121460 386384 121512 386436
rect 124864 386384 124916 386436
rect 128268 386384 128320 386436
rect 182088 386520 182140 386572
rect 233240 386520 233292 386572
rect 350448 386520 350500 386572
rect 401600 386520 401652 386572
rect 462228 386520 462280 386572
rect 513380 386520 513432 386572
rect 149060 386452 149112 386504
rect 154488 386452 154540 386504
rect 205640 386452 205692 386504
rect 238668 386452 238720 386504
rect 289820 386452 289872 386504
rect 293868 386452 293920 386504
rect 345020 386452 345072 386504
rect 378048 386452 378100 386504
rect 429292 386452 429344 386504
rect 434628 386452 434680 386504
rect 485780 386452 485832 386504
rect 518808 386452 518860 386504
rect 569960 386452 570012 386504
rect 178040 386384 178092 386436
rect 209688 386384 209740 386436
rect 262220 386384 262272 386436
rect 266268 386384 266320 386436
rect 317420 386384 317472 386436
rect 322848 386384 322900 386436
rect 374000 386384 374052 386436
rect 405648 386384 405700 386436
rect 458180 386384 458232 386436
rect 489828 386384 489880 386436
rect 542360 386384 542412 386436
rect 544384 386384 544436 386436
rect 548340 386384 548392 386436
rect 120264 386248 120316 386300
rect 122104 386248 122156 386300
rect 204076 385024 204128 385076
rect 212448 385024 212500 385076
rect 204260 384956 204312 385008
rect 204996 384956 205048 385008
rect 568120 378156 568172 378208
rect 580172 378156 580224 378208
rect 15200 365644 15252 365696
rect 35900 365644 35952 365696
rect 36084 365644 36136 365696
rect 63592 365644 63644 365696
rect 64052 365644 64104 365696
rect 91928 365644 91980 365696
rect 92112 365644 92164 365696
rect 119620 365644 119672 365696
rect 122104 365644 122156 365696
rect 147956 365644 148008 365696
rect 148048 365644 148100 365696
rect 175924 365644 175976 365696
rect 176108 365644 176160 365696
rect 203616 365644 203668 365696
rect 204996 365644 205048 365696
rect 231952 365644 232004 365696
rect 232044 365644 232096 365696
rect 259920 365644 259972 365696
rect 260104 365644 260156 365696
rect 287612 365644 287664 365696
rect 288072 365644 288124 365696
rect 315948 365644 316000 365696
rect 316684 365644 316736 365696
rect 343916 365644 343968 365696
rect 344100 365644 344152 365696
rect 371608 365644 371660 365696
rect 372068 365644 372120 365696
rect 399944 365644 399996 365696
rect 400864 365644 400916 365696
rect 427912 365644 427964 365696
rect 428096 365644 428148 365696
rect 455604 365644 455656 365696
rect 456064 365644 456116 365696
rect 483940 365644 483992 365696
rect 484032 365644 484084 365696
rect 511908 365644 511960 365696
rect 512092 365644 512144 365696
rect 539600 365644 539652 365696
rect 540060 365644 540112 365696
rect 567936 365644 567988 365696
rect 16580 365576 16632 365628
rect 36636 365576 36688 365628
rect 44916 365576 44968 365628
rect 71136 365576 71188 365628
rect 82268 365576 82320 365628
rect 93124 365576 93176 365628
rect 110236 365576 110288 365628
rect 124864 365576 124916 365628
rect 128636 365576 128688 365628
rect 149704 365576 149756 365628
rect 156604 365576 156656 365628
rect 182824 365576 182876 365628
rect 194508 365576 194560 365628
rect 204076 365576 204128 365628
rect 212632 365576 212684 365628
rect 232504 365576 232556 365628
rect 240600 365576 240652 365628
rect 267004 365576 267056 365628
rect 278596 365576 278648 365628
rect 289084 365576 289136 365628
rect 306288 365576 306340 365628
rect 318064 365576 318116 365628
rect 324596 365576 324648 365628
rect 345664 365576 345716 365628
rect 362592 365576 362644 365628
rect 373264 365576 373316 365628
rect 390284 365576 390336 365628
rect 400956 365576 401008 365628
rect 408592 365576 408644 365628
rect 428464 365576 428516 365628
rect 436928 365576 436980 365628
rect 462964 365576 463016 365628
rect 474280 365576 474332 365628
rect 485044 365576 485096 365628
rect 502248 365576 502300 365628
rect 514024 365576 514076 365628
rect 520924 365576 520976 365628
rect 541624 365576 541676 365628
rect 26240 365508 26292 365560
rect 43536 365508 43588 365560
rect 54576 365508 54628 365560
rect 66904 365508 66956 365560
rect 138296 365508 138348 365560
rect 151084 365508 151136 365560
rect 166264 365508 166316 365560
rect 177304 365508 177356 365560
rect 222292 365508 222344 365560
rect 233976 365508 234028 365560
rect 250260 365508 250312 365560
rect 261484 365508 261536 365560
rect 334256 365508 334308 365560
rect 347044 365508 347096 365560
rect 418252 365508 418304 365560
rect 429844 365508 429896 365560
rect 446588 365508 446640 365560
rect 457444 365508 457496 365560
rect 530584 365508 530636 365560
rect 544384 365508 544436 365560
rect 558276 364964 558328 365016
rect 567476 364964 567528 365016
rect 548340 362176 548392 362228
rect 568120 362176 568172 362228
rect 148416 361700 148468 361752
rect 165712 361700 165764 361752
rect 175464 361700 175516 361752
rect 193680 361700 193732 361752
rect 203524 361700 203576 361752
rect 221372 361700 221424 361752
rect 232596 361700 232648 361752
rect 249708 361700 249760 361752
rect 260104 361700 260156 361752
rect 277676 361700 277728 361752
rect 296352 361700 296404 361752
rect 316776 361700 316828 361752
rect 345664 361700 345716 361752
rect 361672 361700 361724 361752
rect 371516 361700 371568 361752
rect 389364 361700 389416 361752
rect 399484 361700 399536 361752
rect 417700 361700 417752 361752
rect 428464 361700 428516 361752
rect 445668 361700 445720 361752
rect 456064 361700 456116 361752
rect 473360 361700 473412 361752
rect 483480 361700 483532 361752
rect 501696 361700 501748 361752
rect 511448 361700 511500 361752
rect 529664 361700 529716 361752
rect 36636 361632 36688 361684
rect 53656 361632 53708 361684
rect 64420 361632 64472 361684
rect 81440 361632 81492 361684
rect 119436 361632 119488 361684
rect 137652 361632 137704 361684
rect 156328 361632 156380 361684
rect 178684 361632 178736 361684
rect 212356 361632 212408 361684
rect 232688 361632 232740 361684
rect 268016 361632 268068 361684
rect 287704 361632 287756 361684
rect 315488 361632 315540 361684
rect 333704 361632 333756 361684
rect 352012 361632 352064 361684
rect 374644 361632 374696 361684
rect 408040 361632 408092 361684
rect 428648 361632 428700 361684
rect 464344 361632 464396 361684
rect 483664 361632 483716 361684
rect 492036 361632 492088 361684
rect 512736 361632 512788 361684
rect 541624 361632 541676 361684
rect 557540 361632 557592 361684
rect 15108 361564 15160 361616
rect 25688 361564 25740 361616
rect 36728 361564 36780 361616
rect 63316 361564 63368 361616
rect 66904 361564 66956 361616
rect 91100 361564 91152 361616
rect 93124 361564 93176 361616
rect 119344 361564 119396 361616
rect 122104 361564 122156 361616
rect 147312 361564 147364 361616
rect 148324 361564 148376 361616
rect 175372 361564 175424 361616
rect 177304 361564 177356 361616
rect 203340 361564 203392 361616
rect 204996 361564 205048 361616
rect 231032 361564 231084 361616
rect 232504 361564 232556 361616
rect 259368 361564 259420 361616
rect 260196 361564 260248 361616
rect 287336 361564 287388 361616
rect 289084 361564 289136 361616
rect 315028 361564 315080 361616
rect 316684 361564 316736 361616
rect 343364 361564 343416 361616
rect 344284 361564 344336 361616
rect 371332 361564 371384 361616
rect 373264 361564 373316 361616
rect 399024 361564 399076 361616
rect 400864 361564 400916 361616
rect 427360 361564 427412 361616
rect 428556 361564 428608 361616
rect 455328 361564 455380 361616
rect 456156 361564 456208 361616
rect 483020 361564 483072 361616
rect 485044 361564 485096 361616
rect 511356 361564 511408 361616
rect 512644 361564 512696 361616
rect 539324 361564 539376 361616
rect 540244 361564 540296 361616
rect 567200 361564 567252 361616
rect 109316 359252 109368 359304
rect 91468 358776 91520 358828
rect 287520 358776 287572 358828
rect 305368 359252 305420 359304
rect 42892 356940 42944 356992
rect 43628 356940 43680 356992
rect 2780 345176 2832 345228
rect 4988 345176 5040 345228
rect 63592 342524 63644 342576
rect 64420 342524 64472 342576
rect 147680 342524 147732 342576
rect 148416 342524 148468 342576
rect 512736 341912 512788 341964
rect 519636 341912 519688 341964
rect 287704 341504 287756 341556
rect 295708 341504 295760 341556
rect 428648 341504 428700 341556
rect 435732 341504 435784 341556
rect 232688 341368 232740 341420
rect 239772 341368 239824 341420
rect 483664 341368 483716 341420
rect 491668 341368 491720 341420
rect 316776 341232 316828 341284
rect 323676 341232 323728 341284
rect 13544 340824 13596 340876
rect 66260 340824 66312 340876
rect 70308 340824 70360 340876
rect 121460 340824 121512 340876
rect 126888 340824 126940 340876
rect 178040 340824 178092 340876
rect 209688 340824 209740 340876
rect 262220 340824 262272 340876
rect 266268 340824 266320 340876
rect 317420 340824 317472 340876
rect 322848 340824 322900 340876
rect 374000 340824 374052 340876
rect 405648 340824 405700 340876
rect 458180 340824 458232 340876
rect 489828 340824 489880 340876
rect 42708 340756 42760 340808
rect 93860 340756 93912 340808
rect 97908 340756 97960 340808
rect 149060 340756 149112 340808
rect 154488 340756 154540 340808
rect 205640 340756 205692 340808
rect 231676 340756 231728 340808
rect 232596 340756 232648 340808
rect 238668 340756 238720 340808
rect 289820 340756 289872 340808
rect 293868 340756 293920 340808
rect 345020 340756 345072 340808
rect 378048 340756 378100 340808
rect 429292 340756 429344 340808
rect 434628 340756 434680 340808
rect 485780 340756 485832 340808
rect 518808 340756 518860 340808
rect 35256 340688 35308 340740
rect 36636 340688 36688 340740
rect 182088 340688 182140 340740
rect 233240 340688 233292 340740
rect 343640 340688 343692 340740
rect 345664 340688 345716 340740
rect 350448 340688 350500 340740
rect 401600 340688 401652 340740
rect 462228 340688 462280 340740
rect 513380 340688 513432 340740
rect 539508 340824 539560 340876
rect 541624 340824 541676 340876
rect 542360 340688 542412 340740
rect 569960 340756 570012 340808
rect 547880 340552 547932 340604
rect 548156 340552 548208 340604
rect 71872 338036 71924 338088
rect 100024 338036 100076 338088
rect 25688 337968 25740 338020
rect 36728 337968 36780 338020
rect 42892 337968 42944 338020
rect 15292 337900 15344 337952
rect 43996 337900 44048 337952
rect 53656 337968 53708 338020
rect 66904 337968 66956 338020
rect 81992 337968 82044 338020
rect 93124 337968 93176 338020
rect 99472 337968 99524 338020
rect 127992 338036 128044 338088
rect 165988 338036 166040 338088
rect 177304 338036 177356 338088
rect 178684 338036 178736 338088
rect 184020 338036 184072 338088
rect 109684 337968 109736 338020
rect 122104 337968 122156 338020
rect 137652 337968 137704 338020
rect 148324 337968 148376 338020
rect 183652 337968 183704 338020
rect 211712 338036 211764 338088
rect 277676 338036 277728 338088
rect 289084 338036 289136 338088
rect 306012 338036 306064 338088
rect 316684 338036 316736 338088
rect 361672 338036 361724 338088
rect 373264 338036 373316 338088
rect 374644 338036 374696 338088
rect 379704 338036 379756 338088
rect 193680 337968 193732 338020
rect 204996 337968 205048 338020
rect 222016 337968 222068 338020
rect 232504 337968 232556 338020
rect 249708 337968 249760 338020
rect 260196 337968 260248 338020
rect 333704 337968 333756 338020
rect 344284 337968 344336 338020
rect 379612 337968 379664 338020
rect 408040 338036 408092 338088
rect 474004 338036 474056 338088
rect 485044 338036 485096 338088
rect 501696 338036 501748 338088
rect 512644 338036 512696 338088
rect 548156 338036 548208 338088
rect 557540 338036 557592 338088
rect 390008 337968 390060 338020
rect 400864 337968 400916 338020
rect 417700 337968 417752 338020
rect 428556 337968 428608 338020
rect 445668 337968 445720 338020
rect 456156 337968 456208 338020
rect 529664 337968 529716 338020
rect 540244 337968 540296 338020
rect 72056 337900 72108 337952
rect 127072 337900 127124 337952
rect 156052 337900 156104 337952
rect 238852 337900 238904 337952
rect 268016 337900 268068 337952
rect 323032 337900 323084 337952
rect 352012 337900 352064 337952
rect 434812 337900 434864 337952
rect 463700 337900 463752 337952
rect 518992 337900 519044 337952
rect 547880 337900 547932 337952
rect 26240 335724 26292 335776
rect 35440 335724 35492 335776
rect 71136 335452 71188 335504
rect 82268 335452 82320 335504
rect 99380 335452 99432 335504
rect 100300 335452 100352 335504
rect 183652 335452 183704 335504
rect 222292 335452 222344 335504
rect 261484 335452 261536 335504
rect 268292 335452 268344 335504
rect 295432 335452 295484 335504
rect 334256 335452 334308 335504
rect 379612 335452 379664 335504
rect 418252 335452 418304 335504
rect 463792 335452 463844 335504
rect 36636 335384 36688 335436
rect 53932 335384 53984 335436
rect 71872 335384 71924 335436
rect 109960 335384 110012 335436
rect 124864 335384 124916 335436
rect 128636 335384 128688 335436
rect 151084 335384 151136 335436
rect 156604 335384 156656 335436
rect 182824 335384 182876 335436
rect 193956 335384 194008 335436
rect 232504 335384 232556 335436
rect 15108 335316 15160 335368
rect 16580 335316 16632 335368
rect 66904 335316 66956 335368
rect 72608 335316 72660 335368
rect 93124 335316 93176 335368
rect 99380 335316 99432 335368
rect 99472 335316 99524 335368
rect 138296 335316 138348 335368
rect 149704 335316 149756 335368
rect 166264 335316 166316 335368
rect 177304 335316 177356 335368
rect 184296 335316 184348 335368
rect 233976 335316 234028 335368
rect 240600 335316 240652 335368
rect 267832 335384 267884 335436
rect 306288 335384 306340 335436
rect 352012 335384 352064 335436
rect 390284 335384 390336 335436
rect 400864 335384 400916 335436
rect 408592 335384 408644 335436
rect 429844 335384 429896 335436
rect 436284 335384 436336 335436
rect 457444 335384 457496 335436
rect 464620 335384 464672 335436
rect 491392 335452 491444 335504
rect 529940 335452 529992 335504
rect 502248 335384 502300 335436
rect 512644 335384 512696 335436
rect 520280 335384 520332 335436
rect 250260 335316 250312 335368
rect 267004 335316 267056 335368
rect 277952 335316 278004 335368
rect 289084 335316 289136 335368
rect 296536 335316 296588 335368
rect 318064 335316 318116 335368
rect 324596 335316 324648 335368
rect 347044 335316 347096 335368
rect 361948 335316 362000 335368
rect 373264 335316 373316 335368
rect 380624 335316 380676 335368
rect 428464 335316 428516 335368
rect 445944 335316 445996 335368
rect 462964 335316 463016 335368
rect 474280 335316 474332 335368
rect 485044 335316 485096 335368
rect 492588 335316 492640 335368
rect 511816 335316 511868 335368
rect 514024 335316 514076 335368
rect 541624 335316 541676 335368
rect 558276 335316 558328 335368
rect 348424 332528 348476 332580
rect 352288 332528 352340 332580
rect 544384 332528 544436 332580
rect 548340 332528 548392 332580
rect 568028 332392 568080 332444
rect 120172 332256 120224 332308
rect 122104 332256 122156 332308
rect 568028 332188 568080 332240
rect 209688 331304 209740 331356
rect 262220 331304 262272 331356
rect 204076 331236 204128 331288
rect 212448 331236 212500 331288
rect 293868 331236 293920 331288
rect 345020 331236 345072 331288
rect 405648 331236 405700 331288
rect 458180 331236 458232 331288
rect 489828 331236 489880 331288
rect 542360 331236 542412 331288
rect 204260 328992 204312 329044
rect 204996 328992 205048 329044
rect 400312 328992 400364 329044
rect 400956 328992 401008 329044
rect 570604 324300 570656 324352
rect 579988 324300 580040 324352
rect 13544 314576 13596 314628
rect 66260 314576 66312 314628
rect 70308 314576 70360 314628
rect 121460 314576 121512 314628
rect 126888 314576 126940 314628
rect 178040 314576 178092 314628
rect 182088 314576 182140 314628
rect 233240 314576 233292 314628
rect 238668 314576 238720 314628
rect 289820 314576 289872 314628
rect 322848 314576 322900 314628
rect 374000 314576 374052 314628
rect 378048 314576 378100 314628
rect 429292 314576 429344 314628
rect 434628 314576 434680 314628
rect 485780 314576 485832 314628
rect 518808 314576 518860 314628
rect 569960 314576 570012 314628
rect 42708 314508 42760 314560
rect 93860 314508 93912 314560
rect 97908 314508 97960 314560
rect 149060 314508 149112 314560
rect 154488 314508 154540 314560
rect 205640 314508 205692 314560
rect 266268 314508 266320 314560
rect 317420 314508 317472 314560
rect 350448 314508 350500 314560
rect 401600 314508 401652 314560
rect 462228 314508 462280 314560
rect 513380 314508 513432 314560
rect 15200 311788 15252 311840
rect 35900 311788 35952 311840
rect 36084 311788 36136 311840
rect 63592 311788 63644 311840
rect 64052 311788 64104 311840
rect 91928 311788 91980 311840
rect 92112 311788 92164 311840
rect 119620 311788 119672 311840
rect 122104 311788 122156 311840
rect 147956 311788 148008 311840
rect 148048 311788 148100 311840
rect 175924 311788 175976 311840
rect 176108 311788 176160 311840
rect 203616 311788 203668 311840
rect 204996 311788 205048 311840
rect 231952 311788 232004 311840
rect 232044 311788 232096 311840
rect 259920 311788 259972 311840
rect 260104 311788 260156 311840
rect 287612 311788 287664 311840
rect 288072 311788 288124 311840
rect 315948 311788 316000 311840
rect 316684 311788 316736 311840
rect 343916 311788 343968 311840
rect 344100 311788 344152 311840
rect 371608 311788 371660 311840
rect 372068 311788 372120 311840
rect 399944 311788 399996 311840
rect 400956 311788 401008 311840
rect 427912 311788 427964 311840
rect 428096 311788 428148 311840
rect 455604 311788 455656 311840
rect 456064 311788 456116 311840
rect 483940 311788 483992 311840
rect 484032 311788 484084 311840
rect 511908 311788 511960 311840
rect 514024 311788 514076 311840
rect 539600 311788 539652 311840
rect 540060 311788 540112 311840
rect 567936 311788 567988 311840
rect 16580 311720 16632 311772
rect 36636 311720 36688 311772
rect 44916 311720 44968 311772
rect 71136 311720 71188 311772
rect 82268 311720 82320 311772
rect 93124 311720 93176 311772
rect 110236 311720 110288 311772
rect 124864 311720 124916 311772
rect 128636 311720 128688 311772
rect 149704 311720 149756 311772
rect 156604 311720 156656 311772
rect 182824 311720 182876 311772
rect 194508 311720 194560 311772
rect 204076 311720 204128 311772
rect 212632 311720 212684 311772
rect 232504 311720 232556 311772
rect 240600 311720 240652 311772
rect 267004 311720 267056 311772
rect 278596 311720 278648 311772
rect 289084 311720 289136 311772
rect 306288 311720 306340 311772
rect 318064 311720 318116 311772
rect 324596 311720 324648 311772
rect 347044 311720 347096 311772
rect 362592 311720 362644 311772
rect 373264 311720 373316 311772
rect 390284 311720 390336 311772
rect 400864 311720 400916 311772
rect 408592 311720 408644 311772
rect 428464 311720 428516 311772
rect 436928 311720 436980 311772
rect 462964 311720 463016 311772
rect 474280 311720 474332 311772
rect 485044 311720 485096 311772
rect 502248 311720 502300 311772
rect 512644 311720 512696 311772
rect 520924 311720 520976 311772
rect 541624 311720 541676 311772
rect 26240 311652 26292 311704
rect 43536 311652 43588 311704
rect 54576 311652 54628 311704
rect 66904 311652 66956 311704
rect 138296 311652 138348 311704
rect 151084 311652 151136 311704
rect 166264 311652 166316 311704
rect 177304 311652 177356 311704
rect 222292 311652 222344 311704
rect 233976 311652 234028 311704
rect 250260 311652 250312 311704
rect 261484 311652 261536 311704
rect 334256 311652 334308 311704
rect 348424 311652 348476 311704
rect 418252 311652 418304 311704
rect 429844 311652 429896 311704
rect 446588 311652 446640 311704
rect 457444 311652 457496 311704
rect 530584 311652 530636 311704
rect 544384 311652 544436 311704
rect 558276 311108 558328 311160
rect 567476 311108 567528 311160
rect 548340 308388 548392 308440
rect 568120 308388 568172 308440
rect 212264 307980 212316 308032
rect 232688 307980 232740 308032
rect 296352 307980 296404 308032
rect 316776 307980 316828 308032
rect 408040 307980 408092 308032
rect 428648 307980 428700 308032
rect 148324 307912 148376 307964
rect 165620 307912 165672 307964
rect 175464 307912 175516 307964
rect 193680 307912 193732 307964
rect 203524 307912 203576 307964
rect 221372 307912 221424 307964
rect 260196 307912 260248 307964
rect 277676 307912 277728 307964
rect 287520 307912 287572 307964
rect 305368 307912 305420 307964
rect 345664 307912 345716 307964
rect 361672 307912 361724 307964
rect 371516 307912 371568 307964
rect 389364 307912 389416 307964
rect 399484 307912 399536 307964
rect 417700 307912 417752 307964
rect 456156 307912 456208 307964
rect 473544 307912 473596 307964
rect 483480 307912 483532 307964
rect 501696 307912 501748 307964
rect 511448 307912 511500 307964
rect 529664 307912 529716 307964
rect 36728 307844 36780 307896
rect 53656 307844 53708 307896
rect 64420 307844 64472 307896
rect 81440 307844 81492 307896
rect 91468 307844 91520 307896
rect 109684 307844 109736 307896
rect 119436 307844 119488 307896
rect 137652 307844 137704 307896
rect 156328 307844 156380 307896
rect 178684 307844 178736 307896
rect 232504 307844 232556 307896
rect 249708 307844 249760 307896
rect 268016 307844 268068 307896
rect 287704 307844 287756 307896
rect 315488 307844 315540 307896
rect 333704 307844 333756 307896
rect 352012 307844 352064 307896
rect 374644 307844 374696 307896
rect 428556 307844 428608 307896
rect 445668 307844 445720 307896
rect 464344 307844 464396 307896
rect 483664 307844 483716 307896
rect 492036 307844 492088 307896
rect 512736 307844 512788 307896
rect 541624 307844 541676 307896
rect 557540 307844 557592 307896
rect 15108 307776 15160 307828
rect 25688 307776 25740 307828
rect 36636 307776 36688 307828
rect 63316 307776 63368 307828
rect 66904 307776 66956 307828
rect 91100 307776 91152 307828
rect 93124 307776 93176 307828
rect 119344 307776 119396 307828
rect 122104 307776 122156 307828
rect 147312 307776 147364 307828
rect 148416 307776 148468 307828
rect 175280 307776 175332 307828
rect 177304 307776 177356 307828
rect 203340 307776 203392 307828
rect 204996 307776 205048 307828
rect 231032 307776 231084 307828
rect 232596 307776 232648 307828
rect 259368 307776 259420 307828
rect 260104 307776 260156 307828
rect 287336 307776 287388 307828
rect 289084 307776 289136 307828
rect 315028 307776 315080 307828
rect 316684 307776 316736 307828
rect 343364 307776 343416 307828
rect 344284 307776 344336 307828
rect 371332 307776 371384 307828
rect 373264 307776 373316 307828
rect 399024 307776 399076 307828
rect 400864 307776 400916 307828
rect 427360 307776 427412 307828
rect 428464 307776 428516 307828
rect 455328 307776 455380 307828
rect 456064 307776 456116 307828
rect 483204 307776 483256 307828
rect 485044 307776 485096 307828
rect 511356 307776 511408 307828
rect 512644 307776 512696 307828
rect 539324 307776 539376 307828
rect 540244 307776 540296 307828
rect 567200 307776 567252 307828
rect 42892 300976 42944 301028
rect 43628 300976 43680 301028
rect 3332 293088 3384 293140
rect 7564 293088 7616 293140
rect 63592 291864 63644 291916
rect 64420 291864 64472 291916
rect 259736 291864 259788 291916
rect 260196 291864 260248 291916
rect 455696 291864 455748 291916
rect 456156 291864 456208 291916
rect 287704 288328 287756 288380
rect 295708 288328 295760 288380
rect 316776 288328 316828 288380
rect 323676 288328 323728 288380
rect 232688 287920 232740 287972
rect 239772 287920 239824 287972
rect 428648 287648 428700 287700
rect 435732 287648 435784 287700
rect 512736 287512 512788 287564
rect 519636 287512 519688 287564
rect 483664 287376 483716 287428
rect 491668 287376 491720 287428
rect 13544 286968 13596 287020
rect 66260 286968 66312 287020
rect 70308 286968 70360 287020
rect 121460 286968 121512 287020
rect 154488 286968 154540 287020
rect 205640 286968 205692 287020
rect 209688 286968 209740 287020
rect 262220 286968 262272 287020
rect 266268 286968 266320 287020
rect 317420 286968 317472 287020
rect 322848 286968 322900 287020
rect 374000 286968 374052 287020
rect 405648 286968 405700 287020
rect 458180 286968 458232 287020
rect 489828 286968 489880 287020
rect 542360 286968 542412 287020
rect 42708 286900 42760 286952
rect 93860 286900 93912 286952
rect 97908 286900 97960 286952
rect 149060 286900 149112 286952
rect 182088 286900 182140 286952
rect 233240 286900 233292 286952
rect 238668 286900 238720 286952
rect 289820 286900 289872 286952
rect 293868 286900 293920 286952
rect 126888 286832 126940 286884
rect 178040 286832 178092 286884
rect 343548 286900 343600 286952
rect 345664 286900 345716 286952
rect 378048 286900 378100 286952
rect 429292 286900 429344 286952
rect 434628 286900 434680 286952
rect 485780 286900 485832 286952
rect 518808 286900 518860 286952
rect 569960 286900 570012 286952
rect 345020 286832 345072 286884
rect 350448 286832 350500 286884
rect 401600 286832 401652 286884
rect 462228 286832 462280 286884
rect 513380 286832 513432 286884
rect 427728 286764 427780 286816
rect 428556 286764 428608 286816
rect 539508 286764 539560 286816
rect 541624 286764 541676 286816
rect 35256 286696 35308 286748
rect 36728 286696 36780 286748
rect 547880 286152 547932 286204
rect 548156 286152 548208 286204
rect 15108 285676 15160 285728
rect 16580 285676 16632 285728
rect 71872 284248 71924 284300
rect 100024 284248 100076 284300
rect 25688 284180 25740 284232
rect 36636 284180 36688 284232
rect 42892 284180 42944 284232
rect 15292 284112 15344 284164
rect 43996 284112 44048 284164
rect 53656 284180 53708 284232
rect 66904 284180 66956 284232
rect 81992 284180 82044 284232
rect 93124 284180 93176 284232
rect 99472 284180 99524 284232
rect 127992 284248 128044 284300
rect 165988 284248 166040 284300
rect 177304 284248 177356 284300
rect 178684 284248 178736 284300
rect 184020 284248 184072 284300
rect 109684 284180 109736 284232
rect 122104 284180 122156 284232
rect 137652 284180 137704 284232
rect 148416 284180 148468 284232
rect 183652 284180 183704 284232
rect 211712 284248 211764 284300
rect 277676 284248 277728 284300
rect 289084 284248 289136 284300
rect 306012 284248 306064 284300
rect 316684 284248 316736 284300
rect 361672 284248 361724 284300
rect 373264 284248 373316 284300
rect 374644 284248 374696 284300
rect 379704 284248 379756 284300
rect 193680 284180 193732 284232
rect 204996 284180 205048 284232
rect 222016 284180 222068 284232
rect 232596 284180 232648 284232
rect 249708 284180 249760 284232
rect 260104 284180 260156 284232
rect 333704 284180 333756 284232
rect 344284 284180 344336 284232
rect 379612 284180 379664 284232
rect 408040 284248 408092 284300
rect 474004 284248 474056 284300
rect 485044 284248 485096 284300
rect 501696 284248 501748 284300
rect 512644 284248 512696 284300
rect 548156 284248 548208 284300
rect 557540 284248 557592 284300
rect 390008 284180 390060 284232
rect 400864 284180 400916 284232
rect 417700 284180 417752 284232
rect 428464 284180 428516 284232
rect 445668 284180 445720 284232
rect 456064 284180 456116 284232
rect 529664 284180 529716 284232
rect 540244 284180 540296 284232
rect 72056 284112 72108 284164
rect 127072 284112 127124 284164
rect 156052 284112 156104 284164
rect 238852 284112 238904 284164
rect 268016 284112 268068 284164
rect 323032 284112 323084 284164
rect 352012 284112 352064 284164
rect 434812 284112 434864 284164
rect 463700 284112 463752 284164
rect 518992 284112 519044 284164
rect 547880 284112 547932 284164
rect 26240 280372 26292 280424
rect 35440 280372 35492 280424
rect 71872 280372 71924 280424
rect 71136 280304 71188 280356
rect 36636 280236 36688 280288
rect 53932 280236 53984 280288
rect 39304 280168 39356 280220
rect 44272 280168 44324 280220
rect 66904 280168 66956 280220
rect 72608 280168 72660 280220
rect 352012 280372 352064 280424
rect 99472 280304 99524 280356
rect 100392 280304 100444 280356
rect 183652 280304 183704 280356
rect 222292 280304 222344 280356
rect 267004 280304 267056 280356
rect 277952 280304 278004 280356
rect 295432 280304 295484 280356
rect 334256 280304 334308 280356
rect 347044 280304 347096 280356
rect 109960 280236 110012 280288
rect 124864 280236 124916 280288
rect 128636 280236 128688 280288
rect 151084 280236 151136 280288
rect 156604 280236 156656 280288
rect 182824 280236 182876 280288
rect 193956 280236 194008 280288
rect 232504 280236 232556 280288
rect 82268 280168 82320 280220
rect 93124 280168 93176 280220
rect 100300 280168 100352 280220
rect 100392 280168 100444 280220
rect 138296 280168 138348 280220
rect 149704 280168 149756 280220
rect 166264 280168 166316 280220
rect 177304 280168 177356 280220
rect 184296 280168 184348 280220
rect 233976 280168 234028 280220
rect 240600 280168 240652 280220
rect 267832 280236 267884 280288
rect 306288 280236 306340 280288
rect 250260 280168 250312 280220
rect 261484 280168 261536 280220
rect 268292 280168 268344 280220
rect 289084 280168 289136 280220
rect 296628 280168 296680 280220
rect 318064 280168 318116 280220
rect 324596 280168 324648 280220
rect 348424 280168 348476 280220
rect 352288 280168 352340 280220
rect 463792 280372 463844 280424
rect 379612 280304 379664 280356
rect 418252 280304 418304 280356
rect 390284 280236 390336 280288
rect 400864 280236 400916 280288
rect 408592 280236 408644 280288
rect 429844 280236 429896 280288
rect 436284 280236 436336 280288
rect 457444 280236 457496 280288
rect 464620 280236 464672 280288
rect 491392 280304 491444 280356
rect 529940 280304 529992 280356
rect 502248 280236 502300 280288
rect 541624 280236 541676 280288
rect 361948 280168 362000 280220
rect 373264 280168 373316 280220
rect 380624 280168 380676 280220
rect 428464 280168 428516 280220
rect 445944 280168 445996 280220
rect 462964 280168 463016 280220
rect 474280 280168 474332 280220
rect 485044 280168 485096 280220
rect 492588 280168 492640 280220
rect 512644 280168 512696 280220
rect 520280 280168 520332 280220
rect 544384 280168 544436 280220
rect 548616 280168 548668 280220
rect 558276 280168 558328 280220
rect 568028 278400 568080 278452
rect 120172 278264 120224 278316
rect 122104 278264 122156 278316
rect 512092 278264 512144 278316
rect 514024 278264 514076 278316
rect 568028 278196 568080 278248
rect 126888 277516 126940 277568
rect 178040 277516 178092 277568
rect 182088 277516 182140 277568
rect 233240 277516 233292 277568
rect 462228 277516 462280 277568
rect 513380 277516 513432 277568
rect 42708 277448 42760 277500
rect 93860 277448 93912 277500
rect 97908 277448 97960 277500
rect 149060 277448 149112 277500
rect 154488 277448 154540 277500
rect 205640 277448 205692 277500
rect 209688 277448 209740 277500
rect 262220 277448 262272 277500
rect 266268 277448 266320 277500
rect 317420 277448 317472 277500
rect 322848 277448 322900 277500
rect 374000 277448 374052 277500
rect 378048 277448 378100 277500
rect 429292 277448 429344 277500
rect 434628 277448 434680 277500
rect 485780 277448 485832 277500
rect 518808 277448 518860 277500
rect 569960 277448 570012 277500
rect 13544 277380 13596 277432
rect 66260 277380 66312 277432
rect 70308 277380 70360 277432
rect 121460 277380 121512 277432
rect 204076 277380 204128 277432
rect 212448 277380 212500 277432
rect 238668 277380 238720 277432
rect 289820 277380 289872 277432
rect 293868 277380 293920 277432
rect 345020 277380 345072 277432
rect 350448 277380 350500 277432
rect 401600 277380 401652 277432
rect 405648 277380 405700 277432
rect 458180 277380 458232 277432
rect 489828 277380 489880 277432
rect 542360 277380 542412 277432
rect 204260 272552 204312 272604
rect 204996 272552 205048 272604
rect 400312 272552 400364 272604
rect 400956 272552 401008 272604
rect 15200 256640 15252 256692
rect 35900 256640 35952 256692
rect 36084 256640 36136 256692
rect 63592 256640 63644 256692
rect 64052 256640 64104 256692
rect 91928 256640 91980 256692
rect 92112 256640 92164 256692
rect 119620 256640 119672 256692
rect 122104 256640 122156 256692
rect 147956 256640 148008 256692
rect 148048 256640 148100 256692
rect 175924 256640 175976 256692
rect 176108 256640 176160 256692
rect 203616 256640 203668 256692
rect 204996 256640 205048 256692
rect 231952 256640 232004 256692
rect 232044 256640 232096 256692
rect 259920 256640 259972 256692
rect 260104 256640 260156 256692
rect 287612 256640 287664 256692
rect 288072 256640 288124 256692
rect 315948 256640 316000 256692
rect 316684 256640 316736 256692
rect 343916 256640 343968 256692
rect 344100 256640 344152 256692
rect 371608 256640 371660 256692
rect 372068 256640 372120 256692
rect 399944 256640 399996 256692
rect 400956 256640 401008 256692
rect 427912 256640 427964 256692
rect 428096 256640 428148 256692
rect 455604 256640 455656 256692
rect 456064 256640 456116 256692
rect 483940 256640 483992 256692
rect 484032 256640 484084 256692
rect 511908 256640 511960 256692
rect 514024 256640 514076 256692
rect 539600 256640 539652 256692
rect 540060 256640 540112 256692
rect 567936 256640 567988 256692
rect 16580 256572 16632 256624
rect 36636 256572 36688 256624
rect 44916 256572 44968 256624
rect 71136 256572 71188 256624
rect 82268 256572 82320 256624
rect 93124 256572 93176 256624
rect 110328 256572 110380 256624
rect 124864 256572 124916 256624
rect 128636 256572 128688 256624
rect 149704 256572 149756 256624
rect 156604 256572 156656 256624
rect 182824 256572 182876 256624
rect 194508 256572 194560 256624
rect 204076 256572 204128 256624
rect 212632 256572 212684 256624
rect 232504 256572 232556 256624
rect 240600 256572 240652 256624
rect 267004 256572 267056 256624
rect 278596 256572 278648 256624
rect 289084 256572 289136 256624
rect 306288 256572 306340 256624
rect 318064 256572 318116 256624
rect 324596 256572 324648 256624
rect 347044 256572 347096 256624
rect 362592 256572 362644 256624
rect 373264 256572 373316 256624
rect 390284 256572 390336 256624
rect 400864 256572 400916 256624
rect 408592 256572 408644 256624
rect 428464 256572 428516 256624
rect 436928 256572 436980 256624
rect 462964 256572 463016 256624
rect 474280 256572 474332 256624
rect 485044 256572 485096 256624
rect 502248 256572 502300 256624
rect 512644 256572 512696 256624
rect 520924 256572 520976 256624
rect 541624 256572 541676 256624
rect 26240 256504 26292 256556
rect 39304 256504 39356 256556
rect 54576 256504 54628 256556
rect 66904 256504 66956 256556
rect 138296 256504 138348 256556
rect 151084 256504 151136 256556
rect 166264 256504 166316 256556
rect 177304 256504 177356 256556
rect 222292 256504 222344 256556
rect 233976 256504 234028 256556
rect 250260 256504 250312 256556
rect 261484 256504 261536 256556
rect 334256 256504 334308 256556
rect 348424 256504 348476 256556
rect 418252 256504 418304 256556
rect 429844 256504 429896 256556
rect 446588 256504 446640 256556
rect 457444 256504 457496 256556
rect 530584 256504 530636 256556
rect 544384 256504 544436 256556
rect 558276 255960 558328 256012
rect 567476 255960 567528 256012
rect 548340 254532 548392 254584
rect 568120 254532 568172 254584
rect 212356 254124 212408 254176
rect 232688 254124 232740 254176
rect 296352 254124 296404 254176
rect 316776 254124 316828 254176
rect 408040 254124 408092 254176
rect 428648 254124 428700 254176
rect 492036 254124 492088 254176
rect 512736 254124 512788 254176
rect 2780 254056 2832 254108
rect 5080 254056 5132 254108
rect 148416 254056 148468 254108
rect 165712 254056 165764 254108
rect 175464 254056 175516 254108
rect 193680 254056 193732 254108
rect 203524 254056 203576 254108
rect 221372 254056 221424 254108
rect 260104 254056 260156 254108
rect 277676 254056 277728 254108
rect 287520 254056 287572 254108
rect 305368 254056 305420 254108
rect 345664 254056 345716 254108
rect 361672 254056 361724 254108
rect 371516 254056 371568 254108
rect 389364 254056 389416 254108
rect 399484 254056 399536 254108
rect 417700 254056 417752 254108
rect 456064 254056 456116 254108
rect 473360 254056 473412 254108
rect 483480 254056 483532 254108
rect 501696 254056 501748 254108
rect 36728 253988 36780 254040
rect 53656 253988 53708 254040
rect 64420 253988 64472 254040
rect 81440 253988 81492 254040
rect 91468 253988 91520 254040
rect 109684 253988 109736 254040
rect 119436 253988 119488 254040
rect 137652 253988 137704 254040
rect 156328 253988 156380 254040
rect 178684 253988 178736 254040
rect 232504 253988 232556 254040
rect 249708 253988 249760 254040
rect 268016 253988 268068 254040
rect 287704 253988 287756 254040
rect 315488 253988 315540 254040
rect 333704 253988 333756 254040
rect 352012 253988 352064 254040
rect 374644 253988 374696 254040
rect 428556 253988 428608 254040
rect 445668 253988 445720 254040
rect 464344 253988 464396 254040
rect 483664 253988 483716 254040
rect 511448 253988 511500 254040
rect 529664 253988 529716 254040
rect 541624 253988 541676 254040
rect 557540 253988 557592 254040
rect 15108 253920 15160 253972
rect 25688 253920 25740 253972
rect 36636 253920 36688 253972
rect 63316 253920 63368 253972
rect 66904 253920 66956 253972
rect 91100 253920 91152 253972
rect 93124 253920 93176 253972
rect 119344 253920 119396 253972
rect 122104 253920 122156 253972
rect 147312 253920 147364 253972
rect 148324 253920 148376 253972
rect 175372 253920 175424 253972
rect 177304 253920 177356 253972
rect 203340 253920 203392 253972
rect 204996 253920 205048 253972
rect 231032 253920 231084 253972
rect 232596 253920 232648 253972
rect 259368 253920 259420 253972
rect 260196 253920 260248 253972
rect 287336 253920 287388 253972
rect 289084 253920 289136 253972
rect 315028 253920 315080 253972
rect 316684 253920 316736 253972
rect 343364 253920 343416 253972
rect 344284 253920 344336 253972
rect 371332 253920 371384 253972
rect 373264 253920 373316 253972
rect 399024 253920 399076 253972
rect 400864 253920 400916 253972
rect 427360 253920 427412 253972
rect 428464 253920 428516 253972
rect 455328 253920 455380 253972
rect 456156 253920 456208 253972
rect 483020 253920 483072 253972
rect 485044 253920 485096 253972
rect 511356 253920 511408 253972
rect 512644 253920 512696 253972
rect 539324 253920 539376 253972
rect 540244 253920 540296 253972
rect 567200 253920 567252 253972
rect 350448 251336 350500 251388
rect 401600 251336 401652 251388
rect 462228 251336 462280 251388
rect 513380 251336 513432 251388
rect 42708 251268 42760 251320
rect 126888 251268 126940 251320
rect 178040 251268 178092 251320
rect 182088 251268 182140 251320
rect 233240 251268 233292 251320
rect 238668 251268 238720 251320
rect 289820 251268 289872 251320
rect 293868 251268 293920 251320
rect 345020 251268 345072 251320
rect 378048 251268 378100 251320
rect 429292 251268 429344 251320
rect 434628 251268 434680 251320
rect 485780 251268 485832 251320
rect 518808 251268 518860 251320
rect 569960 251268 570012 251320
rect 93860 251200 93912 251252
rect 97908 251200 97960 251252
rect 149060 251200 149112 251252
rect 154488 251200 154540 251252
rect 205640 251200 205692 251252
rect 209688 251200 209740 251252
rect 262220 251200 262272 251252
rect 266268 251200 266320 251252
rect 317420 251200 317472 251252
rect 322848 251200 322900 251252
rect 374000 251200 374052 251252
rect 405648 251200 405700 251252
rect 458180 251200 458232 251252
rect 489828 251200 489880 251252
rect 542360 251200 542412 251252
rect 42892 249772 42944 249824
rect 43628 249772 43680 249824
rect 2780 240184 2832 240236
rect 5172 240184 5224 240236
rect 63592 235356 63644 235408
rect 64420 235356 64472 235408
rect 147680 235356 147732 235408
rect 148416 235356 148468 235408
rect 512736 234200 512788 234252
rect 519636 234200 519688 234252
rect 428648 233860 428700 233912
rect 435732 233860 435784 233912
rect 232688 233520 232740 233572
rect 239772 233520 239824 233572
rect 287704 233520 287756 233572
rect 295708 233520 295760 233572
rect 316776 233384 316828 233436
rect 323676 233384 323728 233436
rect 483664 233384 483716 233436
rect 491668 233384 491720 233436
rect 13544 233180 13596 233232
rect 66260 233180 66312 233232
rect 70308 233180 70360 233232
rect 121460 233180 121512 233232
rect 427728 233180 427780 233232
rect 428556 233180 428608 233232
rect 539508 233180 539560 233232
rect 541624 233180 541676 233232
rect 15108 232704 15160 232756
rect 16580 232704 16632 232756
rect 343640 232704 343692 232756
rect 345664 232704 345716 232756
rect 547880 232704 547932 232756
rect 548156 232704 548208 232756
rect 35348 231888 35400 231940
rect 36728 231888 36780 231940
rect 149704 231820 149756 231872
rect 579804 231820 579856 231872
rect 71872 230392 71924 230444
rect 100024 230392 100076 230444
rect 25688 230324 25740 230376
rect 36636 230324 36688 230376
rect 42892 230324 42944 230376
rect 15292 230256 15344 230308
rect 43996 230256 44048 230308
rect 53656 230324 53708 230376
rect 66904 230324 66956 230376
rect 81992 230324 82044 230376
rect 93124 230324 93176 230376
rect 99472 230324 99524 230376
rect 127992 230392 128044 230444
rect 165988 230392 166040 230444
rect 177304 230392 177356 230444
rect 178684 230392 178736 230444
rect 184020 230392 184072 230444
rect 109684 230324 109736 230376
rect 122104 230324 122156 230376
rect 137652 230324 137704 230376
rect 148324 230324 148376 230376
rect 183652 230324 183704 230376
rect 211712 230392 211764 230444
rect 277676 230392 277728 230444
rect 289084 230392 289136 230444
rect 306012 230392 306064 230444
rect 316684 230392 316736 230444
rect 361672 230392 361724 230444
rect 373264 230392 373316 230444
rect 379612 230392 379664 230444
rect 408040 230392 408092 230444
rect 474004 230392 474056 230444
rect 485044 230392 485096 230444
rect 501696 230392 501748 230444
rect 512644 230392 512696 230444
rect 548156 230392 548208 230444
rect 557540 230392 557592 230444
rect 193680 230324 193732 230376
rect 204996 230324 205048 230376
rect 222016 230324 222068 230376
rect 232596 230324 232648 230376
rect 249708 230324 249760 230376
rect 260196 230324 260248 230376
rect 333704 230324 333756 230376
rect 344284 230324 344336 230376
rect 374644 230324 374696 230376
rect 379704 230324 379756 230376
rect 390008 230324 390060 230376
rect 400864 230324 400916 230376
rect 417700 230324 417752 230376
rect 428464 230324 428516 230376
rect 445668 230324 445720 230376
rect 456156 230324 456208 230376
rect 529664 230324 529716 230376
rect 540244 230324 540296 230376
rect 72056 230256 72108 230308
rect 127072 230256 127124 230308
rect 156052 230256 156104 230308
rect 238852 230256 238904 230308
rect 268016 230256 268068 230308
rect 323032 230256 323084 230308
rect 352012 230256 352064 230308
rect 434812 230256 434864 230308
rect 463700 230256 463752 230308
rect 518992 230256 519044 230308
rect 547880 230256 547932 230308
rect 26240 226448 26292 226500
rect 35440 226448 35492 226500
rect 71136 226448 71188 226500
rect 82268 226448 82320 226500
rect 184204 226448 184256 226500
rect 222292 226448 222344 226500
rect 261484 226448 261536 226500
rect 268292 226448 268344 226500
rect 296168 226448 296220 226500
rect 334256 226448 334308 226500
rect 352196 226448 352248 226500
rect 36636 226380 36688 226432
rect 53932 226380 53984 226432
rect 72240 226380 72292 226432
rect 109960 226380 110012 226432
rect 124864 226380 124916 226432
rect 128636 226380 128688 226432
rect 152464 226380 152516 226432
rect 156604 226380 156656 226432
rect 182824 226380 182876 226432
rect 193956 226380 194008 226432
rect 232504 226380 232556 226432
rect 39304 226312 39356 226364
rect 44272 226312 44324 226364
rect 66904 226312 66956 226364
rect 72608 226312 72660 226364
rect 93124 226312 93176 226364
rect 100300 226312 100352 226364
rect 100208 226244 100260 226296
rect 138296 226312 138348 226364
rect 151084 226312 151136 226364
rect 166264 226312 166316 226364
rect 177304 226312 177356 226364
rect 184296 226312 184348 226364
rect 233976 226312 234028 226364
rect 240600 226312 240652 226364
rect 268200 226380 268252 226432
rect 306288 226380 306340 226432
rect 347044 226380 347096 226432
rect 361948 226380 362000 226432
rect 380256 226448 380308 226500
rect 418252 226448 418304 226500
rect 462964 226448 463016 226500
rect 474280 226448 474332 226500
rect 492128 226448 492180 226500
rect 529940 226448 529992 226500
rect 390284 226380 390336 226432
rect 400956 226380 401008 226432
rect 408592 226380 408644 226432
rect 429844 226380 429896 226432
rect 436284 226380 436336 226432
rect 464160 226380 464212 226432
rect 502248 226380 502300 226432
rect 512644 226380 512696 226432
rect 520280 226380 520332 226432
rect 541624 226380 541676 226432
rect 250260 226312 250312 226364
rect 267004 226312 267056 226364
rect 277952 226312 278004 226364
rect 289084 226312 289136 226364
rect 296628 226312 296680 226364
rect 318064 226312 318116 226364
rect 324596 226312 324648 226364
rect 348424 226312 348476 226364
rect 352288 226312 352340 226364
rect 373264 226312 373316 226364
rect 380624 226312 380676 226364
rect 428464 226312 428516 226364
rect 445944 226312 445996 226364
rect 457444 226312 457496 226364
rect 464620 226312 464672 226364
rect 485044 226312 485096 226364
rect 492588 226312 492640 226364
rect 544384 226312 544436 226364
rect 548616 226312 548668 226364
rect 558276 226312 558328 226364
rect 568028 224408 568080 224460
rect 120172 224272 120224 224324
rect 122104 224272 122156 224324
rect 210424 224272 210476 224324
rect 212448 224272 212500 224324
rect 512184 224272 512236 224324
rect 514024 224272 514076 224324
rect 568028 224204 568080 224256
rect 182088 223728 182140 223780
rect 233240 223728 233292 223780
rect 350448 223728 350500 223780
rect 401600 223728 401652 223780
rect 462228 223728 462280 223780
rect 513380 223728 513432 223780
rect 42708 223660 42760 223712
rect 93860 223660 93912 223712
rect 97908 223660 97960 223712
rect 149060 223660 149112 223712
rect 154488 223660 154540 223712
rect 205640 223660 205692 223712
rect 238668 223660 238720 223712
rect 289820 223660 289872 223712
rect 293868 223660 293920 223712
rect 345020 223660 345072 223712
rect 378048 223660 378100 223712
rect 429292 223660 429344 223712
rect 434628 223660 434680 223712
rect 485780 223660 485832 223712
rect 518808 223660 518860 223712
rect 569960 223660 570012 223712
rect 13544 223592 13596 223644
rect 66260 223592 66312 223644
rect 70308 223592 70360 223644
rect 121460 223592 121512 223644
rect 126888 223592 126940 223644
rect 178040 223592 178092 223644
rect 209688 223592 209740 223644
rect 262220 223592 262272 223644
rect 266268 223592 266320 223644
rect 317420 223592 317472 223644
rect 322848 223592 322900 223644
rect 374000 223592 374052 223644
rect 405648 223592 405700 223644
rect 458180 223592 458232 223644
rect 489828 223592 489880 223644
rect 542360 223592 542412 223644
rect 204260 221824 204312 221876
rect 204996 221824 205048 221876
rect 64052 219716 64104 219768
rect 64420 219716 64472 219768
rect 231860 203940 231912 203992
rect 232136 203940 232188 203992
rect 15200 202784 15252 202836
rect 35900 202784 35952 202836
rect 36084 202784 36136 202836
rect 63592 202784 63644 202836
rect 64420 202784 64472 202836
rect 91928 202784 91980 202836
rect 92112 202784 92164 202836
rect 119620 202784 119672 202836
rect 122104 202784 122156 202836
rect 147680 202784 147732 202836
rect 148048 202784 148100 202836
rect 175924 202784 175976 202836
rect 176108 202784 176160 202836
rect 203616 202784 203668 202836
rect 204996 202784 205048 202836
rect 231860 202784 231912 202836
rect 232044 202784 232096 202836
rect 259920 202784 259972 202836
rect 260104 202784 260156 202836
rect 287612 202784 287664 202836
rect 288072 202784 288124 202836
rect 315948 202784 316000 202836
rect 316684 202784 316736 202836
rect 343916 202784 343968 202836
rect 344100 202784 344152 202836
rect 371608 202784 371660 202836
rect 372068 202784 372120 202836
rect 399944 202784 399996 202836
rect 400864 202784 400916 202836
rect 427912 202784 427964 202836
rect 428096 202784 428148 202836
rect 455604 202784 455656 202836
rect 456064 202784 456116 202836
rect 483940 202784 483992 202836
rect 484032 202784 484084 202836
rect 511908 202784 511960 202836
rect 514024 202784 514076 202836
rect 539600 202784 539652 202836
rect 540060 202784 540112 202836
rect 567936 202784 567988 202836
rect 16856 202716 16908 202768
rect 36636 202716 36688 202768
rect 44916 202716 44968 202768
rect 71136 202716 71188 202768
rect 82268 202716 82320 202768
rect 93124 202716 93176 202768
rect 110236 202716 110288 202768
rect 124864 202716 124916 202768
rect 128912 202716 128964 202768
rect 151084 202716 151136 202768
rect 156604 202716 156656 202768
rect 182824 202716 182876 202768
rect 194508 202716 194560 202768
rect 210424 202716 210476 202768
rect 213000 202716 213052 202768
rect 232504 202716 232556 202768
rect 240600 202716 240652 202768
rect 267004 202716 267056 202768
rect 278596 202716 278648 202768
rect 289084 202716 289136 202768
rect 306288 202716 306340 202768
rect 318064 202716 318116 202768
rect 324596 202716 324648 202768
rect 347044 202716 347096 202768
rect 362592 202716 362644 202768
rect 373264 202716 373316 202768
rect 390284 202716 390336 202768
rect 400956 202716 401008 202768
rect 408592 202716 408644 202768
rect 428464 202716 428516 202768
rect 436928 202716 436980 202768
rect 462964 202716 463016 202768
rect 474280 202716 474332 202768
rect 485044 202716 485096 202768
rect 502248 202716 502300 202768
rect 512644 202716 512696 202768
rect 520924 202716 520976 202768
rect 541624 202716 541676 202768
rect 26608 202648 26660 202700
rect 39304 202648 39356 202700
rect 54576 202648 54628 202700
rect 66904 202648 66956 202700
rect 138664 202648 138716 202700
rect 152464 202648 152516 202700
rect 166264 202648 166316 202700
rect 177304 202648 177356 202700
rect 222568 202648 222620 202700
rect 233976 202648 234028 202700
rect 250260 202648 250312 202700
rect 261484 202648 261536 202700
rect 334256 202648 334308 202700
rect 348424 202648 348476 202700
rect 418252 202648 418304 202700
rect 429844 202648 429896 202700
rect 446588 202648 446640 202700
rect 457444 202648 457496 202700
rect 530584 202648 530636 202700
rect 544384 202648 544436 202700
rect 558276 202104 558328 202156
rect 567476 202104 567528 202156
rect 3056 201492 3108 201544
rect 64052 201492 64104 201544
rect 548340 200744 548392 200796
rect 568120 200744 568172 200796
rect 296352 200336 296404 200388
rect 316776 200336 316828 200388
rect 408040 200336 408092 200388
rect 428648 200336 428700 200388
rect 492036 200336 492088 200388
rect 512736 200336 512788 200388
rect 148416 200268 148468 200320
rect 165620 200268 165672 200320
rect 175464 200268 175516 200320
rect 193680 200268 193732 200320
rect 203524 200268 203576 200320
rect 221372 200268 221424 200320
rect 232504 200268 232556 200320
rect 249708 200268 249760 200320
rect 260196 200268 260248 200320
rect 277676 200268 277728 200320
rect 287520 200268 287572 200320
rect 305368 200268 305420 200320
rect 345664 200268 345716 200320
rect 361672 200268 361724 200320
rect 371516 200268 371568 200320
rect 389364 200268 389416 200320
rect 399484 200268 399536 200320
rect 417700 200268 417752 200320
rect 456156 200268 456208 200320
rect 473544 200268 473596 200320
rect 483480 200268 483532 200320
rect 501696 200268 501748 200320
rect 36728 200200 36780 200252
rect 53656 200200 53708 200252
rect 64420 200200 64472 200252
rect 81440 200200 81492 200252
rect 91468 200200 91520 200252
rect 109684 200200 109736 200252
rect 119436 200200 119488 200252
rect 137652 200200 137704 200252
rect 156328 200200 156380 200252
rect 178684 200200 178736 200252
rect 212264 200200 212316 200252
rect 232688 200200 232740 200252
rect 268016 200200 268068 200252
rect 287704 200200 287756 200252
rect 315488 200200 315540 200252
rect 333704 200200 333756 200252
rect 352012 200200 352064 200252
rect 374644 200200 374696 200252
rect 428464 200200 428516 200252
rect 445668 200200 445720 200252
rect 464344 200200 464396 200252
rect 483664 200200 483716 200252
rect 511448 200200 511500 200252
rect 529664 200200 529716 200252
rect 541624 200200 541676 200252
rect 557540 200200 557592 200252
rect 15108 200132 15160 200184
rect 25688 200132 25740 200184
rect 36636 200132 36688 200184
rect 63316 200132 63368 200184
rect 66904 200132 66956 200184
rect 91100 200132 91152 200184
rect 93124 200132 93176 200184
rect 119344 200132 119396 200184
rect 124864 200132 124916 200184
rect 147312 200132 147364 200184
rect 148324 200132 148376 200184
rect 175280 200132 175332 200184
rect 177304 200132 177356 200184
rect 203340 200132 203392 200184
rect 204996 200132 205048 200184
rect 231032 200132 231084 200184
rect 232596 200132 232648 200184
rect 259368 200132 259420 200184
rect 260104 200132 260156 200184
rect 287336 200132 287388 200184
rect 289084 200132 289136 200184
rect 315028 200132 315080 200184
rect 316684 200132 316736 200184
rect 343364 200132 343416 200184
rect 344284 200132 344336 200184
rect 371332 200132 371384 200184
rect 373264 200132 373316 200184
rect 399024 200132 399076 200184
rect 400864 200132 400916 200184
rect 427360 200132 427412 200184
rect 428556 200132 428608 200184
rect 455328 200132 455380 200184
rect 456064 200132 456116 200184
rect 483204 200132 483256 200184
rect 485044 200132 485096 200184
rect 511356 200132 511408 200184
rect 512644 200132 512696 200184
rect 539324 200132 539376 200184
rect 540244 200132 540296 200184
rect 567200 200132 567252 200184
rect 42892 193808 42944 193860
rect 43628 193808 43680 193860
rect 570696 191836 570748 191888
rect 580172 191836 580224 191888
rect 2964 187688 3016 187740
rect 11796 187688 11848 187740
rect 147680 185580 147732 185632
rect 148416 185580 148468 185632
rect 259736 185580 259788 185632
rect 260196 185580 260248 185632
rect 455696 185580 455748 185632
rect 456156 185580 456208 185632
rect 63592 181432 63644 181484
rect 64420 181432 64472 181484
rect 512736 180208 512788 180260
rect 519636 180208 519688 180260
rect 428648 180072 428700 180124
rect 435732 180072 435784 180124
rect 232688 179868 232740 179920
rect 239772 179868 239824 179920
rect 483664 179664 483716 179716
rect 491668 179664 491720 179716
rect 316776 179460 316828 179512
rect 323676 179460 323728 179512
rect 287704 179392 287756 179444
rect 295708 179392 295760 179444
rect 13544 179324 13596 179376
rect 66260 179324 66312 179376
rect 70308 179324 70360 179376
rect 121460 179324 121512 179376
rect 126888 179324 126940 179376
rect 178040 179324 178092 179376
rect 209688 179324 209740 179376
rect 262220 179324 262272 179376
rect 266268 179324 266320 179376
rect 317420 179324 317472 179376
rect 322848 179324 322900 179376
rect 374000 179324 374052 179376
rect 405648 179324 405700 179376
rect 458180 179324 458232 179376
rect 489828 179324 489880 179376
rect 42708 179256 42760 179308
rect 93860 179256 93912 179308
rect 97908 179256 97960 179308
rect 149060 179256 149112 179308
rect 154488 179256 154540 179308
rect 205640 179256 205692 179308
rect 238668 179256 238720 179308
rect 289820 179256 289872 179308
rect 293868 179256 293920 179308
rect 182088 179188 182140 179240
rect 233240 179188 233292 179240
rect 343548 179256 343600 179308
rect 345664 179256 345716 179308
rect 378048 179256 378100 179308
rect 429292 179256 429344 179308
rect 434628 179256 434680 179308
rect 485780 179256 485832 179308
rect 518808 179256 518860 179308
rect 345020 179188 345072 179240
rect 350448 179188 350500 179240
rect 401600 179188 401652 179240
rect 462228 179188 462280 179240
rect 513380 179188 513432 179240
rect 539508 179324 539560 179376
rect 541624 179324 541676 179376
rect 542360 179188 542412 179240
rect 569960 179256 570012 179308
rect 15108 178712 15160 178764
rect 16580 178712 16632 178764
rect 35256 178712 35308 178764
rect 36728 178712 36780 178764
rect 547880 178712 547932 178764
rect 548156 178712 548208 178764
rect 71872 176604 71924 176656
rect 100024 176604 100076 176656
rect 25688 176536 25740 176588
rect 36636 176536 36688 176588
rect 42892 176536 42944 176588
rect 15292 176468 15344 176520
rect 43996 176468 44048 176520
rect 53656 176536 53708 176588
rect 66904 176536 66956 176588
rect 81992 176536 82044 176588
rect 93124 176536 93176 176588
rect 99472 176536 99524 176588
rect 127992 176604 128044 176656
rect 165988 176604 166040 176656
rect 177304 176604 177356 176656
rect 178684 176604 178736 176656
rect 184020 176604 184072 176656
rect 109684 176536 109736 176588
rect 124864 176536 124916 176588
rect 137652 176536 137704 176588
rect 148324 176536 148376 176588
rect 183652 176536 183704 176588
rect 211712 176604 211764 176656
rect 277676 176604 277728 176656
rect 289084 176604 289136 176656
rect 306012 176604 306064 176656
rect 316684 176604 316736 176656
rect 361672 176604 361724 176656
rect 373264 176604 373316 176656
rect 374644 176604 374696 176656
rect 379704 176604 379756 176656
rect 193680 176536 193732 176588
rect 204996 176536 205048 176588
rect 222016 176536 222068 176588
rect 232596 176536 232648 176588
rect 249708 176536 249760 176588
rect 260104 176536 260156 176588
rect 333704 176536 333756 176588
rect 344284 176536 344336 176588
rect 379612 176536 379664 176588
rect 408040 176604 408092 176656
rect 474004 176604 474056 176656
rect 485044 176604 485096 176656
rect 501696 176604 501748 176656
rect 512644 176604 512696 176656
rect 548156 176604 548208 176656
rect 557540 176604 557592 176656
rect 390008 176536 390060 176588
rect 400864 176536 400916 176588
rect 417700 176536 417752 176588
rect 428556 176536 428608 176588
rect 445668 176536 445720 176588
rect 456064 176536 456116 176588
rect 529664 176536 529716 176588
rect 540244 176536 540296 176588
rect 72056 176468 72108 176520
rect 127072 176468 127124 176520
rect 156052 176468 156104 176520
rect 238852 176468 238904 176520
rect 268016 176468 268068 176520
rect 323032 176468 323084 176520
rect 352012 176468 352064 176520
rect 434812 176468 434864 176520
rect 463700 176468 463752 176520
rect 518992 176468 519044 176520
rect 547880 176468 547932 176520
rect 26240 172796 26292 172848
rect 35440 172796 35492 172848
rect 71136 172660 71188 172712
rect 82268 172660 82320 172712
rect 99380 172660 99432 172712
rect 100300 172660 100352 172712
rect 183652 172660 183704 172712
rect 222292 172660 222344 172712
rect 261484 172660 261536 172712
rect 268292 172660 268344 172712
rect 295432 172660 295484 172712
rect 334256 172660 334308 172712
rect 352012 172660 352064 172712
rect 36636 172592 36688 172644
rect 53932 172592 53984 172644
rect 71872 172592 71924 172644
rect 109960 172592 110012 172644
rect 124864 172592 124916 172644
rect 128636 172592 128688 172644
rect 152464 172592 152516 172644
rect 156604 172592 156656 172644
rect 182824 172592 182876 172644
rect 193956 172592 194008 172644
rect 232504 172592 232556 172644
rect 39304 172524 39356 172576
rect 44272 172524 44324 172576
rect 66904 172524 66956 172576
rect 72608 172524 72660 172576
rect 93124 172524 93176 172576
rect 99380 172524 99432 172576
rect 99472 172524 99524 172576
rect 138296 172524 138348 172576
rect 151084 172524 151136 172576
rect 166264 172524 166316 172576
rect 177304 172524 177356 172576
rect 184296 172524 184348 172576
rect 233976 172524 234028 172576
rect 240600 172524 240652 172576
rect 267832 172592 267884 172644
rect 306288 172592 306340 172644
rect 345664 172592 345716 172644
rect 361948 172592 362000 172644
rect 379612 172660 379664 172712
rect 418252 172660 418304 172712
rect 463792 172660 463844 172712
rect 390284 172592 390336 172644
rect 400956 172592 401008 172644
rect 408592 172592 408644 172644
rect 429844 172592 429896 172644
rect 436284 172592 436336 172644
rect 457444 172592 457496 172644
rect 464620 172592 464672 172644
rect 485044 172660 485096 172712
rect 492588 172660 492640 172712
rect 502248 172592 502300 172644
rect 514024 172592 514076 172644
rect 520280 172592 520332 172644
rect 541624 172592 541676 172644
rect 250260 172524 250312 172576
rect 267004 172524 267056 172576
rect 277952 172524 278004 172576
rect 289084 172524 289136 172576
rect 296628 172524 296680 172576
rect 318064 172524 318116 172576
rect 324596 172524 324648 172576
rect 347044 172524 347096 172576
rect 352288 172524 352340 172576
rect 373264 172524 373316 172576
rect 380624 172524 380676 172576
rect 428464 172524 428516 172576
rect 445944 172524 445996 172576
rect 462964 172524 463016 172576
rect 474280 172524 474332 172576
rect 491392 172524 491444 172576
rect 529940 172524 529992 172576
rect 544384 172524 544436 172576
rect 548616 172524 548668 172576
rect 558276 172524 558328 172576
rect 210424 171096 210476 171148
rect 212632 171096 212684 171148
rect 568028 170416 568080 170468
rect 63776 170280 63828 170332
rect 65800 170280 65852 170332
rect 120172 170280 120224 170332
rect 122104 170280 122156 170332
rect 568028 170212 568080 170264
rect 204260 165860 204312 165912
rect 204996 165860 205048 165912
rect 13544 151716 13596 151768
rect 66260 151716 66312 151768
rect 70308 151716 70360 151768
rect 121460 151716 121512 151768
rect 126888 151716 126940 151768
rect 178040 151716 178092 151768
rect 209688 151716 209740 151768
rect 262220 151716 262272 151768
rect 266268 151716 266320 151768
rect 317420 151716 317472 151768
rect 322848 151716 322900 151768
rect 374000 151716 374052 151768
rect 405648 151716 405700 151768
rect 458180 151716 458232 151768
rect 489828 151716 489880 151768
rect 542360 151716 542412 151768
rect 42708 151648 42760 151700
rect 93860 151648 93912 151700
rect 97908 151648 97960 151700
rect 149060 151648 149112 151700
rect 154488 151648 154540 151700
rect 205640 151648 205692 151700
rect 238668 151648 238720 151700
rect 289820 151648 289872 151700
rect 293868 151648 293920 151700
rect 345020 151648 345072 151700
rect 378048 151648 378100 151700
rect 429292 151648 429344 151700
rect 434628 151648 434680 151700
rect 485780 151648 485832 151700
rect 518808 151648 518860 151700
rect 569960 151648 570012 151700
rect 182088 151580 182140 151632
rect 233240 151580 233292 151632
rect 350448 151580 350500 151632
rect 401600 151580 401652 151632
rect 462228 151580 462280 151632
rect 513380 151580 513432 151632
rect 15200 148996 15252 149048
rect 35900 148996 35952 149048
rect 36084 148996 36136 149048
rect 63592 148996 63644 149048
rect 65800 148996 65852 149048
rect 91928 148996 91980 149048
rect 92112 148996 92164 149048
rect 119620 148996 119672 149048
rect 122104 148996 122156 149048
rect 147956 148996 148008 149048
rect 148048 148996 148100 149048
rect 175924 148996 175976 149048
rect 176108 148996 176160 149048
rect 203616 148996 203668 149048
rect 204996 148996 205048 149048
rect 231952 148996 232004 149048
rect 232044 148996 232096 149048
rect 259920 148996 259972 149048
rect 260104 148996 260156 149048
rect 287612 148996 287664 149048
rect 288072 148996 288124 149048
rect 315948 148996 316000 149048
rect 316684 148996 316736 149048
rect 343916 148996 343968 149048
rect 344100 148996 344152 149048
rect 371608 148996 371660 149048
rect 372068 148996 372120 149048
rect 399944 148996 399996 149048
rect 400864 148996 400916 149048
rect 427912 148996 427964 149048
rect 428096 148996 428148 149048
rect 455604 148996 455656 149048
rect 456064 148996 456116 149048
rect 483940 148996 483992 149048
rect 484032 148996 484084 149048
rect 511908 148996 511960 149048
rect 512092 148996 512144 149048
rect 539600 148996 539652 149048
rect 540060 148996 540112 149048
rect 567936 148996 567988 149048
rect 16580 148928 16632 148980
rect 36636 148928 36688 148980
rect 44916 148928 44968 148980
rect 71136 148928 71188 148980
rect 82268 148928 82320 148980
rect 93124 148928 93176 148980
rect 110236 148928 110288 148980
rect 124864 148928 124916 148980
rect 128636 148928 128688 148980
rect 151084 148928 151136 148980
rect 156604 148928 156656 148980
rect 182824 148928 182876 148980
rect 194508 148928 194560 148980
rect 210424 148928 210476 148980
rect 212632 148928 212684 148980
rect 232504 148928 232556 148980
rect 240600 148928 240652 148980
rect 267004 148928 267056 148980
rect 278596 148928 278648 148980
rect 289084 148928 289136 148980
rect 306288 148928 306340 148980
rect 318064 148928 318116 148980
rect 324596 148928 324648 148980
rect 345664 148928 345716 148980
rect 362592 148928 362644 148980
rect 373264 148928 373316 148980
rect 390284 148928 390336 148980
rect 400956 148928 401008 148980
rect 408592 148928 408644 148980
rect 428464 148928 428516 148980
rect 436928 148928 436980 148980
rect 462964 148928 463016 148980
rect 474280 148928 474332 148980
rect 485044 148928 485096 148980
rect 502248 148928 502300 148980
rect 514024 148928 514076 148980
rect 520924 148928 520976 148980
rect 541624 148928 541676 148980
rect 26240 148860 26292 148912
rect 39304 148860 39356 148912
rect 54576 148860 54628 148912
rect 66904 148860 66956 148912
rect 138296 148860 138348 148912
rect 152464 148860 152516 148912
rect 166264 148860 166316 148912
rect 177304 148860 177356 148912
rect 222292 148860 222344 148912
rect 233976 148860 234028 148912
rect 250260 148860 250312 148912
rect 261484 148860 261536 148912
rect 334256 148860 334308 148912
rect 347044 148860 347096 148912
rect 418252 148860 418304 148912
rect 429844 148860 429896 148912
rect 446588 148860 446640 148912
rect 457444 148860 457496 148912
rect 530584 148860 530636 148912
rect 544384 148860 544436 148912
rect 558276 148316 558328 148368
rect 567476 148316 567528 148368
rect 548340 146888 548392 146940
rect 568120 146888 568172 146940
rect 212356 146480 212408 146532
rect 232688 146480 232740 146532
rect 296352 146480 296404 146532
rect 316776 146480 316828 146532
rect 408040 146480 408092 146532
rect 428648 146480 428700 146532
rect 492036 146480 492088 146532
rect 512736 146480 512788 146532
rect 148324 146412 148376 146464
rect 165712 146412 165764 146464
rect 175464 146412 175516 146464
rect 193680 146412 193732 146464
rect 203524 146412 203576 146464
rect 221372 146412 221424 146464
rect 260196 146412 260248 146464
rect 277676 146412 277728 146464
rect 287520 146412 287572 146464
rect 305368 146412 305420 146464
rect 345664 146412 345716 146464
rect 361672 146412 361724 146464
rect 371516 146412 371568 146464
rect 389364 146412 389416 146464
rect 399484 146412 399536 146464
rect 417700 146412 417752 146464
rect 456156 146412 456208 146464
rect 473360 146412 473412 146464
rect 483480 146412 483532 146464
rect 501696 146412 501748 146464
rect 36636 146344 36688 146396
rect 53656 146344 53708 146396
rect 64420 146344 64472 146396
rect 81440 146344 81492 146396
rect 91468 146344 91520 146396
rect 109684 146344 109736 146396
rect 119436 146344 119488 146396
rect 137652 146344 137704 146396
rect 156328 146344 156380 146396
rect 178684 146344 178736 146396
rect 232504 146344 232556 146396
rect 249708 146344 249760 146396
rect 268016 146344 268068 146396
rect 287704 146344 287756 146396
rect 315488 146344 315540 146396
rect 333704 146344 333756 146396
rect 352012 146344 352064 146396
rect 374644 146344 374696 146396
rect 428464 146344 428516 146396
rect 445668 146344 445720 146396
rect 464344 146344 464396 146396
rect 483664 146344 483716 146396
rect 511448 146344 511500 146396
rect 529664 146344 529716 146396
rect 541624 146344 541676 146396
rect 557540 146344 557592 146396
rect 15108 146276 15160 146328
rect 25688 146276 25740 146328
rect 36728 146276 36780 146328
rect 63316 146276 63368 146328
rect 66904 146276 66956 146328
rect 91100 146276 91152 146328
rect 93124 146276 93176 146328
rect 119344 146276 119396 146328
rect 124864 146276 124916 146328
rect 147312 146276 147364 146328
rect 148416 146276 148468 146328
rect 175372 146276 175424 146328
rect 177304 146276 177356 146328
rect 203340 146276 203392 146328
rect 204996 146276 205048 146328
rect 231032 146276 231084 146328
rect 232596 146276 232648 146328
rect 259368 146276 259420 146328
rect 260104 146276 260156 146328
rect 287336 146276 287388 146328
rect 289084 146276 289136 146328
rect 315028 146276 315080 146328
rect 316684 146276 316736 146328
rect 343364 146276 343416 146328
rect 344284 146276 344336 146328
rect 371332 146276 371384 146328
rect 373264 146276 373316 146328
rect 399024 146276 399076 146328
rect 400864 146276 400916 146328
rect 427360 146276 427412 146328
rect 428556 146276 428608 146328
rect 455328 146276 455380 146328
rect 456064 146276 456116 146328
rect 483020 146276 483072 146328
rect 485044 146276 485096 146328
rect 511356 146276 511408 146328
rect 512644 146276 512696 146328
rect 539324 146276 539376 146328
rect 540244 146276 540296 146328
rect 567200 146276 567252 146328
rect 3332 136688 3384 136740
rect 9036 136688 9088 136740
rect 42892 135464 42944 135516
rect 43628 135464 43680 135516
rect 63592 128256 63644 128308
rect 64420 128256 64472 128308
rect 259736 128256 259788 128308
rect 260196 128256 260248 128308
rect 455696 128256 455748 128308
rect 456156 128256 456208 128308
rect 232688 126896 232740 126948
rect 239772 126896 239824 126948
rect 483664 126896 483716 126948
rect 491668 126896 491720 126948
rect 512736 126896 512788 126948
rect 519636 126896 519688 126948
rect 428648 126216 428700 126268
rect 435732 126216 435784 126268
rect 287704 126080 287756 126132
rect 295708 126080 295760 126132
rect 316776 126080 316828 126132
rect 323676 126080 323728 126132
rect 13544 125536 13596 125588
rect 66260 125536 66312 125588
rect 70308 125536 70360 125588
rect 121460 125536 121512 125588
rect 126888 125536 126940 125588
rect 178040 125536 178092 125588
rect 209688 125536 209740 125588
rect 262220 125536 262272 125588
rect 266268 125536 266320 125588
rect 317420 125536 317472 125588
rect 322848 125536 322900 125588
rect 374000 125536 374052 125588
rect 405648 125536 405700 125588
rect 458180 125536 458232 125588
rect 489828 125536 489880 125588
rect 542360 125536 542412 125588
rect 42708 125468 42760 125520
rect 93860 125468 93912 125520
rect 97908 125468 97960 125520
rect 149060 125468 149112 125520
rect 154488 125468 154540 125520
rect 205640 125468 205692 125520
rect 238668 125468 238720 125520
rect 289820 125468 289872 125520
rect 293868 125468 293920 125520
rect 345020 125468 345072 125520
rect 378048 125468 378100 125520
rect 429292 125468 429344 125520
rect 434628 125468 434680 125520
rect 485780 125468 485832 125520
rect 518808 125468 518860 125520
rect 569960 125468 570012 125520
rect 182088 125400 182140 125452
rect 233240 125400 233292 125452
rect 350448 125400 350500 125452
rect 401600 125400 401652 125452
rect 462228 125400 462280 125452
rect 513380 125400 513432 125452
rect 343548 124788 343600 124840
rect 345664 124788 345716 124840
rect 35256 124652 35308 124704
rect 36636 124652 36688 124704
rect 547880 124652 547932 124704
rect 548156 124652 548208 124704
rect 15108 124176 15160 124228
rect 16580 124176 16632 124228
rect 71872 122748 71924 122800
rect 100024 122748 100076 122800
rect 25688 122680 25740 122732
rect 36728 122680 36780 122732
rect 42892 122680 42944 122732
rect 15292 122612 15344 122664
rect 43996 122612 44048 122664
rect 53656 122680 53708 122732
rect 66904 122680 66956 122732
rect 81992 122680 82044 122732
rect 93124 122680 93176 122732
rect 99472 122680 99524 122732
rect 127992 122748 128044 122800
rect 165988 122748 166040 122800
rect 177304 122748 177356 122800
rect 178684 122748 178736 122800
rect 184020 122748 184072 122800
rect 109684 122680 109736 122732
rect 124864 122680 124916 122732
rect 137652 122680 137704 122732
rect 148416 122680 148468 122732
rect 183652 122680 183704 122732
rect 211712 122748 211764 122800
rect 231584 122748 231636 122800
rect 232504 122748 232556 122800
rect 277676 122748 277728 122800
rect 289084 122748 289136 122800
rect 306012 122748 306064 122800
rect 316684 122748 316736 122800
rect 361672 122748 361724 122800
rect 373264 122748 373316 122800
rect 379612 122748 379664 122800
rect 408040 122748 408092 122800
rect 474004 122748 474056 122800
rect 485044 122748 485096 122800
rect 501696 122748 501748 122800
rect 512644 122748 512696 122800
rect 539324 122748 539376 122800
rect 541624 122748 541676 122800
rect 548156 122748 548208 122800
rect 557540 122748 557592 122800
rect 193680 122680 193732 122732
rect 204996 122680 205048 122732
rect 221924 122680 221976 122732
rect 232596 122680 232648 122732
rect 249708 122680 249760 122732
rect 260104 122680 260156 122732
rect 333704 122680 333756 122732
rect 344284 122680 344336 122732
rect 374644 122680 374696 122732
rect 379704 122680 379756 122732
rect 390008 122680 390060 122732
rect 400864 122680 400916 122732
rect 417700 122680 417752 122732
rect 428556 122680 428608 122732
rect 445668 122680 445720 122732
rect 456064 122680 456116 122732
rect 529664 122680 529716 122732
rect 540244 122680 540296 122732
rect 71964 122612 72016 122664
rect 127072 122612 127124 122664
rect 155960 122612 156012 122664
rect 238852 122612 238904 122664
rect 268016 122612 268068 122664
rect 323032 122612 323084 122664
rect 352012 122612 352064 122664
rect 434812 122612 434864 122664
rect 463792 122612 463844 122664
rect 518992 122612 519044 122664
rect 547880 122612 547932 122664
rect 71136 118804 71188 118856
rect 82268 118804 82320 118856
rect 99472 118804 99524 118856
rect 138296 118804 138348 118856
rect 183652 118804 183704 118856
rect 222292 118804 222344 118856
rect 267004 118804 267056 118856
rect 277952 118804 278004 118856
rect 295432 118804 295484 118856
rect 334256 118804 334308 118856
rect 352012 118804 352064 118856
rect 26240 118736 26292 118788
rect 35440 118736 35492 118788
rect 36636 118736 36688 118788
rect 53932 118736 53984 118788
rect 71872 118736 71924 118788
rect 109960 118736 110012 118788
rect 120724 118736 120776 118788
rect 128636 118736 128688 118788
rect 151084 118736 151136 118788
rect 156604 118736 156656 118788
rect 182824 118736 182876 118788
rect 193956 118736 194008 118788
rect 232504 118736 232556 118788
rect 39304 118668 39356 118720
rect 44272 118668 44324 118720
rect 66904 118668 66956 118720
rect 72608 118668 72660 118720
rect 93124 118668 93176 118720
rect 100300 118668 100352 118720
rect 148324 118668 148376 118720
rect 166264 118668 166316 118720
rect 177304 118668 177356 118720
rect 184296 118668 184348 118720
rect 233976 118668 234028 118720
rect 240600 118668 240652 118720
rect 267832 118736 267884 118788
rect 306288 118736 306340 118788
rect 345664 118736 345716 118788
rect 361948 118736 362000 118788
rect 379612 118804 379664 118856
rect 418252 118804 418304 118856
rect 463792 118804 463844 118856
rect 390284 118736 390336 118788
rect 400956 118736 401008 118788
rect 408592 118736 408644 118788
rect 429844 118736 429896 118788
rect 436284 118736 436336 118788
rect 457444 118736 457496 118788
rect 464620 118736 464672 118788
rect 491392 118804 491444 118856
rect 250260 118668 250312 118720
rect 261484 118668 261536 118720
rect 268292 118668 268344 118720
rect 289084 118668 289136 118720
rect 296628 118668 296680 118720
rect 318064 118668 318116 118720
rect 324596 118668 324648 118720
rect 347044 118668 347096 118720
rect 352288 118668 352340 118720
rect 373264 118668 373316 118720
rect 380624 118668 380676 118720
rect 428464 118668 428516 118720
rect 445944 118668 445996 118720
rect 462964 118668 463016 118720
rect 474280 118668 474332 118720
rect 485044 118668 485096 118720
rect 492588 118668 492640 118720
rect 541624 118804 541676 118856
rect 502248 118736 502300 118788
rect 514024 118736 514076 118788
rect 520280 118736 520332 118788
rect 558276 118736 558328 118788
rect 529940 118668 529992 118720
rect 544384 118668 544436 118720
rect 548616 118668 548668 118720
rect 547972 118600 548024 118652
rect 567936 118668 567988 118720
rect 63776 116288 63828 116340
rect 65800 116288 65852 116340
rect 120080 116288 120132 116340
rect 122104 116288 122156 116340
rect 210424 116288 210476 116340
rect 212356 116288 212408 116340
rect 204260 114724 204312 114776
rect 204996 114724 205048 114776
rect 13544 97928 13596 97980
rect 66260 97928 66312 97980
rect 97908 97928 97960 97980
rect 149060 97928 149112 97980
rect 154488 97928 154540 97980
rect 205640 97928 205692 97980
rect 209688 97928 209740 97980
rect 262220 97928 262272 97980
rect 266268 97928 266320 97980
rect 317420 97928 317472 97980
rect 322848 97928 322900 97980
rect 374000 97928 374052 97980
rect 405648 97928 405700 97980
rect 458180 97928 458232 97980
rect 489828 97928 489880 97980
rect 542360 97928 542412 97980
rect 70308 97860 70360 97912
rect 121460 97860 121512 97912
rect 126888 97860 126940 97912
rect 178040 97860 178092 97912
rect 182088 97860 182140 97912
rect 233240 97860 233292 97912
rect 238668 97860 238720 97912
rect 289820 97860 289872 97912
rect 293868 97860 293920 97912
rect 345020 97860 345072 97912
rect 378048 97860 378100 97912
rect 429292 97860 429344 97912
rect 434628 97860 434680 97912
rect 485780 97860 485832 97912
rect 518808 97860 518860 97912
rect 569960 97860 570012 97912
rect 42708 97792 42760 97844
rect 93860 97792 93912 97844
rect 350448 97792 350500 97844
rect 401600 97792 401652 97844
rect 462228 97792 462280 97844
rect 513380 97792 513432 97844
rect 547880 95412 547932 95464
rect 548340 95412 548392 95464
rect 15200 95140 15252 95192
rect 35900 95140 35952 95192
rect 36084 95140 36136 95192
rect 63592 95140 63644 95192
rect 65800 95140 65852 95192
rect 91928 95140 91980 95192
rect 92112 95140 92164 95192
rect 119620 95140 119672 95192
rect 122104 95140 122156 95192
rect 147956 95140 148008 95192
rect 148048 95140 148100 95192
rect 175924 95140 175976 95192
rect 176108 95140 176160 95192
rect 203616 95140 203668 95192
rect 204996 95140 205048 95192
rect 231952 95140 232004 95192
rect 232044 95140 232096 95192
rect 259920 95140 259972 95192
rect 260104 95140 260156 95192
rect 287612 95140 287664 95192
rect 288072 95140 288124 95192
rect 315948 95140 316000 95192
rect 316684 95140 316736 95192
rect 343916 95140 343968 95192
rect 344100 95140 344152 95192
rect 371608 95140 371660 95192
rect 372068 95140 372120 95192
rect 399944 95140 399996 95192
rect 400864 95140 400916 95192
rect 427912 95140 427964 95192
rect 428096 95140 428148 95192
rect 455604 95140 455656 95192
rect 456064 95140 456116 95192
rect 483940 95140 483992 95192
rect 484032 95140 484084 95192
rect 511908 95140 511960 95192
rect 512092 95140 512144 95192
rect 539600 95140 539652 95192
rect 540060 95140 540112 95192
rect 567936 95140 567988 95192
rect 16580 95072 16632 95124
rect 36636 95072 36688 95124
rect 44916 95072 44968 95124
rect 71136 95072 71188 95124
rect 82268 95072 82320 95124
rect 93124 95072 93176 95124
rect 110236 95072 110288 95124
rect 120724 95072 120776 95124
rect 128636 95072 128688 95124
rect 148324 95072 148376 95124
rect 156604 95072 156656 95124
rect 182824 95072 182876 95124
rect 194508 95072 194560 95124
rect 210424 95072 210476 95124
rect 212632 95072 212684 95124
rect 232504 95072 232556 95124
rect 240600 95072 240652 95124
rect 267004 95072 267056 95124
rect 278596 95072 278648 95124
rect 289084 95072 289136 95124
rect 306288 95072 306340 95124
rect 318064 95072 318116 95124
rect 324596 95072 324648 95124
rect 345664 95072 345716 95124
rect 362592 95072 362644 95124
rect 373264 95072 373316 95124
rect 390284 95072 390336 95124
rect 400956 95072 401008 95124
rect 408592 95072 408644 95124
rect 428464 95072 428516 95124
rect 436928 95072 436980 95124
rect 462964 95072 463016 95124
rect 474280 95072 474332 95124
rect 485044 95072 485096 95124
rect 502248 95072 502300 95124
rect 514024 95072 514076 95124
rect 520924 95072 520976 95124
rect 541624 95072 541676 95124
rect 26240 95004 26292 95056
rect 39304 95004 39356 95056
rect 54576 95004 54628 95056
rect 66904 95004 66956 95056
rect 138296 95004 138348 95056
rect 151084 95004 151136 95056
rect 166264 95004 166316 95056
rect 177304 95004 177356 95056
rect 222292 95004 222344 95056
rect 233976 95004 234028 95056
rect 250260 95004 250312 95056
rect 261484 95004 261536 95056
rect 334256 95004 334308 95056
rect 347044 95004 347096 95056
rect 418252 95004 418304 95056
rect 429844 95004 429896 95056
rect 446588 95004 446640 95056
rect 457444 95004 457496 95056
rect 530584 95004 530636 95056
rect 544384 95004 544436 95056
rect 558276 94460 558328 94512
rect 567476 94460 567528 94512
rect 408040 91264 408092 91316
rect 428648 91264 428700 91316
rect 148416 91196 148468 91248
rect 165712 91196 165764 91248
rect 175464 91196 175516 91248
rect 193680 91196 193732 91248
rect 203524 91196 203576 91248
rect 221372 91196 221424 91248
rect 232596 91196 232648 91248
rect 249708 91196 249760 91248
rect 260196 91196 260248 91248
rect 277676 91196 277728 91248
rect 287520 91196 287572 91248
rect 305368 91196 305420 91248
rect 315488 91196 315540 91248
rect 333704 91196 333756 91248
rect 345664 91196 345716 91248
rect 361672 91196 361724 91248
rect 371516 91196 371568 91248
rect 389364 91196 389416 91248
rect 399484 91196 399536 91248
rect 417700 91196 417752 91248
rect 456156 91196 456208 91248
rect 473360 91196 473412 91248
rect 483480 91196 483532 91248
rect 501696 91196 501748 91248
rect 511448 91196 511500 91248
rect 529664 91196 529716 91248
rect 36728 91128 36780 91180
rect 53656 91128 53708 91180
rect 64420 91128 64472 91180
rect 81440 91128 81492 91180
rect 91468 91128 91520 91180
rect 109684 91128 109736 91180
rect 119436 91128 119488 91180
rect 137652 91128 137704 91180
rect 156328 91128 156380 91180
rect 178684 91128 178736 91180
rect 212356 91128 212408 91180
rect 232688 91128 232740 91180
rect 268016 91128 268068 91180
rect 287704 91128 287756 91180
rect 296352 91128 296404 91180
rect 316776 91128 316828 91180
rect 352012 91128 352064 91180
rect 374644 91128 374696 91180
rect 428464 91128 428516 91180
rect 445668 91128 445720 91180
rect 464344 91128 464396 91180
rect 483664 91128 483716 91180
rect 492036 91128 492088 91180
rect 512736 91128 512788 91180
rect 541624 91128 541676 91180
rect 557540 91128 557592 91180
rect 15108 91060 15160 91112
rect 25688 91060 25740 91112
rect 36636 91060 36688 91112
rect 63316 91060 63368 91112
rect 66904 91060 66956 91112
rect 91100 91060 91152 91112
rect 93124 91060 93176 91112
rect 119344 91060 119396 91112
rect 124864 91060 124916 91112
rect 147312 91060 147364 91112
rect 148324 91060 148376 91112
rect 175372 91060 175424 91112
rect 177304 91060 177356 91112
rect 203340 91060 203392 91112
rect 204996 91060 205048 91112
rect 231032 91060 231084 91112
rect 232504 91060 232556 91112
rect 259368 91060 259420 91112
rect 260104 91060 260156 91112
rect 287336 91060 287388 91112
rect 289084 91060 289136 91112
rect 315028 91060 315080 91112
rect 316684 91060 316736 91112
rect 343364 91060 343416 91112
rect 344284 91060 344336 91112
rect 371332 91060 371384 91112
rect 373264 91060 373316 91112
rect 399024 91060 399076 91112
rect 400864 91060 400916 91112
rect 427360 91060 427412 91112
rect 428556 91060 428608 91112
rect 455328 91060 455380 91112
rect 456064 91060 456116 91112
rect 483020 91060 483072 91112
rect 485044 91060 485096 91112
rect 511356 91060 511408 91112
rect 512644 91060 512696 91112
rect 539324 91060 539376 91112
rect 540244 91060 540296 91112
rect 567200 91060 567252 91112
rect 434628 88816 434680 88868
rect 485780 88816 485832 88868
rect 405648 88748 405700 88800
rect 458180 88748 458232 88800
rect 42708 88340 42760 88392
rect 93860 88340 93912 88392
rect 97908 88340 97960 88392
rect 149060 88340 149112 88392
rect 154488 88340 154540 88392
rect 205640 88340 205692 88392
rect 209688 88340 209740 88392
rect 262220 88340 262272 88392
rect 266268 88340 266320 88392
rect 317420 88340 317472 88392
rect 322848 88340 322900 88392
rect 374000 88340 374052 88392
rect 378048 88340 378100 88392
rect 429292 88340 429344 88392
rect 489828 88340 489880 88392
rect 542360 88340 542412 88392
rect 42892 85892 42944 85944
rect 43628 85892 43680 85944
rect 3148 84192 3200 84244
rect 14556 84192 14608 84244
rect 428648 72428 428700 72480
rect 435732 72428 435784 72480
rect 63592 72292 63644 72344
rect 64420 72292 64472 72344
rect 147680 72292 147732 72344
rect 148416 72292 148468 72344
rect 232688 72292 232740 72344
rect 239772 72292 239824 72344
rect 259736 72292 259788 72344
rect 260196 72292 260248 72344
rect 316776 72292 316828 72344
rect 323676 72292 323728 72344
rect 455696 72292 455748 72344
rect 456156 72292 456208 72344
rect 483664 72224 483716 72276
rect 491668 72224 491720 72276
rect 287704 72088 287756 72140
rect 295708 72088 295760 72140
rect 512736 72088 512788 72140
rect 519636 72088 519688 72140
rect 13544 71680 13596 71732
rect 66260 71680 66312 71732
rect 70308 71680 70360 71732
rect 121460 71680 121512 71732
rect 126888 71680 126940 71732
rect 178040 71680 178092 71732
rect 182088 71680 182140 71732
rect 233240 71680 233292 71732
rect 238668 71680 238720 71732
rect 289820 71680 289872 71732
rect 293868 71680 293920 71732
rect 345020 71680 345072 71732
rect 350448 71680 350500 71732
rect 401600 71680 401652 71732
rect 462228 71680 462280 71732
rect 513380 71680 513432 71732
rect 518808 71680 518860 71732
rect 569960 71680 570012 71732
rect 231676 71612 231728 71664
rect 232596 71612 232648 71664
rect 343548 71612 343600 71664
rect 345664 71612 345716 71664
rect 539508 71612 539560 71664
rect 541624 71612 541676 71664
rect 15108 70660 15160 70712
rect 16580 70660 16632 70712
rect 35256 70660 35308 70712
rect 36728 70660 36780 70712
rect 547880 70660 547932 70712
rect 548156 70660 548208 70712
rect 71872 68960 71924 69012
rect 100024 68960 100076 69012
rect 25688 68892 25740 68944
rect 36636 68892 36688 68944
rect 42892 68892 42944 68944
rect 15292 68824 15344 68876
rect 43996 68824 44048 68876
rect 53656 68892 53708 68944
rect 66904 68892 66956 68944
rect 81992 68892 82044 68944
rect 93124 68892 93176 68944
rect 99472 68892 99524 68944
rect 127992 68960 128044 69012
rect 165988 68960 166040 69012
rect 177304 68960 177356 69012
rect 178684 68960 178736 69012
rect 184020 68960 184072 69012
rect 109684 68892 109736 68944
rect 124864 68892 124916 68944
rect 137652 68892 137704 68944
rect 148324 68892 148376 68944
rect 183652 68892 183704 68944
rect 211712 68960 211764 69012
rect 222016 68960 222068 69012
rect 232504 68960 232556 69012
rect 277676 68960 277728 69012
rect 289084 68960 289136 69012
rect 306012 68960 306064 69012
rect 316684 68960 316736 69012
rect 361672 68960 361724 69012
rect 373264 68960 373316 69012
rect 379612 68960 379664 69012
rect 408040 68960 408092 69012
rect 474004 68960 474056 69012
rect 485044 68960 485096 69012
rect 501696 68960 501748 69012
rect 512644 68960 512696 69012
rect 548156 68960 548208 69012
rect 557540 68960 557592 69012
rect 193680 68892 193732 68944
rect 204996 68892 205048 68944
rect 249708 68892 249760 68944
rect 260104 68892 260156 68944
rect 333704 68892 333756 68944
rect 344284 68892 344336 68944
rect 374644 68892 374696 68944
rect 379704 68892 379756 68944
rect 390008 68892 390060 68944
rect 400864 68892 400916 68944
rect 417700 68892 417752 68944
rect 428556 68892 428608 68944
rect 445668 68892 445720 68944
rect 456064 68892 456116 68944
rect 529664 68892 529716 68944
rect 540244 68892 540296 68944
rect 72056 68824 72108 68876
rect 127072 68824 127124 68876
rect 156052 68824 156104 68876
rect 238852 68824 238904 68876
rect 268016 68824 268068 68876
rect 323032 68824 323084 68876
rect 352012 68824 352064 68876
rect 434812 68824 434864 68876
rect 463700 68824 463752 68876
rect 518992 68824 519044 68876
rect 547880 68824 547932 68876
rect 26240 65288 26292 65340
rect 35440 65288 35492 65340
rect 71136 65016 71188 65068
rect 82268 65016 82320 65068
rect 99380 65016 99432 65068
rect 100300 65016 100352 65068
rect 183652 65016 183704 65068
rect 222292 65016 222344 65068
rect 261484 65016 261536 65068
rect 268292 65016 268344 65068
rect 295432 65016 295484 65068
rect 334256 65016 334308 65068
rect 352012 65016 352064 65068
rect 36636 64948 36688 65000
rect 53932 64948 53984 65000
rect 71872 64948 71924 65000
rect 109960 64948 110012 65000
rect 124864 64948 124916 65000
rect 128636 64948 128688 65000
rect 152464 64948 152516 65000
rect 156604 64948 156656 65000
rect 182824 64948 182876 65000
rect 193956 64948 194008 65000
rect 232504 64948 232556 65000
rect 39304 64880 39356 64932
rect 44272 64880 44324 64932
rect 66904 64880 66956 64932
rect 72608 64880 72660 64932
rect 93124 64880 93176 64932
rect 99380 64880 99432 64932
rect 99472 64880 99524 64932
rect 138296 64880 138348 64932
rect 151084 64880 151136 64932
rect 166264 64880 166316 64932
rect 177304 64880 177356 64932
rect 184296 64880 184348 64932
rect 210424 64880 210476 64932
rect 212632 64880 212684 64932
rect 233976 64880 234028 64932
rect 240600 64880 240652 64932
rect 267832 64948 267884 65000
rect 306288 64948 306340 65000
rect 345664 64948 345716 65000
rect 361948 64948 362000 65000
rect 379612 65016 379664 65068
rect 418252 65016 418304 65068
rect 463792 65016 463844 65068
rect 390284 64948 390336 65000
rect 400864 64948 400916 65000
rect 408592 64948 408644 65000
rect 429844 64948 429896 65000
rect 436284 64948 436336 65000
rect 457444 64948 457496 65000
rect 464620 64948 464672 65000
rect 485044 65016 485096 65068
rect 492588 65016 492640 65068
rect 502248 64948 502300 65000
rect 514024 64948 514076 65000
rect 520280 64948 520332 65000
rect 541624 64948 541676 65000
rect 558276 64948 558328 65000
rect 250260 64880 250312 64932
rect 267004 64880 267056 64932
rect 277952 64880 278004 64932
rect 289084 64880 289136 64932
rect 296628 64880 296680 64932
rect 318064 64880 318116 64932
rect 324596 64880 324648 64932
rect 347044 64880 347096 64932
rect 352288 64880 352340 64932
rect 373264 64880 373316 64932
rect 380624 64880 380676 64932
rect 428464 64880 428516 64932
rect 445944 64880 445996 64932
rect 462964 64880 463016 64932
rect 474280 64880 474332 64932
rect 491392 64880 491444 64932
rect 529940 64880 529992 64932
rect 547972 64880 548024 64932
rect 567936 64880 567988 64932
rect 63776 62296 63828 62348
rect 65800 62296 65852 62348
rect 120264 62160 120316 62212
rect 122104 62160 122156 62212
rect 42708 62092 42760 62144
rect 93860 62092 93912 62144
rect 97908 62092 97960 62144
rect 149060 62092 149112 62144
rect 154488 62092 154540 62144
rect 205640 62092 205692 62144
rect 209688 62092 209740 62144
rect 262220 62092 262272 62144
rect 266268 62092 266320 62144
rect 317420 62092 317472 62144
rect 322848 62092 322900 62144
rect 374000 62092 374052 62144
rect 378048 62092 378100 62144
rect 429292 62092 429344 62144
rect 434628 62092 434680 62144
rect 485780 62092 485832 62144
rect 489828 62092 489880 62144
rect 542360 62092 542412 62144
rect 544384 62092 544436 62144
rect 548340 62092 548392 62144
rect 400312 58692 400364 58744
rect 400956 58692 401008 58744
rect 204260 57876 204312 57928
rect 204996 57876 205048 57928
rect 2964 44140 3016 44192
rect 11888 44140 11940 44192
rect 13544 44072 13596 44124
rect 66260 44072 66312 44124
rect 70308 44072 70360 44124
rect 121460 44072 121512 44124
rect 126888 44072 126940 44124
rect 178040 44072 178092 44124
rect 182088 44072 182140 44124
rect 233240 44072 233292 44124
rect 238668 44072 238720 44124
rect 289820 44072 289872 44124
rect 293868 44072 293920 44124
rect 345020 44072 345072 44124
rect 350448 44072 350500 44124
rect 401600 44072 401652 44124
rect 405648 44072 405700 44124
rect 458180 44072 458232 44124
rect 462228 44072 462280 44124
rect 513380 44072 513432 44124
rect 518808 44072 518860 44124
rect 569960 44072 570012 44124
rect 15200 41352 15252 41404
rect 35900 41352 35952 41404
rect 36084 41352 36136 41404
rect 63592 41352 63644 41404
rect 65800 41352 65852 41404
rect 91928 41352 91980 41404
rect 92112 41352 92164 41404
rect 119620 41352 119672 41404
rect 122104 41352 122156 41404
rect 147956 41352 148008 41404
rect 148048 41352 148100 41404
rect 175924 41352 175976 41404
rect 176108 41352 176160 41404
rect 203616 41352 203668 41404
rect 204996 41352 205048 41404
rect 231952 41352 232004 41404
rect 232044 41352 232096 41404
rect 259920 41352 259972 41404
rect 260104 41352 260156 41404
rect 287612 41352 287664 41404
rect 288072 41352 288124 41404
rect 315948 41352 316000 41404
rect 316684 41352 316736 41404
rect 343916 41352 343968 41404
rect 344100 41352 344152 41404
rect 371608 41352 371660 41404
rect 372068 41352 372120 41404
rect 399944 41352 399996 41404
rect 400956 41352 401008 41404
rect 427912 41352 427964 41404
rect 428096 41352 428148 41404
rect 455604 41352 455656 41404
rect 456064 41352 456116 41404
rect 483940 41352 483992 41404
rect 484032 41352 484084 41404
rect 511908 41352 511960 41404
rect 512092 41352 512144 41404
rect 539600 41352 539652 41404
rect 540060 41352 540112 41404
rect 567936 41352 567988 41404
rect 16580 41284 16632 41336
rect 36636 41284 36688 41336
rect 44916 41284 44968 41336
rect 71136 41284 71188 41336
rect 82268 41284 82320 41336
rect 93124 41284 93176 41336
rect 110236 41284 110288 41336
rect 124864 41284 124916 41336
rect 128636 41284 128688 41336
rect 151084 41284 151136 41336
rect 156604 41284 156656 41336
rect 182824 41284 182876 41336
rect 194508 41284 194560 41336
rect 210424 41284 210476 41336
rect 212632 41284 212684 41336
rect 232504 41284 232556 41336
rect 240600 41284 240652 41336
rect 267004 41284 267056 41336
rect 278596 41284 278648 41336
rect 289084 41284 289136 41336
rect 306288 41284 306340 41336
rect 318064 41284 318116 41336
rect 324596 41284 324648 41336
rect 345664 41284 345716 41336
rect 362592 41284 362644 41336
rect 373264 41284 373316 41336
rect 390284 41284 390336 41336
rect 400864 41284 400916 41336
rect 408592 41284 408644 41336
rect 428464 41284 428516 41336
rect 436928 41284 436980 41336
rect 462964 41284 463016 41336
rect 474280 41284 474332 41336
rect 485044 41284 485096 41336
rect 502248 41284 502300 41336
rect 514024 41284 514076 41336
rect 520924 41284 520976 41336
rect 541624 41284 541676 41336
rect 26240 41216 26292 41268
rect 39304 41216 39356 41268
rect 54576 41216 54628 41268
rect 66904 41216 66956 41268
rect 138296 41216 138348 41268
rect 152464 41216 152516 41268
rect 166264 41216 166316 41268
rect 177304 41216 177356 41268
rect 222292 41216 222344 41268
rect 233976 41216 234028 41268
rect 250260 41216 250312 41268
rect 261484 41216 261536 41268
rect 334256 41216 334308 41268
rect 347044 41216 347096 41268
rect 418252 41216 418304 41268
rect 429844 41216 429896 41268
rect 446588 41216 446640 41268
rect 457444 41216 457496 41268
rect 530584 41216 530636 41268
rect 544384 41216 544436 41268
rect 558276 40672 558328 40724
rect 567476 40672 567528 40724
rect 46940 39380 46992 39432
rect 204904 39380 204956 39432
rect 19248 39312 19300 39364
rect 234620 39312 234672 39364
rect 547880 38496 547932 38548
rect 548340 38496 548392 38548
rect 26976 38428 27028 38480
rect 36544 38428 36596 38480
rect 53380 38428 53432 38480
rect 65708 38428 65760 38480
rect 5080 38360 5132 38412
rect 33416 38360 33468 38412
rect 35348 38360 35400 38412
rect 149704 38360 149756 38412
rect 5172 38292 5224 38344
rect 38568 38292 38620 38344
rect 43444 38292 43496 38344
rect 54668 38292 54720 38344
rect 59820 38292 59872 38344
rect 322204 38292 322256 38344
rect 14464 38224 14516 38276
rect 20536 38224 20588 38276
rect 23756 38224 23808 38276
rect 462320 38224 462372 38276
rect 11796 38156 11848 38208
rect 45008 38156 45060 38208
rect 61108 38156 61160 38208
rect 570696 38156 570748 38208
rect 10324 38088 10376 38140
rect 30196 38088 30248 38140
rect 32128 38088 32180 38140
rect 543004 38088 543056 38140
rect 4896 38020 4948 38072
rect 41788 38020 41840 38072
rect 51448 38020 51500 38072
rect 580908 38020 580960 38072
rect 6184 37952 6236 38004
rect 22468 37952 22520 38004
rect 25688 37952 25740 38004
rect 580448 37952 580500 38004
rect 16028 37884 16080 37936
rect 580724 37884 580776 37936
rect 57888 37816 57940 37868
rect 64236 37816 64288 37868
rect 50160 37408 50212 37460
rect 61384 37408 61436 37460
rect 149796 37408 149848 37460
rect 165712 37408 165764 37460
rect 175464 37408 175516 37460
rect 193680 37408 193732 37460
rect 203524 37408 203576 37460
rect 221372 37408 221424 37460
rect 232504 37408 232556 37460
rect 249708 37408 249760 37460
rect 260196 37408 260248 37460
rect 277676 37408 277728 37460
rect 287520 37408 287572 37460
rect 305368 37408 305420 37460
rect 345664 37408 345716 37460
rect 361672 37408 361724 37460
rect 371516 37408 371568 37460
rect 389364 37408 389416 37460
rect 399484 37408 399536 37460
rect 417700 37408 417752 37460
rect 456064 37408 456116 37460
rect 473360 37408 473412 37460
rect 483480 37408 483532 37460
rect 501696 37408 501748 37460
rect 42064 37340 42116 37392
rect 48228 37340 48280 37392
rect 56600 37340 56652 37392
rect 91100 37340 91152 37392
rect 91468 37340 91520 37392
rect 109684 37340 109736 37392
rect 122104 37340 122156 37392
rect 137652 37340 137704 37392
rect 156328 37340 156380 37392
rect 178684 37340 178736 37392
rect 212356 37340 212408 37392
rect 232596 37340 232648 37392
rect 268016 37340 268068 37392
rect 287704 37340 287756 37392
rect 296168 37340 296220 37392
rect 316776 37340 316828 37392
rect 322296 37340 322348 37392
rect 333704 37340 333756 37392
rect 352012 37340 352064 37392
rect 374644 37340 374696 37392
rect 408040 37340 408092 37392
rect 428556 37340 428608 37392
rect 429844 37340 429896 37392
rect 445668 37340 445720 37392
rect 464344 37340 464396 37392
rect 483664 37340 483716 37392
rect 492036 37340 492088 37392
rect 512736 37340 512788 37392
rect 518256 37340 518308 37392
rect 529664 37340 529716 37392
rect 541624 37340 541676 37392
rect 557540 37340 557592 37392
rect 13544 37272 13596 37324
rect 81440 37272 81492 37324
rect 93124 37272 93176 37324
rect 119344 37272 119396 37324
rect 120724 37272 120776 37324
rect 147312 37272 147364 37324
rect 148324 37272 148376 37324
rect 175372 37272 175424 37324
rect 177304 37272 177356 37324
rect 203340 37272 203392 37324
rect 204904 37272 204956 37324
rect 231032 37272 231084 37324
rect 239404 37272 239456 37324
rect 259368 37272 259420 37324
rect 260104 37272 260156 37324
rect 287336 37272 287388 37324
rect 289084 37272 289136 37324
rect 315028 37272 315080 37324
rect 316684 37272 316736 37324
rect 343364 37272 343416 37324
rect 344284 37272 344336 37324
rect 371332 37272 371384 37324
rect 373264 37272 373316 37324
rect 399024 37272 399076 37324
rect 400864 37272 400916 37324
rect 427360 37272 427412 37324
rect 428464 37272 428516 37324
rect 455328 37272 455380 37324
rect 456156 37272 456208 37324
rect 483020 37272 483072 37324
rect 485044 37272 485096 37324
rect 511356 37272 511408 37324
rect 512644 37272 512696 37324
rect 539324 37272 539376 37324
rect 540244 37272 540296 37324
rect 567200 37272 567252 37324
rect 64236 36728 64288 36780
rect 568028 36728 568080 36780
rect 64604 36660 64656 36712
rect 580172 36660 580224 36712
rect 64512 36592 64564 36644
rect 580264 36592 580316 36644
rect 13728 36524 13780 36576
rect 580632 36524 580684 36576
rect 39856 36048 39908 36100
rect 61476 36048 61528 36100
rect 36912 35980 36964 36032
rect 93860 35980 93912 36032
rect 28724 35912 28776 35964
rect 579988 35912 580040 35964
rect 3792 35164 3844 35216
rect 61292 35164 61344 35216
rect 63500 35164 63552 35216
rect 580356 35164 580408 35216
rect 266268 34620 266320 34672
rect 317420 34620 317472 34672
rect 434628 34620 434680 34672
rect 485780 34620 485832 34672
rect 70308 34552 70360 34604
rect 121460 34552 121512 34604
rect 126888 34552 126940 34604
rect 178040 34552 178092 34604
rect 182088 34552 182140 34604
rect 233240 34552 233292 34604
rect 238668 34552 238720 34604
rect 289820 34552 289872 34604
rect 322848 34552 322900 34604
rect 374000 34552 374052 34604
rect 378048 34552 378100 34604
rect 429292 34552 429344 34604
rect 462228 34552 462280 34604
rect 513380 34552 513432 34604
rect 518808 34552 518860 34604
rect 569960 34552 570012 34604
rect 97908 34484 97960 34536
rect 149060 34484 149112 34536
rect 154488 34484 154540 34536
rect 205640 34484 205692 34536
rect 209688 34484 209740 34536
rect 262220 34484 262272 34536
rect 293868 34484 293920 34536
rect 345020 34484 345072 34536
rect 350448 34484 350500 34536
rect 401600 34484 401652 34536
rect 405648 34484 405700 34536
rect 458180 34484 458232 34536
rect 489828 34484 489880 34536
rect 542360 34484 542412 34536
rect 3332 31696 3384 31748
rect 12440 31696 12492 31748
rect 238852 30744 238904 30796
rect 239772 30744 239824 30796
rect 63500 27548 63552 27600
rect 71044 27548 71096 27600
rect 4988 23400 5040 23452
rect 12440 23400 12492 23452
rect 4804 22040 4856 22092
rect 12440 22040 12492 22092
rect 259736 21428 259788 21480
rect 260196 21428 260248 21480
rect 9036 20612 9088 20664
rect 12624 20612 12676 20664
rect 428556 18572 428608 18624
rect 435732 18572 435784 18624
rect 287704 18232 287756 18284
rect 295708 18232 295760 18284
rect 316776 18096 316828 18148
rect 323676 18096 323728 18148
rect 232596 17960 232648 18012
rect 239772 17960 239824 18012
rect 483664 17960 483716 18012
rect 491668 17960 491720 18012
rect 512736 17960 512788 18012
rect 519636 17960 519688 18012
rect 7564 17892 7616 17944
rect 12440 17892 12492 17944
rect 3792 16532 3844 16584
rect 63500 16532 63552 16584
rect 119712 16532 119764 16584
rect 122104 16532 122156 16584
rect 147588 16532 147640 16584
rect 149796 16532 149848 16584
rect 343548 16532 343600 16584
rect 345664 16532 345716 16584
rect 427728 16532 427780 16584
rect 429844 16532 429896 16584
rect 539508 16532 539560 16584
rect 541624 16532 541676 16584
rect 41788 15104 41840 15156
rect 429200 15104 429252 15156
rect 52736 15036 52788 15088
rect 233884 15036 233936 15088
rect 39856 13744 39908 13796
rect 65616 13744 65668 13796
rect 81992 13744 82044 13796
rect 93124 13744 93176 13796
rect 165988 13744 166040 13796
rect 177304 13744 177356 13796
rect 178684 13744 178736 13796
rect 184020 13744 184072 13796
rect 193680 13744 193732 13796
rect 204904 13744 204956 13796
rect 249708 13744 249760 13796
rect 260104 13744 260156 13796
rect 277676 13744 277728 13796
rect 289084 13744 289136 13796
rect 306012 13744 306064 13796
rect 316684 13744 316736 13796
rect 361672 13744 361724 13796
rect 373264 13744 373316 13796
rect 374644 13744 374696 13796
rect 379704 13744 379756 13796
rect 390008 13744 390060 13796
rect 400864 13744 400916 13796
rect 474004 13744 474056 13796
rect 485044 13744 485096 13796
rect 501696 13744 501748 13796
rect 512644 13744 512696 13796
rect 529664 13744 529716 13796
rect 540244 13744 540296 13796
rect 547880 13744 547932 13796
rect 557540 13744 557592 13796
rect 17316 13676 17368 13728
rect 570604 13676 570656 13728
rect 3424 13608 3476 13660
rect 28908 13608 28960 13660
rect 32128 13608 32180 13660
rect 580080 13608 580132 13660
rect 4068 13540 4120 13592
rect 25688 13540 25740 13592
rect 36636 13540 36688 13592
rect 580540 13540 580592 13592
rect 8944 13472 8996 13524
rect 30196 13472 30248 13524
rect 43076 13472 43128 13524
rect 580816 13472 580868 13524
rect 26976 13404 27028 13456
rect 378784 13404 378836 13456
rect 379612 13404 379664 13456
rect 408040 13404 408092 13456
rect 417700 13404 417752 13456
rect 428464 13404 428516 13456
rect 434812 13404 434864 13456
rect 463700 13404 463752 13456
rect 511356 13404 511408 13456
rect 518256 13404 518308 13456
rect 518992 13404 519044 13456
rect 547972 13404 548024 13456
rect 3608 13336 3660 13388
rect 57888 13336 57940 13388
rect 71872 13336 71924 13388
rect 100024 13336 100076 13388
rect 3700 13268 3752 13320
rect 54668 13268 54720 13320
rect 99472 13268 99524 13320
rect 127992 13336 128044 13388
rect 109684 13268 109736 13320
rect 120724 13268 120776 13320
rect 127072 13268 127124 13320
rect 156052 13336 156104 13388
rect 183652 13336 183704 13388
rect 211712 13336 211764 13388
rect 222016 13336 222068 13388
rect 239404 13336 239456 13388
rect 315672 13336 315724 13388
rect 322296 13336 322348 13388
rect 323032 13336 323084 13388
rect 352012 13336 352064 13388
rect 445668 13336 445720 13388
rect 456156 13336 456208 13388
rect 137652 13268 137704 13320
rect 148324 13268 148376 13320
rect 333704 13268 333756 13320
rect 344284 13268 344336 13320
rect 6920 13200 6972 13252
rect 55956 13200 56008 13252
rect 238852 13200 238904 13252
rect 268016 13200 268068 13252
rect 3976 13132 4028 13184
rect 22468 13132 22520 13184
rect 23756 13132 23808 13184
rect 65524 13132 65576 13184
rect 1400 13064 1452 13116
rect 33416 13064 33468 13116
rect 38568 13064 38620 13116
rect 72056 13064 72108 13116
rect 20536 12996 20588 13048
rect 578884 12996 578936 13048
rect 3516 12928 3568 12980
rect 46296 12928 46348 12980
rect 3884 12860 3936 12912
rect 51448 12860 51500 12912
rect 11704 12792 11756 12844
rect 35348 12792 35400 12844
rect 64420 3680 64472 3732
rect 125876 3680 125928 3732
rect 64236 3612 64288 3664
rect 126980 3612 127032 3664
rect 61384 3544 61436 3596
rect 132960 3544 133012 3596
rect 13728 3476 13780 3528
rect 129372 3476 129424 3528
rect 572 3408 624 3460
rect 48320 3408 48372 3460
rect 61476 3408 61528 3460
rect 136456 3408 136508 3460
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 2778 658200 2834 658209
rect 2778 658135 2834 658144
rect 2792 657558 2820 658135
rect 2780 657552 2832 657558
rect 2780 657494 2832 657500
rect 6184 657552 6236 657558
rect 6184 657494 6236 657500
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 2778 527912 2834 527921
rect 2778 527847 2834 527856
rect 2792 527202 2820 527847
rect 2780 527196 2832 527202
rect 2780 527138 2832 527144
rect 2778 449576 2834 449585
rect 2778 449511 2834 449520
rect 2792 448662 2820 449511
rect 2780 448656 2832 448662
rect 2780 448598 2832 448604
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 410378 3188 410479
rect 3148 410372 3200 410378
rect 3148 410314 3200 410320
rect 2778 345400 2834 345409
rect 2778 345335 2834 345344
rect 2792 345234 2820 345335
rect 2780 345228 2832 345234
rect 2780 345170 2832 345176
rect 3330 293176 3386 293185
rect 3330 293111 3332 293120
rect 3384 293111 3386 293120
rect 3332 293082 3384 293088
rect 2778 254144 2834 254153
rect 2778 254079 2780 254088
rect 2832 254079 2834 254088
rect 2780 254050 2832 254056
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 2792 240242 2820 241023
rect 2780 240236 2832 240242
rect 2780 240178 2832 240184
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3068 201550 3096 201855
rect 3056 201544 3108 201550
rect 3056 201486 3108 201492
rect 2962 188864 3018 188873
rect 2962 188799 3018 188808
rect 2976 187746 3004 188799
rect 2964 187740 3016 187746
rect 2964 187682 3016 187688
rect 3330 136776 3386 136785
rect 3330 136711 3332 136720
rect 3384 136711 3386 136720
rect 3332 136682 3384 136688
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3160 84250 3188 84623
rect 3148 84244 3200 84250
rect 3148 84186 3200 84192
rect 3330 58576 3386 58585
rect 3330 58511 3386 58520
rect 2962 45520 3018 45529
rect 2962 45455 3018 45464
rect 2976 44198 3004 45455
rect 2964 44192 3016 44198
rect 2964 44134 3016 44140
rect 3344 31754 3372 58511
rect 3332 31748 3384 31754
rect 3332 31690 3384 31696
rect 3436 13666 3464 579935
rect 4804 527196 4856 527202
rect 4804 527138 4856 527144
rect 3514 501800 3570 501809
rect 3514 501735 3570 501744
rect 3424 13660 3476 13666
rect 3424 13602 3476 13608
rect 1400 13116 1452 13122
rect 1400 13058 1452 13064
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 542 -960 654 480
rect 1412 354 1440 13058
rect 3528 12986 3556 501735
rect 3606 475688 3662 475697
rect 3606 475623 3662 475632
rect 3620 13394 3648 475623
rect 3698 397488 3754 397497
rect 3698 397423 3754 397432
rect 3608 13388 3660 13394
rect 3608 13330 3660 13336
rect 3712 13326 3740 397423
rect 3790 358456 3846 358465
rect 3790 358391 3846 358400
rect 3804 35222 3832 358391
rect 3882 306232 3938 306241
rect 3882 306167 3938 306176
rect 3792 35216 3844 35222
rect 3792 35158 3844 35164
rect 3790 19408 3846 19417
rect 3790 19343 3846 19352
rect 3804 16590 3832 19343
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3700 13320 3752 13326
rect 3700 13262 3752 13268
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3896 12918 3924 306167
rect 3974 149832 4030 149841
rect 3974 149767 4030 149776
rect 3988 13190 4016 149767
rect 4066 97608 4122 97617
rect 4066 97543 4122 97552
rect 4080 13598 4108 97543
rect 4816 22098 4844 527138
rect 4896 448656 4948 448662
rect 4896 448598 4948 448604
rect 4908 38078 4936 448598
rect 4988 345228 5040 345234
rect 4988 345170 5040 345176
rect 4896 38072 4948 38078
rect 4896 38014 4948 38020
rect 5000 23458 5028 345170
rect 5080 254108 5132 254114
rect 5080 254050 5132 254056
rect 5092 38418 5120 254050
rect 5172 240236 5224 240242
rect 5172 240178 5224 240184
rect 5080 38412 5132 38418
rect 5080 38354 5132 38360
rect 5184 38350 5212 240178
rect 5172 38344 5224 38350
rect 5172 38286 5224 38292
rect 6196 38010 6224 657494
rect 6184 38004 6236 38010
rect 6184 37946 6236 37952
rect 4988 23452 5040 23458
rect 4988 23394 5040 23400
rect 4804 22092 4856 22098
rect 4804 22034 4856 22040
rect 4068 13592 4120 13598
rect 4068 13534 4120 13540
rect 6932 13258 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 36544 700664 36596 700670
rect 36544 700606 36596 700612
rect 13452 700528 13504 700534
rect 13452 700470 13504 700476
rect 11704 605872 11756 605878
rect 11704 605814 11756 605820
rect 10324 553444 10376 553450
rect 10324 553386 10376 553392
rect 8944 410372 8996 410378
rect 8944 410314 8996 410320
rect 7564 293140 7616 293146
rect 7564 293082 7616 293088
rect 7576 17950 7604 293082
rect 7564 17944 7616 17950
rect 7564 17886 7616 17892
rect 8956 13530 8984 410314
rect 9036 136740 9088 136746
rect 9036 136682 9088 136688
rect 9048 20670 9076 136682
rect 10336 38146 10364 553386
rect 10324 38140 10376 38146
rect 10324 38082 10376 38088
rect 9036 20664 9088 20670
rect 9036 20606 9088 20612
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3884 12912 3936 12918
rect 3884 12854 3936 12860
rect 11716 12850 11744 605814
rect 11796 187740 11848 187746
rect 11796 187682 11848 187688
rect 11808 38214 11836 187682
rect 11888 44192 11940 44198
rect 11888 44134 11940 44140
rect 11796 38208 11848 38214
rect 11796 38150 11848 38156
rect 11900 34513 11928 44134
rect 11886 34504 11942 34513
rect 11886 34439 11942 34448
rect 13464 33153 13492 700470
rect 16120 685908 16172 685914
rect 16120 685850 16172 685856
rect 25688 685908 25740 685914
rect 25688 685850 25740 685856
rect 15304 683590 16054 683618
rect 13634 674248 13690 674257
rect 13634 674183 13690 674192
rect 13648 665174 13676 674183
rect 13636 665168 13688 665174
rect 13636 665110 13688 665116
rect 15304 662250 15332 683590
rect 16132 683330 16160 685850
rect 25700 683876 25728 685850
rect 15844 683324 15896 683330
rect 15844 683266 15896 683272
rect 16120 683324 16172 683330
rect 35374 683318 35480 683346
rect 16120 683266 16172 683272
rect 15856 664154 15884 683266
rect 35256 664760 35308 664766
rect 35308 664708 35374 664714
rect 35256 664702 35374 664708
rect 35268 664686 35374 664702
rect 15844 664148 15896 664154
rect 15844 664090 15896 664096
rect 16580 664148 16632 664154
rect 16580 664090 16632 664096
rect 15488 664006 16054 664034
rect 15292 662244 15344 662250
rect 15292 662186 15344 662192
rect 13636 661700 13688 661706
rect 13636 661642 13688 661648
rect 13542 620256 13598 620265
rect 13542 620191 13598 620200
rect 13556 611318 13584 620191
rect 13544 611312 13596 611318
rect 13544 611254 13596 611260
rect 13544 601724 13596 601730
rect 13544 601666 13596 601672
rect 13556 593473 13584 601666
rect 13542 593464 13598 593473
rect 13542 593399 13598 593408
rect 13542 566264 13598 566273
rect 13542 566199 13598 566208
rect 13556 557530 13584 566199
rect 13544 557524 13596 557530
rect 13544 557466 13596 557472
rect 13542 539472 13598 539481
rect 13542 539407 13598 539416
rect 13556 529922 13584 539407
rect 13544 529916 13596 529922
rect 13544 529858 13596 529864
rect 13542 512272 13598 512281
rect 13542 512207 13598 512216
rect 13556 503674 13584 512207
rect 13544 503668 13596 503674
rect 13544 503610 13596 503616
rect 13542 485480 13598 485489
rect 13542 485415 13598 485424
rect 13556 476066 13584 485415
rect 13544 476060 13596 476066
rect 13544 476002 13596 476008
rect 13544 466472 13596 466478
rect 13544 466414 13596 466420
rect 13556 458289 13584 466414
rect 13542 458280 13598 458289
rect 13542 458215 13598 458224
rect 13542 431488 13598 431497
rect 13542 431423 13598 431432
rect 13556 422278 13584 431423
rect 13544 422272 13596 422278
rect 13544 422214 13596 422220
rect 13542 404288 13598 404297
rect 13542 404223 13598 404232
rect 13556 394670 13584 404223
rect 13544 394664 13596 394670
rect 13544 394606 13596 394612
rect 13544 386436 13596 386442
rect 13544 386378 13596 386384
rect 13556 377505 13584 386378
rect 13542 377496 13598 377505
rect 13542 377431 13598 377440
rect 13542 350296 13598 350305
rect 13542 350231 13598 350240
rect 13556 340882 13584 350231
rect 13544 340876 13596 340882
rect 13544 340818 13596 340824
rect 13542 322960 13598 322969
rect 13542 322895 13598 322904
rect 13556 314634 13584 322895
rect 13544 314628 13596 314634
rect 13544 314570 13596 314576
rect 13542 296304 13598 296313
rect 13542 296239 13598 296248
rect 13556 287026 13584 296239
rect 13544 287020 13596 287026
rect 13544 286962 13596 286968
rect 13544 277432 13596 277438
rect 13544 277374 13596 277380
rect 13556 270065 13584 277374
rect 13542 270056 13598 270065
rect 13542 269991 13598 270000
rect 13542 242312 13598 242321
rect 13542 242247 13598 242256
rect 13556 233238 13584 242247
rect 13544 233232 13596 233238
rect 13544 233174 13596 233180
rect 13544 223644 13596 223650
rect 13544 223586 13596 223592
rect 13556 215393 13584 223586
rect 13542 215384 13598 215393
rect 13542 215319 13598 215328
rect 13542 188320 13598 188329
rect 13542 188255 13598 188264
rect 13556 179382 13584 188255
rect 13544 179376 13596 179382
rect 13544 179318 13596 179324
rect 13542 161392 13598 161401
rect 13542 161327 13598 161336
rect 13556 151774 13584 161327
rect 13544 151768 13596 151774
rect 13544 151710 13596 151716
rect 13542 134328 13598 134337
rect 13542 134263 13598 134272
rect 13556 125594 13584 134263
rect 13544 125588 13596 125594
rect 13544 125530 13596 125536
rect 13542 107400 13598 107409
rect 13542 107335 13598 107344
rect 13556 97986 13584 107335
rect 13544 97980 13596 97986
rect 13544 97922 13596 97928
rect 13542 80336 13598 80345
rect 13542 80271 13598 80280
rect 13556 71738 13584 80271
rect 13544 71732 13596 71738
rect 13544 71674 13596 71680
rect 13542 53408 13598 53417
rect 13542 53343 13598 53352
rect 13556 44130 13584 53343
rect 13544 44124 13596 44130
rect 13544 44066 13596 44072
rect 13544 37324 13596 37330
rect 13544 37266 13596 37272
rect 13450 33144 13506 33153
rect 13450 33079 13506 33088
rect 12440 31748 12492 31754
rect 12440 31690 12492 31696
rect 12452 31113 12480 31690
rect 12438 31104 12494 31113
rect 12438 31039 12494 31048
rect 13556 26353 13584 37266
rect 13648 27713 13676 661642
rect 13728 655580 13780 655586
rect 13728 655522 13780 655528
rect 13740 647465 13768 655522
rect 13726 647456 13782 647465
rect 13726 647391 13782 647400
rect 15488 644474 15516 664006
rect 16592 656948 16620 664090
rect 25700 662318 25728 664020
rect 25688 662312 25740 662318
rect 25688 662254 25740 662260
rect 35452 658374 35480 683318
rect 26240 658368 26292 658374
rect 26240 658310 26292 658316
rect 35440 658368 35492 658374
rect 35440 658310 35492 658316
rect 26252 656948 26280 658310
rect 35926 656254 36124 656282
rect 15212 644446 15516 644474
rect 15212 634778 15240 644446
rect 15200 634772 15252 634778
rect 15200 634714 15252 634720
rect 16592 634710 16620 637092
rect 16580 634704 16632 634710
rect 16580 634646 16632 634652
rect 26252 634642 26280 637092
rect 35912 634778 35940 637092
rect 36096 634778 36124 656254
rect 35900 634772 35952 634778
rect 35900 634714 35952 634720
rect 36084 634772 36136 634778
rect 36084 634714 36136 634720
rect 26240 634636 26292 634642
rect 26240 634578 26292 634584
rect 14464 632120 14516 632126
rect 14464 632062 14516 632068
rect 16120 632120 16172 632126
rect 16120 632062 16172 632068
rect 25688 632120 25740 632126
rect 25688 632062 25740 632068
rect 14476 38282 14504 632062
rect 15304 629598 16054 629626
rect 15304 608462 15332 629598
rect 16132 629338 16160 632062
rect 25700 629884 25728 632062
rect 15844 629332 15896 629338
rect 15844 629274 15896 629280
rect 16120 629332 16172 629338
rect 35374 629326 35480 629354
rect 16120 629274 16172 629280
rect 15856 610706 15884 629274
rect 35268 610706 35374 610722
rect 15844 610700 15896 610706
rect 15844 610642 15896 610648
rect 16580 610700 16632 610706
rect 16580 610642 16632 610648
rect 35256 610700 35374 610706
rect 35308 610694 35374 610700
rect 35256 610642 35308 610648
rect 15488 610014 16054 610042
rect 15292 608456 15344 608462
rect 15292 608398 15344 608404
rect 15488 605834 15516 610014
rect 15212 605806 15516 605834
rect 15212 580990 15240 605806
rect 16592 602956 16620 610642
rect 25700 608530 25728 610028
rect 25688 608524 25740 608530
rect 25688 608466 25740 608472
rect 35452 604518 35480 629326
rect 26240 604512 26292 604518
rect 26240 604454 26292 604460
rect 35440 604512 35492 604518
rect 35440 604454 35492 604460
rect 26252 602956 26280 604454
rect 35926 602262 36124 602290
rect 15200 580984 15252 580990
rect 15200 580926 15252 580932
rect 16592 580922 16620 583100
rect 16580 580916 16632 580922
rect 16580 580858 16632 580864
rect 26252 580854 26280 583100
rect 35912 580990 35940 583100
rect 36096 580990 36124 602262
rect 35900 580984 35952 580990
rect 35900 580926 35952 580932
rect 36084 580984 36136 580990
rect 36084 580926 36136 580932
rect 26240 580848 26292 580854
rect 26240 580790 26292 580796
rect 15844 578264 15896 578270
rect 15844 578206 15896 578212
rect 25688 578264 25740 578270
rect 25688 578206 25740 578212
rect 15292 575272 15344 575278
rect 15292 575214 15344 575220
rect 15304 554606 15332 575214
rect 15856 556238 15884 578206
rect 25700 575892 25728 578206
rect 15948 575334 16054 575362
rect 35374 575334 35480 575362
rect 15948 575278 15976 575334
rect 15936 575272 15988 575278
rect 15936 575214 15988 575220
rect 35268 556714 35374 556730
rect 35256 556708 35374 556714
rect 35308 556702 35374 556708
rect 35256 556650 35308 556656
rect 15844 556232 15896 556238
rect 15844 556174 15896 556180
rect 16580 556232 16632 556238
rect 16580 556174 16632 556180
rect 15488 556022 16054 556050
rect 15292 554600 15344 554606
rect 15292 554542 15344 554548
rect 15488 547874 15516 556022
rect 16592 548964 16620 556174
rect 25700 554674 25728 556036
rect 25688 554668 25740 554674
rect 25688 554610 25740 554616
rect 35452 550934 35480 575334
rect 26240 550928 26292 550934
rect 26240 550870 26292 550876
rect 35440 550928 35492 550934
rect 35440 550870 35492 550876
rect 26252 548964 26280 550870
rect 35926 548270 36124 548298
rect 15212 547846 15516 547874
rect 15212 527134 15240 547846
rect 15200 527128 15252 527134
rect 15200 527070 15252 527076
rect 16592 527066 16620 529108
rect 16580 527060 16632 527066
rect 16580 527002 16632 527008
rect 26252 526998 26280 529108
rect 35912 527134 35940 529108
rect 36096 527134 36124 548270
rect 35900 527128 35952 527134
rect 35900 527070 35952 527076
rect 36084 527128 36136 527134
rect 36084 527070 36136 527076
rect 26240 526992 26292 526998
rect 26240 526934 26292 526940
rect 15108 523048 15160 523054
rect 15108 522990 15160 522996
rect 25688 523048 25740 523054
rect 25688 522990 25740 522996
rect 15120 502722 15148 522990
rect 25700 521900 25728 522990
rect 15304 521206 16054 521234
rect 35374 521206 35480 521234
rect 15108 502716 15160 502722
rect 15108 502658 15160 502664
rect 15304 500818 15332 521206
rect 16580 502716 16632 502722
rect 16580 502658 16632 502664
rect 15488 502030 16054 502058
rect 15292 500812 15344 500818
rect 15292 500754 15344 500760
rect 15488 489914 15516 502030
rect 16592 494972 16620 502658
rect 35268 502314 35374 502330
rect 35256 502308 35374 502314
rect 35308 502302 35374 502308
rect 35256 502250 35308 502256
rect 25700 500886 25728 502044
rect 25688 500880 25740 500886
rect 25688 500822 25740 500828
rect 35452 496942 35480 521206
rect 26240 496936 26292 496942
rect 26240 496878 26292 496884
rect 35440 496936 35492 496942
rect 35440 496878 35492 496884
rect 26252 494972 26280 496878
rect 35926 494278 36124 494306
rect 15212 489886 15516 489914
rect 15212 473346 15240 489886
rect 15200 473340 15252 473346
rect 15200 473282 15252 473288
rect 16592 473278 16620 475116
rect 16580 473272 16632 473278
rect 16580 473214 16632 473220
rect 26252 473210 26280 475116
rect 35912 473346 35940 475116
rect 36096 473346 36124 494278
rect 35900 473340 35952 473346
rect 35900 473282 35952 473288
rect 36084 473340 36136 473346
rect 36084 473282 36136 473288
rect 26240 473204 26292 473210
rect 26240 473146 26292 473152
rect 15660 469260 15712 469266
rect 15660 469202 15712 469208
rect 25688 469260 25740 469266
rect 25688 469202 25740 469208
rect 15292 467288 15344 467294
rect 15292 467230 15344 467236
rect 15304 445602 15332 467230
rect 15672 460934 15700 469202
rect 25700 467908 25728 469202
rect 15936 467288 15988 467294
rect 15988 467236 16054 467242
rect 15936 467230 16054 467236
rect 15948 467214 16054 467230
rect 35374 467214 35480 467242
rect 15672 460906 15884 460934
rect 15856 448730 15884 460906
rect 15844 448724 15896 448730
rect 15844 448666 15896 448672
rect 16672 448724 16724 448730
rect 16672 448666 16724 448672
rect 15672 448038 16054 448066
rect 15292 445596 15344 445602
rect 15292 445538 15344 445544
rect 15672 431954 15700 448038
rect 16684 441614 16712 448666
rect 35256 448520 35308 448526
rect 35308 448468 35374 448474
rect 35256 448462 35374 448468
rect 35268 448446 35374 448462
rect 25700 445670 25728 448052
rect 25688 445664 25740 445670
rect 25688 445606 25740 445612
rect 35452 443426 35480 467214
rect 26608 443420 26660 443426
rect 26608 443362 26660 443368
rect 35440 443420 35492 443426
rect 35440 443362 35492 443368
rect 16684 441586 16804 441614
rect 16776 440858 16804 441586
rect 26620 440994 26648 443362
rect 26266 440966 26648 440994
rect 16606 440830 16804 440858
rect 35926 440286 36124 440314
rect 15212 431926 15700 431954
rect 15212 419490 15240 431926
rect 15200 419484 15252 419490
rect 15200 419426 15252 419432
rect 16592 419422 16620 421124
rect 16580 419416 16632 419422
rect 16580 419358 16632 419364
rect 26252 419354 26280 421124
rect 35912 419490 35940 421124
rect 36096 419490 36124 440286
rect 35900 419484 35952 419490
rect 35900 419426 35952 419432
rect 36084 419484 36136 419490
rect 36084 419426 36136 419432
rect 26240 419348 26292 419354
rect 26240 419290 26292 419296
rect 15108 415472 15160 415478
rect 15108 415414 15160 415420
rect 25688 415472 25740 415478
rect 25688 415414 25740 415420
rect 15120 390454 15148 415414
rect 25700 413916 25728 415414
rect 15304 413222 16054 413250
rect 35374 413222 35480 413250
rect 15304 391814 15332 413222
rect 35268 394602 35374 394618
rect 35256 394596 35374 394602
rect 35308 394590 35374 394596
rect 35256 394538 35308 394544
rect 15672 394046 16054 394074
rect 15292 391808 15344 391814
rect 15292 391750 15344 391756
rect 15108 390448 15160 390454
rect 15108 390390 15160 390396
rect 15672 373994 15700 394046
rect 25700 391882 25728 394060
rect 25688 391876 25740 391882
rect 25688 391818 25740 391824
rect 16580 390448 16632 390454
rect 16580 390390 16632 390396
rect 16592 386852 16620 390390
rect 35452 389842 35480 413222
rect 26240 389836 26292 389842
rect 26240 389778 26292 389784
rect 35440 389836 35492 389842
rect 35440 389778 35492 389784
rect 26252 386852 26280 389778
rect 35926 386294 36124 386322
rect 15212 373966 15700 373994
rect 15212 365702 15240 373966
rect 15200 365696 15252 365702
rect 15200 365638 15252 365644
rect 16592 365634 16620 367132
rect 16580 365628 16632 365634
rect 16580 365570 16632 365576
rect 26252 365566 26280 367132
rect 35912 365702 35940 367132
rect 36096 365702 36124 386294
rect 35900 365696 35952 365702
rect 35900 365638 35952 365644
rect 36084 365696 36136 365702
rect 36084 365638 36136 365644
rect 26240 365560 26292 365566
rect 26240 365502 26292 365508
rect 15108 361616 15160 361622
rect 15108 361558 15160 361564
rect 25688 361616 25740 361622
rect 25688 361558 25740 361564
rect 15120 335374 15148 361558
rect 25700 359924 25728 361558
rect 15304 359230 16054 359258
rect 35374 359230 35480 359258
rect 15304 337958 15332 359230
rect 35268 340746 35374 340762
rect 35256 340740 35374 340746
rect 35308 340734 35374 340740
rect 35256 340682 35308 340688
rect 15488 340054 16054 340082
rect 15292 337952 15344 337958
rect 15292 337894 15344 337900
rect 15108 335368 15160 335374
rect 15488 335354 15516 340054
rect 25700 338026 25728 340068
rect 25688 338020 25740 338026
rect 25688 337962 25740 337968
rect 35452 335782 35480 359230
rect 26240 335776 26292 335782
rect 26240 335718 26292 335724
rect 35440 335776 35492 335782
rect 35440 335718 35492 335724
rect 15108 335310 15160 335316
rect 15212 335326 15516 335354
rect 16580 335368 16632 335374
rect 15212 311846 15240 335326
rect 16580 335310 16632 335316
rect 16592 332860 16620 335310
rect 26252 332860 26280 335718
rect 35926 332302 36124 332330
rect 15200 311840 15252 311846
rect 15200 311782 15252 311788
rect 16592 311778 16620 313140
rect 16580 311772 16632 311778
rect 16580 311714 16632 311720
rect 26252 311710 26280 313140
rect 35912 311846 35940 313140
rect 36096 311846 36124 332302
rect 35900 311840 35952 311846
rect 35900 311782 35952 311788
rect 36084 311840 36136 311846
rect 36084 311782 36136 311788
rect 26240 311704 26292 311710
rect 26240 311646 26292 311652
rect 15108 307828 15160 307834
rect 15108 307770 15160 307776
rect 25688 307828 25740 307834
rect 25688 307770 25740 307776
rect 15120 285734 15148 307770
rect 25700 305932 25728 307770
rect 15304 305238 16054 305266
rect 35374 305238 35480 305266
rect 15108 285728 15160 285734
rect 15108 285670 15160 285676
rect 15304 284170 15332 305238
rect 35268 286754 35374 286770
rect 35256 286748 35374 286754
rect 35308 286742 35374 286748
rect 35256 286690 35308 286696
rect 15672 286062 16054 286090
rect 15292 284164 15344 284170
rect 15292 284106 15344 284112
rect 15672 277394 15700 286062
rect 16580 285728 16632 285734
rect 16580 285670 16632 285676
rect 16592 278868 16620 285670
rect 25700 284238 25728 286076
rect 25688 284232 25740 284238
rect 25688 284174 25740 284180
rect 35452 280430 35480 305238
rect 26240 280424 26292 280430
rect 26240 280366 26292 280372
rect 35440 280424 35492 280430
rect 35440 280366 35492 280372
rect 26252 278868 26280 280366
rect 35926 278310 36124 278338
rect 15212 277366 15700 277394
rect 15212 256698 15240 277366
rect 15200 256692 15252 256698
rect 15200 256634 15252 256640
rect 16592 256630 16620 259148
rect 16580 256624 16632 256630
rect 16580 256566 16632 256572
rect 26252 256562 26280 259148
rect 35912 256698 35940 259148
rect 36096 256698 36124 278310
rect 35900 256692 35952 256698
rect 35900 256634 35952 256640
rect 36084 256692 36136 256698
rect 36084 256634 36136 256640
rect 26240 256556 26292 256562
rect 26240 256498 26292 256504
rect 15108 253972 15160 253978
rect 15108 253914 15160 253920
rect 25688 253972 25740 253978
rect 25688 253914 25740 253920
rect 15120 232762 15148 253914
rect 25700 251940 25728 253914
rect 15304 251246 16054 251274
rect 35374 251246 35480 251274
rect 15108 232756 15160 232762
rect 15108 232698 15160 232704
rect 15304 230314 15332 251246
rect 16580 232756 16632 232762
rect 16580 232698 16632 232704
rect 15672 232070 16054 232098
rect 15292 230308 15344 230314
rect 15292 230250 15344 230256
rect 15672 219434 15700 232070
rect 16592 224876 16620 232698
rect 25700 230382 25728 232084
rect 35360 231946 35388 232084
rect 35348 231940 35400 231946
rect 35348 231882 35400 231888
rect 25688 230376 25740 230382
rect 25688 230318 25740 230324
rect 35452 226506 35480 251246
rect 26240 226500 26292 226506
rect 26240 226442 26292 226448
rect 35440 226500 35492 226506
rect 35440 226442 35492 226448
rect 26252 224876 26280 226442
rect 35926 224318 36124 224346
rect 15212 219406 15700 219434
rect 15212 202842 15240 219406
rect 16606 205006 16896 205034
rect 26266 205006 26648 205034
rect 15200 202836 15252 202842
rect 15200 202778 15252 202784
rect 16868 202774 16896 205006
rect 16856 202768 16908 202774
rect 16856 202710 16908 202716
rect 26620 202706 26648 205006
rect 35820 205006 35926 205034
rect 35820 204898 35848 205006
rect 35820 204870 35940 204898
rect 35912 202842 35940 204870
rect 36096 202842 36124 224318
rect 35900 202836 35952 202842
rect 35900 202778 35952 202784
rect 36084 202836 36136 202842
rect 36084 202778 36136 202784
rect 26608 202700 26660 202706
rect 26608 202642 26660 202648
rect 15108 200184 15160 200190
rect 15108 200126 15160 200132
rect 25688 200184 25740 200190
rect 25688 200126 25740 200132
rect 15120 178770 15148 200126
rect 25700 197948 25728 200126
rect 15304 197254 16054 197282
rect 35374 197254 35480 197282
rect 15108 178764 15160 178770
rect 15108 178706 15160 178712
rect 15304 176526 15332 197254
rect 16580 178764 16632 178770
rect 16580 178706 16632 178712
rect 35256 178764 35308 178770
rect 35256 178706 35308 178712
rect 15488 178078 16054 178106
rect 15292 176520 15344 176526
rect 15292 176462 15344 176468
rect 15488 161474 15516 178078
rect 16592 170884 16620 178706
rect 35268 178650 35296 178706
rect 35268 178622 35374 178650
rect 25700 176594 25728 178092
rect 25688 176588 25740 176594
rect 25688 176530 25740 176536
rect 35452 172854 35480 197254
rect 26240 172848 26292 172854
rect 26240 172790 26292 172796
rect 35440 172848 35492 172854
rect 35440 172790 35492 172796
rect 26252 170884 26280 172790
rect 35926 170326 36124 170354
rect 15212 161446 15516 161474
rect 15212 149054 15240 161446
rect 15200 149048 15252 149054
rect 15200 148990 15252 148996
rect 16592 148986 16620 151028
rect 16580 148980 16632 148986
rect 16580 148922 16632 148928
rect 26252 148918 26280 151028
rect 35912 149054 35940 151028
rect 36096 149054 36124 170326
rect 35900 149048 35952 149054
rect 35900 148990 35952 148996
rect 36084 149048 36136 149054
rect 36084 148990 36136 148996
rect 26240 148912 26292 148918
rect 26240 148854 26292 148860
rect 15108 146328 15160 146334
rect 15108 146270 15160 146276
rect 25688 146328 25740 146334
rect 25688 146270 25740 146276
rect 15120 124234 15148 146270
rect 25700 143956 25728 146270
rect 15304 143262 16054 143290
rect 35374 143262 35480 143290
rect 15108 124228 15160 124234
rect 15108 124170 15160 124176
rect 15304 122670 15332 143262
rect 35256 124704 35308 124710
rect 35308 124652 35374 124658
rect 35256 124646 35374 124652
rect 35268 124630 35374 124646
rect 16580 124228 16632 124234
rect 16580 124170 16632 124176
rect 15488 124086 16054 124114
rect 15292 122664 15344 122670
rect 15292 122606 15344 122612
rect 15488 103514 15516 124086
rect 16592 116892 16620 124170
rect 25700 122738 25728 124100
rect 25688 122732 25740 122738
rect 25688 122674 25740 122680
rect 35452 118794 35480 143262
rect 26240 118788 26292 118794
rect 26240 118730 26292 118736
rect 35440 118788 35492 118794
rect 35440 118730 35492 118736
rect 26252 116892 26280 118730
rect 35926 116334 36124 116362
rect 15212 103486 15516 103514
rect 15212 95198 15240 103486
rect 15200 95192 15252 95198
rect 15200 95134 15252 95140
rect 16592 95130 16620 97036
rect 16580 95124 16632 95130
rect 16580 95066 16632 95072
rect 26252 95062 26280 97036
rect 35912 95198 35940 97036
rect 36096 95198 36124 116334
rect 35900 95192 35952 95198
rect 35900 95134 35952 95140
rect 36084 95192 36136 95198
rect 36084 95134 36136 95140
rect 26240 95056 26292 95062
rect 26240 94998 26292 95004
rect 15108 91112 15160 91118
rect 15108 91054 15160 91060
rect 25688 91112 25740 91118
rect 25688 91054 25740 91060
rect 14556 84244 14608 84250
rect 14556 84186 14608 84192
rect 14464 38276 14516 38282
rect 14464 38218 14516 38224
rect 13728 36576 13780 36582
rect 13728 36518 13780 36524
rect 13740 29753 13768 36518
rect 14568 35894 14596 84186
rect 15120 70718 15148 91054
rect 25700 89964 25728 91054
rect 15304 89270 16054 89298
rect 35374 89270 35480 89298
rect 15108 70712 15160 70718
rect 15108 70654 15160 70660
rect 15304 68882 15332 89270
rect 16580 70712 16632 70718
rect 16580 70654 16632 70660
rect 35256 70712 35308 70718
rect 35308 70660 35374 70666
rect 35256 70654 35374 70660
rect 15488 70094 16054 70122
rect 15292 68876 15344 68882
rect 15292 68818 15344 68824
rect 15488 64874 15516 70094
rect 15212 64846 15516 64874
rect 15212 41410 15240 64846
rect 16592 62900 16620 70654
rect 35268 70638 35374 70654
rect 25700 68950 25728 70108
rect 25688 68944 25740 68950
rect 25688 68886 25740 68892
rect 35452 65346 35480 89270
rect 26240 65340 26292 65346
rect 26240 65282 26292 65288
rect 35440 65340 35492 65346
rect 35440 65282 35492 65288
rect 26252 62900 26280 65282
rect 35926 62206 36124 62234
rect 15200 41404 15252 41410
rect 15200 41346 15252 41352
rect 16592 41342 16620 43044
rect 16580 41336 16632 41342
rect 16580 41278 16632 41284
rect 26252 41274 26280 43044
rect 35912 41410 35940 43044
rect 36096 41410 36124 62206
rect 35900 41404 35952 41410
rect 35900 41346 35952 41352
rect 36084 41404 36136 41410
rect 36084 41346 36136 41352
rect 26240 41268 26292 41274
rect 26240 41210 26292 41216
rect 19248 39364 19300 39370
rect 19248 39306 19300 39312
rect 16028 37936 16080 37942
rect 16028 37878 16080 37884
rect 17314 37904 17370 37913
rect 16040 35972 16068 37878
rect 17314 37839 17370 37848
rect 17328 35972 17356 37839
rect 19260 35972 19288 39306
rect 36556 38486 36584 700606
rect 40512 699990 40540 703520
rect 71044 700596 71096 700602
rect 71044 700538 71096 700544
rect 65524 700460 65576 700466
rect 65524 700402 65576 700408
rect 64144 700392 64196 700398
rect 64144 700334 64196 700340
rect 40500 699984 40552 699990
rect 40500 699926 40552 699932
rect 42064 699984 42116 699990
rect 42064 699926 42116 699932
rect 36728 685976 36780 685982
rect 36728 685918 36780 685924
rect 36636 685908 36688 685914
rect 36636 685850 36688 685856
rect 36648 662318 36676 685850
rect 36740 664766 36768 685918
rect 37278 673568 37334 673577
rect 37278 673503 37334 673512
rect 36728 664760 36780 664766
rect 36728 664702 36780 664708
rect 36636 662312 36688 662318
rect 36636 662254 36688 662260
rect 36636 658368 36688 658374
rect 36636 658310 36688 658316
rect 36648 634710 36676 658310
rect 37292 646785 37320 673503
rect 37278 646776 37334 646785
rect 37278 646711 37334 646720
rect 36636 634704 36688 634710
rect 36636 634646 36688 634652
rect 36728 632188 36780 632194
rect 36728 632130 36780 632136
rect 36636 632120 36688 632126
rect 36636 632062 36688 632068
rect 36648 608530 36676 632062
rect 36740 610706 36768 632130
rect 37278 619576 37334 619585
rect 37278 619511 37334 619520
rect 36728 610700 36780 610706
rect 36728 610642 36780 610648
rect 36636 608524 36688 608530
rect 36636 608466 36688 608472
rect 36636 604580 36688 604586
rect 36636 604522 36688 604528
rect 36648 580922 36676 604522
rect 37292 592793 37320 619511
rect 37278 592784 37334 592793
rect 37278 592719 37334 592728
rect 36636 580916 36688 580922
rect 36636 580858 36688 580864
rect 36728 578332 36780 578338
rect 36728 578274 36780 578280
rect 36636 578264 36688 578270
rect 36636 578206 36688 578212
rect 36648 554674 36676 578206
rect 36740 556714 36768 578274
rect 37278 565584 37334 565593
rect 37278 565519 37334 565528
rect 36728 556708 36780 556714
rect 36728 556650 36780 556656
rect 36636 554668 36688 554674
rect 36636 554610 36688 554616
rect 36636 550724 36688 550730
rect 36636 550666 36688 550672
rect 36648 527066 36676 550666
rect 37292 538801 37320 565519
rect 37278 538792 37334 538801
rect 37278 538727 37334 538736
rect 36636 527060 36688 527066
rect 36636 527002 36688 527008
rect 36636 523116 36688 523122
rect 36636 523058 36688 523064
rect 36648 502314 36676 523058
rect 36728 523048 36780 523054
rect 36728 522990 36780 522996
rect 36636 502308 36688 502314
rect 36636 502250 36688 502256
rect 36740 500886 36768 522990
rect 37278 511592 37334 511601
rect 37278 511527 37334 511536
rect 36728 500880 36780 500886
rect 36728 500822 36780 500828
rect 36636 496936 36688 496942
rect 36636 496878 36688 496884
rect 36648 473278 36676 496878
rect 37292 484809 37320 511527
rect 37278 484800 37334 484809
rect 37278 484735 37334 484744
rect 36636 473272 36688 473278
rect 36636 473214 36688 473220
rect 36728 469328 36780 469334
rect 36728 469270 36780 469276
rect 36636 469260 36688 469266
rect 36636 469202 36688 469208
rect 36648 445670 36676 469202
rect 36740 448526 36768 469270
rect 37278 457600 37334 457609
rect 37278 457535 37334 457544
rect 36728 448520 36780 448526
rect 36728 448462 36780 448468
rect 36636 445664 36688 445670
rect 36636 445606 36688 445612
rect 36636 443080 36688 443086
rect 36636 443022 36688 443028
rect 36648 419422 36676 443022
rect 37292 430817 37320 457535
rect 37278 430808 37334 430817
rect 37278 430743 37334 430752
rect 36636 419416 36688 419422
rect 36636 419358 36688 419364
rect 36728 415540 36780 415546
rect 36728 415482 36780 415488
rect 36636 415472 36688 415478
rect 36636 415414 36688 415420
rect 36648 391882 36676 415414
rect 36740 394602 36768 415482
rect 37278 403608 37334 403617
rect 37278 403543 37334 403552
rect 36728 394596 36780 394602
rect 36728 394538 36780 394544
rect 36636 391876 36688 391882
rect 36636 391818 36688 391824
rect 36636 389292 36688 389298
rect 36636 389234 36688 389240
rect 36648 365634 36676 389234
rect 37292 376825 37320 403543
rect 37278 376816 37334 376825
rect 37278 376751 37334 376760
rect 36636 365628 36688 365634
rect 36636 365570 36688 365576
rect 36636 361684 36688 361690
rect 36636 361626 36688 361632
rect 36648 340746 36676 361626
rect 36728 361616 36780 361622
rect 36728 361558 36780 361564
rect 36636 340740 36688 340746
rect 36636 340682 36688 340688
rect 36740 338026 36768 361558
rect 37278 349616 37334 349625
rect 37278 349551 37334 349560
rect 36728 338020 36780 338026
rect 36728 337962 36780 337968
rect 36636 335436 36688 335442
rect 36636 335378 36688 335384
rect 36648 311778 36676 335378
rect 37292 322833 37320 349551
rect 37278 322824 37334 322833
rect 37278 322759 37334 322768
rect 36636 311772 36688 311778
rect 36636 311714 36688 311720
rect 36728 307896 36780 307902
rect 36728 307838 36780 307844
rect 36636 307828 36688 307834
rect 36636 307770 36688 307776
rect 36648 284238 36676 307770
rect 36740 286754 36768 307838
rect 37278 295624 37334 295633
rect 37278 295559 37334 295568
rect 36728 286748 36780 286754
rect 36728 286690 36780 286696
rect 36636 284232 36688 284238
rect 36636 284174 36688 284180
rect 36636 280288 36688 280294
rect 36636 280230 36688 280236
rect 36648 256630 36676 280230
rect 37292 269113 37320 295559
rect 39304 280220 39356 280226
rect 39304 280162 39356 280168
rect 37278 269104 37334 269113
rect 37278 269039 37334 269048
rect 36636 256624 36688 256630
rect 36636 256566 36688 256572
rect 39316 256562 39344 280162
rect 39304 256556 39356 256562
rect 39304 256498 39356 256504
rect 36728 254040 36780 254046
rect 36728 253982 36780 253988
rect 36636 253972 36688 253978
rect 36636 253914 36688 253920
rect 36648 230382 36676 253914
rect 36740 231946 36768 253982
rect 37278 241632 37334 241641
rect 37278 241567 37334 241576
rect 36728 231940 36780 231946
rect 36728 231882 36780 231888
rect 36636 230376 36688 230382
rect 36636 230318 36688 230324
rect 36636 226432 36688 226438
rect 36636 226374 36688 226380
rect 36648 202774 36676 226374
rect 37292 214713 37320 241567
rect 39304 226364 39356 226370
rect 39304 226306 39356 226312
rect 37278 214704 37334 214713
rect 37278 214639 37334 214648
rect 36636 202768 36688 202774
rect 36636 202710 36688 202716
rect 39316 202706 39344 226306
rect 39304 202700 39356 202706
rect 39304 202642 39356 202648
rect 36728 200252 36780 200258
rect 36728 200194 36780 200200
rect 36636 200184 36688 200190
rect 36636 200126 36688 200132
rect 36648 176594 36676 200126
rect 36740 178770 36768 200194
rect 37278 187640 37334 187649
rect 37278 187575 37334 187584
rect 36728 178764 36780 178770
rect 36728 178706 36780 178712
rect 36636 176588 36688 176594
rect 36636 176530 36688 176536
rect 36636 172644 36688 172650
rect 36636 172586 36688 172592
rect 36648 148986 36676 172586
rect 37292 160721 37320 187575
rect 39304 172576 39356 172582
rect 39304 172518 39356 172524
rect 37278 160712 37334 160721
rect 37278 160647 37334 160656
rect 36636 148980 36688 148986
rect 36636 148922 36688 148928
rect 39316 148918 39344 172518
rect 39304 148912 39356 148918
rect 39304 148854 39356 148860
rect 36636 146396 36688 146402
rect 36636 146338 36688 146344
rect 36648 124710 36676 146338
rect 36728 146328 36780 146334
rect 36728 146270 36780 146276
rect 36636 124704 36688 124710
rect 36636 124646 36688 124652
rect 36740 122738 36768 146270
rect 37278 133648 37334 133657
rect 37278 133583 37334 133592
rect 36728 122732 36780 122738
rect 36728 122674 36780 122680
rect 36636 118788 36688 118794
rect 36636 118730 36688 118736
rect 36648 95130 36676 118730
rect 37292 106729 37320 133583
rect 39304 118720 39356 118726
rect 39304 118662 39356 118668
rect 37278 106720 37334 106729
rect 37278 106655 37334 106664
rect 36636 95124 36688 95130
rect 36636 95066 36688 95072
rect 39316 95062 39344 118662
rect 39304 95056 39356 95062
rect 39304 94998 39356 95004
rect 36728 91180 36780 91186
rect 36728 91122 36780 91128
rect 36636 91112 36688 91118
rect 36636 91054 36688 91060
rect 36648 68950 36676 91054
rect 36740 70718 36768 91122
rect 37278 79656 37334 79665
rect 37278 79591 37334 79600
rect 36728 70712 36780 70718
rect 36728 70654 36780 70660
rect 36636 68944 36688 68950
rect 36636 68886 36688 68892
rect 36636 65000 36688 65006
rect 36636 64942 36688 64948
rect 36648 41342 36676 64942
rect 37292 52737 37320 79591
rect 39304 64932 39356 64938
rect 39304 64874 39356 64880
rect 37278 52728 37334 52737
rect 37278 52663 37334 52672
rect 36636 41336 36688 41342
rect 36636 41278 36688 41284
rect 39316 41274 39344 64874
rect 39304 41268 39356 41274
rect 39304 41210 39356 41216
rect 26976 38480 27028 38486
rect 26976 38422 27028 38428
rect 36544 38480 36596 38486
rect 36544 38422 36596 38428
rect 20536 38276 20588 38282
rect 20536 38218 20588 38224
rect 23756 38276 23808 38282
rect 23756 38218 23808 38224
rect 20548 35972 20576 38218
rect 22468 38004 22520 38010
rect 22468 37946 22520 37952
rect 22480 35972 22508 37946
rect 23768 35972 23796 38218
rect 25688 38004 25740 38010
rect 25688 37946 25740 37952
rect 25700 35972 25728 37946
rect 26988 35972 27016 38422
rect 33416 38412 33468 38418
rect 33416 38354 33468 38360
rect 35348 38412 35400 38418
rect 35348 38354 35400 38360
rect 30196 38140 30248 38146
rect 30196 38082 30248 38088
rect 32128 38140 32180 38146
rect 32128 38082 32180 38088
rect 28736 35970 28934 35986
rect 30208 35972 30236 38082
rect 32140 35972 32168 38082
rect 33428 35972 33456 38354
rect 35360 35972 35388 38354
rect 38568 38344 38620 38350
rect 38568 38286 38620 38292
rect 36912 36032 36964 36038
rect 36662 35980 36912 35986
rect 36662 35974 36964 35980
rect 28724 35964 28934 35970
rect 28776 35958 28934 35964
rect 36662 35958 36952 35974
rect 38580 35972 38608 38286
rect 41788 38072 41840 38078
rect 41788 38014 41840 38020
rect 39856 36100 39908 36106
rect 39856 36042 39908 36048
rect 39868 35972 39896 36042
rect 41800 35972 41828 38014
rect 42076 37398 42104 699926
rect 53656 685976 53708 685982
rect 53656 685918 53708 685924
rect 53668 683876 53696 685918
rect 63316 685908 63368 685914
rect 63316 685850 63368 685856
rect 63328 683876 63356 685850
rect 42904 683318 44022 683346
rect 42708 683188 42760 683194
rect 42708 683130 42760 683136
rect 42720 674257 42748 683130
rect 42706 674248 42762 674257
rect 42706 674183 42762 674192
rect 42904 662318 42932 683318
rect 43444 683256 43496 683262
rect 43444 683198 43496 683204
rect 42892 662312 42944 662318
rect 42892 662254 42944 662260
rect 42708 655648 42760 655654
rect 42708 655590 42760 655596
rect 42720 647465 42748 655590
rect 42706 647456 42762 647465
rect 42706 647391 42762 647400
rect 42892 627292 42944 627298
rect 42892 627234 42944 627240
rect 42706 620256 42762 620265
rect 42706 620191 42762 620200
rect 42720 611250 42748 620191
rect 42708 611244 42760 611250
rect 42708 611186 42760 611192
rect 42904 608530 42932 627234
rect 42892 608524 42944 608530
rect 42892 608466 42944 608472
rect 42708 601792 42760 601798
rect 42708 601734 42760 601740
rect 42720 593473 42748 601734
rect 42706 593464 42762 593473
rect 42706 593399 42762 593408
rect 42892 571260 42944 571266
rect 42892 571202 42944 571208
rect 42706 566264 42762 566273
rect 42706 566199 42762 566208
rect 42720 557462 42748 566199
rect 42708 557456 42760 557462
rect 42708 557398 42760 557404
rect 42904 554674 42932 571202
rect 42892 554668 42944 554674
rect 42892 554610 42944 554616
rect 42706 539472 42762 539481
rect 42706 539407 42762 539416
rect 42720 529854 42748 539407
rect 42708 529848 42760 529854
rect 42708 529790 42760 529796
rect 42708 520328 42760 520334
rect 42708 520270 42760 520276
rect 42720 512281 42748 520270
rect 42892 514072 42944 514078
rect 42892 514014 42944 514020
rect 42706 512272 42762 512281
rect 42706 512207 42762 512216
rect 42904 500886 42932 514014
rect 42892 500880 42944 500886
rect 42892 500822 42944 500828
rect 42706 485480 42762 485489
rect 42706 485415 42762 485424
rect 42720 475998 42748 485415
rect 42708 475992 42760 475998
rect 42708 475934 42760 475940
rect 42708 466540 42760 466546
rect 42708 466482 42760 466488
rect 42720 458289 42748 466482
rect 42892 464092 42944 464098
rect 42892 464034 42944 464040
rect 42706 458280 42762 458289
rect 42706 458215 42762 458224
rect 42904 445670 42932 464034
rect 42892 445664 42944 445670
rect 42892 445606 42944 445612
rect 42708 440292 42760 440298
rect 42708 440234 42760 440240
rect 42720 431497 42748 440234
rect 42706 431488 42762 431497
rect 42706 431423 42762 431432
rect 42892 405952 42944 405958
rect 42892 405894 42944 405900
rect 42706 404288 42762 404297
rect 42706 404223 42762 404232
rect 42720 394602 42748 404223
rect 42708 394596 42760 394602
rect 42708 394538 42760 394544
rect 42904 391882 42932 405894
rect 42892 391876 42944 391882
rect 42892 391818 42944 391824
rect 42708 386504 42760 386510
rect 42708 386446 42760 386452
rect 42720 377505 42748 386446
rect 42706 377496 42762 377505
rect 42706 377431 42762 377440
rect 42892 356992 42944 356998
rect 42892 356934 42944 356940
rect 42706 350296 42762 350305
rect 42706 350231 42762 350240
rect 42720 340814 42748 350231
rect 42708 340808 42760 340814
rect 42708 340750 42760 340756
rect 42904 338026 42932 356934
rect 42892 338020 42944 338026
rect 42892 337962 42944 337968
rect 42706 322960 42762 322969
rect 42706 322895 42762 322904
rect 42720 314566 42748 322895
rect 42708 314560 42760 314566
rect 42708 314502 42760 314508
rect 42892 301028 42944 301034
rect 42892 300970 42944 300976
rect 42706 296304 42762 296313
rect 42706 296239 42762 296248
rect 42720 286958 42748 296239
rect 42708 286952 42760 286958
rect 42708 286894 42760 286900
rect 42904 284238 42932 300970
rect 42892 284232 42944 284238
rect 42892 284174 42944 284180
rect 42708 277500 42760 277506
rect 42708 277442 42760 277448
rect 42720 270065 42748 277442
rect 42706 270056 42762 270065
rect 42706 269991 42762 270000
rect 42708 251320 42760 251326
rect 42708 251262 42760 251268
rect 42720 242321 42748 251262
rect 42892 249824 42944 249830
rect 42892 249766 42944 249772
rect 42706 242312 42762 242321
rect 42706 242247 42762 242256
rect 42904 230382 42932 249766
rect 42892 230376 42944 230382
rect 42892 230318 42944 230324
rect 42708 223712 42760 223718
rect 42708 223654 42760 223660
rect 42720 215393 42748 223654
rect 42706 215384 42762 215393
rect 42706 215319 42762 215328
rect 42892 193860 42944 193866
rect 42892 193802 42944 193808
rect 42706 188320 42762 188329
rect 42706 188255 42762 188264
rect 42720 179314 42748 188255
rect 42708 179308 42760 179314
rect 42708 179250 42760 179256
rect 42904 176594 42932 193802
rect 42892 176588 42944 176594
rect 42892 176530 42944 176536
rect 42706 161392 42762 161401
rect 42706 161327 42762 161336
rect 42720 151706 42748 161327
rect 42708 151700 42760 151706
rect 42708 151642 42760 151648
rect 42892 135516 42944 135522
rect 42892 135458 42944 135464
rect 42706 134328 42762 134337
rect 42706 134263 42762 134272
rect 42720 125526 42748 134263
rect 42708 125520 42760 125526
rect 42708 125462 42760 125468
rect 42904 122738 42932 135458
rect 42892 122732 42944 122738
rect 42892 122674 42944 122680
rect 42706 107400 42762 107409
rect 42706 107335 42762 107344
rect 42720 97850 42748 107335
rect 42708 97844 42760 97850
rect 42708 97786 42760 97792
rect 42708 88392 42760 88398
rect 42708 88334 42760 88340
rect 42720 80345 42748 88334
rect 42892 85944 42944 85950
rect 42892 85886 42944 85892
rect 42706 80336 42762 80345
rect 42706 80271 42762 80280
rect 42904 68950 42932 85886
rect 42892 68944 42944 68950
rect 42892 68886 42944 68892
rect 42708 62144 42760 62150
rect 42708 62086 42760 62092
rect 42720 53417 42748 62086
rect 42706 53408 42762 53417
rect 42706 53343 42762 53352
rect 43456 38350 43484 683198
rect 63592 668772 63644 668778
rect 63592 668714 63644 668720
rect 63604 664714 63632 668714
rect 63342 664686 63632 664714
rect 43640 664006 44022 664034
rect 53576 664006 53682 664034
rect 43640 662250 43668 664006
rect 53576 663794 53604 664006
rect 53576 663766 53788 663794
rect 53760 662318 53788 663766
rect 53748 662312 53800 662318
rect 53748 662254 53800 662260
rect 43628 662244 43680 662250
rect 43628 662186 43680 662192
rect 53932 658368 53984 658374
rect 53932 658310 53984 658316
rect 53944 656962 53972 658310
rect 53944 656934 54280 656962
rect 43548 656254 44620 656282
rect 63940 656254 64092 656282
rect 43548 634642 43576 656254
rect 44620 637078 44956 637106
rect 54280 637078 54616 637106
rect 44928 634710 44956 637078
rect 44916 634704 44968 634710
rect 44916 634646 44968 634652
rect 54588 634642 54616 637078
rect 63604 637078 63940 637106
rect 63604 634778 63632 637078
rect 64064 634778 64092 656254
rect 63592 634772 63644 634778
rect 63592 634714 63644 634720
rect 64052 634772 64104 634778
rect 64052 634714 64104 634720
rect 43536 634636 43588 634642
rect 43536 634578 43588 634584
rect 54576 634636 54628 634642
rect 54576 634578 54628 634584
rect 53656 632188 53708 632194
rect 53656 632130 53708 632136
rect 53668 629884 53696 632130
rect 63316 632120 63368 632126
rect 63316 632062 63368 632068
rect 63328 629884 63356 632062
rect 43640 629326 44022 629354
rect 43640 627298 43668 629326
rect 43628 627292 43680 627298
rect 43628 627234 43680 627240
rect 63592 612808 63644 612814
rect 63592 612750 63644 612756
rect 63604 610722 63632 612750
rect 63342 610694 63632 610722
rect 44008 608462 44036 610028
rect 53668 608530 53696 610028
rect 53656 608524 53708 608530
rect 53656 608466 53708 608472
rect 43996 608456 44048 608462
rect 43996 608398 44048 608404
rect 53932 604580 53984 604586
rect 53932 604522 53984 604528
rect 53944 602970 53972 604522
rect 53944 602942 54280 602970
rect 43548 602262 44620 602290
rect 63940 602262 64092 602290
rect 43548 580854 43576 602262
rect 44620 583086 44956 583114
rect 54280 583086 54616 583114
rect 44928 580922 44956 583086
rect 44916 580916 44968 580922
rect 44916 580858 44968 580864
rect 54588 580854 54616 583086
rect 63604 583086 63940 583114
rect 63604 580990 63632 583086
rect 64064 580990 64092 602262
rect 63592 580984 63644 580990
rect 63592 580926 63644 580932
rect 64052 580984 64104 580990
rect 64052 580926 64104 580932
rect 43536 580848 43588 580854
rect 43536 580790 43588 580796
rect 54576 580848 54628 580854
rect 54576 580790 54628 580796
rect 53656 578332 53708 578338
rect 53656 578274 53708 578280
rect 53668 575892 53696 578274
rect 63316 578264 63368 578270
rect 63316 578206 63368 578212
rect 63328 575892 63356 578206
rect 43640 575334 44022 575362
rect 43640 571266 43668 575334
rect 43628 571260 43680 571266
rect 43628 571202 43680 571208
rect 63592 558340 63644 558346
rect 63592 558282 63644 558288
rect 63604 556730 63632 558282
rect 63342 556702 63632 556730
rect 44008 554606 44036 556036
rect 53668 554674 53696 556036
rect 53656 554668 53708 554674
rect 53656 554610 53708 554616
rect 43996 554600 44048 554606
rect 43996 554542 44048 554548
rect 53932 550724 53984 550730
rect 53932 550666 53984 550672
rect 53944 548978 53972 550666
rect 53944 548950 54280 548978
rect 44100 548270 44620 548298
rect 63940 548270 64092 548298
rect 44100 528554 44128 548270
rect 44620 529094 44956 529122
rect 54280 529094 54616 529122
rect 43548 528526 44128 528554
rect 43548 526998 43576 528526
rect 44928 527066 44956 529094
rect 44916 527060 44968 527066
rect 44916 527002 44968 527008
rect 54588 526998 54616 529094
rect 63604 529094 63940 529122
rect 63604 527134 63632 529094
rect 64064 527134 64092 548270
rect 63592 527128 63644 527134
rect 63592 527070 63644 527076
rect 64052 527128 64104 527134
rect 64052 527070 64104 527076
rect 43536 526992 43588 526998
rect 43536 526934 43588 526940
rect 54576 526992 54628 526998
rect 54576 526934 54628 526940
rect 53656 523116 53708 523122
rect 53656 523058 53708 523064
rect 53668 521900 53696 523058
rect 63316 523048 63368 523054
rect 63316 522990 63368 522996
rect 63328 521900 63356 522990
rect 43640 521206 44022 521234
rect 43640 514078 43668 521206
rect 43628 514072 43680 514078
rect 43628 514014 43680 514020
rect 63592 505640 63644 505646
rect 63592 505582 63644 505588
rect 63604 502738 63632 505582
rect 63342 502710 63632 502738
rect 44008 500818 44036 502044
rect 53668 500886 53696 502044
rect 53656 500880 53708 500886
rect 53656 500822 53708 500828
rect 43996 500812 44048 500818
rect 43996 500754 44048 500760
rect 53932 496936 53984 496942
rect 53932 496878 53984 496884
rect 53944 494986 53972 496878
rect 53944 494958 54280 494986
rect 43548 494278 44620 494306
rect 63940 494278 64092 494306
rect 43548 473210 43576 494278
rect 44620 475102 44956 475130
rect 54280 475102 54616 475130
rect 44928 473278 44956 475102
rect 44916 473272 44968 473278
rect 44916 473214 44968 473220
rect 54588 473210 54616 475102
rect 63604 475102 63940 475130
rect 63604 473346 63632 475102
rect 64064 473346 64092 494278
rect 63592 473340 63644 473346
rect 63592 473282 63644 473288
rect 64052 473340 64104 473346
rect 64052 473282 64104 473288
rect 43536 473204 43588 473210
rect 43536 473146 43588 473152
rect 54576 473204 54628 473210
rect 54576 473146 54628 473152
rect 53656 469328 53708 469334
rect 53656 469270 53708 469276
rect 53668 467908 53696 469270
rect 63316 469260 63368 469266
rect 63316 469202 63368 469208
rect 63328 467908 63356 469202
rect 43640 467214 44022 467242
rect 43640 464098 43668 467214
rect 43628 464092 43680 464098
rect 43628 464034 43680 464040
rect 63592 449676 63644 449682
rect 63592 449618 63644 449624
rect 63604 448746 63632 449618
rect 63342 448718 63632 448746
rect 44008 445602 44036 448052
rect 53668 445670 53696 448052
rect 53656 445664 53708 445670
rect 53656 445606 53708 445612
rect 43996 445596 44048 445602
rect 43996 445538 44048 445544
rect 53932 443080 53984 443086
rect 53932 443022 53984 443028
rect 53944 440994 53972 443022
rect 53944 440966 54280 440994
rect 43548 440286 44620 440314
rect 63940 440286 64092 440314
rect 43548 419354 43576 440286
rect 44620 421110 44956 421138
rect 54280 421110 54616 421138
rect 44928 419422 44956 421110
rect 44916 419416 44968 419422
rect 44916 419358 44968 419364
rect 54588 419354 54616 421110
rect 63604 421110 63940 421138
rect 63604 419490 63632 421110
rect 64064 419490 64092 440286
rect 63592 419484 63644 419490
rect 63592 419426 63644 419432
rect 64052 419484 64104 419490
rect 64052 419426 64104 419432
rect 43536 419348 43588 419354
rect 43536 419290 43588 419296
rect 54576 419348 54628 419354
rect 54576 419290 54628 419296
rect 53656 415540 53708 415546
rect 53656 415482 53708 415488
rect 53668 413916 53696 415482
rect 63316 415472 63368 415478
rect 63316 415414 63368 415420
rect 63328 413916 63356 415414
rect 43640 413222 44022 413250
rect 43640 405958 43668 413222
rect 43628 405952 43680 405958
rect 43628 405894 43680 405900
rect 63592 394664 63644 394670
rect 63342 394612 63592 394618
rect 63342 394606 63644 394612
rect 63342 394590 63632 394606
rect 44008 391814 44036 394060
rect 53668 391882 53696 394060
rect 53656 391876 53708 391882
rect 53656 391818 53708 391824
rect 43996 391808 44048 391814
rect 43996 391750 44048 391756
rect 53932 389292 53984 389298
rect 53932 389234 53984 389240
rect 53944 386866 53972 389234
rect 53944 386838 54280 386866
rect 43548 386430 44620 386458
rect 43548 365566 43576 386430
rect 63940 386294 64092 386322
rect 44620 367118 44956 367146
rect 54280 367118 54616 367146
rect 44928 365634 44956 367118
rect 44916 365628 44968 365634
rect 44916 365570 44968 365576
rect 54588 365566 54616 367118
rect 63604 367118 63940 367146
rect 63604 365702 63632 367118
rect 64064 365702 64092 386294
rect 63592 365696 63644 365702
rect 63592 365638 63644 365644
rect 64052 365696 64104 365702
rect 64052 365638 64104 365644
rect 43536 365560 43588 365566
rect 43536 365502 43588 365508
rect 54576 365560 54628 365566
rect 54576 365502 54628 365508
rect 53656 361684 53708 361690
rect 53656 361626 53708 361632
rect 53668 359924 53696 361626
rect 63316 361616 63368 361622
rect 63316 361558 63368 361564
rect 63328 359924 63356 361558
rect 43640 359230 44022 359258
rect 43640 356998 43668 359230
rect 43628 356992 43680 356998
rect 43628 356934 43680 356940
rect 63592 342576 63644 342582
rect 63592 342518 63644 342524
rect 63604 340762 63632 342518
rect 63342 340734 63632 340762
rect 44008 337958 44036 340068
rect 53668 338026 53696 340068
rect 53656 338020 53708 338026
rect 53656 337962 53708 337968
rect 43996 337952 44048 337958
rect 43996 337894 44048 337900
rect 53932 335436 53984 335442
rect 53932 335378 53984 335384
rect 53944 332874 53972 335378
rect 53944 332846 54280 332874
rect 43548 332574 44620 332602
rect 43548 311710 43576 332574
rect 63940 332302 64092 332330
rect 44620 313126 44956 313154
rect 54280 313126 54616 313154
rect 44928 311778 44956 313126
rect 44916 311772 44968 311778
rect 44916 311714 44968 311720
rect 54588 311710 54616 313126
rect 63604 313126 63940 313154
rect 63604 311846 63632 313126
rect 64064 311846 64092 332302
rect 63592 311840 63644 311846
rect 63592 311782 63644 311788
rect 64052 311840 64104 311846
rect 64052 311782 64104 311788
rect 43536 311704 43588 311710
rect 43536 311646 43588 311652
rect 54576 311704 54628 311710
rect 54576 311646 54628 311652
rect 53656 307896 53708 307902
rect 53656 307838 53708 307844
rect 53668 305932 53696 307838
rect 63316 307828 63368 307834
rect 63316 307770 63368 307776
rect 63328 305932 63356 307770
rect 43640 305238 44022 305266
rect 43640 301034 43668 305238
rect 43628 301028 43680 301034
rect 43628 300970 43680 300976
rect 63592 291916 63644 291922
rect 63592 291858 63644 291864
rect 63604 286770 63632 291858
rect 63342 286742 63632 286770
rect 44008 284170 44036 286076
rect 53668 284238 53696 286076
rect 53656 284232 53708 284238
rect 53656 284174 53708 284180
rect 43996 284164 44048 284170
rect 43996 284106 44048 284112
rect 53932 280288 53984 280294
rect 53932 280230 53984 280236
rect 44272 280220 44324 280226
rect 44272 280162 44324 280168
rect 44284 278882 44312 280162
rect 53944 278882 53972 280230
rect 44284 278854 44620 278882
rect 53944 278854 54280 278882
rect 63940 278310 64092 278338
rect 44620 259134 44956 259162
rect 54280 259134 54616 259162
rect 44928 256630 44956 259134
rect 44916 256624 44968 256630
rect 44916 256566 44968 256572
rect 54588 256562 54616 259134
rect 63604 259134 63940 259162
rect 63604 256698 63632 259134
rect 64064 256698 64092 278310
rect 63592 256692 63644 256698
rect 63592 256634 63644 256640
rect 64052 256692 64104 256698
rect 64052 256634 64104 256640
rect 54576 256556 54628 256562
rect 54576 256498 54628 256504
rect 53656 254040 53708 254046
rect 53656 253982 53708 253988
rect 53668 251940 53696 253982
rect 63316 253972 63368 253978
rect 63316 253914 63368 253920
rect 63328 251940 63356 253914
rect 43640 251246 44022 251274
rect 43640 249830 43668 251246
rect 43628 249824 43680 249830
rect 43628 249766 43680 249772
rect 63592 235408 63644 235414
rect 63592 235350 63644 235356
rect 63604 232778 63632 235350
rect 63342 232750 63632 232778
rect 44008 230314 44036 232084
rect 53668 230382 53696 232084
rect 53656 230376 53708 230382
rect 53656 230318 53708 230324
rect 43996 230308 44048 230314
rect 43996 230250 44048 230256
rect 53932 226432 53984 226438
rect 53932 226374 53984 226380
rect 44272 226364 44324 226370
rect 44272 226306 44324 226312
rect 44284 224890 44312 226306
rect 53944 224890 53972 226374
rect 44284 224862 44620 224890
rect 53944 224862 54280 224890
rect 63940 224318 64092 224346
rect 64064 219774 64092 224318
rect 64052 219768 64104 219774
rect 64052 219710 64104 219716
rect 44620 205006 44956 205034
rect 54280 205006 54616 205034
rect 44928 202774 44956 205006
rect 44916 202768 44968 202774
rect 44916 202710 44968 202716
rect 54588 202706 54616 205006
rect 63604 205006 63940 205034
rect 63604 202842 63632 205006
rect 63592 202836 63644 202842
rect 63592 202778 63644 202784
rect 54576 202700 54628 202706
rect 54576 202642 54628 202648
rect 64052 201544 64104 201550
rect 64052 201486 64104 201492
rect 53656 200252 53708 200258
rect 53656 200194 53708 200200
rect 53668 197948 53696 200194
rect 63316 200184 63368 200190
rect 63316 200126 63368 200132
rect 63328 197948 63356 200126
rect 43640 197254 44022 197282
rect 43640 193866 43668 197254
rect 43628 193860 43680 193866
rect 43628 193802 43680 193808
rect 63592 181484 63644 181490
rect 63592 181426 63644 181432
rect 63604 178786 63632 181426
rect 63342 178758 63632 178786
rect 44008 176526 44036 178092
rect 53668 176594 53696 178092
rect 53656 176588 53708 176594
rect 53656 176530 53708 176536
rect 43996 176520 44048 176526
rect 43996 176462 44048 176468
rect 53932 172644 53984 172650
rect 53932 172586 53984 172592
rect 44272 172576 44324 172582
rect 44272 172518 44324 172524
rect 44284 170898 44312 172518
rect 53944 170898 53972 172586
rect 44284 170870 44620 170898
rect 53944 170870 54280 170898
rect 63788 170338 63940 170354
rect 63776 170332 63940 170338
rect 63828 170326 63940 170332
rect 63776 170274 63828 170280
rect 44620 151014 44956 151042
rect 54280 151014 54616 151042
rect 44928 148986 44956 151014
rect 44916 148980 44968 148986
rect 44916 148922 44968 148928
rect 54588 148918 54616 151014
rect 63604 151014 63940 151042
rect 63604 149054 63632 151014
rect 63592 149048 63644 149054
rect 63592 148990 63644 148996
rect 54576 148912 54628 148918
rect 54576 148854 54628 148860
rect 53656 146396 53708 146402
rect 53656 146338 53708 146344
rect 53668 143956 53696 146338
rect 63316 146328 63368 146334
rect 63316 146270 63368 146276
rect 63328 143956 63356 146270
rect 43640 143262 44022 143290
rect 43640 135522 43668 143262
rect 43628 135516 43680 135522
rect 43628 135458 43680 135464
rect 63592 128308 63644 128314
rect 63592 128250 63644 128256
rect 63604 124794 63632 128250
rect 63342 124766 63632 124794
rect 44008 122670 44036 124100
rect 53668 122738 53696 124100
rect 53656 122732 53708 122738
rect 53656 122674 53708 122680
rect 43996 122664 44048 122670
rect 43996 122606 44048 122612
rect 53932 118788 53984 118794
rect 53932 118730 53984 118736
rect 44272 118720 44324 118726
rect 44272 118662 44324 118668
rect 44284 116906 44312 118662
rect 53944 116906 53972 118730
rect 44284 116878 44620 116906
rect 53944 116878 54280 116906
rect 63788 116346 63940 116362
rect 63776 116340 63940 116346
rect 63828 116334 63940 116340
rect 63776 116282 63828 116288
rect 44620 97022 44956 97050
rect 54280 97022 54616 97050
rect 44928 95130 44956 97022
rect 44916 95124 44968 95130
rect 44916 95066 44968 95072
rect 54588 95062 54616 97022
rect 63604 97022 63940 97050
rect 63604 95198 63632 97022
rect 63592 95192 63644 95198
rect 63592 95134 63644 95140
rect 54576 95056 54628 95062
rect 54576 94998 54628 95004
rect 53656 91180 53708 91186
rect 53656 91122 53708 91128
rect 53668 89964 53696 91122
rect 63316 91112 63368 91118
rect 63316 91054 63368 91060
rect 63328 89964 63356 91054
rect 43640 89270 44022 89298
rect 43640 85950 43668 89270
rect 43628 85944 43680 85950
rect 43628 85886 43680 85892
rect 63592 72344 63644 72350
rect 63592 72286 63644 72292
rect 63604 70666 63632 72286
rect 63342 70638 63632 70666
rect 44008 68882 44036 70108
rect 53668 68950 53696 70108
rect 53656 68944 53708 68950
rect 53656 68886 53708 68892
rect 43996 68876 44048 68882
rect 43996 68818 44048 68824
rect 53932 65000 53984 65006
rect 53932 64942 53984 64948
rect 44272 64932 44324 64938
rect 44272 64874 44324 64880
rect 44284 62914 44312 64874
rect 53944 62914 53972 64942
rect 44284 62886 44620 62914
rect 53944 62886 54280 62914
rect 63788 62354 63940 62370
rect 63776 62348 63940 62354
rect 63828 62342 63940 62348
rect 63776 62290 63828 62296
rect 44620 43030 44956 43058
rect 54280 43030 54616 43058
rect 44928 41342 44956 43030
rect 44916 41336 44968 41342
rect 44916 41278 44968 41284
rect 54588 41274 54616 43030
rect 63604 43030 63940 43058
rect 63604 41410 63632 43030
rect 63592 41404 63644 41410
rect 63592 41346 63644 41352
rect 54576 41268 54628 41274
rect 54576 41210 54628 41216
rect 46940 39432 46992 39438
rect 46940 39374 46992 39380
rect 43444 38344 43496 38350
rect 43444 38286 43496 38292
rect 45008 38208 45060 38214
rect 45008 38150 45060 38156
rect 42064 37392 42116 37398
rect 42064 37334 42116 37340
rect 45020 35972 45048 38150
rect 46952 35972 46980 39374
rect 53380 38480 53432 38486
rect 53380 38422 53432 38428
rect 51448 38072 51500 38078
rect 51448 38014 51500 38020
rect 50160 37460 50212 37466
rect 50160 37402 50212 37408
rect 48228 37392 48280 37398
rect 48228 37334 48280 37340
rect 48240 35972 48268 37334
rect 50172 35972 50200 37402
rect 51460 35972 51488 38014
rect 53392 35972 53420 38422
rect 54668 38344 54720 38350
rect 54668 38286 54720 38292
rect 59820 38344 59872 38350
rect 59820 38286 59872 38292
rect 54680 35972 54708 38286
rect 57888 37868 57940 37874
rect 57888 37810 57940 37816
rect 56600 37392 56652 37398
rect 56600 37334 56652 37340
rect 56612 35972 56640 37334
rect 57900 35972 57928 37810
rect 59832 35972 59860 38286
rect 61108 38208 61160 38214
rect 61108 38150 61160 38156
rect 61120 35972 61148 38150
rect 61384 37460 61436 37466
rect 61384 37402 61436 37408
rect 28724 35906 28776 35912
rect 14568 35866 15148 35894
rect 13726 29744 13782 29753
rect 13726 29679 13782 29688
rect 13634 27704 13690 27713
rect 13634 27639 13690 27648
rect 13542 26344 13598 26353
rect 13542 26279 13598 26288
rect 13726 24168 13782 24177
rect 13726 24103 13782 24112
rect 12440 23452 12492 23458
rect 12440 23394 12492 23400
rect 12452 22953 12480 23394
rect 12438 22944 12494 22953
rect 12438 22879 12494 22888
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 12452 20913 12480 22034
rect 12438 20904 12494 20913
rect 12438 20839 12494 20848
rect 12624 20664 12676 20670
rect 12624 20606 12676 20612
rect 12636 19553 12664 20606
rect 12622 19544 12678 19553
rect 12622 19479 12678 19488
rect 12440 17944 12492 17950
rect 12440 17886 12492 17892
rect 12452 17513 12480 17886
rect 12438 17504 12494 17513
rect 12438 17439 12494 17448
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 13740 3534 13768 24103
rect 15120 16574 15148 35866
rect 43442 35320 43498 35329
rect 43498 35278 43746 35306
rect 43442 35255 43498 35264
rect 61292 35216 61344 35222
rect 61292 35158 61344 35164
rect 61304 34377 61332 35158
rect 61290 34368 61346 34377
rect 61290 34303 61346 34312
rect 15120 16546 15608 16574
rect 15580 16538 15608 16546
rect 48042 16552 48098 16561
rect 15580 16510 16054 16538
rect 48098 16510 48254 16538
rect 48042 16487 48098 16496
rect 17328 13734 17356 16116
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 19260 13297 19288 16116
rect 19246 13288 19302 13297
rect 19246 13223 19302 13232
rect 20548 13054 20576 16116
rect 22480 13190 22508 16116
rect 23768 13190 23796 16116
rect 25700 13598 25728 16116
rect 25688 13592 25740 13598
rect 25688 13534 25740 13540
rect 26988 13462 27016 16116
rect 28920 13666 28948 16116
rect 28908 13660 28960 13666
rect 28908 13602 28960 13608
rect 30208 13530 30236 16116
rect 32140 13666 32168 16116
rect 32128 13660 32180 13666
rect 32128 13602 32180 13608
rect 30196 13524 30248 13530
rect 30196 13466 30248 13472
rect 26976 13456 27028 13462
rect 26976 13398 27028 13404
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 33428 13122 33456 16116
rect 33416 13116 33468 13122
rect 33416 13058 33468 13064
rect 20536 13048 20588 13054
rect 20536 12990 20588 12996
rect 35360 12850 35388 16116
rect 36648 13598 36676 16116
rect 36636 13592 36688 13598
rect 36636 13534 36688 13540
rect 38580 13122 38608 16116
rect 39868 13802 39896 16116
rect 41800 15162 41828 16116
rect 41788 15156 41840 15162
rect 41788 15098 41840 15104
rect 39856 13796 39908 13802
rect 39856 13738 39908 13744
rect 43088 13530 43116 16116
rect 43076 13524 43128 13530
rect 43076 13466 43128 13472
rect 45020 13161 45048 16116
rect 45006 13152 45062 13161
rect 38568 13116 38620 13122
rect 45006 13087 45062 13096
rect 38568 13058 38620 13064
rect 46308 12986 46336 16116
rect 48332 16102 49542 16130
rect 46296 12980 46348 12986
rect 46296 12922 46348 12928
rect 35348 12844 35400 12850
rect 35348 12786 35400 12792
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 48332 3466 48360 16102
rect 51460 12918 51488 16116
rect 52748 15094 52776 16116
rect 52736 15088 52788 15094
rect 52736 15030 52788 15036
rect 54680 13326 54708 16116
rect 54668 13320 54720 13326
rect 54668 13262 54720 13268
rect 55968 13258 55996 16116
rect 57900 13394 57928 16116
rect 59832 13569 59860 16116
rect 59818 13560 59874 13569
rect 59818 13495 59874 13504
rect 61120 13433 61148 16116
rect 61106 13424 61162 13433
rect 57888 13388 57940 13394
rect 61106 13359 61162 13368
rect 57888 13330 57940 13336
rect 55956 13252 56008 13258
rect 55956 13194 56008 13200
rect 51448 12912 51500 12918
rect 51448 12854 51500 12860
rect 61396 3602 61424 37402
rect 61476 36100 61528 36106
rect 61476 36042 61528 36048
rect 61384 3596 61436 3602
rect 61384 3538 61436 3544
rect 61488 3466 61516 36042
rect 63500 35216 63552 35222
rect 63500 35158 63552 35164
rect 63512 28393 63540 35158
rect 63498 28384 63554 28393
rect 63498 28319 63554 28328
rect 63500 27600 63552 27606
rect 63500 27542 63552 27548
rect 63512 27033 63540 27542
rect 63498 27024 63554 27033
rect 63498 26959 63554 26968
rect 63498 21448 63554 21457
rect 63498 21383 63554 21392
rect 63512 16590 63540 21383
rect 64064 20233 64092 201486
rect 64156 23633 64184 700334
rect 64236 700324 64288 700330
rect 64236 700266 64288 700272
rect 64248 37874 64276 700266
rect 64328 685976 64380 685982
rect 64328 685918 64380 685924
rect 64340 668778 64368 685918
rect 64328 668772 64380 668778
rect 64328 668714 64380 668720
rect 64328 632188 64380 632194
rect 64328 632130 64380 632136
rect 64340 612814 64368 632130
rect 64328 612808 64380 612814
rect 64328 612750 64380 612756
rect 64328 578332 64380 578338
rect 64328 578274 64380 578280
rect 64340 558346 64368 578274
rect 64328 558340 64380 558346
rect 64328 558282 64380 558288
rect 64328 523116 64380 523122
rect 64328 523058 64380 523064
rect 64340 505646 64368 523058
rect 64328 505640 64380 505646
rect 64328 505582 64380 505588
rect 64328 470620 64380 470626
rect 64328 470562 64380 470568
rect 64236 37868 64288 37874
rect 64236 37810 64288 37816
rect 64236 36780 64288 36786
rect 64236 36722 64288 36728
rect 64248 35193 64276 36722
rect 64234 35184 64290 35193
rect 64234 35119 64290 35128
rect 64234 30288 64290 30297
rect 64234 30223 64290 30232
rect 64142 23624 64198 23633
rect 64142 23559 64198 23568
rect 64050 20224 64106 20233
rect 64050 20159 64106 20168
rect 63500 16584 63552 16590
rect 63500 16526 63552 16532
rect 64248 3670 64276 30223
rect 64340 18193 64368 470562
rect 64420 469328 64472 469334
rect 64420 469270 64472 469276
rect 64432 449682 64460 469270
rect 64420 449676 64472 449682
rect 64420 449618 64472 449624
rect 64420 415540 64472 415546
rect 64420 415482 64472 415488
rect 64432 394670 64460 415482
rect 64420 394664 64472 394670
rect 64420 394606 64472 394612
rect 64420 361684 64472 361690
rect 64420 361626 64472 361632
rect 64432 342582 64460 361626
rect 64420 342576 64472 342582
rect 64420 342518 64472 342524
rect 64420 307896 64472 307902
rect 64420 307838 64472 307844
rect 64432 291922 64460 307838
rect 64420 291916 64472 291922
rect 64420 291858 64472 291864
rect 64420 254040 64472 254046
rect 64420 253982 64472 253988
rect 64432 235414 64460 253982
rect 64420 235408 64472 235414
rect 64420 235350 64472 235356
rect 64420 219768 64472 219774
rect 64420 219710 64472 219716
rect 64432 202842 64460 219710
rect 64420 202836 64472 202842
rect 64420 202778 64472 202784
rect 64420 200252 64472 200258
rect 64420 200194 64472 200200
rect 64432 181490 64460 200194
rect 64420 181484 64472 181490
rect 64420 181426 64472 181432
rect 64420 146396 64472 146402
rect 64420 146338 64472 146344
rect 64432 128314 64460 146338
rect 64420 128308 64472 128314
rect 64420 128250 64472 128256
rect 64420 91180 64472 91186
rect 64420 91122 64472 91128
rect 64432 72350 64460 91122
rect 64420 72344 64472 72350
rect 64420 72286 64472 72292
rect 64604 36712 64656 36718
rect 64604 36654 64656 36660
rect 64512 36644 64564 36650
rect 64512 36586 64564 36592
rect 64524 31657 64552 36586
rect 64510 31648 64566 31657
rect 64510 31583 64566 31592
rect 64616 26234 64644 36654
rect 64524 26206 64644 26234
rect 64418 24984 64474 24993
rect 64418 24919 64474 24928
rect 64326 18184 64382 18193
rect 64326 18119 64382 18128
rect 64432 3738 64460 24919
rect 64524 16833 64552 26206
rect 64510 16824 64566 16833
rect 64510 16759 64566 16768
rect 65536 13190 65564 700402
rect 65616 699712 65668 699718
rect 65616 699654 65668 699660
rect 65628 13802 65656 699654
rect 65708 696992 65760 696998
rect 65708 696934 65760 696940
rect 65720 38486 65748 696934
rect 66904 685908 66956 685914
rect 66904 685850 66956 685856
rect 66258 673568 66314 673577
rect 66258 673503 66314 673512
rect 66272 665174 66300 673503
rect 66260 665168 66312 665174
rect 66260 665110 66312 665116
rect 66916 662318 66944 685850
rect 70306 673840 70362 673849
rect 70306 673775 70362 673784
rect 70320 665174 70348 673775
rect 70308 665168 70360 665174
rect 70308 665110 70360 665116
rect 66904 662312 66956 662318
rect 66904 662254 66956 662260
rect 66904 658300 66956 658306
rect 66904 658242 66956 658248
rect 66260 655580 66312 655586
rect 66260 655522 66312 655528
rect 66272 646785 66300 655522
rect 66258 646776 66314 646785
rect 66258 646711 66314 646720
rect 66916 634642 66944 658242
rect 70308 655580 70360 655586
rect 70308 655522 70360 655528
rect 70320 647465 70348 655522
rect 70306 647456 70362 647465
rect 70306 647391 70362 647400
rect 66904 634636 66956 634642
rect 66904 634578 66956 634584
rect 66904 632120 66956 632126
rect 66904 632062 66956 632068
rect 66258 619576 66314 619585
rect 66258 619511 66314 619520
rect 66272 611318 66300 619511
rect 66260 611312 66312 611318
rect 66260 611254 66312 611260
rect 66916 608530 66944 632062
rect 70306 620256 70362 620265
rect 70306 620191 70362 620200
rect 70320 611318 70348 620191
rect 70308 611312 70360 611318
rect 70308 611254 70360 611260
rect 66904 608524 66956 608530
rect 66904 608466 66956 608472
rect 66904 604512 66956 604518
rect 66904 604454 66956 604460
rect 66260 601724 66312 601730
rect 66260 601666 66312 601672
rect 66272 592793 66300 601666
rect 66258 592784 66314 592793
rect 66258 592719 66314 592728
rect 66916 580854 66944 604454
rect 70308 601724 70360 601730
rect 70308 601666 70360 601672
rect 70320 593473 70348 601666
rect 70306 593464 70362 593473
rect 70306 593399 70362 593408
rect 66904 580848 66956 580854
rect 66904 580790 66956 580796
rect 66904 578264 66956 578270
rect 66904 578206 66956 578212
rect 66258 565584 66314 565593
rect 66258 565519 66314 565528
rect 66272 557530 66300 565519
rect 66260 557524 66312 557530
rect 66260 557466 66312 557472
rect 66916 554674 66944 578206
rect 70306 566264 70362 566273
rect 70306 566199 70362 566208
rect 70320 557530 70348 566199
rect 70308 557524 70360 557530
rect 70308 557466 70360 557472
rect 66904 554668 66956 554674
rect 66904 554610 66956 554616
rect 66904 550656 66956 550662
rect 66904 550598 66956 550604
rect 66258 538792 66314 538801
rect 66258 538727 66314 538736
rect 66272 529922 66300 538727
rect 66260 529916 66312 529922
rect 66260 529858 66312 529864
rect 66916 526998 66944 550598
rect 70306 539472 70362 539481
rect 70306 539407 70362 539416
rect 70320 529922 70348 539407
rect 70308 529916 70360 529922
rect 70308 529858 70360 529864
rect 66904 526992 66956 526998
rect 66904 526934 66956 526940
rect 66904 523048 66956 523054
rect 66904 522990 66956 522996
rect 66258 511592 66314 511601
rect 66258 511527 66314 511536
rect 66272 503674 66300 511527
rect 66260 503668 66312 503674
rect 66260 503610 66312 503616
rect 66916 500886 66944 522990
rect 70306 512272 70362 512281
rect 70306 512207 70362 512216
rect 70320 503674 70348 512207
rect 70308 503668 70360 503674
rect 70308 503610 70360 503616
rect 66904 500880 66956 500886
rect 66904 500822 66956 500828
rect 66904 496868 66956 496874
rect 66904 496810 66956 496816
rect 66258 484800 66314 484809
rect 66258 484735 66314 484744
rect 66272 476066 66300 484735
rect 66260 476060 66312 476066
rect 66260 476002 66312 476008
rect 66916 473210 66944 496810
rect 70306 485480 70362 485489
rect 70306 485415 70362 485424
rect 70320 476066 70348 485415
rect 70308 476060 70360 476066
rect 70308 476002 70360 476008
rect 66904 473204 66956 473210
rect 66904 473146 66956 473152
rect 66904 469260 66956 469266
rect 66904 469202 66956 469208
rect 66260 466472 66312 466478
rect 66260 466414 66312 466420
rect 66272 457609 66300 466414
rect 66258 457600 66314 457609
rect 66258 457535 66314 457544
rect 66916 445670 66944 469202
rect 70308 466472 70360 466478
rect 70308 466414 70360 466420
rect 70320 458289 70348 466414
rect 70306 458280 70362 458289
rect 70306 458215 70362 458224
rect 66904 445664 66956 445670
rect 66904 445606 66956 445612
rect 66904 443012 66956 443018
rect 66904 442954 66956 442960
rect 66258 430808 66314 430817
rect 66258 430743 66314 430752
rect 66272 422278 66300 430743
rect 66260 422272 66312 422278
rect 66260 422214 66312 422220
rect 66916 419354 66944 442954
rect 70306 430944 70362 430953
rect 70306 430879 70362 430888
rect 70320 422278 70348 430879
rect 70308 422272 70360 422278
rect 70308 422214 70360 422220
rect 66904 419348 66956 419354
rect 66904 419290 66956 419296
rect 66904 415472 66956 415478
rect 66904 415414 66956 415420
rect 66258 403608 66314 403617
rect 66258 403543 66314 403552
rect 66272 394534 66300 403543
rect 66260 394528 66312 394534
rect 66260 394470 66312 394476
rect 66916 391882 66944 415414
rect 70306 404288 70362 404297
rect 70306 404223 70362 404232
rect 70320 394670 70348 404223
rect 70308 394664 70360 394670
rect 70308 394606 70360 394612
rect 66904 391876 66956 391882
rect 66904 391818 66956 391824
rect 66904 389224 66956 389230
rect 66904 389166 66956 389172
rect 66260 386436 66312 386442
rect 66260 386378 66312 386384
rect 66272 376825 66300 386378
rect 66258 376816 66314 376825
rect 66258 376751 66314 376760
rect 66916 365566 66944 389166
rect 70308 386436 70360 386442
rect 70308 386378 70360 386384
rect 70320 378049 70348 386378
rect 70306 378040 70362 378049
rect 70306 377975 70362 377984
rect 66904 365560 66956 365566
rect 66904 365502 66956 365508
rect 66904 361616 66956 361622
rect 66904 361558 66956 361564
rect 66258 349616 66314 349625
rect 66258 349551 66314 349560
rect 66272 340882 66300 349551
rect 66260 340876 66312 340882
rect 66260 340818 66312 340824
rect 66916 338026 66944 361558
rect 70306 350296 70362 350305
rect 70306 350231 70362 350240
rect 70320 340882 70348 350231
rect 70308 340876 70360 340882
rect 70308 340818 70360 340824
rect 66904 338020 66956 338026
rect 66904 337962 66956 337968
rect 66904 335368 66956 335374
rect 66904 335310 66956 335316
rect 66258 322144 66314 322153
rect 66258 322079 66314 322088
rect 66272 314634 66300 322079
rect 66260 314628 66312 314634
rect 66260 314570 66312 314576
rect 66916 311710 66944 335310
rect 70306 322960 70362 322969
rect 70306 322895 70362 322904
rect 70320 314634 70348 322895
rect 70308 314628 70360 314634
rect 70308 314570 70360 314576
rect 66904 311704 66956 311710
rect 66904 311646 66956 311652
rect 66904 307828 66956 307834
rect 66904 307770 66956 307776
rect 66258 295624 66314 295633
rect 66258 295559 66314 295568
rect 66272 287026 66300 295559
rect 66260 287020 66312 287026
rect 66260 286962 66312 286968
rect 66916 284238 66944 307770
rect 70306 296304 70362 296313
rect 70306 296239 70362 296248
rect 70320 287026 70348 296239
rect 70308 287020 70360 287026
rect 70308 286962 70360 286968
rect 66904 284232 66956 284238
rect 66904 284174 66956 284180
rect 66904 280220 66956 280226
rect 66904 280162 66956 280168
rect 66260 277432 66312 277438
rect 66260 277374 66312 277380
rect 66272 269113 66300 277374
rect 66258 269104 66314 269113
rect 66258 269039 66314 269048
rect 66916 256562 66944 280162
rect 70308 277432 70360 277438
rect 70308 277374 70360 277380
rect 70320 270065 70348 277374
rect 70306 270056 70362 270065
rect 70306 269991 70362 270000
rect 66904 256556 66956 256562
rect 66904 256498 66956 256504
rect 66904 253972 66956 253978
rect 66904 253914 66956 253920
rect 66258 241632 66314 241641
rect 66258 241567 66314 241576
rect 66272 233238 66300 241567
rect 66260 233232 66312 233238
rect 66260 233174 66312 233180
rect 66916 230382 66944 253914
rect 70306 242312 70362 242321
rect 70306 242247 70362 242256
rect 70320 233238 70348 242247
rect 70308 233232 70360 233238
rect 70308 233174 70360 233180
rect 66904 230376 66956 230382
rect 66904 230318 66956 230324
rect 66904 226364 66956 226370
rect 66904 226306 66956 226312
rect 66260 223644 66312 223650
rect 66260 223586 66312 223592
rect 66272 214713 66300 223586
rect 66258 214704 66314 214713
rect 66258 214639 66314 214648
rect 66916 202706 66944 226306
rect 70308 223644 70360 223650
rect 70308 223586 70360 223592
rect 70320 215937 70348 223586
rect 70306 215928 70362 215937
rect 70306 215863 70362 215872
rect 66904 202700 66956 202706
rect 66904 202642 66956 202648
rect 66904 200184 66956 200190
rect 66904 200126 66956 200132
rect 66258 187640 66314 187649
rect 66258 187575 66314 187584
rect 66272 179382 66300 187575
rect 66260 179376 66312 179382
rect 66260 179318 66312 179324
rect 66916 176594 66944 200126
rect 70306 188320 70362 188329
rect 70306 188255 70362 188264
rect 70320 179382 70348 188255
rect 70308 179376 70360 179382
rect 70308 179318 70360 179324
rect 66904 176588 66956 176594
rect 66904 176530 66956 176536
rect 66904 172576 66956 172582
rect 66904 172518 66956 172524
rect 65800 170332 65852 170338
rect 65800 170274 65852 170280
rect 65812 149054 65840 170274
rect 66258 160712 66314 160721
rect 66258 160647 66314 160656
rect 66272 151774 66300 160647
rect 66260 151768 66312 151774
rect 66260 151710 66312 151716
rect 65800 149048 65852 149054
rect 65800 148990 65852 148996
rect 66916 148918 66944 172518
rect 70306 160848 70362 160857
rect 70306 160783 70362 160792
rect 70320 151774 70348 160783
rect 70308 151768 70360 151774
rect 70308 151710 70360 151716
rect 66904 148912 66956 148918
rect 66904 148854 66956 148860
rect 66904 146328 66956 146334
rect 66904 146270 66956 146276
rect 66258 133648 66314 133657
rect 66258 133583 66314 133592
rect 66272 125594 66300 133583
rect 66260 125588 66312 125594
rect 66260 125530 66312 125536
rect 66916 122738 66944 146270
rect 70306 134328 70362 134337
rect 70306 134263 70362 134272
rect 70320 125594 70348 134263
rect 70308 125588 70360 125594
rect 70308 125530 70360 125536
rect 66904 122732 66956 122738
rect 66904 122674 66956 122680
rect 66904 118720 66956 118726
rect 66904 118662 66956 118668
rect 65800 116340 65852 116346
rect 65800 116282 65852 116288
rect 65812 95198 65840 116282
rect 66258 106720 66314 106729
rect 66258 106655 66314 106664
rect 66272 97986 66300 106655
rect 66260 97980 66312 97986
rect 66260 97922 66312 97928
rect 65800 95192 65852 95198
rect 65800 95134 65852 95140
rect 66916 95062 66944 118662
rect 70306 107400 70362 107409
rect 70306 107335 70362 107344
rect 70320 97918 70348 107335
rect 70308 97912 70360 97918
rect 70308 97854 70360 97860
rect 66904 95056 66956 95062
rect 66904 94998 66956 95004
rect 66904 91112 66956 91118
rect 66904 91054 66956 91060
rect 66258 79656 66314 79665
rect 66258 79591 66314 79600
rect 66272 71738 66300 79591
rect 66260 71732 66312 71738
rect 66260 71674 66312 71680
rect 66916 68950 66944 91054
rect 70306 80336 70362 80345
rect 70306 80271 70362 80280
rect 70320 71738 70348 80271
rect 70308 71732 70360 71738
rect 70308 71674 70360 71680
rect 66904 68944 66956 68950
rect 66904 68886 66956 68892
rect 66904 64932 66956 64938
rect 66904 64874 66956 64880
rect 65800 62348 65852 62354
rect 65800 62290 65852 62296
rect 65812 41410 65840 62290
rect 66258 52728 66314 52737
rect 66258 52663 66314 52672
rect 66272 44130 66300 52663
rect 66260 44124 66312 44130
rect 66260 44066 66312 44072
rect 65800 41404 65852 41410
rect 65800 41346 65852 41352
rect 66916 41274 66944 64874
rect 70306 53408 70362 53417
rect 70306 53343 70362 53352
rect 70320 44130 70348 53343
rect 70308 44124 70360 44130
rect 70308 44066 70360 44072
rect 66904 41268 66956 41274
rect 66904 41210 66956 41216
rect 65708 38480 65760 38486
rect 65708 38422 65760 38428
rect 70308 34604 70360 34610
rect 70308 34546 70360 34552
rect 70320 26897 70348 34546
rect 71056 27606 71084 700538
rect 72988 699718 73016 703520
rect 105464 700670 105492 703520
rect 105452 700664 105504 700670
rect 105452 700606 105504 700612
rect 137848 700466 137876 703520
rect 170324 700466 170352 703520
rect 137836 700460 137888 700466
rect 137836 700402 137888 700408
rect 153844 700460 153896 700466
rect 153844 700402 153896 700408
rect 170312 700460 170364 700466
rect 170312 700402 170364 700408
rect 72976 699712 73028 699718
rect 72976 699654 73028 699660
rect 148324 686044 148376 686050
rect 148324 685986 148376 685992
rect 81440 685976 81492 685982
rect 81440 685918 81492 685924
rect 91468 685976 91520 685982
rect 91468 685918 91520 685924
rect 109684 685976 109736 685982
rect 109684 685918 109736 685924
rect 119436 685976 119488 685982
rect 119436 685918 119488 685924
rect 137652 685976 137704 685982
rect 137652 685918 137704 685924
rect 81452 683890 81480 685918
rect 91100 685908 91152 685914
rect 91100 685850 91152 685856
rect 91112 683890 91140 685850
rect 81452 683862 81696 683890
rect 91112 683862 91356 683890
rect 71884 683318 72036 683346
rect 71884 662386 71912 683318
rect 91480 664714 91508 685918
rect 93124 685908 93176 685914
rect 93124 685850 93176 685856
rect 91356 664686 91508 664714
rect 72022 663794 72050 664020
rect 81696 664006 82032 664034
rect 71976 663766 72050 663794
rect 71872 662380 71924 662386
rect 71872 662322 71924 662328
rect 71976 662250 72004 663766
rect 82004 662318 82032 664006
rect 93136 662318 93164 685850
rect 109696 683876 109724 685918
rect 119344 685908 119396 685914
rect 119344 685850 119396 685856
rect 119356 683876 119384 685850
rect 99484 683318 100050 683346
rect 93860 683188 93912 683194
rect 93860 683130 93912 683136
rect 97908 683188 97960 683194
rect 97908 683130 97960 683136
rect 93872 673577 93900 683130
rect 97920 674257 97948 683130
rect 97906 674248 97962 674257
rect 97906 674183 97962 674192
rect 93858 673568 93914 673577
rect 93858 673503 93914 673512
rect 99484 662318 99512 683318
rect 119448 664714 119476 685918
rect 122104 685908 122156 685914
rect 122104 685850 122156 685856
rect 121458 673568 121514 673577
rect 121458 673503 121514 673512
rect 121472 665174 121500 673503
rect 121460 665168 121512 665174
rect 121460 665110 121512 665116
rect 119370 664686 119476 664714
rect 100036 662386 100064 664020
rect 100024 662380 100076 662386
rect 100024 662322 100076 662328
rect 109696 662318 109724 664020
rect 122116 662318 122144 685850
rect 137664 683876 137692 685918
rect 147312 685908 147364 685914
rect 147312 685850 147364 685856
rect 147324 683876 147352 685850
rect 127084 683318 128018 683346
rect 126886 674248 126942 674257
rect 126886 674183 126942 674192
rect 126900 665174 126928 674183
rect 126888 665168 126940 665174
rect 126888 665110 126940 665116
rect 81992 662312 82044 662318
rect 81992 662254 82044 662260
rect 93124 662312 93176 662318
rect 93124 662254 93176 662260
rect 99472 662312 99524 662318
rect 99472 662254 99524 662260
rect 109684 662312 109736 662318
rect 109684 662254 109736 662260
rect 122104 662312 122156 662318
rect 122104 662254 122156 662260
rect 127084 662250 127112 683318
rect 148336 673454 148364 685986
rect 148416 685908 148468 685914
rect 148416 685850 148468 685856
rect 147784 673426 148364 673454
rect 147784 664714 147812 673426
rect 147338 664686 147812 664714
rect 127728 664006 128018 664034
rect 137678 664006 137968 664034
rect 127728 662386 127756 664006
rect 127716 662380 127768 662386
rect 127716 662322 127768 662328
rect 137940 662318 137968 664006
rect 148428 662318 148456 685850
rect 149060 683188 149112 683194
rect 149060 683130 149112 683136
rect 149072 673577 149100 683130
rect 149058 673568 149114 673577
rect 149058 673503 149114 673512
rect 137928 662312 137980 662318
rect 137928 662254 137980 662260
rect 148416 662312 148468 662318
rect 148416 662254 148468 662260
rect 71964 662244 72016 662250
rect 71964 662186 72016 662192
rect 127072 662244 127124 662250
rect 127072 662186 127124 662192
rect 71136 658436 71188 658442
rect 71136 658378 71188 658384
rect 82268 658436 82320 658442
rect 82268 658378 82320 658384
rect 99472 658436 99524 658442
rect 99472 658378 99524 658384
rect 100392 658436 100444 658442
rect 100392 658378 100444 658384
rect 71148 634710 71176 658378
rect 71872 658368 71924 658374
rect 71872 658310 71924 658316
rect 71884 654134 71912 658310
rect 72608 658300 72660 658306
rect 72608 658242 72660 658248
rect 72620 656948 72648 658242
rect 82280 656948 82308 658378
rect 93124 658300 93176 658306
rect 93124 658242 93176 658248
rect 91954 656254 92152 656282
rect 71884 654106 72280 654134
rect 72252 637786 72280 654106
rect 72252 637758 72634 637786
rect 82280 634710 82308 637092
rect 91940 634778 91968 637092
rect 92124 634778 92152 656254
rect 91928 634772 91980 634778
rect 91928 634714 91980 634720
rect 92112 634772 92164 634778
rect 92112 634714 92164 634720
rect 93136 634710 93164 658242
rect 93860 655648 93912 655654
rect 93860 655590 93912 655596
rect 97908 655648 97960 655654
rect 97908 655590 97960 655596
rect 93872 646785 93900 655590
rect 97920 647465 97948 655590
rect 99484 654134 99512 658378
rect 100404 658306 100432 658378
rect 109960 658368 110012 658374
rect 109960 658310 110012 658316
rect 124864 658368 124916 658374
rect 124864 658310 124916 658316
rect 128636 658368 128688 658374
rect 128636 658310 128688 658316
rect 151084 658368 151136 658374
rect 151084 658310 151136 658316
rect 100300 658300 100352 658306
rect 100300 658242 100352 658248
rect 100392 658300 100444 658306
rect 100392 658242 100444 658248
rect 100312 656962 100340 658242
rect 109972 656962 110000 658310
rect 100312 656934 100648 656962
rect 109972 656934 110308 656962
rect 119968 656266 120212 656282
rect 119968 656260 120224 656266
rect 119968 656254 120172 656260
rect 120172 656202 120224 656208
rect 122104 656260 122156 656266
rect 122104 656202 122156 656208
rect 121460 655580 121512 655586
rect 121460 655522 121512 655528
rect 99484 654106 100248 654134
rect 97906 647456 97962 647465
rect 97906 647391 97962 647400
rect 93858 646776 93914 646785
rect 93858 646711 93914 646720
rect 100220 637786 100248 654106
rect 121472 646785 121500 655522
rect 121458 646776 121514 646785
rect 121458 646711 121514 646720
rect 100220 637758 100648 637786
rect 110294 636834 110322 637092
rect 119632 637078 119968 637106
rect 110294 636806 110368 636834
rect 110340 634710 110368 636806
rect 119632 634778 119660 637078
rect 122116 634778 122144 656202
rect 119620 634772 119672 634778
rect 119620 634714 119672 634720
rect 122104 634772 122156 634778
rect 122104 634714 122156 634720
rect 124876 634710 124904 658310
rect 128648 656948 128676 658310
rect 138296 658300 138348 658306
rect 138296 658242 138348 658248
rect 149704 658300 149756 658306
rect 149704 658242 149756 658248
rect 138308 656948 138336 658242
rect 147982 656254 148088 656282
rect 126888 655580 126940 655586
rect 126888 655522 126940 655528
rect 126900 647465 126928 655522
rect 126886 647456 126942 647465
rect 126886 647391 126942 647400
rect 128648 634710 128676 637092
rect 71136 634704 71188 634710
rect 71136 634646 71188 634652
rect 82268 634704 82320 634710
rect 82268 634646 82320 634652
rect 93124 634704 93176 634710
rect 93124 634646 93176 634652
rect 110328 634704 110380 634710
rect 110328 634646 110380 634652
rect 124864 634704 124916 634710
rect 124864 634646 124916 634652
rect 128636 634704 128688 634710
rect 128636 634646 128688 634652
rect 138308 634642 138336 637092
rect 147968 634778 147996 637092
rect 148060 634778 148088 656254
rect 149060 655648 149112 655654
rect 149060 655590 149112 655596
rect 149072 646785 149100 655590
rect 149058 646776 149114 646785
rect 149058 646711 149114 646720
rect 147956 634772 148008 634778
rect 147956 634714 148008 634720
rect 148048 634772 148100 634778
rect 148048 634714 148100 634720
rect 149716 634710 149744 658242
rect 149704 634704 149756 634710
rect 149704 634646 149756 634652
rect 151096 634642 151124 658310
rect 138296 634636 138348 634642
rect 138296 634578 138348 634584
rect 151084 634636 151136 634642
rect 151084 634578 151136 634584
rect 148324 632256 148376 632262
rect 148324 632198 148376 632204
rect 81440 632188 81492 632194
rect 81440 632130 81492 632136
rect 91468 632188 91520 632194
rect 91468 632130 91520 632136
rect 109684 632188 109736 632194
rect 109684 632130 109736 632136
rect 119436 632188 119488 632194
rect 119436 632130 119488 632136
rect 137652 632188 137704 632194
rect 137652 632130 137704 632136
rect 81452 629898 81480 632130
rect 91100 632120 91152 632126
rect 91100 632062 91152 632068
rect 91112 629898 91140 632062
rect 81452 629870 81696 629898
rect 91112 629870 91356 629898
rect 71884 629326 72036 629354
rect 71884 608598 71912 629326
rect 91480 610722 91508 632130
rect 93124 632120 93176 632126
rect 93124 632062 93176 632068
rect 91356 610694 91508 610722
rect 72036 610014 72096 610042
rect 81696 610014 82032 610042
rect 71872 608592 71924 608598
rect 71872 608534 71924 608540
rect 72068 608462 72096 610014
rect 82004 608530 82032 610014
rect 93136 608530 93164 632062
rect 109696 629884 109724 632130
rect 119344 632120 119396 632126
rect 119344 632062 119396 632068
rect 119356 629884 119384 632062
rect 99484 629326 100050 629354
rect 97906 620256 97962 620265
rect 97906 620191 97962 620200
rect 93858 619576 93914 619585
rect 93858 619511 93914 619520
rect 93872 611250 93900 619511
rect 97920 611250 97948 620191
rect 93860 611244 93912 611250
rect 93860 611186 93912 611192
rect 97908 611244 97960 611250
rect 97908 611186 97960 611192
rect 99484 608530 99512 629326
rect 119448 610722 119476 632130
rect 124864 632120 124916 632126
rect 124864 632062 124916 632068
rect 121458 619576 121514 619585
rect 121458 619511 121514 619520
rect 121472 611318 121500 619511
rect 121460 611312 121512 611318
rect 121460 611254 121512 611260
rect 119370 610694 119476 610722
rect 100036 608598 100064 610028
rect 100024 608592 100076 608598
rect 100024 608534 100076 608540
rect 109696 608530 109724 610028
rect 124876 608530 124904 632062
rect 137664 629884 137692 632130
rect 147312 632120 147364 632126
rect 147312 632062 147364 632068
rect 147324 629884 147352 632062
rect 127084 629326 128018 629354
rect 126886 620256 126942 620265
rect 126886 620191 126942 620200
rect 126900 611318 126928 620191
rect 126888 611312 126940 611318
rect 126888 611254 126940 611260
rect 81992 608524 82044 608530
rect 81992 608466 82044 608472
rect 93124 608524 93176 608530
rect 93124 608466 93176 608472
rect 99472 608524 99524 608530
rect 99472 608466 99524 608472
rect 109684 608524 109736 608530
rect 109684 608466 109736 608472
rect 124864 608524 124916 608530
rect 124864 608466 124916 608472
rect 127084 608462 127112 629326
rect 148336 615494 148364 632198
rect 148416 632120 148468 632126
rect 148416 632062 148468 632068
rect 147784 615466 148364 615494
rect 147784 610722 147812 615466
rect 147338 610694 147812 610722
rect 128004 608598 128032 610028
rect 127992 608592 128044 608598
rect 127992 608534 128044 608540
rect 137664 608530 137692 610028
rect 148428 608530 148456 632062
rect 149058 619576 149114 619585
rect 149058 619511 149114 619520
rect 149072 611250 149100 619511
rect 149060 611244 149112 611250
rect 149060 611186 149112 611192
rect 137652 608524 137704 608530
rect 137652 608466 137704 608472
rect 148416 608524 148468 608530
rect 148416 608466 148468 608472
rect 72056 608456 72108 608462
rect 72056 608398 72108 608404
rect 127072 608456 127124 608462
rect 127072 608398 127124 608404
rect 71136 604648 71188 604654
rect 71136 604590 71188 604596
rect 82268 604648 82320 604654
rect 82268 604590 82320 604596
rect 99472 604648 99524 604654
rect 99472 604590 99524 604596
rect 100392 604648 100444 604654
rect 100392 604590 100444 604596
rect 71148 580922 71176 604590
rect 71872 604580 71924 604586
rect 71872 604522 71924 604528
rect 71884 596174 71912 604522
rect 72608 604512 72660 604518
rect 72608 604454 72660 604460
rect 72620 602956 72648 604454
rect 82280 602956 82308 604590
rect 93124 604512 93176 604518
rect 93124 604454 93176 604460
rect 91954 602262 92152 602290
rect 71884 596146 72280 596174
rect 72252 583794 72280 596146
rect 72252 583766 72634 583794
rect 82280 580922 82308 583100
rect 91940 580990 91968 583100
rect 92124 580990 92152 602262
rect 91928 580984 91980 580990
rect 91928 580926 91980 580932
rect 92112 580984 92164 580990
rect 92112 580926 92164 580932
rect 93136 580922 93164 604454
rect 93860 601792 93912 601798
rect 93860 601734 93912 601740
rect 97908 601792 97960 601798
rect 97908 601734 97960 601740
rect 93872 592793 93900 601734
rect 97920 593473 97948 601734
rect 99484 596174 99512 604590
rect 100404 604518 100432 604590
rect 109960 604580 110012 604586
rect 109960 604522 110012 604528
rect 151084 604580 151136 604586
rect 151084 604522 151136 604528
rect 100300 604512 100352 604518
rect 100300 604454 100352 604460
rect 100392 604512 100444 604518
rect 100392 604454 100444 604460
rect 100312 602970 100340 604454
rect 109972 602970 110000 604522
rect 138296 604512 138348 604518
rect 138296 604454 138348 604460
rect 149704 604512 149756 604518
rect 149704 604454 149756 604460
rect 100312 602942 100648 602970
rect 109972 602942 110308 602970
rect 138308 602956 138336 604454
rect 119968 602274 120212 602290
rect 128280 602274 128662 602290
rect 119968 602268 120224 602274
rect 119968 602262 120172 602268
rect 120172 602210 120224 602216
rect 122104 602268 122156 602274
rect 122104 602210 122156 602216
rect 124864 602268 124916 602274
rect 124864 602210 124916 602216
rect 128268 602268 128662 602274
rect 128320 602262 128662 602268
rect 147982 602262 148088 602290
rect 128268 602210 128320 602216
rect 121460 601724 121512 601730
rect 121460 601666 121512 601672
rect 99484 596146 100248 596174
rect 97906 593464 97962 593473
rect 97906 593399 97962 593408
rect 93858 592784 93914 592793
rect 93858 592719 93914 592728
rect 100220 583794 100248 596146
rect 121472 592793 121500 601666
rect 121458 592784 121514 592793
rect 121458 592719 121514 592728
rect 100220 583766 100648 583794
rect 110248 583086 110308 583114
rect 119632 583086 119968 583114
rect 110248 580922 110276 583086
rect 119632 580990 119660 583086
rect 122116 580990 122144 602210
rect 119620 580984 119672 580990
rect 119620 580926 119672 580932
rect 122104 580984 122156 580990
rect 122104 580926 122156 580932
rect 124876 580922 124904 602210
rect 126888 601724 126940 601730
rect 126888 601666 126940 601672
rect 126900 593473 126928 601666
rect 126886 593464 126942 593473
rect 126886 593399 126942 593408
rect 128648 580922 128676 583100
rect 71136 580916 71188 580922
rect 71136 580858 71188 580864
rect 82268 580916 82320 580922
rect 82268 580858 82320 580864
rect 93124 580916 93176 580922
rect 93124 580858 93176 580864
rect 110236 580916 110288 580922
rect 110236 580858 110288 580864
rect 124864 580916 124916 580922
rect 124864 580858 124916 580864
rect 128636 580916 128688 580922
rect 128636 580858 128688 580864
rect 138308 580854 138336 583100
rect 147968 580990 147996 583100
rect 148060 580990 148088 602262
rect 149060 601792 149112 601798
rect 149060 601734 149112 601740
rect 149072 592793 149100 601734
rect 149058 592784 149114 592793
rect 149058 592719 149114 592728
rect 147956 580984 148008 580990
rect 147956 580926 148008 580932
rect 148048 580984 148100 580990
rect 148048 580926 148100 580932
rect 149716 580922 149744 604454
rect 149704 580916 149756 580922
rect 149704 580858 149756 580864
rect 151096 580854 151124 604522
rect 138296 580848 138348 580854
rect 138296 580790 138348 580796
rect 151084 580848 151136 580854
rect 151084 580790 151136 580796
rect 148416 578400 148468 578406
rect 148416 578342 148468 578348
rect 81440 578332 81492 578338
rect 81440 578274 81492 578280
rect 91468 578332 91520 578338
rect 91468 578274 91520 578280
rect 109684 578332 109736 578338
rect 109684 578274 109736 578280
rect 119436 578332 119488 578338
rect 119436 578274 119488 578280
rect 137652 578332 137704 578338
rect 137652 578274 137704 578280
rect 81452 575906 81480 578274
rect 91100 578264 91152 578270
rect 91100 578206 91152 578212
rect 91112 575906 91140 578206
rect 81452 575878 81696 575906
rect 91112 575878 91356 575906
rect 71884 575334 72036 575362
rect 71884 554742 71912 575334
rect 91480 556730 91508 578274
rect 93124 578264 93176 578270
rect 93124 578206 93176 578212
rect 91356 556702 91508 556730
rect 72036 556022 72096 556050
rect 81696 556022 82032 556050
rect 71872 554736 71924 554742
rect 71872 554678 71924 554684
rect 72068 554606 72096 556022
rect 82004 554674 82032 556022
rect 93136 554674 93164 578206
rect 109696 575892 109724 578274
rect 119344 578264 119396 578270
rect 119344 578206 119396 578212
rect 119356 575892 119384 578206
rect 99484 575334 100050 575362
rect 97906 566264 97962 566273
rect 97906 566199 97962 566208
rect 93858 565584 93914 565593
rect 93858 565519 93914 565528
rect 93872 557462 93900 565519
rect 97920 557462 97948 566199
rect 93860 557456 93912 557462
rect 93860 557398 93912 557404
rect 97908 557456 97960 557462
rect 97908 557398 97960 557404
rect 99484 554674 99512 575334
rect 119448 556730 119476 578274
rect 124864 578264 124916 578270
rect 124864 578206 124916 578212
rect 121458 565584 121514 565593
rect 121458 565519 121514 565528
rect 121472 557530 121500 565519
rect 121460 557524 121512 557530
rect 121460 557466 121512 557472
rect 119370 556702 119476 556730
rect 100036 554742 100064 556036
rect 100024 554736 100076 554742
rect 100024 554678 100076 554684
rect 109696 554674 109724 556036
rect 124876 554674 124904 578206
rect 137664 575892 137692 578274
rect 147312 578264 147364 578270
rect 147312 578206 147364 578212
rect 148324 578264 148376 578270
rect 148324 578206 148376 578212
rect 147324 575892 147352 578206
rect 127084 575334 128018 575362
rect 126886 566264 126942 566273
rect 126886 566199 126942 566208
rect 126900 557530 126928 566199
rect 126888 557524 126940 557530
rect 126888 557466 126940 557472
rect 81992 554668 82044 554674
rect 81992 554610 82044 554616
rect 93124 554668 93176 554674
rect 93124 554610 93176 554616
rect 99472 554668 99524 554674
rect 99472 554610 99524 554616
rect 109684 554668 109736 554674
rect 109684 554610 109736 554616
rect 124864 554668 124916 554674
rect 124864 554610 124916 554616
rect 127084 554606 127112 575334
rect 147680 562352 147732 562358
rect 147680 562294 147732 562300
rect 147692 556730 147720 562294
rect 147338 556702 147720 556730
rect 128004 554742 128032 556036
rect 127992 554736 128044 554742
rect 127992 554678 128044 554684
rect 137664 554674 137692 556036
rect 148336 554674 148364 578206
rect 148428 562358 148456 578342
rect 149058 565584 149114 565593
rect 149058 565519 149114 565528
rect 148416 562352 148468 562358
rect 148416 562294 148468 562300
rect 149072 557462 149100 565519
rect 149060 557456 149112 557462
rect 149060 557398 149112 557404
rect 137652 554668 137704 554674
rect 137652 554610 137704 554616
rect 148324 554668 148376 554674
rect 148324 554610 148376 554616
rect 72056 554600 72108 554606
rect 72056 554542 72108 554548
rect 127072 554600 127124 554606
rect 127072 554542 127124 554548
rect 71136 550792 71188 550798
rect 71136 550734 71188 550740
rect 82268 550792 82320 550798
rect 82268 550734 82320 550740
rect 99472 550792 99524 550798
rect 99472 550734 99524 550740
rect 100392 550792 100444 550798
rect 100392 550734 100444 550740
rect 71148 527066 71176 550734
rect 71872 550724 71924 550730
rect 71872 550666 71924 550672
rect 71884 538214 71912 550666
rect 72608 550656 72660 550662
rect 72608 550598 72660 550604
rect 72620 548964 72648 550598
rect 82280 548964 82308 550734
rect 93124 550656 93176 550662
rect 93124 550598 93176 550604
rect 91954 548270 92152 548298
rect 71884 538186 72280 538214
rect 72252 529666 72280 538186
rect 72252 529638 72634 529666
rect 82280 527066 82308 529108
rect 91940 527134 91968 529108
rect 92124 527134 92152 548270
rect 91928 527128 91980 527134
rect 91928 527070 91980 527076
rect 92112 527128 92164 527134
rect 92112 527070 92164 527076
rect 93136 527066 93164 550598
rect 97906 539472 97962 539481
rect 97906 539407 97962 539416
rect 93858 538792 93914 538801
rect 93858 538727 93914 538736
rect 93872 529854 93900 538727
rect 97920 529854 97948 539407
rect 99484 538214 99512 550734
rect 100404 550662 100432 550734
rect 109960 550724 110012 550730
rect 109960 550666 110012 550672
rect 151084 550724 151136 550730
rect 151084 550666 151136 550672
rect 100300 550656 100352 550662
rect 100300 550598 100352 550604
rect 100392 550656 100444 550662
rect 100392 550598 100444 550604
rect 100312 548978 100340 550598
rect 109972 548978 110000 550666
rect 138296 550656 138348 550662
rect 138296 550598 138348 550604
rect 149704 550656 149756 550662
rect 149704 550598 149756 550604
rect 100312 548950 100648 548978
rect 109972 548950 110308 548978
rect 138308 548964 138336 550598
rect 119968 548282 120120 548298
rect 128280 548282 128662 548298
rect 119968 548276 120132 548282
rect 119968 548270 120080 548276
rect 120080 548218 120132 548224
rect 122104 548276 122156 548282
rect 122104 548218 122156 548224
rect 124864 548276 124916 548282
rect 124864 548218 124916 548224
rect 128268 548276 128662 548282
rect 128320 548270 128662 548276
rect 147982 548270 148088 548298
rect 128268 548218 128320 548224
rect 121458 538792 121514 538801
rect 121458 538727 121514 538736
rect 99484 538186 100248 538214
rect 93860 529848 93912 529854
rect 93860 529790 93912 529796
rect 97908 529848 97960 529854
rect 97908 529790 97960 529796
rect 100220 529666 100248 538186
rect 121472 529922 121500 538727
rect 121460 529916 121512 529922
rect 121460 529858 121512 529864
rect 100220 529638 100648 529666
rect 110294 528850 110322 529108
rect 119632 529094 119968 529122
rect 110294 528822 110368 528850
rect 110340 527066 110368 528822
rect 119632 527134 119660 529094
rect 122116 527134 122144 548218
rect 119620 527128 119672 527134
rect 119620 527070 119672 527076
rect 122104 527128 122156 527134
rect 122104 527070 122156 527076
rect 124876 527066 124904 548218
rect 126886 539472 126942 539481
rect 126886 539407 126942 539416
rect 126900 529922 126928 539407
rect 126888 529916 126940 529922
rect 126888 529858 126940 529864
rect 128648 527066 128676 529108
rect 71136 527060 71188 527066
rect 71136 527002 71188 527008
rect 82268 527060 82320 527066
rect 82268 527002 82320 527008
rect 93124 527060 93176 527066
rect 93124 527002 93176 527008
rect 110328 527060 110380 527066
rect 110328 527002 110380 527008
rect 124864 527060 124916 527066
rect 124864 527002 124916 527008
rect 128636 527060 128688 527066
rect 128636 527002 128688 527008
rect 138308 526998 138336 529108
rect 147968 527134 147996 529108
rect 148060 527134 148088 548270
rect 149058 538792 149114 538801
rect 149058 538727 149114 538736
rect 149072 529854 149100 538727
rect 149060 529848 149112 529854
rect 149060 529790 149112 529796
rect 147956 527128 148008 527134
rect 147956 527070 148008 527076
rect 148048 527128 148100 527134
rect 148048 527070 148100 527076
rect 149716 527066 149744 550598
rect 149704 527060 149756 527066
rect 149704 527002 149756 527008
rect 151096 526998 151124 550666
rect 138296 526992 138348 526998
rect 138296 526934 138348 526940
rect 151084 526992 151136 526998
rect 151084 526934 151136 526940
rect 148416 523184 148468 523190
rect 148416 523126 148468 523132
rect 81440 523116 81492 523122
rect 81440 523058 81492 523064
rect 91468 523116 91520 523122
rect 91468 523058 91520 523064
rect 109684 523116 109736 523122
rect 109684 523058 109736 523064
rect 119436 523116 119488 523122
rect 119436 523058 119488 523064
rect 137652 523116 137704 523122
rect 137652 523058 137704 523064
rect 81452 521914 81480 523058
rect 91100 523048 91152 523054
rect 91100 522990 91152 522996
rect 91112 521914 91140 522990
rect 81452 521886 81696 521914
rect 91112 521886 91356 521914
rect 71884 521206 72036 521234
rect 71884 500954 71912 521206
rect 91480 502738 91508 523058
rect 93124 523048 93176 523054
rect 93124 522990 93176 522996
rect 91356 502710 91508 502738
rect 72036 502030 72096 502058
rect 81696 502030 82032 502058
rect 71872 500948 71924 500954
rect 71872 500890 71924 500896
rect 72068 500818 72096 502030
rect 82004 500886 82032 502030
rect 93136 500886 93164 522990
rect 109696 521900 109724 523058
rect 119344 523048 119396 523054
rect 119344 522990 119396 522996
rect 119356 521900 119384 522990
rect 99484 521206 100050 521234
rect 93860 520328 93912 520334
rect 93860 520270 93912 520276
rect 97908 520328 97960 520334
rect 97908 520270 97960 520276
rect 93872 511601 93900 520270
rect 97920 512281 97948 520270
rect 97906 512272 97962 512281
rect 97906 512207 97962 512216
rect 93858 511592 93914 511601
rect 93858 511527 93914 511536
rect 99484 500886 99512 521206
rect 119448 502738 119476 523058
rect 124864 523048 124916 523054
rect 124864 522990 124916 522996
rect 121458 511592 121514 511601
rect 121458 511527 121514 511536
rect 121472 503674 121500 511527
rect 121460 503668 121512 503674
rect 121460 503610 121512 503616
rect 119370 502710 119476 502738
rect 100036 500954 100064 502044
rect 100024 500948 100076 500954
rect 100024 500890 100076 500896
rect 109696 500886 109724 502044
rect 124876 500886 124904 522990
rect 137664 521900 137692 523058
rect 147312 523048 147364 523054
rect 147312 522990 147364 522996
rect 148324 523048 148376 523054
rect 148324 522990 148376 522996
rect 147324 521900 147352 522990
rect 127084 521206 128018 521234
rect 126886 512272 126942 512281
rect 126886 512207 126942 512216
rect 126900 503674 126928 512207
rect 126888 503668 126940 503674
rect 126888 503610 126940 503616
rect 81992 500880 82044 500886
rect 81992 500822 82044 500828
rect 93124 500880 93176 500886
rect 93124 500822 93176 500828
rect 99472 500880 99524 500886
rect 99472 500822 99524 500828
rect 109684 500880 109736 500886
rect 109684 500822 109736 500828
rect 124864 500880 124916 500886
rect 124864 500822 124916 500828
rect 127084 500818 127112 521206
rect 147680 505640 147732 505646
rect 147680 505582 147732 505588
rect 147692 502738 147720 505582
rect 147338 502710 147720 502738
rect 128004 500954 128032 502044
rect 127992 500948 128044 500954
rect 127992 500890 128044 500896
rect 137664 500886 137692 502044
rect 148336 500886 148364 522990
rect 148428 505646 148456 523126
rect 149060 520328 149112 520334
rect 149060 520270 149112 520276
rect 149072 511601 149100 520270
rect 149058 511592 149114 511601
rect 149058 511527 149114 511536
rect 148416 505640 148468 505646
rect 148416 505582 148468 505588
rect 137652 500880 137704 500886
rect 137652 500822 137704 500828
rect 148324 500880 148376 500886
rect 148324 500822 148376 500828
rect 72056 500812 72108 500818
rect 72056 500754 72108 500760
rect 127072 500812 127124 500818
rect 127072 500754 127124 500760
rect 71136 497004 71188 497010
rect 71136 496946 71188 496952
rect 82268 497004 82320 497010
rect 82268 496946 82320 496952
rect 71148 473278 71176 496946
rect 72240 496936 72292 496942
rect 72240 496878 72292 496884
rect 72252 475674 72280 496878
rect 72608 496868 72660 496874
rect 72608 496810 72660 496816
rect 72620 494972 72648 496810
rect 82280 494972 82308 496946
rect 109960 496936 110012 496942
rect 109960 496878 110012 496884
rect 151084 496936 151136 496942
rect 151084 496878 151136 496884
rect 93124 496868 93176 496874
rect 93124 496810 93176 496816
rect 100300 496868 100352 496874
rect 100300 496810 100352 496816
rect 91954 494278 92152 494306
rect 72252 475646 72634 475674
rect 82280 473278 82308 475116
rect 91940 473346 91968 475116
rect 92124 473346 92152 494278
rect 91928 473340 91980 473346
rect 91928 473282 91980 473288
rect 92112 473340 92164 473346
rect 92112 473282 92164 473288
rect 93136 473278 93164 496810
rect 100208 496800 100260 496806
rect 100208 496742 100260 496748
rect 97906 485480 97962 485489
rect 97906 485415 97962 485424
rect 93858 484800 93914 484809
rect 93858 484735 93914 484744
rect 93872 475998 93900 484735
rect 97920 475998 97948 485415
rect 93860 475992 93912 475998
rect 93860 475934 93912 475940
rect 97908 475992 97960 475998
rect 97908 475934 97960 475940
rect 100220 475674 100248 496742
rect 100312 494986 100340 496810
rect 109972 494986 110000 496878
rect 138296 496868 138348 496874
rect 138296 496810 138348 496816
rect 149704 496868 149756 496874
rect 149704 496810 149756 496816
rect 100312 494958 100648 494986
rect 109972 494958 110308 494986
rect 138308 494972 138336 496810
rect 119968 494290 120212 494306
rect 128280 494290 128662 494306
rect 119968 494284 120224 494290
rect 119968 494278 120172 494284
rect 120172 494226 120224 494232
rect 122104 494284 122156 494290
rect 122104 494226 122156 494232
rect 124864 494284 124916 494290
rect 124864 494226 124916 494232
rect 128268 494284 128662 494290
rect 128320 494278 128662 494284
rect 147982 494278 148088 494306
rect 128268 494226 128320 494232
rect 121458 484800 121514 484809
rect 121458 484735 121514 484744
rect 121472 476066 121500 484735
rect 121460 476060 121512 476066
rect 121460 476002 121512 476008
rect 100220 475646 100648 475674
rect 110248 475102 110308 475130
rect 119632 475102 119968 475130
rect 110248 473278 110276 475102
rect 119632 473346 119660 475102
rect 122116 473346 122144 494226
rect 119620 473340 119672 473346
rect 119620 473282 119672 473288
rect 122104 473340 122156 473346
rect 122104 473282 122156 473288
rect 124876 473278 124904 494226
rect 126886 485480 126942 485489
rect 126886 485415 126942 485424
rect 126900 476066 126928 485415
rect 126888 476060 126940 476066
rect 126888 476002 126940 476008
rect 128648 473278 128676 475116
rect 71136 473272 71188 473278
rect 71136 473214 71188 473220
rect 82268 473272 82320 473278
rect 82268 473214 82320 473220
rect 93124 473272 93176 473278
rect 93124 473214 93176 473220
rect 110236 473272 110288 473278
rect 110236 473214 110288 473220
rect 124864 473272 124916 473278
rect 124864 473214 124916 473220
rect 128636 473272 128688 473278
rect 128636 473214 128688 473220
rect 138308 473210 138336 475116
rect 147968 473346 147996 475116
rect 148060 473346 148088 494278
rect 149058 484800 149114 484809
rect 149058 484735 149114 484744
rect 149072 475998 149100 484735
rect 149060 475992 149112 475998
rect 149060 475934 149112 475940
rect 147956 473340 148008 473346
rect 147956 473282 148008 473288
rect 148048 473340 148100 473346
rect 148048 473282 148100 473288
rect 149716 473278 149744 496810
rect 149704 473272 149756 473278
rect 149704 473214 149756 473220
rect 151096 473210 151124 496878
rect 138296 473204 138348 473210
rect 138296 473146 138348 473152
rect 151084 473204 151136 473210
rect 151084 473146 151136 473152
rect 148324 469396 148376 469402
rect 148324 469338 148376 469344
rect 81440 469328 81492 469334
rect 81440 469270 81492 469276
rect 91468 469328 91520 469334
rect 91468 469270 91520 469276
rect 109684 469328 109736 469334
rect 109684 469270 109736 469276
rect 119436 469328 119488 469334
rect 119436 469270 119488 469276
rect 137652 469328 137704 469334
rect 137652 469270 137704 469276
rect 81452 467922 81480 469270
rect 91100 469260 91152 469266
rect 91100 469202 91152 469208
rect 91112 467922 91140 469202
rect 81452 467894 81696 467922
rect 91112 467894 91356 467922
rect 71884 467214 72036 467242
rect 71884 445738 71912 467214
rect 91480 448746 91508 469270
rect 93124 469260 93176 469266
rect 93124 469202 93176 469208
rect 91356 448718 91508 448746
rect 72036 448038 72096 448066
rect 81696 448038 82032 448066
rect 71872 445732 71924 445738
rect 71872 445674 71924 445680
rect 72068 445602 72096 448038
rect 82004 445670 82032 448038
rect 93136 445670 93164 469202
rect 109696 467908 109724 469270
rect 119344 469260 119396 469266
rect 119344 469202 119396 469208
rect 119356 467908 119384 469202
rect 99484 467214 100050 467242
rect 93860 466540 93912 466546
rect 93860 466482 93912 466488
rect 97908 466540 97960 466546
rect 97908 466482 97960 466488
rect 93872 457609 93900 466482
rect 97920 458289 97948 466482
rect 97906 458280 97962 458289
rect 97906 458215 97962 458224
rect 93858 457600 93914 457609
rect 93858 457535 93914 457544
rect 99484 445670 99512 467214
rect 119448 448746 119476 469270
rect 124864 469260 124916 469266
rect 124864 469202 124916 469208
rect 121460 466472 121512 466478
rect 121460 466414 121512 466420
rect 121472 457609 121500 466414
rect 121458 457600 121514 457609
rect 121458 457535 121514 457544
rect 119370 448718 119476 448746
rect 100036 445738 100064 448052
rect 100024 445732 100076 445738
rect 100024 445674 100076 445680
rect 109696 445670 109724 448052
rect 124876 445670 124904 469202
rect 137664 467908 137692 469270
rect 147312 469260 147364 469266
rect 147312 469202 147364 469208
rect 147324 467908 147352 469202
rect 127084 467214 128018 467242
rect 126888 466472 126940 466478
rect 126888 466414 126940 466420
rect 126900 458289 126928 466414
rect 126886 458280 126942 458289
rect 126886 458215 126942 458224
rect 81992 445664 82044 445670
rect 81992 445606 82044 445612
rect 93124 445664 93176 445670
rect 93124 445606 93176 445612
rect 99472 445664 99524 445670
rect 99472 445606 99524 445612
rect 109684 445664 109736 445670
rect 109684 445606 109736 445612
rect 124864 445664 124916 445670
rect 124864 445606 124916 445612
rect 127084 445602 127112 467214
rect 148336 451274 148364 469338
rect 148416 469260 148468 469266
rect 148416 469202 148468 469208
rect 147784 451246 148364 451274
rect 147784 448474 147812 451246
rect 147338 448446 147812 448474
rect 128004 445738 128032 448052
rect 127992 445732 128044 445738
rect 127992 445674 128044 445680
rect 137664 445670 137692 448052
rect 148428 445670 148456 469202
rect 149060 466540 149112 466546
rect 149060 466482 149112 466488
rect 149072 457609 149100 466482
rect 149058 457600 149114 457609
rect 149058 457535 149114 457544
rect 137652 445664 137704 445670
rect 137652 445606 137704 445612
rect 148416 445664 148468 445670
rect 148416 445606 148468 445612
rect 72056 445596 72108 445602
rect 72056 445538 72108 445544
rect 127072 445596 127124 445602
rect 127072 445538 127124 445544
rect 71136 443148 71188 443154
rect 71136 443090 71188 443096
rect 82268 443148 82320 443154
rect 82268 443090 82320 443096
rect 99380 443148 99432 443154
rect 99380 443090 99432 443096
rect 100300 443148 100352 443154
rect 100300 443090 100352 443096
rect 71148 419422 71176 443090
rect 71872 443080 71924 443086
rect 71872 443022 71924 443028
rect 71884 441614 71912 443022
rect 72608 443012 72660 443018
rect 72608 442954 72660 442960
rect 71884 441586 72280 441614
rect 72252 421682 72280 441586
rect 72620 440980 72648 442954
rect 82280 440980 82308 443090
rect 99392 443018 99420 443090
rect 93124 443012 93176 443018
rect 93124 442954 93176 442960
rect 99380 443012 99432 443018
rect 99380 442954 99432 442960
rect 99472 443012 99524 443018
rect 99472 442954 99524 442960
rect 91954 440286 92152 440314
rect 72252 421654 72634 421682
rect 82280 419422 82308 421124
rect 91940 419490 91968 421124
rect 92124 419490 92152 440286
rect 91928 419484 91980 419490
rect 91928 419426 91980 419432
rect 92112 419484 92164 419490
rect 92112 419426 92164 419432
rect 93136 419422 93164 442954
rect 99484 441614 99512 442954
rect 99484 441586 100248 441614
rect 93860 440292 93912 440298
rect 93860 440234 93912 440240
rect 97908 440292 97960 440298
rect 97908 440234 97960 440240
rect 93872 430817 93900 440234
rect 97920 431497 97948 440234
rect 97906 431488 97962 431497
rect 97906 431423 97962 431432
rect 93858 430808 93914 430817
rect 93858 430743 93914 430752
rect 100220 421682 100248 441586
rect 100312 440994 100340 443090
rect 109960 443080 110012 443086
rect 109960 443022 110012 443028
rect 124864 443080 124916 443086
rect 124864 443022 124916 443028
rect 128360 443080 128412 443086
rect 128360 443022 128412 443028
rect 151084 443080 151136 443086
rect 151084 443022 151136 443028
rect 109972 440994 110000 443022
rect 100312 440966 100648 440994
rect 109972 440966 110308 440994
rect 119968 440286 120304 440314
rect 120276 440230 120304 440286
rect 120264 440224 120316 440230
rect 120264 440166 120316 440172
rect 122104 440224 122156 440230
rect 122104 440166 122156 440172
rect 121458 430808 121514 430817
rect 121458 430743 121514 430752
rect 121472 422278 121500 430743
rect 121460 422272 121512 422278
rect 121460 422214 121512 422220
rect 100220 421654 100648 421682
rect 110248 421110 110308 421138
rect 119632 421110 119968 421138
rect 110248 419422 110276 421110
rect 119632 419490 119660 421110
rect 122116 419490 122144 440166
rect 119620 419484 119672 419490
rect 119620 419426 119672 419432
rect 122104 419484 122156 419490
rect 122104 419426 122156 419432
rect 124876 419422 124904 443022
rect 128372 440994 128400 443022
rect 138020 443012 138072 443018
rect 138020 442954 138072 442960
rect 149704 443012 149756 443018
rect 149704 442954 149756 442960
rect 138032 440994 138060 442954
rect 128372 440966 128662 440994
rect 138032 440966 138322 440994
rect 147982 440286 148088 440314
rect 126886 431488 126942 431497
rect 126886 431423 126942 431432
rect 126900 422278 126928 431423
rect 126888 422272 126940 422278
rect 126888 422214 126940 422220
rect 128648 419422 128676 421124
rect 71136 419416 71188 419422
rect 71136 419358 71188 419364
rect 82268 419416 82320 419422
rect 82268 419358 82320 419364
rect 93124 419416 93176 419422
rect 93124 419358 93176 419364
rect 110236 419416 110288 419422
rect 110236 419358 110288 419364
rect 124864 419416 124916 419422
rect 124864 419358 124916 419364
rect 128636 419416 128688 419422
rect 128636 419358 128688 419364
rect 138308 419354 138336 421124
rect 147968 419490 147996 421124
rect 148060 419490 148088 440286
rect 149060 440292 149112 440298
rect 149060 440234 149112 440240
rect 149072 430817 149100 440234
rect 149058 430808 149114 430817
rect 149058 430743 149114 430752
rect 147956 419484 148008 419490
rect 147956 419426 148008 419432
rect 148048 419484 148100 419490
rect 148048 419426 148100 419432
rect 149716 419422 149744 442954
rect 149704 419416 149756 419422
rect 149704 419358 149756 419364
rect 151096 419354 151124 443022
rect 138296 419348 138348 419354
rect 138296 419290 138348 419296
rect 151084 419348 151136 419354
rect 151084 419290 151136 419296
rect 119436 415608 119488 415614
rect 119436 415550 119488 415556
rect 137652 415608 137704 415614
rect 137652 415550 137704 415556
rect 148324 415608 148376 415614
rect 148324 415550 148376 415556
rect 81440 415540 81492 415546
rect 81440 415482 81492 415488
rect 91468 415540 91520 415546
rect 91468 415482 91520 415488
rect 109684 415540 109736 415546
rect 109684 415482 109736 415488
rect 81452 413930 81480 415482
rect 91100 415472 91152 415478
rect 91100 415414 91152 415420
rect 91112 413930 91140 415414
rect 81452 413902 81696 413930
rect 91112 413902 91356 413930
rect 71884 413222 72036 413250
rect 71884 391950 71912 413222
rect 91480 394754 91508 415482
rect 93124 415472 93176 415478
rect 93124 415414 93176 415420
rect 91356 394726 91508 394754
rect 72022 393802 72050 394060
rect 81696 394046 82032 394074
rect 71976 393774 72050 393802
rect 71872 391944 71924 391950
rect 71872 391886 71924 391892
rect 71976 391814 72004 393774
rect 82004 391882 82032 394046
rect 93136 391882 93164 415414
rect 109696 413916 109724 415482
rect 119344 415472 119396 415478
rect 119344 415414 119396 415420
rect 119356 413916 119384 415414
rect 99484 413222 100050 413250
rect 97906 404288 97962 404297
rect 97906 404223 97962 404232
rect 93858 403608 93914 403617
rect 93858 403543 93914 403552
rect 93872 394602 93900 403543
rect 97920 394602 97948 404223
rect 93860 394596 93912 394602
rect 93860 394538 93912 394544
rect 97908 394596 97960 394602
rect 97908 394538 97960 394544
rect 99484 391882 99512 413222
rect 119448 394754 119476 415550
rect 127992 415540 128044 415546
rect 127992 415482 128044 415488
rect 122104 415472 122156 415478
rect 122104 415414 122156 415420
rect 121458 403608 121514 403617
rect 121458 403543 121514 403552
rect 119370 394726 119476 394754
rect 121472 394670 121500 403543
rect 121460 394664 121512 394670
rect 121460 394606 121512 394612
rect 100036 391950 100064 394060
rect 100024 391944 100076 391950
rect 100024 391886 100076 391892
rect 109696 391882 109724 394060
rect 122116 391882 122144 415414
rect 128004 413916 128032 415482
rect 137664 413916 137692 415550
rect 147312 415472 147364 415478
rect 147312 415414 147364 415420
rect 147324 413916 147352 415414
rect 126886 404288 126942 404297
rect 126886 404223 126942 404232
rect 126900 394670 126928 404223
rect 148336 402974 148364 415550
rect 148508 415540 148560 415546
rect 148508 415482 148560 415488
rect 148416 415472 148468 415478
rect 148416 415414 148468 415420
rect 147784 402946 148364 402974
rect 126888 394664 126940 394670
rect 147784 394618 147812 402946
rect 126888 394606 126940 394612
rect 147338 394590 147812 394618
rect 128004 391950 128032 394060
rect 127992 391944 128044 391950
rect 127992 391886 128044 391892
rect 137664 391882 137692 394060
rect 148428 391882 148456 415414
rect 148520 395350 148548 415482
rect 149058 403608 149114 403617
rect 149058 403543 149114 403552
rect 148508 395344 148560 395350
rect 148508 395286 148560 395292
rect 149072 394602 149100 403543
rect 149060 394596 149112 394602
rect 149060 394538 149112 394544
rect 81992 391876 82044 391882
rect 81992 391818 82044 391824
rect 93124 391876 93176 391882
rect 93124 391818 93176 391824
rect 99472 391876 99524 391882
rect 99472 391818 99524 391824
rect 109684 391876 109736 391882
rect 109684 391818 109736 391824
rect 122104 391876 122156 391882
rect 122104 391818 122156 391824
rect 137652 391876 137704 391882
rect 137652 391818 137704 391824
rect 148416 391876 148468 391882
rect 148416 391818 148468 391824
rect 71964 391808 72016 391814
rect 71964 391750 72016 391756
rect 71136 389360 71188 389366
rect 71136 389302 71188 389308
rect 82268 389360 82320 389366
rect 82268 389302 82320 389308
rect 99472 389360 99524 389366
rect 99472 389302 99524 389308
rect 100392 389360 100444 389366
rect 100392 389302 100444 389308
rect 71148 365634 71176 389302
rect 71872 389292 71924 389298
rect 71872 389234 71924 389240
rect 71884 383654 71912 389234
rect 72608 389224 72660 389230
rect 72608 389166 72660 389172
rect 72620 386852 72648 389166
rect 82280 386852 82308 389302
rect 93124 389224 93176 389230
rect 93124 389166 93176 389172
rect 91954 386294 92152 386322
rect 71884 383626 72280 383654
rect 72252 367690 72280 383626
rect 72252 367662 72634 367690
rect 82280 365634 82308 367132
rect 91940 365702 91968 367132
rect 92124 365702 92152 386294
rect 91928 365696 91980 365702
rect 91928 365638 91980 365644
rect 92112 365696 92164 365702
rect 92112 365638 92164 365644
rect 93136 365634 93164 389166
rect 93860 386504 93912 386510
rect 93860 386446 93912 386452
rect 97908 386504 97960 386510
rect 97908 386446 97960 386452
rect 93872 376825 93900 386446
rect 97920 377505 97948 386446
rect 99484 383654 99512 389302
rect 100404 389230 100432 389302
rect 109960 389292 110012 389298
rect 109960 389234 110012 389240
rect 151084 389292 151136 389298
rect 151084 389234 151136 389240
rect 100300 389224 100352 389230
rect 100300 389166 100352 389172
rect 100392 389224 100444 389230
rect 100392 389166 100444 389172
rect 100312 386866 100340 389166
rect 109972 386866 110000 389234
rect 138296 389224 138348 389230
rect 138296 389166 138348 389172
rect 149704 389224 149756 389230
rect 149704 389166 149756 389172
rect 100312 386838 100648 386866
rect 109972 386838 110308 386866
rect 138308 386852 138336 389166
rect 126888 386572 126940 386578
rect 126888 386514 126940 386520
rect 121460 386436 121512 386442
rect 121460 386378 121512 386384
rect 124864 386436 124916 386442
rect 124864 386378 124916 386384
rect 119968 386306 120304 386322
rect 119968 386300 120316 386306
rect 119968 386294 120264 386300
rect 120264 386242 120316 386248
rect 99484 383626 100248 383654
rect 97906 377496 97962 377505
rect 97906 377431 97962 377440
rect 93858 376816 93914 376825
rect 93858 376751 93914 376760
rect 100220 367690 100248 383626
rect 121472 376825 121500 386378
rect 122104 386300 122156 386306
rect 122104 386242 122156 386248
rect 121458 376816 121514 376825
rect 121458 376751 121514 376760
rect 100220 367662 100648 367690
rect 110248 367118 110308 367146
rect 119632 367118 119968 367146
rect 110248 365634 110276 367118
rect 119632 365702 119660 367118
rect 122116 365702 122144 386242
rect 119620 365696 119672 365702
rect 119620 365638 119672 365644
rect 122104 365696 122156 365702
rect 122104 365638 122156 365644
rect 124876 365634 124904 386378
rect 126900 377505 126928 386514
rect 149060 386504 149112 386510
rect 128280 386442 128662 386458
rect 149060 386446 149112 386452
rect 128268 386436 128662 386442
rect 128320 386430 128662 386436
rect 128268 386378 128320 386384
rect 147982 386294 148088 386322
rect 126886 377496 126942 377505
rect 126886 377431 126942 377440
rect 128648 365634 128676 367132
rect 71136 365628 71188 365634
rect 71136 365570 71188 365576
rect 82268 365628 82320 365634
rect 82268 365570 82320 365576
rect 93124 365628 93176 365634
rect 93124 365570 93176 365576
rect 110236 365628 110288 365634
rect 110236 365570 110288 365576
rect 124864 365628 124916 365634
rect 124864 365570 124916 365576
rect 128636 365628 128688 365634
rect 128636 365570 128688 365576
rect 138308 365566 138336 367132
rect 147968 365702 147996 367132
rect 148060 365702 148088 386294
rect 149072 376825 149100 386446
rect 149058 376816 149114 376825
rect 149058 376751 149114 376760
rect 147956 365696 148008 365702
rect 147956 365638 148008 365644
rect 148048 365696 148100 365702
rect 148048 365638 148100 365644
rect 149716 365634 149744 389166
rect 149704 365628 149756 365634
rect 149704 365570 149756 365576
rect 151096 365566 151124 389234
rect 138296 365560 138348 365566
rect 138296 365502 138348 365508
rect 151084 365560 151136 365566
rect 151084 365502 151136 365508
rect 148416 361752 148468 361758
rect 148416 361694 148468 361700
rect 81440 361684 81492 361690
rect 81440 361626 81492 361632
rect 119436 361684 119488 361690
rect 119436 361626 119488 361632
rect 137652 361684 137704 361690
rect 137652 361626 137704 361632
rect 81452 359938 81480 361626
rect 91100 361616 91152 361622
rect 91100 361558 91152 361564
rect 93124 361616 93176 361622
rect 93124 361558 93176 361564
rect 119344 361616 119396 361622
rect 119344 361558 119396 361564
rect 91112 359938 91140 361558
rect 81452 359910 81696 359938
rect 91112 359910 91356 359938
rect 71884 359230 72036 359258
rect 71884 338094 71912 359230
rect 91468 358828 91520 358834
rect 91468 358770 91520 358776
rect 91480 340762 91508 358770
rect 91356 340734 91508 340762
rect 72036 340054 72096 340082
rect 81696 340054 82032 340082
rect 71872 338088 71924 338094
rect 71872 338030 71924 338036
rect 72068 337958 72096 340054
rect 82004 338026 82032 340054
rect 93136 338026 93164 361558
rect 119356 359924 119384 361558
rect 109316 359304 109368 359310
rect 99484 359230 100050 359258
rect 109368 359252 109710 359258
rect 109316 359246 109710 359252
rect 109328 359230 109710 359246
rect 97906 350296 97962 350305
rect 97906 350231 97962 350240
rect 93858 349616 93914 349625
rect 93858 349551 93914 349560
rect 93872 340814 93900 349551
rect 97920 340814 97948 350231
rect 93860 340808 93912 340814
rect 93860 340750 93912 340756
rect 97908 340808 97960 340814
rect 97908 340750 97960 340756
rect 99484 338026 99512 359230
rect 119448 340762 119476 361626
rect 122104 361616 122156 361622
rect 122104 361558 122156 361564
rect 121458 349616 121514 349625
rect 121458 349551 121514 349560
rect 121472 340882 121500 349551
rect 121460 340876 121512 340882
rect 121460 340818 121512 340824
rect 119370 340734 119476 340762
rect 100036 338094 100064 340068
rect 100024 338088 100076 338094
rect 100024 338030 100076 338036
rect 109696 338026 109724 340068
rect 122116 338026 122144 361558
rect 137664 359924 137692 361626
rect 147312 361616 147364 361622
rect 147312 361558 147364 361564
rect 148324 361616 148376 361622
rect 148324 361558 148376 361564
rect 147324 359924 147352 361558
rect 127084 359230 128018 359258
rect 126886 350296 126942 350305
rect 126886 350231 126942 350240
rect 126900 340882 126928 350231
rect 126888 340876 126940 340882
rect 126888 340818 126940 340824
rect 81992 338020 82044 338026
rect 81992 337962 82044 337968
rect 93124 338020 93176 338026
rect 93124 337962 93176 337968
rect 99472 338020 99524 338026
rect 99472 337962 99524 337968
rect 109684 338020 109736 338026
rect 109684 337962 109736 337968
rect 122104 338020 122156 338026
rect 122104 337962 122156 337968
rect 127084 337958 127112 359230
rect 147680 342576 147732 342582
rect 147680 342518 147732 342524
rect 147692 340762 147720 342518
rect 147338 340734 147720 340762
rect 128004 338094 128032 340068
rect 127992 338088 128044 338094
rect 127992 338030 128044 338036
rect 137664 338026 137692 340068
rect 148336 338026 148364 361558
rect 148428 342582 148456 361694
rect 149058 349616 149114 349625
rect 149058 349551 149114 349560
rect 148416 342576 148468 342582
rect 148416 342518 148468 342524
rect 149072 340814 149100 349551
rect 149060 340808 149112 340814
rect 149060 340750 149112 340756
rect 137652 338020 137704 338026
rect 137652 337962 137704 337968
rect 148324 338020 148376 338026
rect 148324 337962 148376 337968
rect 72056 337952 72108 337958
rect 72056 337894 72108 337900
rect 127072 337952 127124 337958
rect 127072 337894 127124 337900
rect 71136 335504 71188 335510
rect 71136 335446 71188 335452
rect 82268 335504 82320 335510
rect 82268 335446 82320 335452
rect 99380 335504 99432 335510
rect 99380 335446 99432 335452
rect 100300 335504 100352 335510
rect 100300 335446 100352 335452
rect 71148 311778 71176 335446
rect 71872 335436 71924 335442
rect 71872 335378 71924 335384
rect 71884 325694 71912 335378
rect 72608 335368 72660 335374
rect 72608 335310 72660 335316
rect 72620 332860 72648 335310
rect 82280 332860 82308 335446
rect 99392 335374 99420 335446
rect 93124 335368 93176 335374
rect 93124 335310 93176 335316
rect 99380 335368 99432 335374
rect 99380 335310 99432 335316
rect 99472 335368 99524 335374
rect 99472 335310 99524 335316
rect 91954 332302 92152 332330
rect 71884 325666 72280 325694
rect 72252 313698 72280 325666
rect 72252 313670 72634 313698
rect 82280 311778 82308 313140
rect 91940 311846 91968 313140
rect 92124 311846 92152 332302
rect 91928 311840 91980 311846
rect 91928 311782 91980 311788
rect 92112 311840 92164 311846
rect 92112 311782 92164 311788
rect 93136 311778 93164 335310
rect 99484 325694 99512 335310
rect 100312 332874 100340 335446
rect 109960 335436 110012 335442
rect 109960 335378 110012 335384
rect 124864 335436 124916 335442
rect 124864 335378 124916 335384
rect 128636 335436 128688 335442
rect 128636 335378 128688 335384
rect 151084 335436 151136 335442
rect 151084 335378 151136 335384
rect 109972 332874 110000 335378
rect 100312 332846 100648 332874
rect 109972 332846 110308 332874
rect 119968 332314 120212 332330
rect 119968 332308 120224 332314
rect 119968 332302 120172 332308
rect 120172 332250 120224 332256
rect 122104 332308 122156 332314
rect 122104 332250 122156 332256
rect 99484 325666 100248 325694
rect 97906 322960 97962 322969
rect 97906 322895 97962 322904
rect 93858 322144 93914 322153
rect 93858 322079 93914 322088
rect 93872 314566 93900 322079
rect 97920 314566 97948 322895
rect 93860 314560 93912 314566
rect 93860 314502 93912 314508
rect 97908 314560 97960 314566
rect 97908 314502 97960 314508
rect 100220 313698 100248 325666
rect 121458 322144 121514 322153
rect 121458 322079 121514 322088
rect 121472 314634 121500 322079
rect 121460 314628 121512 314634
rect 121460 314570 121512 314576
rect 100220 313670 100648 313698
rect 110248 313126 110308 313154
rect 119632 313126 119968 313154
rect 110248 311778 110276 313126
rect 119632 311846 119660 313126
rect 122116 311846 122144 332250
rect 119620 311840 119672 311846
rect 119620 311782 119672 311788
rect 122104 311840 122156 311846
rect 122104 311782 122156 311788
rect 124876 311778 124904 335378
rect 128648 332860 128676 335378
rect 138296 335368 138348 335374
rect 138296 335310 138348 335316
rect 149704 335368 149756 335374
rect 149704 335310 149756 335316
rect 138308 332860 138336 335310
rect 147982 332302 148088 332330
rect 126886 322960 126942 322969
rect 126886 322895 126942 322904
rect 126900 314634 126928 322895
rect 126888 314628 126940 314634
rect 126888 314570 126940 314576
rect 128648 311778 128676 313140
rect 71136 311772 71188 311778
rect 71136 311714 71188 311720
rect 82268 311772 82320 311778
rect 82268 311714 82320 311720
rect 93124 311772 93176 311778
rect 93124 311714 93176 311720
rect 110236 311772 110288 311778
rect 110236 311714 110288 311720
rect 124864 311772 124916 311778
rect 124864 311714 124916 311720
rect 128636 311772 128688 311778
rect 128636 311714 128688 311720
rect 138308 311710 138336 313140
rect 147968 311846 147996 313140
rect 148060 311846 148088 332302
rect 149058 322144 149114 322153
rect 149058 322079 149114 322088
rect 149072 314566 149100 322079
rect 149060 314560 149112 314566
rect 149060 314502 149112 314508
rect 147956 311840 148008 311846
rect 147956 311782 148008 311788
rect 148048 311840 148100 311846
rect 148048 311782 148100 311788
rect 149716 311778 149744 335310
rect 149704 311772 149756 311778
rect 149704 311714 149756 311720
rect 151096 311710 151124 335378
rect 138296 311704 138348 311710
rect 138296 311646 138348 311652
rect 151084 311704 151136 311710
rect 151084 311646 151136 311652
rect 148324 307964 148376 307970
rect 148324 307906 148376 307912
rect 81440 307896 81492 307902
rect 81440 307838 81492 307844
rect 91468 307896 91520 307902
rect 91468 307838 91520 307844
rect 109684 307896 109736 307902
rect 109684 307838 109736 307844
rect 119436 307896 119488 307902
rect 119436 307838 119488 307844
rect 137652 307896 137704 307902
rect 137652 307838 137704 307844
rect 81452 305946 81480 307838
rect 91100 307828 91152 307834
rect 91100 307770 91152 307776
rect 91112 305946 91140 307770
rect 81452 305918 81696 305946
rect 91112 305918 91356 305946
rect 71884 305238 72036 305266
rect 71884 284306 71912 305238
rect 91480 286770 91508 307838
rect 93124 307828 93176 307834
rect 93124 307770 93176 307776
rect 91356 286742 91508 286770
rect 72036 286062 72096 286090
rect 81696 286062 82032 286090
rect 71872 284300 71924 284306
rect 71872 284242 71924 284248
rect 72068 284170 72096 286062
rect 82004 284238 82032 286062
rect 93136 284238 93164 307770
rect 109696 305932 109724 307838
rect 119344 307828 119396 307834
rect 119344 307770 119396 307776
rect 119356 305932 119384 307770
rect 99484 305238 100050 305266
rect 97906 296304 97962 296313
rect 97906 296239 97962 296248
rect 93858 295624 93914 295633
rect 93858 295559 93914 295568
rect 93872 286958 93900 295559
rect 97920 286958 97948 296239
rect 93860 286952 93912 286958
rect 93860 286894 93912 286900
rect 97908 286952 97960 286958
rect 97908 286894 97960 286900
rect 99484 284238 99512 305238
rect 119448 286770 119476 307838
rect 122104 307828 122156 307834
rect 122104 307770 122156 307776
rect 121458 295624 121514 295633
rect 121458 295559 121514 295568
rect 121472 287026 121500 295559
rect 121460 287020 121512 287026
rect 121460 286962 121512 286968
rect 119370 286742 119476 286770
rect 100036 284306 100064 286076
rect 100024 284300 100076 284306
rect 100024 284242 100076 284248
rect 109696 284238 109724 286076
rect 122116 284238 122144 307770
rect 137664 305932 137692 307838
rect 147312 307828 147364 307834
rect 147312 307770 147364 307776
rect 147324 305932 147352 307770
rect 127084 305238 128018 305266
rect 126886 296304 126942 296313
rect 126886 296239 126942 296248
rect 126900 286890 126928 296239
rect 126888 286884 126940 286890
rect 126888 286826 126940 286832
rect 81992 284232 82044 284238
rect 81992 284174 82044 284180
rect 93124 284232 93176 284238
rect 93124 284174 93176 284180
rect 99472 284232 99524 284238
rect 99472 284174 99524 284180
rect 109684 284232 109736 284238
rect 109684 284174 109736 284180
rect 122104 284232 122156 284238
rect 122104 284174 122156 284180
rect 127084 284170 127112 305238
rect 148336 287054 148364 307906
rect 148416 307828 148468 307834
rect 148416 307770 148468 307776
rect 147784 287026 148364 287054
rect 147784 286770 147812 287026
rect 147338 286742 147812 286770
rect 128004 284306 128032 286076
rect 127992 284300 128044 284306
rect 127992 284242 128044 284248
rect 137664 284238 137692 286076
rect 148428 284238 148456 307770
rect 149058 295624 149114 295633
rect 149058 295559 149114 295568
rect 149072 286958 149100 295559
rect 149060 286952 149112 286958
rect 149060 286894 149112 286900
rect 137652 284232 137704 284238
rect 137652 284174 137704 284180
rect 148416 284232 148468 284238
rect 148416 284174 148468 284180
rect 72056 284164 72108 284170
rect 72056 284106 72108 284112
rect 127072 284164 127124 284170
rect 127072 284106 127124 284112
rect 71872 280424 71924 280430
rect 71872 280366 71924 280372
rect 71136 280356 71188 280362
rect 71136 280298 71188 280304
rect 71148 256630 71176 280298
rect 71884 267734 71912 280366
rect 99472 280356 99524 280362
rect 99472 280298 99524 280304
rect 100392 280356 100444 280362
rect 100392 280298 100444 280304
rect 72608 280220 72660 280226
rect 72608 280162 72660 280168
rect 82268 280220 82320 280226
rect 82268 280162 82320 280168
rect 93124 280220 93176 280226
rect 93124 280162 93176 280168
rect 72620 278868 72648 280162
rect 82280 278868 82308 280162
rect 91954 278310 92152 278338
rect 71884 267706 72280 267734
rect 72252 259706 72280 267706
rect 72252 259678 72634 259706
rect 82280 256630 82308 259148
rect 91940 256698 91968 259148
rect 92124 256698 92152 278310
rect 91928 256692 91980 256698
rect 91928 256634 91980 256640
rect 92112 256692 92164 256698
rect 92112 256634 92164 256640
rect 93136 256630 93164 280162
rect 93860 277500 93912 277506
rect 93860 277442 93912 277448
rect 97908 277500 97960 277506
rect 97908 277442 97960 277448
rect 93872 269113 93900 277442
rect 97920 270065 97948 277442
rect 97906 270056 97962 270065
rect 97906 269991 97962 270000
rect 93858 269104 93914 269113
rect 93858 269039 93914 269048
rect 99484 267734 99512 280298
rect 100404 280226 100432 280298
rect 109960 280288 110012 280294
rect 109960 280230 110012 280236
rect 124864 280288 124916 280294
rect 124864 280230 124916 280236
rect 128636 280288 128688 280294
rect 128636 280230 128688 280236
rect 151084 280288 151136 280294
rect 151084 280230 151136 280236
rect 100300 280220 100352 280226
rect 100300 280162 100352 280168
rect 100392 280220 100444 280226
rect 100392 280162 100444 280168
rect 100312 278882 100340 280162
rect 109972 278882 110000 280230
rect 100312 278854 100648 278882
rect 109972 278854 110308 278882
rect 119968 278322 120212 278338
rect 119968 278316 120224 278322
rect 119968 278310 120172 278316
rect 120172 278258 120224 278264
rect 122104 278316 122156 278322
rect 122104 278258 122156 278264
rect 121460 277432 121512 277438
rect 121460 277374 121512 277380
rect 121472 269113 121500 277374
rect 121458 269104 121514 269113
rect 121458 269039 121514 269048
rect 99484 267706 100248 267734
rect 100220 259706 100248 267706
rect 100220 259678 100648 259706
rect 110294 258890 110322 259148
rect 119632 259134 119968 259162
rect 110294 258862 110368 258890
rect 110340 256630 110368 258862
rect 119632 256698 119660 259134
rect 122116 256698 122144 278258
rect 119620 256692 119672 256698
rect 119620 256634 119672 256640
rect 122104 256692 122156 256698
rect 122104 256634 122156 256640
rect 124876 256630 124904 280230
rect 128648 278868 128676 280230
rect 138296 280220 138348 280226
rect 138296 280162 138348 280168
rect 149704 280220 149756 280226
rect 149704 280162 149756 280168
rect 138308 278868 138336 280162
rect 147982 278310 148088 278338
rect 126888 277568 126940 277574
rect 126888 277510 126940 277516
rect 126900 270065 126928 277510
rect 126886 270056 126942 270065
rect 126886 269991 126942 270000
rect 128648 256630 128676 259148
rect 71136 256624 71188 256630
rect 71136 256566 71188 256572
rect 82268 256624 82320 256630
rect 82268 256566 82320 256572
rect 93124 256624 93176 256630
rect 93124 256566 93176 256572
rect 110328 256624 110380 256630
rect 110328 256566 110380 256572
rect 124864 256624 124916 256630
rect 124864 256566 124916 256572
rect 128636 256624 128688 256630
rect 128636 256566 128688 256572
rect 138308 256562 138336 259148
rect 147968 256698 147996 259148
rect 148060 256698 148088 278310
rect 149060 277500 149112 277506
rect 149060 277442 149112 277448
rect 149072 269113 149100 277442
rect 149058 269104 149114 269113
rect 149058 269039 149114 269048
rect 147956 256692 148008 256698
rect 147956 256634 148008 256640
rect 148048 256692 148100 256698
rect 148048 256634 148100 256640
rect 149716 256630 149744 280162
rect 149704 256624 149756 256630
rect 149704 256566 149756 256572
rect 151096 256562 151124 280230
rect 138296 256556 138348 256562
rect 138296 256498 138348 256504
rect 151084 256556 151136 256562
rect 151084 256498 151136 256504
rect 148416 254108 148468 254114
rect 148416 254050 148468 254056
rect 81440 254040 81492 254046
rect 81440 253982 81492 253988
rect 91468 254040 91520 254046
rect 91468 253982 91520 253988
rect 109684 254040 109736 254046
rect 109684 253982 109736 253988
rect 119436 254040 119488 254046
rect 119436 253982 119488 253988
rect 137652 254040 137704 254046
rect 137652 253982 137704 253988
rect 81452 251954 81480 253982
rect 91100 253972 91152 253978
rect 91100 253914 91152 253920
rect 91112 251954 91140 253914
rect 81452 251926 81696 251954
rect 91112 251926 91356 251954
rect 71884 251246 72036 251274
rect 71884 230450 71912 251246
rect 91480 232778 91508 253982
rect 93124 253972 93176 253978
rect 93124 253914 93176 253920
rect 91356 232750 91508 232778
rect 72036 232070 72096 232098
rect 81696 232070 82032 232098
rect 71872 230444 71924 230450
rect 71872 230386 71924 230392
rect 72068 230314 72096 232070
rect 82004 230382 82032 232070
rect 93136 230382 93164 253914
rect 109696 251940 109724 253982
rect 119344 253972 119396 253978
rect 119344 253914 119396 253920
rect 119356 251940 119384 253914
rect 93860 251252 93912 251258
rect 93860 251194 93912 251200
rect 97908 251252 97960 251258
rect 97908 251194 97960 251200
rect 99484 251246 100050 251274
rect 93872 241641 93900 251194
rect 97920 242321 97948 251194
rect 97906 242312 97962 242321
rect 97906 242247 97962 242256
rect 93858 241632 93914 241641
rect 93858 241567 93914 241576
rect 99484 230382 99512 251246
rect 119448 232778 119476 253982
rect 122104 253972 122156 253978
rect 122104 253914 122156 253920
rect 121458 241632 121514 241641
rect 121458 241567 121514 241576
rect 121472 233238 121500 241567
rect 121460 233232 121512 233238
rect 121460 233174 121512 233180
rect 119370 232750 119476 232778
rect 100036 230450 100064 232084
rect 100024 230444 100076 230450
rect 100024 230386 100076 230392
rect 109696 230382 109724 232084
rect 122116 230382 122144 253914
rect 137664 251940 137692 253982
rect 147312 253972 147364 253978
rect 147312 253914 147364 253920
rect 148324 253972 148376 253978
rect 148324 253914 148376 253920
rect 147324 251940 147352 253914
rect 126888 251320 126940 251326
rect 126888 251262 126940 251268
rect 126900 242321 126928 251262
rect 127084 251246 128018 251274
rect 126886 242312 126942 242321
rect 126886 242247 126942 242256
rect 81992 230376 82044 230382
rect 81992 230318 82044 230324
rect 93124 230376 93176 230382
rect 93124 230318 93176 230324
rect 99472 230376 99524 230382
rect 99472 230318 99524 230324
rect 109684 230376 109736 230382
rect 109684 230318 109736 230324
rect 122104 230376 122156 230382
rect 122104 230318 122156 230324
rect 127084 230314 127112 251246
rect 147680 235408 147732 235414
rect 147680 235350 147732 235356
rect 147692 232778 147720 235350
rect 147338 232750 147720 232778
rect 128004 230450 128032 232084
rect 127992 230444 128044 230450
rect 127992 230386 128044 230392
rect 137664 230382 137692 232084
rect 148336 230382 148364 253914
rect 148428 235414 148456 254050
rect 149060 251252 149112 251258
rect 149060 251194 149112 251200
rect 149072 241641 149100 251194
rect 149058 241632 149114 241641
rect 149058 241567 149114 241576
rect 148416 235408 148468 235414
rect 148416 235350 148468 235356
rect 149704 231872 149756 231878
rect 149704 231814 149756 231820
rect 137652 230376 137704 230382
rect 137652 230318 137704 230324
rect 148324 230376 148376 230382
rect 148324 230318 148376 230324
rect 72056 230308 72108 230314
rect 72056 230250 72108 230256
rect 127072 230308 127124 230314
rect 127072 230250 127124 230256
rect 71136 226500 71188 226506
rect 71136 226442 71188 226448
rect 82268 226500 82320 226506
rect 82268 226442 82320 226448
rect 71148 202774 71176 226442
rect 72240 226432 72292 226438
rect 72240 226374 72292 226380
rect 72252 205714 72280 226374
rect 72608 226364 72660 226370
rect 72608 226306 72660 226312
rect 72620 224876 72648 226306
rect 82280 224876 82308 226442
rect 109960 226432 110012 226438
rect 109960 226374 110012 226380
rect 124864 226432 124916 226438
rect 124864 226374 124916 226380
rect 128636 226432 128688 226438
rect 128636 226374 128688 226380
rect 93124 226364 93176 226370
rect 93124 226306 93176 226312
rect 100300 226364 100352 226370
rect 100300 226306 100352 226312
rect 91954 224318 92152 224346
rect 72252 205686 72634 205714
rect 82280 202774 82308 205020
rect 91940 202842 91968 205020
rect 92124 202842 92152 224318
rect 91928 202836 91980 202842
rect 91928 202778 91980 202784
rect 92112 202836 92164 202842
rect 92112 202778 92164 202784
rect 93136 202774 93164 226306
rect 100208 226296 100260 226302
rect 100208 226238 100260 226244
rect 93860 223712 93912 223718
rect 93860 223654 93912 223660
rect 97908 223712 97960 223718
rect 97908 223654 97960 223660
rect 93872 214713 93900 223654
rect 97920 215393 97948 223654
rect 97906 215384 97962 215393
rect 97906 215319 97962 215328
rect 93858 214704 93914 214713
rect 93858 214639 93914 214648
rect 100220 205714 100248 226238
rect 100312 224890 100340 226306
rect 109972 224890 110000 226374
rect 100312 224862 100648 224890
rect 109972 224862 110308 224890
rect 119968 224330 120212 224346
rect 119968 224324 120224 224330
rect 119968 224318 120172 224324
rect 120172 224266 120224 224272
rect 122104 224324 122156 224330
rect 122104 224266 122156 224272
rect 121460 223644 121512 223650
rect 121460 223586 121512 223592
rect 121472 214713 121500 223586
rect 121458 214704 121514 214713
rect 121458 214639 121514 214648
rect 100220 205686 100648 205714
rect 110248 205006 110308 205034
rect 119632 205006 119968 205034
rect 110248 202774 110276 205006
rect 119632 202842 119660 205006
rect 122116 202842 122144 224266
rect 119620 202836 119672 202842
rect 119620 202778 119672 202784
rect 122104 202836 122156 202842
rect 122104 202778 122156 202784
rect 124876 202774 124904 226374
rect 128648 224876 128676 226374
rect 138296 226364 138348 226370
rect 138296 226306 138348 226312
rect 138308 224876 138336 226306
rect 147982 224318 148088 224346
rect 126888 223644 126940 223650
rect 126888 223586 126940 223592
rect 126900 215393 126928 223586
rect 126886 215384 126942 215393
rect 126886 215319 126942 215328
rect 128662 205006 128952 205034
rect 138322 205006 138704 205034
rect 128924 202774 128952 205006
rect 71136 202768 71188 202774
rect 71136 202710 71188 202716
rect 82268 202768 82320 202774
rect 82268 202710 82320 202716
rect 93124 202768 93176 202774
rect 93124 202710 93176 202716
rect 110236 202768 110288 202774
rect 110236 202710 110288 202716
rect 124864 202768 124916 202774
rect 124864 202710 124916 202716
rect 128912 202768 128964 202774
rect 128912 202710 128964 202716
rect 138676 202706 138704 205006
rect 147692 205006 147982 205034
rect 147692 202842 147720 205006
rect 148060 202842 148088 224318
rect 149060 223712 149112 223718
rect 149060 223654 149112 223660
rect 149072 214713 149100 223654
rect 149058 214704 149114 214713
rect 149058 214639 149114 214648
rect 147680 202836 147732 202842
rect 147680 202778 147732 202784
rect 148048 202836 148100 202842
rect 148048 202778 148100 202784
rect 138664 202700 138716 202706
rect 138664 202642 138716 202648
rect 148416 200320 148468 200326
rect 148416 200262 148468 200268
rect 81440 200252 81492 200258
rect 81440 200194 81492 200200
rect 91468 200252 91520 200258
rect 91468 200194 91520 200200
rect 109684 200252 109736 200258
rect 109684 200194 109736 200200
rect 119436 200252 119488 200258
rect 119436 200194 119488 200200
rect 137652 200252 137704 200258
rect 137652 200194 137704 200200
rect 81452 197962 81480 200194
rect 91100 200184 91152 200190
rect 91100 200126 91152 200132
rect 91112 197962 91140 200126
rect 81452 197934 81696 197962
rect 91112 197934 91356 197962
rect 71884 197254 72036 197282
rect 71884 176662 71912 197254
rect 91480 178786 91508 200194
rect 93124 200184 93176 200190
rect 93124 200126 93176 200132
rect 91356 178758 91508 178786
rect 72036 178078 72096 178106
rect 81696 178078 82032 178106
rect 71872 176656 71924 176662
rect 71872 176598 71924 176604
rect 72068 176526 72096 178078
rect 82004 176594 82032 178078
rect 93136 176594 93164 200126
rect 109696 197948 109724 200194
rect 119344 200184 119396 200190
rect 119344 200126 119396 200132
rect 119356 197948 119384 200126
rect 99484 197254 100050 197282
rect 97906 188320 97962 188329
rect 97906 188255 97962 188264
rect 93858 187640 93914 187649
rect 93858 187575 93914 187584
rect 93872 179314 93900 187575
rect 97920 179314 97948 188255
rect 93860 179308 93912 179314
rect 93860 179250 93912 179256
rect 97908 179308 97960 179314
rect 97908 179250 97960 179256
rect 99484 176594 99512 197254
rect 119448 178786 119476 200194
rect 124864 200184 124916 200190
rect 124864 200126 124916 200132
rect 121458 187640 121514 187649
rect 121458 187575 121514 187584
rect 121472 179382 121500 187575
rect 121460 179376 121512 179382
rect 121460 179318 121512 179324
rect 119370 178758 119476 178786
rect 100036 176662 100064 178092
rect 100024 176656 100076 176662
rect 100024 176598 100076 176604
rect 109696 176594 109724 178092
rect 124876 176594 124904 200126
rect 137664 197948 137692 200194
rect 147312 200184 147364 200190
rect 147312 200126 147364 200132
rect 148324 200184 148376 200190
rect 148324 200126 148376 200132
rect 147324 197948 147352 200126
rect 127084 197254 128018 197282
rect 126886 188320 126942 188329
rect 126886 188255 126942 188264
rect 126900 179382 126928 188255
rect 126888 179376 126940 179382
rect 126888 179318 126940 179324
rect 81992 176588 82044 176594
rect 81992 176530 82044 176536
rect 93124 176588 93176 176594
rect 93124 176530 93176 176536
rect 99472 176588 99524 176594
rect 99472 176530 99524 176536
rect 109684 176588 109736 176594
rect 109684 176530 109736 176536
rect 124864 176588 124916 176594
rect 124864 176530 124916 176536
rect 127084 176526 127112 197254
rect 147680 185632 147732 185638
rect 147680 185574 147732 185580
rect 147692 178786 147720 185574
rect 147338 178758 147720 178786
rect 128004 176662 128032 178092
rect 127992 176656 128044 176662
rect 127992 176598 128044 176604
rect 137664 176594 137692 178092
rect 148336 176594 148364 200126
rect 148428 185638 148456 200262
rect 149058 187640 149114 187649
rect 149058 187575 149114 187584
rect 148416 185632 148468 185638
rect 148416 185574 148468 185580
rect 149072 179314 149100 187575
rect 149060 179308 149112 179314
rect 149060 179250 149112 179256
rect 137652 176588 137704 176594
rect 137652 176530 137704 176536
rect 148324 176588 148376 176594
rect 148324 176530 148376 176536
rect 72056 176520 72108 176526
rect 72056 176462 72108 176468
rect 127072 176520 127124 176526
rect 127072 176462 127124 176468
rect 71136 172712 71188 172718
rect 71136 172654 71188 172660
rect 82268 172712 82320 172718
rect 82268 172654 82320 172660
rect 99380 172712 99432 172718
rect 99380 172654 99432 172660
rect 100300 172712 100352 172718
rect 100300 172654 100352 172660
rect 71148 148986 71176 172654
rect 71872 172644 71924 172650
rect 71872 172586 71924 172592
rect 71884 171134 71912 172586
rect 72608 172576 72660 172582
rect 72608 172518 72660 172524
rect 71884 171106 72280 171134
rect 72252 151722 72280 171106
rect 72620 170884 72648 172518
rect 82280 170884 82308 172654
rect 99392 172582 99420 172654
rect 93124 172576 93176 172582
rect 93124 172518 93176 172524
rect 99380 172576 99432 172582
rect 99380 172518 99432 172524
rect 99472 172576 99524 172582
rect 99472 172518 99524 172524
rect 91954 170326 92152 170354
rect 72252 151694 72634 151722
rect 82280 148986 82308 151028
rect 91940 149054 91968 151028
rect 92124 149054 92152 170326
rect 91928 149048 91980 149054
rect 91928 148990 91980 148996
rect 92112 149048 92164 149054
rect 92112 148990 92164 148996
rect 93136 148986 93164 172518
rect 99484 171134 99512 172518
rect 99484 171106 100248 171134
rect 97906 161392 97962 161401
rect 97906 161327 97962 161336
rect 93858 160712 93914 160721
rect 93858 160647 93914 160656
rect 93872 151706 93900 160647
rect 97920 151706 97948 161327
rect 100220 151722 100248 171106
rect 100312 170898 100340 172654
rect 109960 172644 110012 172650
rect 109960 172586 110012 172592
rect 124864 172644 124916 172650
rect 124864 172586 124916 172592
rect 128636 172644 128688 172650
rect 128636 172586 128688 172592
rect 109972 170898 110000 172586
rect 100312 170870 100648 170898
rect 109972 170870 110308 170898
rect 119968 170338 120212 170354
rect 119968 170332 120224 170338
rect 119968 170326 120172 170332
rect 120172 170274 120224 170280
rect 122104 170332 122156 170338
rect 122104 170274 122156 170280
rect 121458 160712 121514 160721
rect 121458 160647 121514 160656
rect 121472 151774 121500 160647
rect 121460 151768 121512 151774
rect 93860 151700 93912 151706
rect 93860 151642 93912 151648
rect 97908 151700 97960 151706
rect 100220 151694 100648 151722
rect 121460 151710 121512 151716
rect 97908 151642 97960 151648
rect 110248 151014 110308 151042
rect 119632 151014 119968 151042
rect 110248 148986 110276 151014
rect 119632 149054 119660 151014
rect 122116 149054 122144 170274
rect 119620 149048 119672 149054
rect 119620 148990 119672 148996
rect 122104 149048 122156 149054
rect 122104 148990 122156 148996
rect 124876 148986 124904 172586
rect 128648 170884 128676 172586
rect 138296 172576 138348 172582
rect 138296 172518 138348 172524
rect 138308 170884 138336 172518
rect 147982 170326 148088 170354
rect 126886 161392 126942 161401
rect 126886 161327 126942 161336
rect 126900 151774 126928 161327
rect 126888 151768 126940 151774
rect 126888 151710 126940 151716
rect 128648 148986 128676 151028
rect 71136 148980 71188 148986
rect 71136 148922 71188 148928
rect 82268 148980 82320 148986
rect 82268 148922 82320 148928
rect 93124 148980 93176 148986
rect 93124 148922 93176 148928
rect 110236 148980 110288 148986
rect 110236 148922 110288 148928
rect 124864 148980 124916 148986
rect 124864 148922 124916 148928
rect 128636 148980 128688 148986
rect 128636 148922 128688 148928
rect 138308 148918 138336 151028
rect 147968 149054 147996 151028
rect 148060 149054 148088 170326
rect 149058 160712 149114 160721
rect 149058 160647 149114 160656
rect 149072 151706 149100 160647
rect 149060 151700 149112 151706
rect 149060 151642 149112 151648
rect 147956 149048 148008 149054
rect 147956 148990 148008 148996
rect 148048 149048 148100 149054
rect 148048 148990 148100 148996
rect 138296 148912 138348 148918
rect 138296 148854 138348 148860
rect 148324 146464 148376 146470
rect 148324 146406 148376 146412
rect 81440 146396 81492 146402
rect 81440 146338 81492 146344
rect 91468 146396 91520 146402
rect 91468 146338 91520 146344
rect 109684 146396 109736 146402
rect 109684 146338 109736 146344
rect 119436 146396 119488 146402
rect 119436 146338 119488 146344
rect 137652 146396 137704 146402
rect 137652 146338 137704 146344
rect 81452 143970 81480 146338
rect 91100 146328 91152 146334
rect 91100 146270 91152 146276
rect 91112 143970 91140 146270
rect 81452 143942 81696 143970
rect 91112 143942 91356 143970
rect 71884 143262 72036 143290
rect 71884 122806 71912 143262
rect 91480 124794 91508 146338
rect 93124 146328 93176 146334
rect 93124 146270 93176 146276
rect 91356 124766 91508 124794
rect 72022 123842 72050 124100
rect 81696 124086 82032 124114
rect 71976 123814 72050 123842
rect 71872 122800 71924 122806
rect 71872 122742 71924 122748
rect 71976 122670 72004 123814
rect 82004 122738 82032 124086
rect 93136 122738 93164 146270
rect 109696 143956 109724 146338
rect 119344 146328 119396 146334
rect 119344 146270 119396 146276
rect 119356 143956 119384 146270
rect 99484 143262 100050 143290
rect 97906 134328 97962 134337
rect 97906 134263 97962 134272
rect 93858 133648 93914 133657
rect 93858 133583 93914 133592
rect 93872 125526 93900 133583
rect 97920 125526 97948 134263
rect 93860 125520 93912 125526
rect 93860 125462 93912 125468
rect 97908 125520 97960 125526
rect 97908 125462 97960 125468
rect 99484 122738 99512 143262
rect 119448 124794 119476 146338
rect 124864 146328 124916 146334
rect 124864 146270 124916 146276
rect 121458 133648 121514 133657
rect 121458 133583 121514 133592
rect 121472 125594 121500 133583
rect 121460 125588 121512 125594
rect 121460 125530 121512 125536
rect 119370 124766 119476 124794
rect 100036 122806 100064 124100
rect 100024 122800 100076 122806
rect 100024 122742 100076 122748
rect 109696 122738 109724 124100
rect 124876 122738 124904 146270
rect 137664 143956 137692 146338
rect 147312 146328 147364 146334
rect 147312 146270 147364 146276
rect 147324 143956 147352 146270
rect 127084 143262 128018 143290
rect 126886 134328 126942 134337
rect 126886 134263 126942 134272
rect 126900 125594 126928 134263
rect 126888 125588 126940 125594
rect 126888 125530 126940 125536
rect 81992 122732 82044 122738
rect 81992 122674 82044 122680
rect 93124 122732 93176 122738
rect 93124 122674 93176 122680
rect 99472 122732 99524 122738
rect 99472 122674 99524 122680
rect 109684 122732 109736 122738
rect 109684 122674 109736 122680
rect 124864 122732 124916 122738
rect 124864 122674 124916 122680
rect 127084 122670 127112 143262
rect 148336 132494 148364 146406
rect 148416 146328 148468 146334
rect 148416 146270 148468 146276
rect 147784 132466 148364 132494
rect 147784 124794 147812 132466
rect 147338 124766 147812 124794
rect 128004 122806 128032 124100
rect 127992 122800 128044 122806
rect 127992 122742 128044 122748
rect 137664 122738 137692 124100
rect 148428 122738 148456 146270
rect 149058 133648 149114 133657
rect 149058 133583 149114 133592
rect 149072 125526 149100 133583
rect 149060 125520 149112 125526
rect 149060 125462 149112 125468
rect 137652 122732 137704 122738
rect 137652 122674 137704 122680
rect 148416 122732 148468 122738
rect 148416 122674 148468 122680
rect 71964 122664 72016 122670
rect 71964 122606 72016 122612
rect 127072 122664 127124 122670
rect 127072 122606 127124 122612
rect 71136 118856 71188 118862
rect 71136 118798 71188 118804
rect 82268 118856 82320 118862
rect 82268 118798 82320 118804
rect 99472 118856 99524 118862
rect 99472 118798 99524 118804
rect 138296 118856 138348 118862
rect 138296 118798 138348 118804
rect 71148 95130 71176 118798
rect 71872 118788 71924 118794
rect 71872 118730 71924 118736
rect 71884 113174 71912 118730
rect 72608 118720 72660 118726
rect 72608 118662 72660 118668
rect 72620 116892 72648 118662
rect 82280 116892 82308 118798
rect 93124 118720 93176 118726
rect 93124 118662 93176 118668
rect 91954 116334 92152 116362
rect 71884 113146 72280 113174
rect 72252 97730 72280 113146
rect 72252 97702 72634 97730
rect 82280 95130 82308 97036
rect 91940 95198 91968 97036
rect 92124 95198 92152 116334
rect 91928 95192 91980 95198
rect 91928 95134 91980 95140
rect 92112 95192 92164 95198
rect 92112 95134 92164 95140
rect 93136 95130 93164 118662
rect 99484 113174 99512 118798
rect 109960 118788 110012 118794
rect 109960 118730 110012 118736
rect 120724 118788 120776 118794
rect 120724 118730 120776 118736
rect 128636 118788 128688 118794
rect 128636 118730 128688 118736
rect 100300 118720 100352 118726
rect 100300 118662 100352 118668
rect 100312 116906 100340 118662
rect 109972 116906 110000 118730
rect 100312 116878 100648 116906
rect 109972 116878 110308 116906
rect 119968 116346 120120 116362
rect 119968 116340 120132 116346
rect 119968 116334 120080 116340
rect 120080 116282 120132 116288
rect 99484 113146 100248 113174
rect 97906 107400 97962 107409
rect 97906 107335 97962 107344
rect 93858 106720 93914 106729
rect 93858 106655 93914 106664
rect 93872 97850 93900 106655
rect 97920 97986 97948 107335
rect 97908 97980 97960 97986
rect 97908 97922 97960 97928
rect 93860 97844 93912 97850
rect 93860 97786 93912 97792
rect 100220 97730 100248 113146
rect 100220 97702 100648 97730
rect 110248 97022 110308 97050
rect 119632 97022 119968 97050
rect 110248 95130 110276 97022
rect 119632 95198 119660 97022
rect 119620 95192 119672 95198
rect 119620 95134 119672 95140
rect 120736 95130 120764 118730
rect 128648 116892 128676 118730
rect 138308 116892 138336 118798
rect 148324 118720 148376 118726
rect 148324 118662 148376 118668
rect 122104 116340 122156 116346
rect 147982 116334 148088 116362
rect 122104 116282 122156 116288
rect 121458 106720 121514 106729
rect 121458 106655 121514 106664
rect 121472 97918 121500 106655
rect 121460 97912 121512 97918
rect 121460 97854 121512 97860
rect 122116 95198 122144 116282
rect 126886 107400 126942 107409
rect 126886 107335 126942 107344
rect 126900 97918 126928 107335
rect 126888 97912 126940 97918
rect 126888 97854 126940 97860
rect 122104 95192 122156 95198
rect 122104 95134 122156 95140
rect 128648 95130 128676 97036
rect 71136 95124 71188 95130
rect 71136 95066 71188 95072
rect 82268 95124 82320 95130
rect 82268 95066 82320 95072
rect 93124 95124 93176 95130
rect 93124 95066 93176 95072
rect 110236 95124 110288 95130
rect 110236 95066 110288 95072
rect 120724 95124 120776 95130
rect 120724 95066 120776 95072
rect 128636 95124 128688 95130
rect 128636 95066 128688 95072
rect 138308 95062 138336 97036
rect 147968 95198 147996 97036
rect 148060 95198 148088 116334
rect 147956 95192 148008 95198
rect 147956 95134 148008 95140
rect 148048 95192 148100 95198
rect 148048 95134 148100 95140
rect 148336 95130 148364 118662
rect 149058 106720 149114 106729
rect 149058 106655 149114 106664
rect 149072 97986 149100 106655
rect 149060 97980 149112 97986
rect 149060 97922 149112 97928
rect 148324 95124 148376 95130
rect 148324 95066 148376 95072
rect 138296 95056 138348 95062
rect 138296 94998 138348 95004
rect 148416 91248 148468 91254
rect 148416 91190 148468 91196
rect 81440 91180 81492 91186
rect 81440 91122 81492 91128
rect 91468 91180 91520 91186
rect 91468 91122 91520 91128
rect 109684 91180 109736 91186
rect 109684 91122 109736 91128
rect 119436 91180 119488 91186
rect 119436 91122 119488 91128
rect 137652 91180 137704 91186
rect 137652 91122 137704 91128
rect 81452 89978 81480 91122
rect 91100 91112 91152 91118
rect 91100 91054 91152 91060
rect 91112 89978 91140 91054
rect 81452 89950 81696 89978
rect 91112 89950 91356 89978
rect 71884 89270 72036 89298
rect 71884 69018 71912 89270
rect 91480 70666 91508 91122
rect 93124 91112 93176 91118
rect 93124 91054 93176 91060
rect 91356 70638 91508 70666
rect 72036 70094 72096 70122
rect 81696 70094 82032 70122
rect 71872 69012 71924 69018
rect 71872 68954 71924 68960
rect 72068 68882 72096 70094
rect 82004 68950 82032 70094
rect 93136 68950 93164 91054
rect 109696 89964 109724 91122
rect 119344 91112 119396 91118
rect 119344 91054 119396 91060
rect 119356 89964 119384 91054
rect 99484 89270 100050 89298
rect 93860 88392 93912 88398
rect 93860 88334 93912 88340
rect 97908 88392 97960 88398
rect 97908 88334 97960 88340
rect 93872 79665 93900 88334
rect 97920 80345 97948 88334
rect 97906 80336 97962 80345
rect 97906 80271 97962 80280
rect 93858 79656 93914 79665
rect 93858 79591 93914 79600
rect 99484 68950 99512 89270
rect 119448 70666 119476 91122
rect 124864 91112 124916 91118
rect 124864 91054 124916 91060
rect 121458 79656 121514 79665
rect 121458 79591 121514 79600
rect 121472 71738 121500 79591
rect 121460 71732 121512 71738
rect 121460 71674 121512 71680
rect 119370 70638 119476 70666
rect 100036 69018 100064 70108
rect 100024 69012 100076 69018
rect 100024 68954 100076 68960
rect 109696 68950 109724 70108
rect 124876 68950 124904 91054
rect 137664 89964 137692 91122
rect 147312 91112 147364 91118
rect 147312 91054 147364 91060
rect 148324 91112 148376 91118
rect 148324 91054 148376 91060
rect 147324 89964 147352 91054
rect 127084 89270 128018 89298
rect 126886 80336 126942 80345
rect 126886 80271 126942 80280
rect 126900 71738 126928 80271
rect 126888 71732 126940 71738
rect 126888 71674 126940 71680
rect 81992 68944 82044 68950
rect 81992 68886 82044 68892
rect 93124 68944 93176 68950
rect 93124 68886 93176 68892
rect 99472 68944 99524 68950
rect 99472 68886 99524 68892
rect 109684 68944 109736 68950
rect 109684 68886 109736 68892
rect 124864 68944 124916 68950
rect 124864 68886 124916 68892
rect 127084 68882 127112 89270
rect 147680 72344 147732 72350
rect 147680 72286 147732 72292
rect 147692 70666 147720 72286
rect 147338 70638 147720 70666
rect 128004 69018 128032 70108
rect 127992 69012 128044 69018
rect 127992 68954 128044 68960
rect 137664 68950 137692 70108
rect 148336 68950 148364 91054
rect 148428 72350 148456 91190
rect 149060 88392 149112 88398
rect 149060 88334 149112 88340
rect 149072 79665 149100 88334
rect 149058 79656 149114 79665
rect 149058 79591 149114 79600
rect 148416 72344 148468 72350
rect 148416 72286 148468 72292
rect 137652 68944 137704 68950
rect 137652 68886 137704 68892
rect 148324 68944 148376 68950
rect 148324 68886 148376 68892
rect 72056 68876 72108 68882
rect 72056 68818 72108 68824
rect 127072 68876 127124 68882
rect 127072 68818 127124 68824
rect 71136 65068 71188 65074
rect 71136 65010 71188 65016
rect 82268 65068 82320 65074
rect 82268 65010 82320 65016
rect 99380 65068 99432 65074
rect 99380 65010 99432 65016
rect 100300 65068 100352 65074
rect 100300 65010 100352 65016
rect 71148 41342 71176 65010
rect 71872 65000 71924 65006
rect 71872 64942 71924 64948
rect 71884 55214 71912 64942
rect 72608 64932 72660 64938
rect 72608 64874 72660 64880
rect 72620 62900 72648 64874
rect 82280 62900 82308 65010
rect 99392 64938 99420 65010
rect 93124 64932 93176 64938
rect 93124 64874 93176 64880
rect 99380 64932 99432 64938
rect 99380 64874 99432 64880
rect 99472 64932 99524 64938
rect 99472 64874 99524 64880
rect 91954 62206 92152 62234
rect 71884 55186 72280 55214
rect 72252 43738 72280 55186
rect 72252 43710 72634 43738
rect 82280 41342 82308 43044
rect 91940 41410 91968 43044
rect 92124 41410 92152 62206
rect 91928 41404 91980 41410
rect 91928 41346 91980 41352
rect 92112 41404 92164 41410
rect 92112 41346 92164 41352
rect 93136 41342 93164 64874
rect 93860 62144 93912 62150
rect 93860 62086 93912 62092
rect 97908 62144 97960 62150
rect 97908 62086 97960 62092
rect 93872 52737 93900 62086
rect 97920 53417 97948 62086
rect 99484 55214 99512 64874
rect 100312 62914 100340 65010
rect 109960 65000 110012 65006
rect 109960 64942 110012 64948
rect 124864 65000 124916 65006
rect 124864 64942 124916 64948
rect 128636 65000 128688 65006
rect 128636 64942 128688 64948
rect 109972 62914 110000 64942
rect 100312 62886 100648 62914
rect 109972 62886 110308 62914
rect 119968 62218 120304 62234
rect 119968 62212 120316 62218
rect 119968 62206 120264 62212
rect 120264 62154 120316 62160
rect 122104 62212 122156 62218
rect 122104 62154 122156 62160
rect 99484 55186 100248 55214
rect 97906 53408 97962 53417
rect 97906 53343 97962 53352
rect 93858 52728 93914 52737
rect 93858 52663 93914 52672
rect 100220 43738 100248 55186
rect 121458 52728 121514 52737
rect 121458 52663 121514 52672
rect 121472 44130 121500 52663
rect 121460 44124 121512 44130
rect 121460 44066 121512 44072
rect 100220 43710 100648 43738
rect 110248 43030 110308 43058
rect 119632 43030 119968 43058
rect 110248 41342 110276 43030
rect 119632 41410 119660 43030
rect 122116 41410 122144 62154
rect 119620 41404 119672 41410
rect 119620 41346 119672 41352
rect 122104 41404 122156 41410
rect 122104 41346 122156 41352
rect 124876 41342 124904 64942
rect 128648 62900 128676 64942
rect 138296 64932 138348 64938
rect 138296 64874 138348 64880
rect 138308 62900 138336 64874
rect 147982 62206 148088 62234
rect 126886 53408 126942 53417
rect 126886 53343 126942 53352
rect 126900 44130 126928 53343
rect 126888 44124 126940 44130
rect 126888 44066 126940 44072
rect 128648 41342 128676 43044
rect 71136 41336 71188 41342
rect 71136 41278 71188 41284
rect 82268 41336 82320 41342
rect 82268 41278 82320 41284
rect 93124 41336 93176 41342
rect 93124 41278 93176 41284
rect 110236 41336 110288 41342
rect 110236 41278 110288 41284
rect 124864 41336 124916 41342
rect 124864 41278 124916 41284
rect 128636 41336 128688 41342
rect 128636 41278 128688 41284
rect 138308 41274 138336 43044
rect 147968 41410 147996 43044
rect 148060 41410 148088 62206
rect 149060 62144 149112 62150
rect 149060 62086 149112 62092
rect 149072 52737 149100 62086
rect 149058 52728 149114 52737
rect 149058 52663 149114 52672
rect 147956 41404 148008 41410
rect 147956 41346 148008 41352
rect 148048 41404 148100 41410
rect 148048 41346 148100 41352
rect 138296 41268 138348 41274
rect 138296 41210 138348 41216
rect 149716 38418 149744 231814
rect 152464 226432 152516 226438
rect 152464 226374 152516 226380
rect 151084 226364 151136 226370
rect 151084 226306 151136 226312
rect 151096 202774 151124 226306
rect 151084 202768 151136 202774
rect 151084 202710 151136 202716
rect 152476 202706 152504 226374
rect 152464 202700 152516 202706
rect 152464 202642 152516 202648
rect 152464 172644 152516 172650
rect 152464 172586 152516 172592
rect 151084 172576 151136 172582
rect 151084 172518 151136 172524
rect 151096 148986 151124 172518
rect 151084 148980 151136 148986
rect 151084 148922 151136 148928
rect 152476 148918 152504 172586
rect 152464 148912 152516 148918
rect 152464 148854 152516 148860
rect 151084 118788 151136 118794
rect 151084 118730 151136 118736
rect 151096 95062 151124 118730
rect 151084 95056 151136 95062
rect 151084 94998 151136 95004
rect 152464 65000 152516 65006
rect 152464 64942 152516 64948
rect 151084 64932 151136 64938
rect 151084 64874 151136 64880
rect 151096 41342 151124 64874
rect 151084 41336 151136 41342
rect 151084 41278 151136 41284
rect 152476 41274 152504 64942
rect 153856 42129 153884 700402
rect 202800 700330 202828 703520
rect 204904 700460 204956 700466
rect 204904 700402 204956 700408
rect 202788 700324 202840 700330
rect 202788 700266 202840 700272
rect 165712 686044 165764 686050
rect 165712 685986 165764 685992
rect 175464 686044 175516 686050
rect 175464 685986 175516 685992
rect 193680 686044 193732 686050
rect 193680 685986 193732 685992
rect 203524 686044 203576 686050
rect 203524 685986 203576 685992
rect 156328 685976 156380 685982
rect 156328 685918 156380 685924
rect 156340 683890 156368 685918
rect 156032 683862 156368 683890
rect 165724 683754 165752 685986
rect 175372 685908 175424 685914
rect 175372 685850 175424 685856
rect 175384 683754 175412 685850
rect 165692 683726 165752 683754
rect 175352 683726 175412 683754
rect 154488 683188 154540 683194
rect 154488 683130 154540 683136
rect 154500 674257 154528 683130
rect 154486 674248 154542 674257
rect 154486 674183 154542 674192
rect 175476 664714 175504 685986
rect 178684 685976 178736 685982
rect 178684 685918 178736 685924
rect 177304 685908 177356 685914
rect 177304 685850 177356 685856
rect 175352 664686 175504 664714
rect 156018 663794 156046 664020
rect 165692 664006 166028 664034
rect 155972 663766 156046 663794
rect 155972 662250 156000 663766
rect 166000 662386 166028 664006
rect 177316 662386 177344 685850
rect 178038 673568 178094 673577
rect 178038 673503 178094 673512
rect 178052 665174 178080 673503
rect 178040 665168 178092 665174
rect 178040 665110 178092 665116
rect 178696 662386 178724 685918
rect 193692 683876 193720 685986
rect 203340 685908 203392 685914
rect 203340 685850 203392 685856
rect 203352 683876 203380 685850
rect 183664 683318 184046 683346
rect 182088 683256 182140 683262
rect 182088 683198 182140 683204
rect 182100 674257 182128 683198
rect 182086 674248 182142 674257
rect 182086 674183 182142 674192
rect 165988 662380 166040 662386
rect 165988 662322 166040 662328
rect 177304 662380 177356 662386
rect 177304 662322 177356 662328
rect 178684 662380 178736 662386
rect 178684 662322 178736 662328
rect 183664 662318 183692 683318
rect 203536 664714 203564 685986
rect 203366 664686 203564 664714
rect 184032 662386 184060 664020
rect 184020 662380 184072 662386
rect 184020 662322 184072 662328
rect 193692 662318 193720 664020
rect 183652 662312 183704 662318
rect 183652 662254 183704 662260
rect 193680 662312 193732 662318
rect 193680 662254 193732 662260
rect 155960 662244 156012 662250
rect 155960 662186 156012 662192
rect 183652 658436 183704 658442
rect 183652 658378 183704 658384
rect 156604 658368 156656 658374
rect 156604 658310 156656 658316
rect 182824 658368 182876 658374
rect 182824 658310 182876 658316
rect 156616 656948 156644 658310
rect 166264 658300 166316 658306
rect 166264 658242 166316 658248
rect 177304 658300 177356 658306
rect 177304 658242 177356 658248
rect 166276 656948 166304 658242
rect 175950 656254 176148 656282
rect 156420 655648 156472 655654
rect 156420 655590 156472 655596
rect 156432 648009 156460 655590
rect 156418 648000 156474 648009
rect 156418 647935 156474 647944
rect 156616 634710 156644 637092
rect 156604 634704 156656 634710
rect 156604 634646 156656 634652
rect 166276 634642 166304 637092
rect 175936 634778 175964 637092
rect 176120 634778 176148 656254
rect 175924 634772 175976 634778
rect 175924 634714 175976 634720
rect 176108 634772 176160 634778
rect 176108 634714 176160 634720
rect 177316 634642 177344 658242
rect 178040 655580 178092 655586
rect 178040 655522 178092 655528
rect 178052 646785 178080 655522
rect 178038 646776 178094 646785
rect 178038 646711 178094 646720
rect 182836 634710 182864 658310
rect 183664 654134 183692 658378
rect 193956 658368 194008 658374
rect 193956 658310 194008 658316
rect 184296 658300 184348 658306
rect 184296 658242 184348 658248
rect 184308 656962 184336 658242
rect 193968 656962 193996 658310
rect 184308 656934 184644 656962
rect 193968 656934 194304 656962
rect 203964 656254 204300 656282
rect 184388 655716 184440 655722
rect 184388 655658 184440 655664
rect 183664 654106 184244 654134
rect 184216 637786 184244 654106
rect 184400 648009 184428 655658
rect 204272 654362 204300 656254
rect 204260 654356 204312 654362
rect 204260 654298 204312 654304
rect 184386 648000 184442 648009
rect 184386 647935 184442 647944
rect 184216 637758 184644 637786
rect 194304 637078 194548 637106
rect 194520 634710 194548 637078
rect 203628 637078 203964 637106
rect 203628 634778 203656 637078
rect 203616 634772 203668 634778
rect 203616 634714 203668 634720
rect 182824 634704 182876 634710
rect 182824 634646 182876 634652
rect 194508 634704 194560 634710
rect 194508 634646 194560 634652
rect 166264 634636 166316 634642
rect 166264 634578 166316 634584
rect 177304 634636 177356 634642
rect 177304 634578 177356 634584
rect 165712 632256 165764 632262
rect 165712 632198 165764 632204
rect 175464 632256 175516 632262
rect 175464 632198 175516 632204
rect 193680 632256 193732 632262
rect 193680 632198 193732 632204
rect 203524 632256 203576 632262
rect 203524 632198 203576 632204
rect 156328 632188 156380 632194
rect 156328 632130 156380 632136
rect 156340 629898 156368 632130
rect 156032 629870 156368 629898
rect 165724 629762 165752 632198
rect 175372 632120 175424 632126
rect 175372 632062 175424 632068
rect 175384 629762 175412 632062
rect 165692 629734 165752 629762
rect 175352 629734 175412 629762
rect 154486 620256 154542 620265
rect 154486 620191 154542 620200
rect 154500 611250 154528 620191
rect 154488 611244 154540 611250
rect 154488 611186 154540 611192
rect 175476 610722 175504 632198
rect 178684 632188 178736 632194
rect 178684 632130 178736 632136
rect 177304 632120 177356 632126
rect 177304 632062 177356 632068
rect 175352 610694 175504 610722
rect 156032 610014 156092 610042
rect 165692 610014 166028 610042
rect 156064 608462 156092 610014
rect 166000 608598 166028 610014
rect 177316 608598 177344 632062
rect 178038 619576 178094 619585
rect 178038 619511 178094 619520
rect 178052 611318 178080 619511
rect 178040 611312 178092 611318
rect 178040 611254 178092 611260
rect 178696 608598 178724 632130
rect 193692 629884 193720 632198
rect 203340 632120 203392 632126
rect 203340 632062 203392 632068
rect 203352 629884 203380 632062
rect 183664 629326 184046 629354
rect 182086 620256 182142 620265
rect 182086 620191 182142 620200
rect 182100 611182 182128 620191
rect 182088 611176 182140 611182
rect 182088 611118 182140 611124
rect 165988 608592 166040 608598
rect 165988 608534 166040 608540
rect 177304 608592 177356 608598
rect 177304 608534 177356 608540
rect 178684 608592 178736 608598
rect 178684 608534 178736 608540
rect 183664 608530 183692 629326
rect 203536 610722 203564 632198
rect 203366 610694 203564 610722
rect 184032 608598 184060 610028
rect 184020 608592 184072 608598
rect 184020 608534 184072 608540
rect 193692 608530 193720 610028
rect 183652 608524 183704 608530
rect 183652 608466 183704 608472
rect 193680 608524 193732 608530
rect 193680 608466 193732 608472
rect 156052 608456 156104 608462
rect 156052 608398 156104 608404
rect 183652 604648 183704 604654
rect 183652 604590 183704 604596
rect 156604 604580 156656 604586
rect 156604 604522 156656 604528
rect 182824 604580 182876 604586
rect 182824 604522 182876 604528
rect 156616 602956 156644 604522
rect 166264 604512 166316 604518
rect 166264 604454 166316 604460
rect 177304 604512 177356 604518
rect 177304 604454 177356 604460
rect 166276 602956 166304 604454
rect 175950 602262 176148 602290
rect 154488 601792 154540 601798
rect 154488 601734 154540 601740
rect 154500 593473 154528 601734
rect 154486 593464 154542 593473
rect 154486 593399 154542 593408
rect 156616 580922 156644 583100
rect 156604 580916 156656 580922
rect 156604 580858 156656 580864
rect 166276 580854 166304 583100
rect 175936 580990 175964 583100
rect 176120 580990 176148 602262
rect 175924 580984 175976 580990
rect 175924 580926 175976 580932
rect 176108 580984 176160 580990
rect 176108 580926 176160 580932
rect 177316 580854 177344 604454
rect 182088 601860 182140 601866
rect 182088 601802 182140 601808
rect 178040 601724 178092 601730
rect 178040 601666 178092 601672
rect 178052 592793 178080 601666
rect 182100 593473 182128 601802
rect 182086 593464 182142 593473
rect 182086 593399 182142 593408
rect 178038 592784 178094 592793
rect 178038 592719 178094 592728
rect 182836 580922 182864 604522
rect 183664 596174 183692 604590
rect 193956 604580 194008 604586
rect 193956 604522 194008 604528
rect 184296 604512 184348 604518
rect 184296 604454 184348 604460
rect 184308 602970 184336 604454
rect 193968 602970 193996 604522
rect 184308 602942 184644 602970
rect 193968 602942 194304 602970
rect 203964 602262 204300 602290
rect 204272 599282 204300 602262
rect 204260 599276 204312 599282
rect 204260 599218 204312 599224
rect 183664 596146 184244 596174
rect 184216 583794 184244 596146
rect 184216 583766 184644 583794
rect 194304 583086 194548 583114
rect 194520 580922 194548 583086
rect 203628 583086 203964 583114
rect 203628 580990 203656 583086
rect 203616 580984 203668 580990
rect 203616 580926 203668 580932
rect 182824 580916 182876 580922
rect 182824 580858 182876 580864
rect 194508 580916 194560 580922
rect 194508 580858 194560 580864
rect 166264 580848 166316 580854
rect 166264 580790 166316 580796
rect 177304 580848 177356 580854
rect 177304 580790 177356 580796
rect 165620 578400 165672 578406
rect 165620 578342 165672 578348
rect 175464 578400 175516 578406
rect 175464 578342 175516 578348
rect 193680 578400 193732 578406
rect 193680 578342 193732 578348
rect 203524 578400 203576 578406
rect 203524 578342 203576 578348
rect 156328 578332 156380 578338
rect 156328 578274 156380 578280
rect 156340 575906 156368 578274
rect 165632 576178 165660 578342
rect 175280 578264 175332 578270
rect 175280 578206 175332 578212
rect 175292 576178 175320 578206
rect 165632 576150 165706 576178
rect 175292 576150 175366 576178
rect 156032 575878 156368 575906
rect 165678 575892 165706 576150
rect 175338 575892 175366 576150
rect 154486 566264 154542 566273
rect 154486 566199 154542 566208
rect 154500 557462 154528 566199
rect 154488 557456 154540 557462
rect 154488 557398 154540 557404
rect 175476 556730 175504 578342
rect 178684 578332 178736 578338
rect 178684 578274 178736 578280
rect 177304 578264 177356 578270
rect 177304 578206 177356 578212
rect 175352 556702 175504 556730
rect 156032 556022 156092 556050
rect 165692 556022 166028 556050
rect 156064 554606 156092 556022
rect 166000 554742 166028 556022
rect 177316 554742 177344 578206
rect 178038 565584 178094 565593
rect 178038 565519 178094 565528
rect 178052 557530 178080 565519
rect 178040 557524 178092 557530
rect 178040 557466 178092 557472
rect 178696 554742 178724 578274
rect 193692 575892 193720 578342
rect 203340 578264 203392 578270
rect 203340 578206 203392 578212
rect 203352 575892 203380 578206
rect 183664 575334 184046 575362
rect 182086 566264 182142 566273
rect 182086 566199 182142 566208
rect 182100 557394 182128 566199
rect 182088 557388 182140 557394
rect 182088 557330 182140 557336
rect 165988 554736 166040 554742
rect 165988 554678 166040 554684
rect 177304 554736 177356 554742
rect 177304 554678 177356 554684
rect 178684 554736 178736 554742
rect 178684 554678 178736 554684
rect 183664 554674 183692 575334
rect 203536 556730 203564 578342
rect 203366 556702 203564 556730
rect 184032 554742 184060 556036
rect 184020 554736 184072 554742
rect 184020 554678 184072 554684
rect 193692 554674 193720 556036
rect 183652 554668 183704 554674
rect 183652 554610 183704 554616
rect 193680 554668 193732 554674
rect 193680 554610 193732 554616
rect 156052 554600 156104 554606
rect 156052 554542 156104 554548
rect 183652 550792 183704 550798
rect 183652 550734 183704 550740
rect 156604 550724 156656 550730
rect 156604 550666 156656 550672
rect 182824 550724 182876 550730
rect 182824 550666 182876 550672
rect 156616 548964 156644 550666
rect 166264 550656 166316 550662
rect 166264 550598 166316 550604
rect 177304 550656 177356 550662
rect 177304 550598 177356 550604
rect 166276 548964 166304 550598
rect 175950 548270 176148 548298
rect 154486 539472 154542 539481
rect 154486 539407 154542 539416
rect 154500 529854 154528 539407
rect 154488 529848 154540 529854
rect 154488 529790 154540 529796
rect 156616 527066 156644 529108
rect 156604 527060 156656 527066
rect 156604 527002 156656 527008
rect 166276 526998 166304 529108
rect 175936 527134 175964 529108
rect 176120 527134 176148 548270
rect 175924 527128 175976 527134
rect 175924 527070 175976 527076
rect 176108 527128 176160 527134
rect 176108 527070 176160 527076
rect 177316 526998 177344 550598
rect 182086 539472 182142 539481
rect 182086 539407 182142 539416
rect 178038 538792 178094 538801
rect 178038 538727 178094 538736
rect 178052 529922 178080 538727
rect 178040 529916 178092 529922
rect 178040 529858 178092 529864
rect 182100 529786 182128 539407
rect 182088 529780 182140 529786
rect 182088 529722 182140 529728
rect 182836 527066 182864 550666
rect 183664 538214 183692 550734
rect 193956 550724 194008 550730
rect 193956 550666 194008 550672
rect 184296 550656 184348 550662
rect 184296 550598 184348 550604
rect 184308 548978 184336 550598
rect 193968 548978 193996 550666
rect 184308 548950 184644 548978
rect 193968 548950 194304 548978
rect 203964 548270 204300 548298
rect 204272 547126 204300 548270
rect 204260 547120 204312 547126
rect 204260 547062 204312 547068
rect 183664 538186 184244 538214
rect 184216 529666 184244 538186
rect 184216 529638 184644 529666
rect 194304 529094 194548 529122
rect 194520 527066 194548 529094
rect 203628 529094 203964 529122
rect 203628 527134 203656 529094
rect 203616 527128 203668 527134
rect 203616 527070 203668 527076
rect 182824 527060 182876 527066
rect 182824 527002 182876 527008
rect 194508 527060 194560 527066
rect 194508 527002 194560 527008
rect 166264 526992 166316 526998
rect 166264 526934 166316 526940
rect 177304 526992 177356 526998
rect 177304 526934 177356 526940
rect 165712 523184 165764 523190
rect 165712 523126 165764 523132
rect 175464 523184 175516 523190
rect 175464 523126 175516 523132
rect 193680 523184 193732 523190
rect 193680 523126 193732 523132
rect 203524 523184 203576 523190
rect 203524 523126 203576 523132
rect 156328 523116 156380 523122
rect 156328 523058 156380 523064
rect 156340 521914 156368 523058
rect 156032 521886 156368 521914
rect 165724 521778 165752 523126
rect 175372 523048 175424 523054
rect 175372 522990 175424 522996
rect 175384 521778 175412 522990
rect 165692 521750 165752 521778
rect 175352 521750 175412 521778
rect 155868 520328 155920 520334
rect 155868 520270 155920 520276
rect 155880 518906 155908 520270
rect 154488 518900 154540 518906
rect 154488 518842 154540 518848
rect 155868 518900 155920 518906
rect 155868 518842 155920 518848
rect 154500 512281 154528 518842
rect 154486 512272 154542 512281
rect 154486 512207 154542 512216
rect 175476 502738 175504 523126
rect 178684 523116 178736 523122
rect 178684 523058 178736 523064
rect 177304 523048 177356 523054
rect 177304 522990 177356 522996
rect 175352 502710 175504 502738
rect 156032 502030 156092 502058
rect 165692 502030 166028 502058
rect 156064 500818 156092 502030
rect 166000 500954 166028 502030
rect 177316 500954 177344 522990
rect 178038 511592 178094 511601
rect 178038 511527 178094 511536
rect 178052 503674 178080 511527
rect 178040 503668 178092 503674
rect 178040 503610 178092 503616
rect 178696 500954 178724 523058
rect 193692 521900 193720 523126
rect 203340 523048 203392 523054
rect 203340 522990 203392 522996
rect 203352 521900 203380 522990
rect 183664 521206 184046 521234
rect 182086 512272 182142 512281
rect 182086 512207 182142 512216
rect 182100 503674 182128 512207
rect 182088 503668 182140 503674
rect 182088 503610 182140 503616
rect 165988 500948 166040 500954
rect 165988 500890 166040 500896
rect 177304 500948 177356 500954
rect 177304 500890 177356 500896
rect 178684 500948 178736 500954
rect 178684 500890 178736 500896
rect 183664 500886 183692 521206
rect 203536 502738 203564 523126
rect 203366 502710 203564 502738
rect 184032 500954 184060 502044
rect 184020 500948 184072 500954
rect 184020 500890 184072 500896
rect 193692 500886 193720 502044
rect 183652 500880 183704 500886
rect 183652 500822 183704 500828
rect 193680 500880 193732 500886
rect 193680 500822 193732 500828
rect 156052 500812 156104 500818
rect 156052 500754 156104 500760
rect 184204 497004 184256 497010
rect 184204 496946 184256 496952
rect 156604 496936 156656 496942
rect 156604 496878 156656 496884
rect 182824 496936 182876 496942
rect 182824 496878 182876 496884
rect 156616 494972 156644 496878
rect 166264 496868 166316 496874
rect 166264 496810 166316 496816
rect 177304 496868 177356 496874
rect 177304 496810 177356 496816
rect 166276 494972 166304 496810
rect 175950 494278 176148 494306
rect 154486 485480 154542 485489
rect 154486 485415 154542 485424
rect 154500 475998 154528 485415
rect 154488 475992 154540 475998
rect 154488 475934 154540 475940
rect 156616 473278 156644 475116
rect 156604 473272 156656 473278
rect 156604 473214 156656 473220
rect 166276 473210 166304 475116
rect 175936 473346 175964 475116
rect 176120 473346 176148 494278
rect 175924 473340 175976 473346
rect 175924 473282 175976 473288
rect 176108 473340 176160 473346
rect 176108 473282 176160 473288
rect 177316 473210 177344 496810
rect 182086 485480 182142 485489
rect 182086 485415 182142 485424
rect 178038 484800 178094 484809
rect 178038 484735 178094 484744
rect 178052 476066 178080 484735
rect 178040 476060 178092 476066
rect 178040 476002 178092 476008
rect 182100 475930 182128 485415
rect 182088 475924 182140 475930
rect 182088 475866 182140 475872
rect 182836 473278 182864 496878
rect 184216 475674 184244 496946
rect 193956 496936 194008 496942
rect 193956 496878 194008 496884
rect 184296 496868 184348 496874
rect 184296 496810 184348 496816
rect 184308 494986 184336 496810
rect 193968 494986 193996 496878
rect 184308 494958 184644 494986
rect 193968 494958 194304 494986
rect 203964 494278 204300 494306
rect 204272 492114 204300 494278
rect 204260 492108 204312 492114
rect 204260 492050 204312 492056
rect 184216 475646 184644 475674
rect 194304 475102 194548 475130
rect 194520 473278 194548 475102
rect 203628 475102 203964 475130
rect 203628 473346 203656 475102
rect 203616 473340 203668 473346
rect 203616 473282 203668 473288
rect 182824 473272 182876 473278
rect 182824 473214 182876 473220
rect 194508 473272 194560 473278
rect 194508 473214 194560 473220
rect 166264 473204 166316 473210
rect 166264 473146 166316 473152
rect 177304 473204 177356 473210
rect 177304 473146 177356 473152
rect 165712 469396 165764 469402
rect 165712 469338 165764 469344
rect 175464 469396 175516 469402
rect 175464 469338 175516 469344
rect 193680 469396 193732 469402
rect 193680 469338 193732 469344
rect 203524 469396 203576 469402
rect 203524 469338 203576 469344
rect 156328 469328 156380 469334
rect 156328 469270 156380 469276
rect 156340 467922 156368 469270
rect 156032 467894 156368 467922
rect 165724 467786 165752 469338
rect 175372 469260 175424 469266
rect 175372 469202 175424 469208
rect 175384 467786 175412 469202
rect 165692 467758 165752 467786
rect 175352 467758 175412 467786
rect 154488 466540 154540 466546
rect 154488 466482 154540 466488
rect 154500 458289 154528 466482
rect 154486 458280 154542 458289
rect 154486 458215 154542 458224
rect 175476 448746 175504 469338
rect 178684 469328 178736 469334
rect 178684 469270 178736 469276
rect 177304 469260 177356 469266
rect 177304 469202 177356 469208
rect 175352 448718 175504 448746
rect 156032 448038 156092 448066
rect 165692 448038 166028 448066
rect 156064 445602 156092 448038
rect 166000 445738 166028 448038
rect 177316 445738 177344 469202
rect 178040 466472 178092 466478
rect 178040 466414 178092 466420
rect 178052 457609 178080 466414
rect 178038 457600 178094 457609
rect 178038 457535 178094 457544
rect 178696 445738 178724 469270
rect 193692 467908 193720 469338
rect 203340 469260 203392 469266
rect 203340 469202 203392 469208
rect 203352 467908 203380 469202
rect 183664 467214 184046 467242
rect 182088 466608 182140 466614
rect 182088 466550 182140 466556
rect 182100 458289 182128 466550
rect 182086 458280 182142 458289
rect 182086 458215 182142 458224
rect 165988 445732 166040 445738
rect 165988 445674 166040 445680
rect 177304 445732 177356 445738
rect 177304 445674 177356 445680
rect 178684 445732 178736 445738
rect 178684 445674 178736 445680
rect 183664 445670 183692 467214
rect 203536 448746 203564 469338
rect 203366 448718 203564 448746
rect 184032 445738 184060 448052
rect 184020 445732 184072 445738
rect 184020 445674 184072 445680
rect 193692 445670 193720 448052
rect 183652 445664 183704 445670
rect 183652 445606 183704 445612
rect 193680 445664 193732 445670
rect 193680 445606 193732 445612
rect 156052 445596 156104 445602
rect 156052 445538 156104 445544
rect 183652 443148 183704 443154
rect 183652 443090 183704 443096
rect 156604 443080 156656 443086
rect 156604 443022 156656 443028
rect 182824 443080 182876 443086
rect 182824 443022 182876 443028
rect 156616 440980 156644 443022
rect 166264 443012 166316 443018
rect 166264 442954 166316 442960
rect 177304 443012 177356 443018
rect 177304 442954 177356 442960
rect 166276 440980 166304 442954
rect 154488 440292 154540 440298
rect 175950 440286 176148 440314
rect 154488 440234 154540 440240
rect 154500 431497 154528 440234
rect 154486 431488 154542 431497
rect 154486 431423 154542 431432
rect 156616 419422 156644 421124
rect 156604 419416 156656 419422
rect 156604 419358 156656 419364
rect 166276 419354 166304 421124
rect 175936 419490 175964 421124
rect 176120 419490 176148 440286
rect 175924 419484 175976 419490
rect 175924 419426 175976 419432
rect 176108 419484 176160 419490
rect 176108 419426 176160 419432
rect 177316 419354 177344 442954
rect 182086 431488 182142 431497
rect 182086 431423 182142 431432
rect 178038 430808 178094 430817
rect 178038 430743 178094 430752
rect 178052 422278 178080 430743
rect 182100 422278 182128 431423
rect 178040 422272 178092 422278
rect 178040 422214 178092 422220
rect 182088 422272 182140 422278
rect 182088 422214 182140 422220
rect 182836 419422 182864 443022
rect 183664 441614 183692 443090
rect 193956 443080 194008 443086
rect 193956 443022 194008 443028
rect 184296 443012 184348 443018
rect 184296 442954 184348 442960
rect 183664 441586 184244 441614
rect 184216 421682 184244 441586
rect 184308 440994 184336 442954
rect 193968 440994 193996 443022
rect 184308 440966 184644 440994
rect 193968 440966 194304 440994
rect 203964 440286 204300 440314
rect 204272 436150 204300 440286
rect 204260 436144 204312 436150
rect 204260 436086 204312 436092
rect 184216 421654 184644 421682
rect 194304 421110 194548 421138
rect 194520 419422 194548 421110
rect 203628 421110 203964 421138
rect 203628 419490 203656 421110
rect 203616 419484 203668 419490
rect 203616 419426 203668 419432
rect 182824 419416 182876 419422
rect 182824 419358 182876 419364
rect 194508 419416 194560 419422
rect 194508 419358 194560 419364
rect 166264 419348 166316 419354
rect 166264 419290 166316 419296
rect 177304 419348 177356 419354
rect 177304 419290 177356 419296
rect 165712 415608 165764 415614
rect 165712 415550 165764 415556
rect 175464 415608 175516 415614
rect 175464 415550 175516 415556
rect 193680 415608 193732 415614
rect 193680 415550 193732 415556
rect 203524 415608 203576 415614
rect 203524 415550 203576 415556
rect 156328 415540 156380 415546
rect 156328 415482 156380 415488
rect 156340 413930 156368 415482
rect 156032 413902 156368 413930
rect 165724 413794 165752 415550
rect 175372 415472 175424 415478
rect 175372 415414 175424 415420
rect 175384 413794 175412 415414
rect 165692 413766 165752 413794
rect 175352 413766 175412 413794
rect 154486 404288 154542 404297
rect 154486 404223 154542 404232
rect 154500 394534 154528 404223
rect 155868 395344 155920 395350
rect 155868 395286 155920 395292
rect 155880 394754 155908 395286
rect 175476 394754 175504 415550
rect 178684 415540 178736 415546
rect 178684 415482 178736 415488
rect 177304 415472 177356 415478
rect 177304 415414 177356 415420
rect 155880 394726 156032 394754
rect 175352 394726 175504 394754
rect 154488 394528 154540 394534
rect 154488 394470 154540 394476
rect 165692 394046 166028 394074
rect 166000 391950 166028 394046
rect 177316 391950 177344 415414
rect 178038 403608 178094 403617
rect 178038 403543 178094 403552
rect 178052 394670 178080 403543
rect 178040 394664 178092 394670
rect 178040 394606 178092 394612
rect 178696 391950 178724 415482
rect 193692 413916 193720 415550
rect 203340 415472 203392 415478
rect 203340 415414 203392 415420
rect 203352 413916 203380 415414
rect 183664 413222 184046 413250
rect 182086 404288 182142 404297
rect 182086 404223 182142 404232
rect 182100 394602 182128 404223
rect 182088 394596 182140 394602
rect 182088 394538 182140 394544
rect 165988 391944 166040 391950
rect 165988 391886 166040 391892
rect 177304 391944 177356 391950
rect 177304 391886 177356 391892
rect 178684 391944 178736 391950
rect 178684 391886 178736 391892
rect 183664 391882 183692 413222
rect 203536 394754 203564 415550
rect 203366 394726 203564 394754
rect 184032 391950 184060 394060
rect 184020 391944 184072 391950
rect 184020 391886 184072 391892
rect 193692 391882 193720 394060
rect 183652 391876 183704 391882
rect 183652 391818 183704 391824
rect 193680 391876 193732 391882
rect 193680 391818 193732 391824
rect 183652 389360 183704 389366
rect 183652 389302 183704 389308
rect 156604 389292 156656 389298
rect 156604 389234 156656 389240
rect 182824 389292 182876 389298
rect 182824 389234 182876 389240
rect 156616 386852 156644 389234
rect 166264 389224 166316 389230
rect 166264 389166 166316 389172
rect 177304 389224 177356 389230
rect 177304 389166 177356 389172
rect 166276 386852 166304 389166
rect 154488 386504 154540 386510
rect 154488 386446 154540 386452
rect 154500 377505 154528 386446
rect 175950 386294 176148 386322
rect 154486 377496 154542 377505
rect 154486 377431 154542 377440
rect 156616 365634 156644 367132
rect 156604 365628 156656 365634
rect 156604 365570 156656 365576
rect 166276 365566 166304 367132
rect 175936 365702 175964 367132
rect 176120 365702 176148 386294
rect 175924 365696 175976 365702
rect 175924 365638 175976 365644
rect 176108 365696 176160 365702
rect 176108 365638 176160 365644
rect 177316 365566 177344 389166
rect 182088 386572 182140 386578
rect 182088 386514 182140 386520
rect 178040 386436 178092 386442
rect 178040 386378 178092 386384
rect 178052 376825 178080 386378
rect 182100 377505 182128 386514
rect 182086 377496 182142 377505
rect 182086 377431 182142 377440
rect 178038 376816 178094 376825
rect 178038 376751 178094 376760
rect 182836 365634 182864 389234
rect 183664 383654 183692 389302
rect 193956 389292 194008 389298
rect 193956 389234 194008 389240
rect 184296 389224 184348 389230
rect 184296 389166 184348 389172
rect 184308 386866 184336 389166
rect 193968 386866 193996 389234
rect 184308 386838 184644 386866
rect 193968 386838 194304 386866
rect 203964 386430 204300 386458
rect 204076 385076 204128 385082
rect 204076 385018 204128 385024
rect 183664 383626 184244 383654
rect 184216 367690 184244 383626
rect 184216 367662 184644 367690
rect 194304 367118 194548 367146
rect 194520 365634 194548 367118
rect 203628 367118 203964 367146
rect 203628 365702 203656 367118
rect 203616 365696 203668 365702
rect 203616 365638 203668 365644
rect 204088 365634 204116 385018
rect 204272 385014 204300 386430
rect 204260 385008 204312 385014
rect 204260 384950 204312 384956
rect 182824 365628 182876 365634
rect 182824 365570 182876 365576
rect 194508 365628 194560 365634
rect 194508 365570 194560 365576
rect 204076 365628 204128 365634
rect 204076 365570 204128 365576
rect 166264 365560 166316 365566
rect 166264 365502 166316 365508
rect 177304 365560 177356 365566
rect 177304 365502 177356 365508
rect 165712 361752 165764 361758
rect 165712 361694 165764 361700
rect 175464 361752 175516 361758
rect 175464 361694 175516 361700
rect 193680 361752 193732 361758
rect 193680 361694 193732 361700
rect 203524 361752 203576 361758
rect 203524 361694 203576 361700
rect 156328 361684 156380 361690
rect 156328 361626 156380 361632
rect 156340 359938 156368 361626
rect 156032 359910 156368 359938
rect 165724 359802 165752 361694
rect 175372 361616 175424 361622
rect 175372 361558 175424 361564
rect 175384 359802 175412 361558
rect 165692 359774 165752 359802
rect 175352 359774 175412 359802
rect 154486 350296 154542 350305
rect 154486 350231 154542 350240
rect 154500 340814 154528 350231
rect 154488 340808 154540 340814
rect 175476 340762 175504 361694
rect 178684 361684 178736 361690
rect 178684 361626 178736 361632
rect 177304 361616 177356 361622
rect 177304 361558 177356 361564
rect 154488 340750 154540 340756
rect 175352 340734 175504 340762
rect 156032 340054 156092 340082
rect 165692 340054 166028 340082
rect 156064 337958 156092 340054
rect 166000 338094 166028 340054
rect 177316 338094 177344 361558
rect 178038 349616 178094 349625
rect 178038 349551 178094 349560
rect 178052 340882 178080 349551
rect 178040 340876 178092 340882
rect 178040 340818 178092 340824
rect 178696 338094 178724 361626
rect 193692 359924 193720 361694
rect 203340 361616 203392 361622
rect 203340 361558 203392 361564
rect 203352 359924 203380 361558
rect 183664 359230 184046 359258
rect 182086 350296 182142 350305
rect 182086 350231 182142 350240
rect 182100 340746 182128 350231
rect 182088 340740 182140 340746
rect 182088 340682 182140 340688
rect 165988 338088 166040 338094
rect 165988 338030 166040 338036
rect 177304 338088 177356 338094
rect 177304 338030 177356 338036
rect 178684 338088 178736 338094
rect 178684 338030 178736 338036
rect 183664 338026 183692 359230
rect 203536 340762 203564 361694
rect 203366 340734 203564 340762
rect 184032 338094 184060 340068
rect 184020 338088 184072 338094
rect 184020 338030 184072 338036
rect 193692 338026 193720 340068
rect 183652 338020 183704 338026
rect 183652 337962 183704 337968
rect 193680 338020 193732 338026
rect 193680 337962 193732 337968
rect 156052 337952 156104 337958
rect 156052 337894 156104 337900
rect 183652 335504 183704 335510
rect 183652 335446 183704 335452
rect 156604 335436 156656 335442
rect 156604 335378 156656 335384
rect 182824 335436 182876 335442
rect 182824 335378 182876 335384
rect 156616 332860 156644 335378
rect 166264 335368 166316 335374
rect 166264 335310 166316 335316
rect 177304 335368 177356 335374
rect 177304 335310 177356 335316
rect 166276 332860 166304 335310
rect 175950 332302 176148 332330
rect 154486 322960 154542 322969
rect 154486 322895 154542 322904
rect 154500 314566 154528 322895
rect 154488 314560 154540 314566
rect 154488 314502 154540 314508
rect 156616 311778 156644 313140
rect 156604 311772 156656 311778
rect 156604 311714 156656 311720
rect 166276 311710 166304 313140
rect 175936 311846 175964 313140
rect 176120 311846 176148 332302
rect 175924 311840 175976 311846
rect 175924 311782 175976 311788
rect 176108 311840 176160 311846
rect 176108 311782 176160 311788
rect 177316 311710 177344 335310
rect 182086 322960 182142 322969
rect 182086 322895 182142 322904
rect 178038 322144 178094 322153
rect 178038 322079 178094 322088
rect 178052 314634 178080 322079
rect 182100 314634 182128 322895
rect 178040 314628 178092 314634
rect 178040 314570 178092 314576
rect 182088 314628 182140 314634
rect 182088 314570 182140 314576
rect 182836 311778 182864 335378
rect 183664 325694 183692 335446
rect 193956 335436 194008 335442
rect 193956 335378 194008 335384
rect 184296 335368 184348 335374
rect 184296 335310 184348 335316
rect 184308 332874 184336 335310
rect 193968 332874 193996 335378
rect 184308 332846 184644 332874
rect 193968 332846 194304 332874
rect 203964 332302 204300 332330
rect 204076 331288 204128 331294
rect 204076 331230 204128 331236
rect 183664 325666 184244 325694
rect 184216 313698 184244 325666
rect 184216 313670 184644 313698
rect 194304 313126 194548 313154
rect 194520 311778 194548 313126
rect 203628 313126 203964 313154
rect 203628 311846 203656 313126
rect 203616 311840 203668 311846
rect 203616 311782 203668 311788
rect 204088 311778 204116 331230
rect 204272 329050 204300 332302
rect 204260 329044 204312 329050
rect 204260 328986 204312 328992
rect 182824 311772 182876 311778
rect 182824 311714 182876 311720
rect 194508 311772 194560 311778
rect 194508 311714 194560 311720
rect 204076 311772 204128 311778
rect 204076 311714 204128 311720
rect 166264 311704 166316 311710
rect 166264 311646 166316 311652
rect 177304 311704 177356 311710
rect 177304 311646 177356 311652
rect 165620 307964 165672 307970
rect 165620 307906 165672 307912
rect 175464 307964 175516 307970
rect 175464 307906 175516 307912
rect 193680 307964 193732 307970
rect 193680 307906 193732 307912
rect 203524 307964 203576 307970
rect 203524 307906 203576 307912
rect 156328 307896 156380 307902
rect 156328 307838 156380 307844
rect 156340 305946 156368 307838
rect 165632 306082 165660 307906
rect 175280 307828 175332 307834
rect 175280 307770 175332 307776
rect 175292 306082 175320 307770
rect 165632 306054 165706 306082
rect 175292 306054 175366 306082
rect 156032 305918 156368 305946
rect 165678 305932 165706 306054
rect 175338 305932 175366 306054
rect 154486 296304 154542 296313
rect 154486 296239 154542 296248
rect 154500 287026 154528 296239
rect 154488 287020 154540 287026
rect 154488 286962 154540 286968
rect 175476 286770 175504 307906
rect 178684 307896 178736 307902
rect 178684 307838 178736 307844
rect 177304 307828 177356 307834
rect 177304 307770 177356 307776
rect 175352 286742 175504 286770
rect 156032 286062 156092 286090
rect 165692 286062 166028 286090
rect 156064 284170 156092 286062
rect 166000 284306 166028 286062
rect 177316 284306 177344 307770
rect 178038 295624 178094 295633
rect 178038 295559 178094 295568
rect 178052 286890 178080 295559
rect 178040 286884 178092 286890
rect 178040 286826 178092 286832
rect 178696 284306 178724 307838
rect 193692 305932 193720 307906
rect 203340 307828 203392 307834
rect 203340 307770 203392 307776
rect 203352 305932 203380 307770
rect 183664 305238 184046 305266
rect 182086 296304 182142 296313
rect 182086 296239 182142 296248
rect 182100 286958 182128 296239
rect 182088 286952 182140 286958
rect 182088 286894 182140 286900
rect 165988 284300 166040 284306
rect 165988 284242 166040 284248
rect 177304 284300 177356 284306
rect 177304 284242 177356 284248
rect 178684 284300 178736 284306
rect 178684 284242 178736 284248
rect 183664 284238 183692 305238
rect 203536 286770 203564 307906
rect 203366 286742 203564 286770
rect 184032 284306 184060 286076
rect 184020 284300 184072 284306
rect 184020 284242 184072 284248
rect 193692 284238 193720 286076
rect 183652 284232 183704 284238
rect 183652 284174 183704 284180
rect 193680 284232 193732 284238
rect 193680 284174 193732 284180
rect 156052 284164 156104 284170
rect 156052 284106 156104 284112
rect 183652 280356 183704 280362
rect 183652 280298 183704 280304
rect 156604 280288 156656 280294
rect 156604 280230 156656 280236
rect 182824 280288 182876 280294
rect 182824 280230 182876 280236
rect 156616 278868 156644 280230
rect 166264 280220 166316 280226
rect 166264 280162 166316 280168
rect 177304 280220 177356 280226
rect 177304 280162 177356 280168
rect 166276 278868 166304 280162
rect 175950 278310 176148 278338
rect 154488 277500 154540 277506
rect 154488 277442 154540 277448
rect 154500 270065 154528 277442
rect 154486 270056 154542 270065
rect 154486 269991 154542 270000
rect 156616 256630 156644 259148
rect 156604 256624 156656 256630
rect 156604 256566 156656 256572
rect 166276 256562 166304 259148
rect 175936 256698 175964 259148
rect 176120 256698 176148 278310
rect 175924 256692 175976 256698
rect 175924 256634 175976 256640
rect 176108 256692 176160 256698
rect 176108 256634 176160 256640
rect 177316 256562 177344 280162
rect 178040 277568 178092 277574
rect 178040 277510 178092 277516
rect 182088 277568 182140 277574
rect 182088 277510 182140 277516
rect 178052 269113 178080 277510
rect 182100 270065 182128 277510
rect 182086 270056 182142 270065
rect 182086 269991 182142 270000
rect 178038 269104 178094 269113
rect 178038 269039 178094 269048
rect 182836 256630 182864 280230
rect 183664 267734 183692 280298
rect 193956 280288 194008 280294
rect 193956 280230 194008 280236
rect 184296 280220 184348 280226
rect 184296 280162 184348 280168
rect 184308 278882 184336 280162
rect 193968 278882 193996 280230
rect 184308 278854 184644 278882
rect 193968 278854 194304 278882
rect 203964 278310 204300 278338
rect 204076 277432 204128 277438
rect 204076 277374 204128 277380
rect 183664 267706 184244 267734
rect 184216 259706 184244 267706
rect 184216 259678 184644 259706
rect 194304 259134 194548 259162
rect 194520 256630 194548 259134
rect 203628 259134 203964 259162
rect 203628 256698 203656 259134
rect 203616 256692 203668 256698
rect 203616 256634 203668 256640
rect 204088 256630 204116 277374
rect 204272 272610 204300 278310
rect 204260 272604 204312 272610
rect 204260 272546 204312 272552
rect 182824 256624 182876 256630
rect 182824 256566 182876 256572
rect 194508 256624 194560 256630
rect 194508 256566 194560 256572
rect 204076 256624 204128 256630
rect 204076 256566 204128 256572
rect 166264 256556 166316 256562
rect 166264 256498 166316 256504
rect 177304 256556 177356 256562
rect 177304 256498 177356 256504
rect 165712 254108 165764 254114
rect 165712 254050 165764 254056
rect 175464 254108 175516 254114
rect 175464 254050 175516 254056
rect 193680 254108 193732 254114
rect 193680 254050 193732 254056
rect 203524 254108 203576 254114
rect 203524 254050 203576 254056
rect 156328 254040 156380 254046
rect 156328 253982 156380 253988
rect 156340 251954 156368 253982
rect 156032 251926 156368 251954
rect 165724 251818 165752 254050
rect 175372 253972 175424 253978
rect 175372 253914 175424 253920
rect 175384 251818 175412 253914
rect 165692 251790 165752 251818
rect 175352 251790 175412 251818
rect 154488 251252 154540 251258
rect 154488 251194 154540 251200
rect 154500 242321 154528 251194
rect 154486 242312 154542 242321
rect 154486 242247 154542 242256
rect 175476 232778 175504 254050
rect 178684 254040 178736 254046
rect 178684 253982 178736 253988
rect 177304 253972 177356 253978
rect 177304 253914 177356 253920
rect 175352 232750 175504 232778
rect 156032 232070 156092 232098
rect 165692 232070 166028 232098
rect 156064 230314 156092 232070
rect 166000 230450 166028 232070
rect 177316 230450 177344 253914
rect 178040 251320 178092 251326
rect 178040 251262 178092 251268
rect 178052 241641 178080 251262
rect 178038 241632 178094 241641
rect 178038 241567 178094 241576
rect 178696 230450 178724 253982
rect 193692 251940 193720 254050
rect 203340 253972 203392 253978
rect 203340 253914 203392 253920
rect 203352 251940 203380 253914
rect 182088 251320 182140 251326
rect 182088 251262 182140 251268
rect 182100 242321 182128 251262
rect 183664 251246 184046 251274
rect 182086 242312 182142 242321
rect 182086 242247 182142 242256
rect 165988 230444 166040 230450
rect 165988 230386 166040 230392
rect 177304 230444 177356 230450
rect 177304 230386 177356 230392
rect 178684 230444 178736 230450
rect 178684 230386 178736 230392
rect 183664 230382 183692 251246
rect 203536 232778 203564 254050
rect 203366 232750 203564 232778
rect 184032 230450 184060 232084
rect 184020 230444 184072 230450
rect 184020 230386 184072 230392
rect 193692 230382 193720 232084
rect 183652 230376 183704 230382
rect 183652 230318 183704 230324
rect 193680 230376 193732 230382
rect 193680 230318 193732 230324
rect 156052 230308 156104 230314
rect 156052 230250 156104 230256
rect 184204 226500 184256 226506
rect 184204 226442 184256 226448
rect 156604 226432 156656 226438
rect 156604 226374 156656 226380
rect 182824 226432 182876 226438
rect 182824 226374 182876 226380
rect 156616 224876 156644 226374
rect 166264 226364 166316 226370
rect 166264 226306 166316 226312
rect 177304 226364 177356 226370
rect 177304 226306 177356 226312
rect 166276 224876 166304 226306
rect 175950 224318 176148 224346
rect 154488 223712 154540 223718
rect 154488 223654 154540 223660
rect 154500 215393 154528 223654
rect 154486 215384 154542 215393
rect 154486 215319 154542 215328
rect 156616 202774 156644 205020
rect 156604 202768 156656 202774
rect 156604 202710 156656 202716
rect 166276 202706 166304 205020
rect 175936 202842 175964 205020
rect 176120 202842 176148 224318
rect 175924 202836 175976 202842
rect 175924 202778 175976 202784
rect 176108 202836 176160 202842
rect 176108 202778 176160 202784
rect 177316 202706 177344 226306
rect 182088 223780 182140 223786
rect 182088 223722 182140 223728
rect 178040 223644 178092 223650
rect 178040 223586 178092 223592
rect 178052 214713 178080 223586
rect 182100 215393 182128 223722
rect 182086 215384 182142 215393
rect 182086 215319 182142 215328
rect 178038 214704 178094 214713
rect 178038 214639 178094 214648
rect 182836 202774 182864 226374
rect 184216 205714 184244 226442
rect 193956 226432 194008 226438
rect 193956 226374 194008 226380
rect 184296 226364 184348 226370
rect 184296 226306 184348 226312
rect 184308 224890 184336 226306
rect 193968 224890 193996 226374
rect 184308 224862 184644 224890
rect 193968 224862 194304 224890
rect 203964 224318 204300 224346
rect 204272 221882 204300 224318
rect 204260 221876 204312 221882
rect 204260 221818 204312 221824
rect 184216 205686 184644 205714
rect 194304 205006 194548 205034
rect 194520 202774 194548 205006
rect 203628 205006 203964 205034
rect 203628 202842 203656 205006
rect 203616 202836 203668 202842
rect 203616 202778 203668 202784
rect 182824 202768 182876 202774
rect 182824 202710 182876 202716
rect 194508 202768 194560 202774
rect 194508 202710 194560 202716
rect 166264 202700 166316 202706
rect 166264 202642 166316 202648
rect 177304 202700 177356 202706
rect 177304 202642 177356 202648
rect 165620 200320 165672 200326
rect 165620 200262 165672 200268
rect 175464 200320 175516 200326
rect 175464 200262 175516 200268
rect 193680 200320 193732 200326
rect 193680 200262 193732 200268
rect 203524 200320 203576 200326
rect 203524 200262 203576 200268
rect 156328 200252 156380 200258
rect 156328 200194 156380 200200
rect 156340 197962 156368 200194
rect 165632 198234 165660 200262
rect 175280 200184 175332 200190
rect 175280 200126 175332 200132
rect 175292 198234 175320 200126
rect 165632 198206 165706 198234
rect 175292 198206 175366 198234
rect 156032 197934 156368 197962
rect 165678 197948 165706 198206
rect 175338 197948 175366 198206
rect 154486 188320 154542 188329
rect 154486 188255 154542 188264
rect 154500 179314 154528 188255
rect 154488 179308 154540 179314
rect 154488 179250 154540 179256
rect 175476 178786 175504 200262
rect 178684 200252 178736 200258
rect 178684 200194 178736 200200
rect 177304 200184 177356 200190
rect 177304 200126 177356 200132
rect 175352 178758 175504 178786
rect 156032 178078 156092 178106
rect 165692 178078 166028 178106
rect 156064 176526 156092 178078
rect 166000 176662 166028 178078
rect 177316 176662 177344 200126
rect 178038 187640 178094 187649
rect 178038 187575 178094 187584
rect 178052 179382 178080 187575
rect 178040 179376 178092 179382
rect 178040 179318 178092 179324
rect 178696 176662 178724 200194
rect 193692 197948 193720 200262
rect 203340 200184 203392 200190
rect 203340 200126 203392 200132
rect 203352 197948 203380 200126
rect 183664 197254 184046 197282
rect 182086 188320 182142 188329
rect 182086 188255 182142 188264
rect 182100 179246 182128 188255
rect 182088 179240 182140 179246
rect 182088 179182 182140 179188
rect 165988 176656 166040 176662
rect 165988 176598 166040 176604
rect 177304 176656 177356 176662
rect 177304 176598 177356 176604
rect 178684 176656 178736 176662
rect 178684 176598 178736 176604
rect 183664 176594 183692 197254
rect 203536 178786 203564 200262
rect 203366 178758 203564 178786
rect 184032 176662 184060 178092
rect 184020 176656 184072 176662
rect 184020 176598 184072 176604
rect 193692 176594 193720 178092
rect 183652 176588 183704 176594
rect 183652 176530 183704 176536
rect 193680 176588 193732 176594
rect 193680 176530 193732 176536
rect 156052 176520 156104 176526
rect 156052 176462 156104 176468
rect 183652 172712 183704 172718
rect 183652 172654 183704 172660
rect 156604 172644 156656 172650
rect 156604 172586 156656 172592
rect 182824 172644 182876 172650
rect 182824 172586 182876 172592
rect 156616 170884 156644 172586
rect 166264 172576 166316 172582
rect 166264 172518 166316 172524
rect 177304 172576 177356 172582
rect 177304 172518 177356 172524
rect 166276 170884 166304 172518
rect 175950 170326 176148 170354
rect 154486 161392 154542 161401
rect 154486 161327 154542 161336
rect 154500 151706 154528 161327
rect 154488 151700 154540 151706
rect 154488 151642 154540 151648
rect 156616 148986 156644 151028
rect 156604 148980 156656 148986
rect 156604 148922 156656 148928
rect 166276 148918 166304 151028
rect 175936 149054 175964 151028
rect 176120 149054 176148 170326
rect 175924 149048 175976 149054
rect 175924 148990 175976 148996
rect 176108 149048 176160 149054
rect 176108 148990 176160 148996
rect 177316 148918 177344 172518
rect 182086 161392 182142 161401
rect 182086 161327 182142 161336
rect 178038 160712 178094 160721
rect 178038 160647 178094 160656
rect 178052 151774 178080 160647
rect 178040 151768 178092 151774
rect 178040 151710 178092 151716
rect 182100 151638 182128 161327
rect 182088 151632 182140 151638
rect 182088 151574 182140 151580
rect 182836 148986 182864 172586
rect 183664 171134 183692 172654
rect 193956 172644 194008 172650
rect 193956 172586 194008 172592
rect 184296 172576 184348 172582
rect 184296 172518 184348 172524
rect 183664 171106 184244 171134
rect 184216 151722 184244 171106
rect 184308 170898 184336 172518
rect 193968 170898 193996 172586
rect 184308 170870 184644 170898
rect 193968 170870 194304 170898
rect 203964 170326 204300 170354
rect 204272 165918 204300 170326
rect 204260 165912 204312 165918
rect 204260 165854 204312 165860
rect 184216 151694 184644 151722
rect 194304 151014 194548 151042
rect 194520 148986 194548 151014
rect 203628 151014 203964 151042
rect 203628 149054 203656 151014
rect 203616 149048 203668 149054
rect 203616 148990 203668 148996
rect 182824 148980 182876 148986
rect 182824 148922 182876 148928
rect 194508 148980 194560 148986
rect 194508 148922 194560 148928
rect 166264 148912 166316 148918
rect 166264 148854 166316 148860
rect 177304 148912 177356 148918
rect 177304 148854 177356 148860
rect 165712 146464 165764 146470
rect 165712 146406 165764 146412
rect 175464 146464 175516 146470
rect 175464 146406 175516 146412
rect 193680 146464 193732 146470
rect 193680 146406 193732 146412
rect 203524 146464 203576 146470
rect 203524 146406 203576 146412
rect 156328 146396 156380 146402
rect 156328 146338 156380 146344
rect 156340 143970 156368 146338
rect 156032 143942 156368 143970
rect 165724 143834 165752 146406
rect 175372 146328 175424 146334
rect 175372 146270 175424 146276
rect 175384 143834 175412 146270
rect 165692 143806 165752 143834
rect 175352 143806 175412 143834
rect 154486 134328 154542 134337
rect 154486 134263 154542 134272
rect 154500 125526 154528 134263
rect 154488 125520 154540 125526
rect 154488 125462 154540 125468
rect 175476 124794 175504 146406
rect 178684 146396 178736 146402
rect 178684 146338 178736 146344
rect 177304 146328 177356 146334
rect 177304 146270 177356 146276
rect 175352 124766 175504 124794
rect 156018 123842 156046 124100
rect 165692 124086 166028 124114
rect 155972 123814 156046 123842
rect 155972 122670 156000 123814
rect 166000 122806 166028 124086
rect 177316 122806 177344 146270
rect 178038 133648 178094 133657
rect 178038 133583 178094 133592
rect 178052 125594 178080 133583
rect 178040 125588 178092 125594
rect 178040 125530 178092 125536
rect 178696 122806 178724 146338
rect 193692 143956 193720 146406
rect 203340 146328 203392 146334
rect 203340 146270 203392 146276
rect 203352 143956 203380 146270
rect 183664 143262 184046 143290
rect 182086 134328 182142 134337
rect 182086 134263 182142 134272
rect 182100 125458 182128 134263
rect 182088 125452 182140 125458
rect 182088 125394 182140 125400
rect 165988 122800 166040 122806
rect 165988 122742 166040 122748
rect 177304 122800 177356 122806
rect 177304 122742 177356 122748
rect 178684 122800 178736 122806
rect 178684 122742 178736 122748
rect 183664 122738 183692 143262
rect 203536 124794 203564 146406
rect 203366 124766 203564 124794
rect 184032 122806 184060 124100
rect 184020 122800 184072 122806
rect 184020 122742 184072 122748
rect 193692 122738 193720 124100
rect 183652 122732 183704 122738
rect 183652 122674 183704 122680
rect 193680 122732 193732 122738
rect 193680 122674 193732 122680
rect 155960 122664 156012 122670
rect 155960 122606 156012 122612
rect 183652 118856 183704 118862
rect 183652 118798 183704 118804
rect 156604 118788 156656 118794
rect 156604 118730 156656 118736
rect 182824 118788 182876 118794
rect 182824 118730 182876 118736
rect 156616 116892 156644 118730
rect 166264 118720 166316 118726
rect 166264 118662 166316 118668
rect 177304 118720 177356 118726
rect 177304 118662 177356 118668
rect 166276 116892 166304 118662
rect 175950 116334 176148 116362
rect 154486 107400 154542 107409
rect 154486 107335 154542 107344
rect 154500 97986 154528 107335
rect 154488 97980 154540 97986
rect 154488 97922 154540 97928
rect 156616 95130 156644 97036
rect 156604 95124 156656 95130
rect 156604 95066 156656 95072
rect 166276 95062 166304 97036
rect 175936 95198 175964 97036
rect 176120 95198 176148 116334
rect 175924 95192 175976 95198
rect 175924 95134 175976 95140
rect 176108 95192 176160 95198
rect 176108 95134 176160 95140
rect 177316 95062 177344 118662
rect 182086 107400 182142 107409
rect 182086 107335 182142 107344
rect 178038 106720 178094 106729
rect 178038 106655 178094 106664
rect 178052 97918 178080 106655
rect 182100 97918 182128 107335
rect 178040 97912 178092 97918
rect 178040 97854 178092 97860
rect 182088 97912 182140 97918
rect 182088 97854 182140 97860
rect 182836 95130 182864 118730
rect 183664 113174 183692 118798
rect 193956 118788 194008 118794
rect 193956 118730 194008 118736
rect 184296 118720 184348 118726
rect 184296 118662 184348 118668
rect 184308 116906 184336 118662
rect 193968 116906 193996 118730
rect 184308 116878 184644 116906
rect 193968 116878 194304 116906
rect 203964 116334 204300 116362
rect 204272 114782 204300 116334
rect 204260 114776 204312 114782
rect 204260 114718 204312 114724
rect 183664 113146 184244 113174
rect 184216 97730 184244 113146
rect 184216 97702 184644 97730
rect 194304 97022 194548 97050
rect 194520 95130 194548 97022
rect 203628 97022 203964 97050
rect 203628 95198 203656 97022
rect 203616 95192 203668 95198
rect 203616 95134 203668 95140
rect 182824 95124 182876 95130
rect 182824 95066 182876 95072
rect 194508 95124 194560 95130
rect 194508 95066 194560 95072
rect 166264 95056 166316 95062
rect 166264 94998 166316 95004
rect 177304 95056 177356 95062
rect 177304 94998 177356 95004
rect 165712 91248 165764 91254
rect 165712 91190 165764 91196
rect 175464 91248 175516 91254
rect 175464 91190 175516 91196
rect 193680 91248 193732 91254
rect 193680 91190 193732 91196
rect 203524 91248 203576 91254
rect 203524 91190 203576 91196
rect 156328 91180 156380 91186
rect 156328 91122 156380 91128
rect 156340 89978 156368 91122
rect 156032 89950 156368 89978
rect 165724 89842 165752 91190
rect 175372 91112 175424 91118
rect 175372 91054 175424 91060
rect 175384 89842 175412 91054
rect 165692 89814 165752 89842
rect 175352 89814 175412 89842
rect 154488 88392 154540 88398
rect 154488 88334 154540 88340
rect 154500 80345 154528 88334
rect 154486 80336 154542 80345
rect 154486 80271 154542 80280
rect 175476 70666 175504 91190
rect 178684 91180 178736 91186
rect 178684 91122 178736 91128
rect 177304 91112 177356 91118
rect 177304 91054 177356 91060
rect 175352 70638 175504 70666
rect 156032 70094 156092 70122
rect 165692 70094 166028 70122
rect 156064 68882 156092 70094
rect 166000 69018 166028 70094
rect 177316 69018 177344 91054
rect 178038 79656 178094 79665
rect 178038 79591 178094 79600
rect 178052 71738 178080 79591
rect 178040 71732 178092 71738
rect 178040 71674 178092 71680
rect 178696 69018 178724 91122
rect 193692 89964 193720 91190
rect 203340 91112 203392 91118
rect 203340 91054 203392 91060
rect 203352 89964 203380 91054
rect 183664 89270 184046 89298
rect 182086 80336 182142 80345
rect 182086 80271 182142 80280
rect 182100 71738 182128 80271
rect 182088 71732 182140 71738
rect 182088 71674 182140 71680
rect 165988 69012 166040 69018
rect 165988 68954 166040 68960
rect 177304 69012 177356 69018
rect 177304 68954 177356 68960
rect 178684 69012 178736 69018
rect 178684 68954 178736 68960
rect 183664 68950 183692 89270
rect 203536 70666 203564 91190
rect 203366 70638 203564 70666
rect 184032 69018 184060 70108
rect 184020 69012 184072 69018
rect 184020 68954 184072 68960
rect 193692 68950 193720 70108
rect 183652 68944 183704 68950
rect 183652 68886 183704 68892
rect 193680 68944 193732 68950
rect 193680 68886 193732 68892
rect 156052 68876 156104 68882
rect 156052 68818 156104 68824
rect 183652 65068 183704 65074
rect 183652 65010 183704 65016
rect 156604 65000 156656 65006
rect 156604 64942 156656 64948
rect 182824 65000 182876 65006
rect 182824 64942 182876 64948
rect 156616 62900 156644 64942
rect 166264 64932 166316 64938
rect 166264 64874 166316 64880
rect 177304 64932 177356 64938
rect 177304 64874 177356 64880
rect 166276 62900 166304 64874
rect 175950 62206 176148 62234
rect 154488 62144 154540 62150
rect 154488 62086 154540 62092
rect 154500 53417 154528 62086
rect 154486 53408 154542 53417
rect 154486 53343 154542 53352
rect 153842 42120 153898 42129
rect 153842 42055 153898 42064
rect 156616 41342 156644 43044
rect 156604 41336 156656 41342
rect 156604 41278 156656 41284
rect 166276 41274 166304 43044
rect 175936 41410 175964 43044
rect 176120 41410 176148 62206
rect 175924 41404 175976 41410
rect 175924 41346 175976 41352
rect 176108 41404 176160 41410
rect 176108 41346 176160 41352
rect 177316 41274 177344 64874
rect 182086 53408 182142 53417
rect 182086 53343 182142 53352
rect 178038 52728 178094 52737
rect 178038 52663 178094 52672
rect 178052 44130 178080 52663
rect 182100 44130 182128 53343
rect 178040 44124 178092 44130
rect 178040 44066 178092 44072
rect 182088 44124 182140 44130
rect 182088 44066 182140 44072
rect 182836 41342 182864 64942
rect 183664 55214 183692 65010
rect 193956 65000 194008 65006
rect 193956 64942 194008 64948
rect 184296 64932 184348 64938
rect 184296 64874 184348 64880
rect 184308 62914 184336 64874
rect 193968 62914 193996 64942
rect 184308 62886 184644 62914
rect 193968 62886 194304 62914
rect 203964 62206 204300 62234
rect 204272 57934 204300 62206
rect 204260 57928 204312 57934
rect 204260 57870 204312 57876
rect 183664 55186 184244 55214
rect 184216 43738 184244 55186
rect 184216 43710 184644 43738
rect 194304 43030 194548 43058
rect 194520 41342 194548 43030
rect 203628 43030 203964 43058
rect 203628 41410 203656 43030
rect 203616 41404 203668 41410
rect 203616 41346 203668 41352
rect 182824 41336 182876 41342
rect 182824 41278 182876 41284
rect 194508 41336 194560 41342
rect 194508 41278 194560 41284
rect 152464 41268 152516 41274
rect 152464 41210 152516 41216
rect 166264 41268 166316 41274
rect 166264 41210 166316 41216
rect 177304 41268 177356 41274
rect 177304 41210 177356 41216
rect 204916 39438 204944 700402
rect 233884 700324 233936 700330
rect 233884 700266 233936 700272
rect 212356 686112 212408 686118
rect 212356 686054 212408 686060
rect 232688 686112 232740 686118
rect 232688 686054 232740 686060
rect 204996 685908 205048 685914
rect 204996 685850 205048 685856
rect 205008 662318 205036 685850
rect 212368 683890 212396 686054
rect 221372 686044 221424 686050
rect 221372 685986 221424 685992
rect 212060 683862 212396 683890
rect 221384 683890 221412 685986
rect 232596 685976 232648 685982
rect 232596 685918 232648 685924
rect 231032 685908 231084 685914
rect 231032 685850 231084 685856
rect 232504 685908 232556 685914
rect 232504 685850 232556 685856
rect 231044 683890 231072 685850
rect 221384 683862 221720 683890
rect 231044 683862 231380 683890
rect 205640 683188 205692 683194
rect 205640 683130 205692 683136
rect 205652 674121 205680 683130
rect 209686 674248 209742 674257
rect 209686 674183 209742 674192
rect 205638 674112 205694 674121
rect 205638 674047 205694 674056
rect 209700 665174 209728 674183
rect 209688 665168 209740 665174
rect 209688 665110 209740 665116
rect 211724 664006 212060 664034
rect 221720 664006 222056 664034
rect 231380 664006 231624 664034
rect 211724 662386 211752 664006
rect 211712 662380 211764 662386
rect 211712 662322 211764 662328
rect 222028 662318 222056 664006
rect 231596 663746 231624 664006
rect 231584 663740 231636 663746
rect 231584 663682 231636 663688
rect 232516 662318 232544 685850
rect 232608 663746 232636 685918
rect 232700 665310 232728 686054
rect 233240 683256 233292 683262
rect 233240 683198 233292 683204
rect 233252 673577 233280 683198
rect 233238 673568 233294 673577
rect 233238 673503 233294 673512
rect 232688 665304 232740 665310
rect 232688 665246 232740 665252
rect 232596 663740 232648 663746
rect 232596 663682 232648 663688
rect 204996 662312 205048 662318
rect 204996 662254 205048 662260
rect 222016 662312 222068 662318
rect 222016 662254 222068 662260
rect 232504 662312 232556 662318
rect 232504 662254 232556 662260
rect 222292 658436 222344 658442
rect 222292 658378 222344 658384
rect 222304 656948 222332 658378
rect 232504 658368 232556 658374
rect 232504 658310 232556 658316
rect 212368 656266 212658 656282
rect 210424 656260 210476 656266
rect 210424 656202 210476 656208
rect 212356 656260 212658 656266
rect 212408 656254 212658 656260
rect 231978 656254 232084 656282
rect 212356 656202 212408 656208
rect 205640 655648 205692 655654
rect 205640 655590 205692 655596
rect 204996 654356 205048 654362
rect 204996 654298 205048 654304
rect 205008 634778 205036 654298
rect 205652 646785 205680 655590
rect 209688 655580 209740 655586
rect 209688 655522 209740 655528
rect 209700 647465 209728 655522
rect 209686 647456 209742 647465
rect 209686 647391 209742 647400
rect 205638 646776 205694 646785
rect 205638 646711 205694 646720
rect 204996 634772 205048 634778
rect 204996 634714 205048 634720
rect 210436 634710 210464 656202
rect 212644 634710 212672 637092
rect 210424 634704 210476 634710
rect 210424 634646 210476 634652
rect 212632 634704 212684 634710
rect 212632 634646 212684 634652
rect 222304 634642 222332 637092
rect 231964 634778 231992 637092
rect 232056 634778 232084 656254
rect 231952 634772 232004 634778
rect 231952 634714 232004 634720
rect 232044 634772 232096 634778
rect 232044 634714 232096 634720
rect 232516 634710 232544 658310
rect 233240 655716 233292 655722
rect 233240 655658 233292 655664
rect 233252 646785 233280 655658
rect 233238 646776 233294 646785
rect 233238 646711 233294 646720
rect 232504 634704 232556 634710
rect 232504 634646 232556 634652
rect 222292 634636 222344 634642
rect 222292 634578 222344 634584
rect 212356 632324 212408 632330
rect 212356 632266 212408 632272
rect 232688 632324 232740 632330
rect 232688 632266 232740 632272
rect 204996 632120 205048 632126
rect 204996 632062 205048 632068
rect 205008 608530 205036 632062
rect 212368 629898 212396 632266
rect 221372 632256 221424 632262
rect 221372 632198 221424 632204
rect 212060 629870 212396 629898
rect 221384 629898 221412 632198
rect 232504 632188 232556 632194
rect 232504 632130 232556 632136
rect 231032 632120 231084 632126
rect 231032 632062 231084 632068
rect 231044 629898 231072 632062
rect 221384 629870 221720 629898
rect 231044 629870 231380 629898
rect 209686 620256 209742 620265
rect 209686 620191 209742 620200
rect 205638 619576 205694 619585
rect 205638 619511 205694 619520
rect 205652 611250 205680 619511
rect 209700 611318 209728 620191
rect 232516 615494 232544 632130
rect 232596 632120 232648 632126
rect 232596 632062 232648 632068
rect 231872 615466 232544 615494
rect 209688 611312 209740 611318
rect 231872 611266 231900 615466
rect 209688 611254 209740 611260
rect 205640 611244 205692 611250
rect 205640 611186 205692 611192
rect 231780 611238 231900 611266
rect 231780 610722 231808 611238
rect 231380 610694 231808 610722
rect 211724 610014 212060 610042
rect 221720 610014 222056 610042
rect 211724 608598 211752 610014
rect 211712 608592 211764 608598
rect 211712 608534 211764 608540
rect 222028 608530 222056 610014
rect 232608 608530 232636 632062
rect 232700 611998 232728 632266
rect 233238 619576 233294 619585
rect 233238 619511 233294 619520
rect 232688 611992 232740 611998
rect 232688 611934 232740 611940
rect 233252 611182 233280 619511
rect 233240 611176 233292 611182
rect 233240 611118 233292 611124
rect 204996 608524 205048 608530
rect 204996 608466 205048 608472
rect 222016 608524 222068 608530
rect 222016 608466 222068 608472
rect 232596 608524 232648 608530
rect 232596 608466 232648 608472
rect 222292 604648 222344 604654
rect 222292 604590 222344 604596
rect 222304 602956 222332 604590
rect 232504 604580 232556 604586
rect 232504 604522 232556 604528
rect 212368 602274 212658 602290
rect 210424 602268 210476 602274
rect 210424 602210 210476 602216
rect 212356 602268 212658 602274
rect 212408 602262 212658 602268
rect 231978 602262 232084 602290
rect 212356 602210 212408 602216
rect 205640 601792 205692 601798
rect 205640 601734 205692 601740
rect 204996 599276 205048 599282
rect 204996 599218 205048 599224
rect 205008 580990 205036 599218
rect 205652 592793 205680 601734
rect 209688 601724 209740 601730
rect 209688 601666 209740 601672
rect 209700 593473 209728 601666
rect 209686 593464 209742 593473
rect 209686 593399 209742 593408
rect 205638 592784 205694 592793
rect 205638 592719 205694 592728
rect 204996 580984 205048 580990
rect 204996 580926 205048 580932
rect 210436 580922 210464 602210
rect 212644 580922 212672 583100
rect 210424 580916 210476 580922
rect 210424 580858 210476 580864
rect 212632 580916 212684 580922
rect 212632 580858 212684 580864
rect 222304 580854 222332 583100
rect 231964 580990 231992 583100
rect 232056 580990 232084 602262
rect 231952 580984 232004 580990
rect 231952 580926 232004 580932
rect 232044 580984 232096 580990
rect 232044 580926 232096 580932
rect 232516 580922 232544 604522
rect 233240 601860 233292 601866
rect 233240 601802 233292 601808
rect 233252 592793 233280 601802
rect 233238 592784 233294 592793
rect 233238 592719 233294 592728
rect 232504 580916 232556 580922
rect 232504 580858 232556 580864
rect 222292 580848 222344 580854
rect 222292 580790 222344 580796
rect 212264 578468 212316 578474
rect 212264 578410 212316 578416
rect 232688 578468 232740 578474
rect 232688 578410 232740 578416
rect 204996 578264 205048 578270
rect 204996 578206 205048 578212
rect 205008 554674 205036 578206
rect 212276 575906 212304 578410
rect 221372 578400 221424 578406
rect 221372 578342 221424 578348
rect 212060 575878 212304 575906
rect 221384 575906 221412 578342
rect 232504 578332 232556 578338
rect 232504 578274 232556 578280
rect 231032 578264 231084 578270
rect 231032 578206 231084 578212
rect 231044 575906 231072 578206
rect 221384 575878 221720 575906
rect 231044 575878 231380 575906
rect 209686 566264 209742 566273
rect 209686 566199 209742 566208
rect 205638 565584 205694 565593
rect 205638 565519 205694 565528
rect 205652 557462 205680 565519
rect 209700 557530 209728 566199
rect 232516 557534 232544 578274
rect 232596 578264 232648 578270
rect 232596 578206 232648 578212
rect 209688 557524 209740 557530
rect 209688 557466 209740 557472
rect 231780 557506 232544 557534
rect 205640 557456 205692 557462
rect 205640 557398 205692 557404
rect 231780 556730 231808 557506
rect 231380 556702 231808 556730
rect 211724 556022 212060 556050
rect 221720 556022 222056 556050
rect 211724 554742 211752 556022
rect 211712 554736 211764 554742
rect 211712 554678 211764 554684
rect 222028 554674 222056 556022
rect 232608 554674 232636 578206
rect 232700 558210 232728 578410
rect 233238 565584 233294 565593
rect 233238 565519 233294 565528
rect 232688 558204 232740 558210
rect 232688 558146 232740 558152
rect 233252 557394 233280 565519
rect 233240 557388 233292 557394
rect 233240 557330 233292 557336
rect 204996 554668 205048 554674
rect 204996 554610 205048 554616
rect 222016 554668 222068 554674
rect 222016 554610 222068 554616
rect 232596 554668 232648 554674
rect 232596 554610 232648 554616
rect 222292 550792 222344 550798
rect 222292 550734 222344 550740
rect 222304 548964 222332 550734
rect 232504 550724 232556 550730
rect 232504 550666 232556 550672
rect 212368 548282 212658 548298
rect 210424 548276 210476 548282
rect 210424 548218 210476 548224
rect 212356 548276 212658 548282
rect 212408 548270 212658 548276
rect 231978 548270 232084 548298
rect 212356 548218 212408 548224
rect 204996 547120 205048 547126
rect 204996 547062 205048 547068
rect 205008 527134 205036 547062
rect 209686 539472 209742 539481
rect 209686 539407 209742 539416
rect 205638 538792 205694 538801
rect 205638 538727 205694 538736
rect 205652 529854 205680 538727
rect 209700 529922 209728 539407
rect 209688 529916 209740 529922
rect 209688 529858 209740 529864
rect 205640 529848 205692 529854
rect 205640 529790 205692 529796
rect 204996 527128 205048 527134
rect 204996 527070 205048 527076
rect 210436 527066 210464 548218
rect 212644 527066 212672 529108
rect 210424 527060 210476 527066
rect 210424 527002 210476 527008
rect 212632 527060 212684 527066
rect 212632 527002 212684 527008
rect 222304 526998 222332 529108
rect 231964 527134 231992 529108
rect 232056 527134 232084 548270
rect 231952 527128 232004 527134
rect 231952 527070 232004 527076
rect 232044 527128 232096 527134
rect 232044 527070 232096 527076
rect 232516 527066 232544 550666
rect 233238 538792 233294 538801
rect 233238 538727 233294 538736
rect 233252 529786 233280 538727
rect 233240 529780 233292 529786
rect 233240 529722 233292 529728
rect 232504 527060 232556 527066
rect 232504 527002 232556 527008
rect 222292 526992 222344 526998
rect 222292 526934 222344 526940
rect 212356 523252 212408 523258
rect 212356 523194 212408 523200
rect 232688 523252 232740 523258
rect 232688 523194 232740 523200
rect 204996 523048 205048 523054
rect 204996 522990 205048 522996
rect 205008 500886 205036 522990
rect 212368 521914 212396 523194
rect 221372 523184 221424 523190
rect 221372 523126 221424 523132
rect 212060 521886 212396 521914
rect 221384 521914 221412 523126
rect 232504 523116 232556 523122
rect 232504 523058 232556 523064
rect 231032 523048 231084 523054
rect 231032 522990 231084 522996
rect 231044 521914 231072 522990
rect 221384 521886 221720 521914
rect 231044 521886 231380 521914
rect 205640 520328 205692 520334
rect 205640 520270 205692 520276
rect 209688 520328 209740 520334
rect 209688 520270 209740 520276
rect 205652 511601 205680 520270
rect 209700 512281 209728 520270
rect 209686 512272 209742 512281
rect 209686 512207 209742 512216
rect 205638 511592 205694 511601
rect 205638 511527 205694 511536
rect 232516 509234 232544 523058
rect 232596 523048 232648 523054
rect 232596 522990 232648 522996
rect 231872 509206 232544 509234
rect 231872 502874 231900 509206
rect 231780 502846 231900 502874
rect 231780 502738 231808 502846
rect 231380 502710 231808 502738
rect 211724 502030 212060 502058
rect 221720 502030 222056 502058
rect 211724 500954 211752 502030
rect 211712 500948 211764 500954
rect 211712 500890 211764 500896
rect 222028 500886 222056 502030
rect 232608 500886 232636 522990
rect 232700 504286 232728 523194
rect 233238 511592 233294 511601
rect 233238 511527 233294 511536
rect 232688 504280 232740 504286
rect 232688 504222 232740 504228
rect 233252 503674 233280 511527
rect 233240 503668 233292 503674
rect 233240 503610 233292 503616
rect 204996 500880 205048 500886
rect 204996 500822 205048 500828
rect 222016 500880 222068 500886
rect 222016 500822 222068 500828
rect 232596 500880 232648 500886
rect 232596 500822 232648 500828
rect 222292 497004 222344 497010
rect 222292 496946 222344 496952
rect 222304 494972 222332 496946
rect 232504 496936 232556 496942
rect 232504 496878 232556 496884
rect 212368 494290 212658 494306
rect 210424 494284 210476 494290
rect 210424 494226 210476 494232
rect 212356 494284 212658 494290
rect 212408 494278 212658 494284
rect 231978 494278 232084 494306
rect 212356 494226 212408 494232
rect 204996 492108 205048 492114
rect 204996 492050 205048 492056
rect 205008 473346 205036 492050
rect 209686 485480 209742 485489
rect 209686 485415 209742 485424
rect 205638 484800 205694 484809
rect 205638 484735 205694 484744
rect 205652 475998 205680 484735
rect 209700 476066 209728 485415
rect 209688 476060 209740 476066
rect 209688 476002 209740 476008
rect 205640 475992 205692 475998
rect 205640 475934 205692 475940
rect 204996 473340 205048 473346
rect 204996 473282 205048 473288
rect 210436 473278 210464 494226
rect 212644 473278 212672 475116
rect 210424 473272 210476 473278
rect 210424 473214 210476 473220
rect 212632 473272 212684 473278
rect 212632 473214 212684 473220
rect 222304 473210 222332 475116
rect 231964 473346 231992 475116
rect 232056 473346 232084 494278
rect 231952 473340 232004 473346
rect 231952 473282 232004 473288
rect 232044 473340 232096 473346
rect 232044 473282 232096 473288
rect 232516 473278 232544 496878
rect 233238 484800 233294 484809
rect 233238 484735 233294 484744
rect 233252 475930 233280 484735
rect 233240 475924 233292 475930
rect 233240 475866 233292 475872
rect 232504 473272 232556 473278
rect 232504 473214 232556 473220
rect 222292 473204 222344 473210
rect 222292 473146 222344 473152
rect 212356 469464 212408 469470
rect 212356 469406 212408 469412
rect 232688 469464 232740 469470
rect 232688 469406 232740 469412
rect 204996 469260 205048 469266
rect 204996 469202 205048 469208
rect 205008 445670 205036 469202
rect 212368 467922 212396 469406
rect 221372 469396 221424 469402
rect 221372 469338 221424 469344
rect 212060 467894 212396 467922
rect 221384 467922 221412 469338
rect 232596 469328 232648 469334
rect 232596 469270 232648 469276
rect 231032 469260 231084 469266
rect 231032 469202 231084 469208
rect 232504 469260 232556 469266
rect 232504 469202 232556 469208
rect 231044 467922 231072 469202
rect 221384 467894 221720 467922
rect 231044 467894 231380 467922
rect 205640 466540 205692 466546
rect 205640 466482 205692 466488
rect 205652 457609 205680 466482
rect 209688 466472 209740 466478
rect 209688 466414 209740 466420
rect 209700 458289 209728 466414
rect 209686 458280 209742 458289
rect 209686 458215 209742 458224
rect 205638 457600 205694 457609
rect 205638 457535 205694 457544
rect 231676 448520 231728 448526
rect 231380 448468 231676 448474
rect 231380 448462 231728 448468
rect 231380 448446 231716 448462
rect 211724 448038 212060 448066
rect 221720 448038 222056 448066
rect 211724 445738 211752 448038
rect 222028 445738 222056 448038
rect 232516 445738 232544 469202
rect 232608 448526 232636 469270
rect 232700 449954 232728 469406
rect 233240 466608 233292 466614
rect 233240 466550 233292 466556
rect 233252 457609 233280 466550
rect 233238 457600 233294 457609
rect 233238 457535 233294 457544
rect 232688 449948 232740 449954
rect 232688 449890 232740 449896
rect 232596 448520 232648 448526
rect 232596 448462 232648 448468
rect 211712 445732 211764 445738
rect 211712 445674 211764 445680
rect 222016 445732 222068 445738
rect 222016 445674 222068 445680
rect 232504 445732 232556 445738
rect 232504 445674 232556 445680
rect 204996 445664 205048 445670
rect 204996 445606 205048 445612
rect 222200 443148 222252 443154
rect 222200 443090 222252 443096
rect 210424 441652 210476 441658
rect 210424 441594 210476 441600
rect 212540 441652 212592 441658
rect 222212 441614 222240 443090
rect 232504 443080 232556 443086
rect 232504 443022 232556 443028
rect 212592 441600 212764 441614
rect 212540 441594 212764 441600
rect 205640 440292 205692 440298
rect 205640 440234 205692 440240
rect 209688 440292 209740 440298
rect 209688 440234 209740 440240
rect 204996 436144 205048 436150
rect 204996 436086 205048 436092
rect 205008 419490 205036 436086
rect 205652 431361 205680 440234
rect 209700 431497 209728 440234
rect 209686 431488 209742 431497
rect 209686 431423 209742 431432
rect 205638 431352 205694 431361
rect 205638 431287 205694 431296
rect 204996 419484 205048 419490
rect 204996 419426 205048 419432
rect 210436 419422 210464 441594
rect 212552 441586 212764 441594
rect 222212 441586 222424 441614
rect 212736 440994 212764 441586
rect 212658 440966 212764 440994
rect 222396 440858 222424 441586
rect 222318 440830 222424 440858
rect 231978 440286 232084 440314
rect 212644 419422 212672 421124
rect 210424 419416 210476 419422
rect 210424 419358 210476 419364
rect 212632 419416 212684 419422
rect 212632 419358 212684 419364
rect 222304 419354 222332 421124
rect 231964 419490 231992 421124
rect 232056 419490 232084 440286
rect 231952 419484 232004 419490
rect 231952 419426 232004 419432
rect 232044 419484 232096 419490
rect 232044 419426 232096 419432
rect 232516 419422 232544 443022
rect 233238 430808 233294 430817
rect 233238 430743 233294 430752
rect 233252 422278 233280 430743
rect 233240 422272 233292 422278
rect 233240 422214 233292 422220
rect 232504 419416 232556 419422
rect 232504 419358 232556 419364
rect 222292 419348 222344 419354
rect 222292 419290 222344 419296
rect 212356 415676 212408 415682
rect 212356 415618 212408 415624
rect 232688 415676 232740 415682
rect 232688 415618 232740 415624
rect 204996 415472 205048 415478
rect 204996 415414 205048 415420
rect 205008 391882 205036 415414
rect 212368 413930 212396 415618
rect 221372 415608 221424 415614
rect 221372 415550 221424 415556
rect 212060 413902 212396 413930
rect 221384 413930 221412 415550
rect 232596 415540 232648 415546
rect 232596 415482 232648 415488
rect 231032 415472 231084 415478
rect 231032 415414 231084 415420
rect 232504 415472 232556 415478
rect 232504 415414 232556 415420
rect 231044 413930 231072 415414
rect 221384 413902 221720 413930
rect 231044 413902 231380 413930
rect 209686 404288 209742 404297
rect 209686 404223 209742 404232
rect 205638 403608 205694 403617
rect 205638 403543 205694 403552
rect 205652 394534 205680 403543
rect 209700 394670 209728 404223
rect 209688 394664 209740 394670
rect 209688 394606 209740 394612
rect 205640 394528 205692 394534
rect 205640 394470 205692 394476
rect 211724 394046 212060 394074
rect 221720 394046 221964 394074
rect 231380 394046 231624 394074
rect 211724 391950 211752 394046
rect 221936 391950 221964 394046
rect 231596 393310 231624 394046
rect 231584 393304 231636 393310
rect 231584 393246 231636 393252
rect 232516 391950 232544 415414
rect 232608 393310 232636 415482
rect 232700 395078 232728 415618
rect 233238 403608 233294 403617
rect 233238 403543 233294 403552
rect 232688 395072 232740 395078
rect 232688 395014 232740 395020
rect 233252 394602 233280 403543
rect 233240 394596 233292 394602
rect 233240 394538 233292 394544
rect 232596 393304 232648 393310
rect 232596 393246 232648 393252
rect 211712 391944 211764 391950
rect 211712 391886 211764 391892
rect 221924 391944 221976 391950
rect 221924 391886 221976 391892
rect 232504 391944 232556 391950
rect 232504 391886 232556 391892
rect 204996 391876 205048 391882
rect 204996 391818 205048 391824
rect 222292 389360 222344 389366
rect 222292 389302 222344 389308
rect 222304 386852 222332 389302
rect 232504 389292 232556 389298
rect 232504 389234 232556 389240
rect 205640 386504 205692 386510
rect 205640 386446 205692 386452
rect 204996 385008 205048 385014
rect 204996 384950 205048 384956
rect 205008 365702 205036 384950
rect 205652 377369 205680 386446
rect 209688 386436 209740 386442
rect 209688 386378 209740 386384
rect 209700 377505 209728 386378
rect 212460 386294 212658 386322
rect 231978 386294 232084 386322
rect 212460 385082 212488 386294
rect 212448 385076 212500 385082
rect 212448 385018 212500 385024
rect 209686 377496 209742 377505
rect 209686 377431 209742 377440
rect 205638 377360 205694 377369
rect 205638 377295 205694 377304
rect 204996 365696 205048 365702
rect 204996 365638 205048 365644
rect 212644 365634 212672 367132
rect 212632 365628 212684 365634
rect 212632 365570 212684 365576
rect 222304 365566 222332 367132
rect 231964 365702 231992 367132
rect 232056 365702 232084 386294
rect 231952 365696 232004 365702
rect 231952 365638 232004 365644
rect 232044 365696 232096 365702
rect 232044 365638 232096 365644
rect 232516 365634 232544 389234
rect 233240 386572 233292 386578
rect 233240 386514 233292 386520
rect 233252 376825 233280 386514
rect 233238 376816 233294 376825
rect 233238 376751 233294 376760
rect 232504 365628 232556 365634
rect 232504 365570 232556 365576
rect 222292 365560 222344 365566
rect 222292 365502 222344 365508
rect 221372 361752 221424 361758
rect 221372 361694 221424 361700
rect 232596 361752 232648 361758
rect 232596 361694 232648 361700
rect 212356 361684 212408 361690
rect 212356 361626 212408 361632
rect 204996 361616 205048 361622
rect 204996 361558 205048 361564
rect 205008 338026 205036 361558
rect 212368 359938 212396 361626
rect 212060 359910 212396 359938
rect 221384 359938 221412 361694
rect 231032 361616 231084 361622
rect 231032 361558 231084 361564
rect 232504 361616 232556 361622
rect 232504 361558 232556 361564
rect 231044 359938 231072 361558
rect 221384 359910 221720 359938
rect 231044 359910 231380 359938
rect 209686 350296 209742 350305
rect 209686 350231 209742 350240
rect 205638 349616 205694 349625
rect 205638 349551 205694 349560
rect 205652 340814 205680 349551
rect 209700 340882 209728 350231
rect 209688 340876 209740 340882
rect 209688 340818 209740 340824
rect 205640 340808 205692 340814
rect 231676 340808 231728 340814
rect 205640 340750 205692 340756
rect 231380 340756 231676 340762
rect 231380 340750 231728 340756
rect 231380 340734 231716 340750
rect 211724 340054 212060 340082
rect 221720 340054 222056 340082
rect 211724 338094 211752 340054
rect 211712 338088 211764 338094
rect 211712 338030 211764 338036
rect 222028 338026 222056 340054
rect 232516 338026 232544 361558
rect 232608 340814 232636 361694
rect 232688 361684 232740 361690
rect 232688 361626 232740 361632
rect 232700 341426 232728 361626
rect 233238 349616 233294 349625
rect 233238 349551 233294 349560
rect 232688 341420 232740 341426
rect 232688 341362 232740 341368
rect 232596 340808 232648 340814
rect 232596 340750 232648 340756
rect 233252 340746 233280 349551
rect 233240 340740 233292 340746
rect 233240 340682 233292 340688
rect 204996 338020 205048 338026
rect 204996 337962 205048 337968
rect 222016 338020 222068 338026
rect 222016 337962 222068 337968
rect 232504 338020 232556 338026
rect 232504 337962 232556 337968
rect 222292 335504 222344 335510
rect 222292 335446 222344 335452
rect 222304 332860 222332 335446
rect 232504 335436 232556 335442
rect 232504 335378 232556 335384
rect 212460 332302 212658 332330
rect 231978 332302 232084 332330
rect 209688 331356 209740 331362
rect 209688 331298 209740 331304
rect 204996 329044 205048 329050
rect 204996 328986 205048 328992
rect 205008 311846 205036 328986
rect 209700 324057 209728 331298
rect 212460 331294 212488 332302
rect 212448 331288 212500 331294
rect 212448 331230 212500 331236
rect 209686 324048 209742 324057
rect 209686 323983 209742 323992
rect 205638 322144 205694 322153
rect 205638 322079 205694 322088
rect 205652 314566 205680 322079
rect 205640 314560 205692 314566
rect 205640 314502 205692 314508
rect 204996 311840 205048 311846
rect 204996 311782 205048 311788
rect 212644 311778 212672 313140
rect 212632 311772 212684 311778
rect 212632 311714 212684 311720
rect 222304 311710 222332 313140
rect 231964 311846 231992 313140
rect 232056 311846 232084 332302
rect 231952 311840 232004 311846
rect 231952 311782 232004 311788
rect 232044 311840 232096 311846
rect 232044 311782 232096 311788
rect 232516 311778 232544 335378
rect 233238 322144 233294 322153
rect 233238 322079 233294 322088
rect 233252 314634 233280 322079
rect 233240 314628 233292 314634
rect 233240 314570 233292 314576
rect 232504 311772 232556 311778
rect 232504 311714 232556 311720
rect 222292 311704 222344 311710
rect 222292 311646 222344 311652
rect 212264 308032 212316 308038
rect 212264 307974 212316 307980
rect 232688 308032 232740 308038
rect 232688 307974 232740 307980
rect 204996 307828 205048 307834
rect 204996 307770 205048 307776
rect 205008 284238 205036 307770
rect 212276 305946 212304 307974
rect 221372 307964 221424 307970
rect 221372 307906 221424 307912
rect 212060 305918 212304 305946
rect 221384 305946 221412 307906
rect 232504 307896 232556 307902
rect 232504 307838 232556 307844
rect 231032 307828 231084 307834
rect 231032 307770 231084 307776
rect 231044 305946 231072 307770
rect 221384 305918 221720 305946
rect 231044 305918 231380 305946
rect 209686 296304 209742 296313
rect 209686 296239 209742 296248
rect 205638 295624 205694 295633
rect 205638 295559 205694 295568
rect 205652 287026 205680 295559
rect 209700 287026 209728 296239
rect 232516 287054 232544 307838
rect 232596 307828 232648 307834
rect 232596 307770 232648 307776
rect 231780 287026 232544 287054
rect 205640 287020 205692 287026
rect 205640 286962 205692 286968
rect 209688 287020 209740 287026
rect 209688 286962 209740 286968
rect 231780 286770 231808 287026
rect 231380 286742 231808 286770
rect 211724 286062 212060 286090
rect 221720 286062 222056 286090
rect 211724 284306 211752 286062
rect 211712 284300 211764 284306
rect 211712 284242 211764 284248
rect 222028 284238 222056 286062
rect 232608 284238 232636 307770
rect 232700 287978 232728 307974
rect 233238 295624 233294 295633
rect 233238 295559 233294 295568
rect 232688 287972 232740 287978
rect 232688 287914 232740 287920
rect 233252 286958 233280 295559
rect 233240 286952 233292 286958
rect 233240 286894 233292 286900
rect 204996 284232 205048 284238
rect 204996 284174 205048 284180
rect 222016 284232 222068 284238
rect 222016 284174 222068 284180
rect 232596 284232 232648 284238
rect 232596 284174 232648 284180
rect 222292 280356 222344 280362
rect 222292 280298 222344 280304
rect 222304 278868 222332 280298
rect 232504 280288 232556 280294
rect 232504 280230 232556 280236
rect 212460 278310 212658 278338
rect 231978 278310 232084 278338
rect 205640 277500 205692 277506
rect 205640 277442 205692 277448
rect 209688 277500 209740 277506
rect 209688 277442 209740 277448
rect 204996 272604 205048 272610
rect 204996 272546 205048 272552
rect 205008 256698 205036 272546
rect 205652 269113 205680 277442
rect 209700 269929 209728 277442
rect 212460 277438 212488 278310
rect 212448 277432 212500 277438
rect 212448 277374 212500 277380
rect 209686 269920 209742 269929
rect 209686 269855 209742 269864
rect 205638 269104 205694 269113
rect 205638 269039 205694 269048
rect 204996 256692 205048 256698
rect 204996 256634 205048 256640
rect 212644 256630 212672 259148
rect 212632 256624 212684 256630
rect 212632 256566 212684 256572
rect 222304 256562 222332 259148
rect 231964 256698 231992 259148
rect 232056 256698 232084 278310
rect 231952 256692 232004 256698
rect 231952 256634 232004 256640
rect 232044 256692 232096 256698
rect 232044 256634 232096 256640
rect 232516 256630 232544 280230
rect 233240 277568 233292 277574
rect 233240 277510 233292 277516
rect 233252 269113 233280 277510
rect 233238 269104 233294 269113
rect 233238 269039 233294 269048
rect 232504 256624 232556 256630
rect 232504 256566 232556 256572
rect 222292 256556 222344 256562
rect 222292 256498 222344 256504
rect 212356 254176 212408 254182
rect 212356 254118 212408 254124
rect 232688 254176 232740 254182
rect 232688 254118 232740 254124
rect 204996 253972 205048 253978
rect 204996 253914 205048 253920
rect 205008 230382 205036 253914
rect 212368 251954 212396 254118
rect 221372 254108 221424 254114
rect 221372 254050 221424 254056
rect 212060 251926 212396 251954
rect 221384 251954 221412 254050
rect 232504 254040 232556 254046
rect 232504 253982 232556 253988
rect 231032 253972 231084 253978
rect 231032 253914 231084 253920
rect 231044 251954 231072 253914
rect 221384 251926 221720 251954
rect 231044 251926 231380 251954
rect 205640 251252 205692 251258
rect 205640 251194 205692 251200
rect 209688 251252 209740 251258
rect 209688 251194 209740 251200
rect 205652 241641 205680 251194
rect 209700 242321 209728 251194
rect 209686 242312 209742 242321
rect 209686 242247 209742 242256
rect 205638 241632 205694 241641
rect 205638 241567 205694 241576
rect 232516 238754 232544 253982
rect 232596 253972 232648 253978
rect 232596 253914 232648 253920
rect 231872 238726 232544 238754
rect 231872 232914 231900 238726
rect 231780 232886 231900 232914
rect 231780 232778 231808 232886
rect 231380 232750 231808 232778
rect 211724 232070 212060 232098
rect 221720 232070 222056 232098
rect 211724 230450 211752 232070
rect 211712 230444 211764 230450
rect 211712 230386 211764 230392
rect 222028 230382 222056 232070
rect 232608 230382 232636 253914
rect 232700 233578 232728 254118
rect 233240 251320 233292 251326
rect 233240 251262 233292 251268
rect 233252 241641 233280 251262
rect 233238 241632 233294 241641
rect 233238 241567 233294 241576
rect 232688 233572 232740 233578
rect 232688 233514 232740 233520
rect 204996 230376 205048 230382
rect 204996 230318 205048 230324
rect 222016 230376 222068 230382
rect 222016 230318 222068 230324
rect 232596 230376 232648 230382
rect 232596 230318 232648 230324
rect 222292 226500 222344 226506
rect 222292 226442 222344 226448
rect 222304 224876 222332 226442
rect 232504 226432 232556 226438
rect 232504 226374 232556 226380
rect 212460 224330 212658 224346
rect 210424 224324 210476 224330
rect 210424 224266 210476 224272
rect 212448 224324 212658 224330
rect 212500 224318 212658 224324
rect 231978 224318 232084 224346
rect 212448 224266 212500 224272
rect 205640 223712 205692 223718
rect 205640 223654 205692 223660
rect 204996 221876 205048 221882
rect 204996 221818 205048 221824
rect 205008 202842 205036 221818
rect 205652 215257 205680 223654
rect 209688 223644 209740 223650
rect 209688 223586 209740 223592
rect 209700 215393 209728 223586
rect 209686 215384 209742 215393
rect 209686 215319 209742 215328
rect 205638 215248 205694 215257
rect 205638 215183 205694 215192
rect 204996 202836 205048 202842
rect 204996 202778 205048 202784
rect 210436 202774 210464 224266
rect 232056 212534 232084 224318
rect 232056 212506 232268 212534
rect 212658 205006 213040 205034
rect 222318 205006 222608 205034
rect 231978 205006 232176 205034
rect 213012 202774 213040 205006
rect 210424 202768 210476 202774
rect 210424 202710 210476 202716
rect 213000 202768 213052 202774
rect 213000 202710 213052 202716
rect 222580 202706 222608 205006
rect 232148 203998 232176 205006
rect 231860 203992 231912 203998
rect 231860 203934 231912 203940
rect 232136 203992 232188 203998
rect 232136 203934 232188 203940
rect 231872 202842 231900 203934
rect 232240 203810 232268 212506
rect 232056 203782 232268 203810
rect 232056 202842 232084 203782
rect 231860 202836 231912 202842
rect 231860 202778 231912 202784
rect 232044 202836 232096 202842
rect 232044 202778 232096 202784
rect 232516 202774 232544 226374
rect 233240 223780 233292 223786
rect 233240 223722 233292 223728
rect 233252 214713 233280 223722
rect 233238 214704 233294 214713
rect 233238 214639 233294 214648
rect 232504 202768 232556 202774
rect 232504 202710 232556 202716
rect 222568 202700 222620 202706
rect 222568 202642 222620 202648
rect 221372 200320 221424 200326
rect 221372 200262 221424 200268
rect 232504 200320 232556 200326
rect 232504 200262 232556 200268
rect 212264 200252 212316 200258
rect 212264 200194 212316 200200
rect 204996 200184 205048 200190
rect 204996 200126 205048 200132
rect 205008 176594 205036 200126
rect 212276 197962 212304 200194
rect 212060 197934 212304 197962
rect 221384 197962 221412 200262
rect 231032 200184 231084 200190
rect 231032 200126 231084 200132
rect 231044 197962 231072 200126
rect 221384 197934 221720 197962
rect 231044 197934 231380 197962
rect 209686 188320 209742 188329
rect 209686 188255 209742 188264
rect 205638 187640 205694 187649
rect 205638 187575 205694 187584
rect 205652 179314 205680 187575
rect 209700 179382 209728 188255
rect 232516 180794 232544 200262
rect 232688 200252 232740 200258
rect 232688 200194 232740 200200
rect 232596 200184 232648 200190
rect 232596 200126 232648 200132
rect 231872 180766 232544 180794
rect 209688 179376 209740 179382
rect 209688 179318 209740 179324
rect 205640 179308 205692 179314
rect 205640 179250 205692 179256
rect 231872 178922 231900 180766
rect 231780 178894 231900 178922
rect 231780 178786 231808 178894
rect 231380 178758 231808 178786
rect 211724 178078 212060 178106
rect 221720 178078 222056 178106
rect 211724 176662 211752 178078
rect 211712 176656 211764 176662
rect 211712 176598 211764 176604
rect 222028 176594 222056 178078
rect 232608 176594 232636 200126
rect 232700 179926 232728 200194
rect 233238 187640 233294 187649
rect 233238 187575 233294 187584
rect 232688 179920 232740 179926
rect 232688 179862 232740 179868
rect 233252 179246 233280 187575
rect 233240 179240 233292 179246
rect 233240 179182 233292 179188
rect 204996 176588 205048 176594
rect 204996 176530 205048 176536
rect 222016 176588 222068 176594
rect 222016 176530 222068 176536
rect 232596 176588 232648 176594
rect 232596 176530 232648 176536
rect 222292 172712 222344 172718
rect 222292 172654 222344 172660
rect 210424 171148 210476 171154
rect 210424 171090 210476 171096
rect 212632 171148 212684 171154
rect 212684 171106 212764 171134
rect 212632 171090 212684 171096
rect 204996 165912 205048 165918
rect 204996 165854 205048 165860
rect 205008 149054 205036 165854
rect 209686 161392 209742 161401
rect 209686 161327 209742 161336
rect 205638 160168 205694 160177
rect 205638 160103 205694 160112
rect 205652 151706 205680 160103
rect 209700 151774 209728 161327
rect 209688 151768 209740 151774
rect 209688 151710 209740 151716
rect 205640 151700 205692 151706
rect 205640 151642 205692 151648
rect 204996 149048 205048 149054
rect 204996 148990 205048 148996
rect 210436 148986 210464 171090
rect 212736 170898 212764 171106
rect 212658 170870 212764 170898
rect 222304 170884 222332 172654
rect 232504 172644 232556 172650
rect 232504 172586 232556 172592
rect 231978 170326 232084 170354
rect 212644 148986 212672 151028
rect 210424 148980 210476 148986
rect 210424 148922 210476 148928
rect 212632 148980 212684 148986
rect 212632 148922 212684 148928
rect 222304 148918 222332 151028
rect 231964 149054 231992 151028
rect 232056 149054 232084 170326
rect 231952 149048 232004 149054
rect 231952 148990 232004 148996
rect 232044 149048 232096 149054
rect 232044 148990 232096 148996
rect 232516 148986 232544 172586
rect 233238 160712 233294 160721
rect 233238 160647 233294 160656
rect 233252 151638 233280 160647
rect 233240 151632 233292 151638
rect 233240 151574 233292 151580
rect 232504 148980 232556 148986
rect 232504 148922 232556 148928
rect 222292 148912 222344 148918
rect 222292 148854 222344 148860
rect 212356 146532 212408 146538
rect 212356 146474 212408 146480
rect 232688 146532 232740 146538
rect 232688 146474 232740 146480
rect 204996 146328 205048 146334
rect 204996 146270 205048 146276
rect 205008 122738 205036 146270
rect 212368 143970 212396 146474
rect 221372 146464 221424 146470
rect 221372 146406 221424 146412
rect 212060 143942 212396 143970
rect 221384 143970 221412 146406
rect 232504 146396 232556 146402
rect 232504 146338 232556 146344
rect 231032 146328 231084 146334
rect 231032 146270 231084 146276
rect 231044 143970 231072 146270
rect 221384 143942 221720 143970
rect 231044 143942 231380 143970
rect 209686 134328 209742 134337
rect 209686 134263 209742 134272
rect 205638 133648 205694 133657
rect 205638 133583 205694 133592
rect 205652 125526 205680 133583
rect 209700 125594 209728 134263
rect 209688 125588 209740 125594
rect 209688 125530 209740 125536
rect 205640 125520 205692 125526
rect 205640 125462 205692 125468
rect 211724 124086 212060 124114
rect 221720 124086 221964 124114
rect 231380 124086 231624 124114
rect 211724 122806 211752 124086
rect 211712 122800 211764 122806
rect 211712 122742 211764 122748
rect 221936 122738 221964 124086
rect 231596 122806 231624 124086
rect 232516 122806 232544 146338
rect 232596 146328 232648 146334
rect 232596 146270 232648 146276
rect 231584 122800 231636 122806
rect 231584 122742 231636 122748
rect 232504 122800 232556 122806
rect 232504 122742 232556 122748
rect 232608 122738 232636 146270
rect 232700 126954 232728 146474
rect 233238 133648 233294 133657
rect 233238 133583 233294 133592
rect 232688 126948 232740 126954
rect 232688 126890 232740 126896
rect 233252 125458 233280 133583
rect 233240 125452 233292 125458
rect 233240 125394 233292 125400
rect 204996 122732 205048 122738
rect 204996 122674 205048 122680
rect 221924 122732 221976 122738
rect 221924 122674 221976 122680
rect 232596 122732 232648 122738
rect 232596 122674 232648 122680
rect 222292 118856 222344 118862
rect 222292 118798 222344 118804
rect 222304 116892 222332 118798
rect 232504 118788 232556 118794
rect 232504 118730 232556 118736
rect 212368 116346 212658 116362
rect 210424 116340 210476 116346
rect 210424 116282 210476 116288
rect 212356 116340 212658 116346
rect 212408 116334 212658 116340
rect 231978 116334 232084 116362
rect 212356 116282 212408 116288
rect 204996 114776 205048 114782
rect 204996 114718 205048 114724
rect 205008 95198 205036 114718
rect 209686 107400 209742 107409
rect 209686 107335 209742 107344
rect 205638 106720 205694 106729
rect 205638 106655 205694 106664
rect 205652 97986 205680 106655
rect 209700 97986 209728 107335
rect 205640 97980 205692 97986
rect 205640 97922 205692 97928
rect 209688 97980 209740 97986
rect 209688 97922 209740 97928
rect 204996 95192 205048 95198
rect 204996 95134 205048 95140
rect 210436 95130 210464 116282
rect 212644 95130 212672 97036
rect 210424 95124 210476 95130
rect 210424 95066 210476 95072
rect 212632 95124 212684 95130
rect 212632 95066 212684 95072
rect 222304 95062 222332 97036
rect 231964 95198 231992 97036
rect 232056 95198 232084 116334
rect 231952 95192 232004 95198
rect 231952 95134 232004 95140
rect 232044 95192 232096 95198
rect 232044 95134 232096 95140
rect 232516 95130 232544 118730
rect 233238 106720 233294 106729
rect 233238 106655 233294 106664
rect 233252 97918 233280 106655
rect 233240 97912 233292 97918
rect 233240 97854 233292 97860
rect 232504 95124 232556 95130
rect 232504 95066 232556 95072
rect 222292 95056 222344 95062
rect 222292 94998 222344 95004
rect 221372 91248 221424 91254
rect 221372 91190 221424 91196
rect 232596 91248 232648 91254
rect 232596 91190 232648 91196
rect 212356 91180 212408 91186
rect 212356 91122 212408 91128
rect 204996 91112 205048 91118
rect 204996 91054 205048 91060
rect 205008 68950 205036 91054
rect 212368 89978 212396 91122
rect 212060 89950 212396 89978
rect 221384 89978 221412 91190
rect 231032 91112 231084 91118
rect 231032 91054 231084 91060
rect 232504 91112 232556 91118
rect 232504 91054 232556 91060
rect 231044 89978 231072 91054
rect 221384 89950 221720 89978
rect 231044 89950 231380 89978
rect 205640 88392 205692 88398
rect 205640 88334 205692 88340
rect 209688 88392 209740 88398
rect 209688 88334 209740 88340
rect 205652 79665 205680 88334
rect 209700 80345 209728 88334
rect 209686 80336 209742 80345
rect 209686 80271 209742 80280
rect 205638 79656 205694 79665
rect 205638 79591 205694 79600
rect 231676 71664 231728 71670
rect 231676 71606 231728 71612
rect 231688 70666 231716 71606
rect 231380 70638 231716 70666
rect 211724 70094 212060 70122
rect 221720 70094 222056 70122
rect 211724 69018 211752 70094
rect 222028 69018 222056 70094
rect 232516 69018 232544 91054
rect 232608 71670 232636 91190
rect 232688 91180 232740 91186
rect 232688 91122 232740 91128
rect 232700 72350 232728 91122
rect 233238 79656 233294 79665
rect 233238 79591 233294 79600
rect 232688 72344 232740 72350
rect 232688 72286 232740 72292
rect 233252 71738 233280 79591
rect 233240 71732 233292 71738
rect 233240 71674 233292 71680
rect 232596 71664 232648 71670
rect 232596 71606 232648 71612
rect 211712 69012 211764 69018
rect 211712 68954 211764 68960
rect 222016 69012 222068 69018
rect 222016 68954 222068 68960
rect 232504 69012 232556 69018
rect 232504 68954 232556 68960
rect 204996 68944 205048 68950
rect 204996 68886 205048 68892
rect 222292 65068 222344 65074
rect 222292 65010 222344 65016
rect 210424 64932 210476 64938
rect 210424 64874 210476 64880
rect 212632 64932 212684 64938
rect 212632 64874 212684 64880
rect 205640 62144 205692 62150
rect 205640 62086 205692 62092
rect 209688 62144 209740 62150
rect 209688 62086 209740 62092
rect 204996 57928 205048 57934
rect 204996 57870 205048 57876
rect 205008 41410 205036 57870
rect 205652 52737 205680 62086
rect 209700 53417 209728 62086
rect 209686 53408 209742 53417
rect 209686 53343 209742 53352
rect 205638 52728 205694 52737
rect 205638 52663 205694 52672
rect 204996 41404 205048 41410
rect 204996 41346 205048 41352
rect 210436 41342 210464 64874
rect 212644 62900 212672 64874
rect 222304 62900 222332 65010
rect 232504 65000 232556 65006
rect 232504 64942 232556 64948
rect 231978 62206 232084 62234
rect 212644 41342 212672 43044
rect 210424 41336 210476 41342
rect 210424 41278 210476 41284
rect 212632 41336 212684 41342
rect 212632 41278 212684 41284
rect 222304 41274 222332 43044
rect 231964 41410 231992 43044
rect 232056 41410 232084 62206
rect 231952 41404 232004 41410
rect 231952 41346 232004 41352
rect 232044 41404 232096 41410
rect 232044 41346 232096 41352
rect 232516 41342 232544 64942
rect 233238 52728 233294 52737
rect 233238 52663 233294 52672
rect 233252 44130 233280 52663
rect 233240 44124 233292 44130
rect 233240 44066 233292 44072
rect 232504 41336 232556 41342
rect 232504 41278 232556 41284
rect 222292 41268 222344 41274
rect 222292 41210 222344 41216
rect 204904 39432 204956 39438
rect 204904 39374 204956 39380
rect 149704 38412 149756 38418
rect 149704 38354 149756 38360
rect 149796 37460 149848 37466
rect 149796 37402 149848 37408
rect 165712 37460 165764 37466
rect 165712 37402 165764 37408
rect 175464 37460 175516 37466
rect 175464 37402 175516 37408
rect 193680 37460 193732 37466
rect 193680 37402 193732 37408
rect 203524 37460 203576 37466
rect 203524 37402 203576 37408
rect 221372 37460 221424 37466
rect 221372 37402 221424 37408
rect 232504 37460 232556 37466
rect 232504 37402 232556 37408
rect 91100 37392 91152 37398
rect 91100 37334 91152 37340
rect 91468 37392 91520 37398
rect 91468 37334 91520 37340
rect 109684 37392 109736 37398
rect 109684 37334 109736 37340
rect 122104 37392 122156 37398
rect 122104 37334 122156 37340
rect 137652 37392 137704 37398
rect 137652 37334 137704 37340
rect 81440 37324 81492 37330
rect 81440 37266 81492 37272
rect 81452 35986 81480 37266
rect 91112 35986 91140 37334
rect 81452 35958 81696 35986
rect 91112 35958 91356 35986
rect 71884 35278 72036 35306
rect 71044 27600 71096 27606
rect 71044 27542 71096 27548
rect 70306 26888 70362 26897
rect 70306 26823 70362 26832
rect 65616 13796 65668 13802
rect 65616 13738 65668 13744
rect 71884 13394 71912 35278
rect 91480 16674 91508 37334
rect 93124 37324 93176 37330
rect 93124 37266 93176 37272
rect 91356 16646 91508 16674
rect 72036 16102 72096 16130
rect 81696 16102 82032 16130
rect 71872 13388 71924 13394
rect 71872 13330 71924 13336
rect 65524 13184 65576 13190
rect 65524 13126 65576 13132
rect 72068 13122 72096 16102
rect 82004 13802 82032 16102
rect 93136 13802 93164 37266
rect 93860 36032 93912 36038
rect 93860 35974 93912 35980
rect 93872 25673 93900 35974
rect 109696 35972 109724 37334
rect 119344 37324 119396 37330
rect 119344 37266 119396 37272
rect 120724 37324 120776 37330
rect 120724 37266 120776 37272
rect 119356 35972 119384 37266
rect 99484 35278 100050 35306
rect 97908 34536 97960 34542
rect 97908 34478 97960 34484
rect 97920 26353 97948 34478
rect 97906 26344 97962 26353
rect 97906 26279 97962 26288
rect 93858 25664 93914 25673
rect 93858 25599 93914 25608
rect 81992 13796 82044 13802
rect 81992 13738 82044 13744
rect 93124 13796 93176 13802
rect 93124 13738 93176 13744
rect 99484 13326 99512 35278
rect 119712 16584 119764 16590
rect 119370 16532 119712 16538
rect 119370 16526 119764 16532
rect 119370 16510 119752 16526
rect 100036 13394 100064 16116
rect 100024 13388 100076 13394
rect 100024 13330 100076 13336
rect 109696 13326 109724 16116
rect 120736 13326 120764 37266
rect 121460 34604 121512 34610
rect 121460 34546 121512 34552
rect 121472 25673 121500 34546
rect 121458 25664 121514 25673
rect 121458 25599 121514 25608
rect 122116 16590 122144 37334
rect 137664 35972 137692 37334
rect 147312 37324 147364 37330
rect 147312 37266 147364 37272
rect 148324 37324 148376 37330
rect 148324 37266 148376 37272
rect 147324 35972 147352 37266
rect 127084 35278 128018 35306
rect 126888 34604 126940 34610
rect 126888 34546 126940 34552
rect 126900 26353 126928 34546
rect 126886 26344 126942 26353
rect 126886 26279 126942 26288
rect 122104 16584 122156 16590
rect 122104 16526 122156 16532
rect 127084 13326 127112 35278
rect 147588 16584 147640 16590
rect 147338 16532 147588 16538
rect 147338 16526 147640 16532
rect 147338 16510 147628 16526
rect 128004 13394 128032 16116
rect 127992 13388 128044 13394
rect 127992 13330 128044 13336
rect 137664 13326 137692 16116
rect 148336 13326 148364 37266
rect 149060 34536 149112 34542
rect 149060 34478 149112 34484
rect 149072 25673 149100 34478
rect 149058 25664 149114 25673
rect 149058 25599 149114 25608
rect 149808 16590 149836 37402
rect 156328 37392 156380 37398
rect 156328 37334 156380 37340
rect 156340 35986 156368 37334
rect 165724 35986 165752 37402
rect 175372 37324 175424 37330
rect 175372 37266 175424 37272
rect 175384 35986 175412 37266
rect 156032 35958 156368 35986
rect 165692 35958 165752 35986
rect 175352 35958 175412 35986
rect 154488 34536 154540 34542
rect 154488 34478 154540 34484
rect 154500 26353 154528 34478
rect 154486 26344 154542 26353
rect 154486 26279 154542 26288
rect 175476 16674 175504 37402
rect 178684 37392 178736 37398
rect 178684 37334 178736 37340
rect 177304 37324 177356 37330
rect 177304 37266 177356 37272
rect 175352 16646 175504 16674
rect 149796 16584 149848 16590
rect 149796 16526 149848 16532
rect 156032 16102 156092 16130
rect 165692 16102 166028 16130
rect 156064 13394 156092 16102
rect 166000 13802 166028 16102
rect 177316 13802 177344 37266
rect 178040 34604 178092 34610
rect 178040 34546 178092 34552
rect 178052 25673 178080 34546
rect 178038 25664 178094 25673
rect 178038 25599 178094 25608
rect 178696 13802 178724 37334
rect 193692 35972 193720 37402
rect 203340 37324 203392 37330
rect 203340 37266 203392 37272
rect 203352 35972 203380 37266
rect 183664 35278 184046 35306
rect 182088 34604 182140 34610
rect 182088 34546 182140 34552
rect 182100 26353 182128 34546
rect 182086 26344 182142 26353
rect 182086 26279 182142 26288
rect 165988 13796 166040 13802
rect 165988 13738 166040 13744
rect 177304 13796 177356 13802
rect 177304 13738 177356 13744
rect 178684 13796 178736 13802
rect 178684 13738 178736 13744
rect 183664 13394 183692 35278
rect 203536 16674 203564 37402
rect 212356 37392 212408 37398
rect 212356 37334 212408 37340
rect 204904 37324 204956 37330
rect 204904 37266 204956 37272
rect 203366 16646 203564 16674
rect 184032 13802 184060 16116
rect 193692 13802 193720 16116
rect 204916 13802 204944 37266
rect 212368 35986 212396 37334
rect 212060 35958 212396 35986
rect 221384 35986 221412 37402
rect 231032 37324 231084 37330
rect 231032 37266 231084 37272
rect 231044 35986 231072 37266
rect 221384 35958 221720 35986
rect 231044 35958 231380 35986
rect 205640 34536 205692 34542
rect 205640 34478 205692 34484
rect 209688 34536 209740 34542
rect 209688 34478 209740 34484
rect 205652 25945 205680 34478
rect 209700 26353 209728 34478
rect 209686 26344 209742 26353
rect 209686 26279 209742 26288
rect 205638 25936 205694 25945
rect 205638 25871 205694 25880
rect 232516 16574 232544 37402
rect 232596 37392 232648 37398
rect 232596 37334 232648 37340
rect 232608 18018 232636 37334
rect 233240 34604 233292 34610
rect 233240 34546 233292 34552
rect 233252 25673 233280 34546
rect 233238 25664 233294 25673
rect 233238 25599 233294 25608
rect 232596 18012 232648 18018
rect 232596 17954 232648 17960
rect 231780 16546 232544 16574
rect 231780 16538 231808 16546
rect 231380 16510 231808 16538
rect 211724 16102 212060 16130
rect 221720 16102 222056 16130
rect 184020 13796 184072 13802
rect 184020 13738 184072 13744
rect 193680 13796 193732 13802
rect 193680 13738 193732 13744
rect 204904 13796 204956 13802
rect 204904 13738 204956 13744
rect 211724 13394 211752 16102
rect 222028 13394 222056 16102
rect 233896 15094 233924 700266
rect 233976 658300 234028 658306
rect 233976 658242 234028 658248
rect 233988 634642 234016 658242
rect 233976 634636 234028 634642
rect 233976 634578 234028 634584
rect 233976 604512 234028 604518
rect 233976 604454 234028 604460
rect 233988 580854 234016 604454
rect 233976 580848 234028 580854
rect 233976 580790 234028 580796
rect 233976 550656 234028 550662
rect 233976 550598 234028 550604
rect 233988 526998 234016 550598
rect 233976 526992 234028 526998
rect 233976 526934 234028 526940
rect 233976 496868 234028 496874
rect 233976 496810 234028 496816
rect 233988 473210 234016 496810
rect 233976 473204 234028 473210
rect 233976 473146 234028 473152
rect 233976 443012 234028 443018
rect 233976 442954 234028 442960
rect 233988 419354 234016 442954
rect 233976 419348 234028 419354
rect 233976 419290 234028 419296
rect 233976 389224 234028 389230
rect 233976 389166 234028 389172
rect 233988 365566 234016 389166
rect 233976 365560 234028 365566
rect 233976 365502 234028 365508
rect 233976 335368 234028 335374
rect 233976 335310 234028 335316
rect 233988 311710 234016 335310
rect 233976 311704 234028 311710
rect 233976 311646 234028 311652
rect 233976 280220 234028 280226
rect 233976 280162 234028 280168
rect 233988 256562 234016 280162
rect 233976 256556 234028 256562
rect 233976 256498 234028 256504
rect 233976 226364 234028 226370
rect 233976 226306 234028 226312
rect 233988 202706 234016 226306
rect 233976 202700 234028 202706
rect 233976 202642 234028 202648
rect 233976 172576 234028 172582
rect 233976 172518 234028 172524
rect 233988 148918 234016 172518
rect 233976 148912 234028 148918
rect 233976 148854 234028 148860
rect 233976 118720 234028 118726
rect 233976 118662 234028 118668
rect 233988 95062 234016 118662
rect 233976 95056 234028 95062
rect 233976 94998 234028 95004
rect 233976 64932 234028 64938
rect 233976 64874 234028 64880
rect 233988 41274 234016 64874
rect 233976 41268 234028 41274
rect 233976 41210 234028 41216
rect 234632 39370 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700602 267688 703520
rect 267648 700596 267700 700602
rect 267648 700538 267700 700544
rect 300136 700534 300164 703520
rect 332520 700534 332548 703520
rect 300124 700528 300176 700534
rect 300124 700470 300176 700476
rect 322204 700528 322256 700534
rect 322204 700470 322256 700476
rect 332508 700528 332560 700534
rect 332508 700470 332560 700476
rect 296352 686112 296404 686118
rect 296352 686054 296404 686060
rect 316776 686112 316828 686118
rect 316776 686054 316828 686060
rect 260104 686044 260156 686050
rect 260104 685986 260156 685992
rect 277676 686044 277728 686050
rect 277676 685986 277728 685992
rect 287520 686044 287572 686050
rect 287520 685986 287572 685992
rect 249708 685976 249760 685982
rect 249708 685918 249760 685924
rect 249720 683876 249748 685918
rect 259368 685908 259420 685914
rect 259368 685850 259420 685856
rect 259380 683876 259408 685850
rect 238864 683318 240074 683346
rect 238668 683188 238720 683194
rect 238668 683130 238720 683136
rect 238680 674257 238708 683130
rect 238666 674248 238722 674257
rect 238666 674183 238722 674192
rect 238864 662250 238892 683318
rect 260116 673454 260144 685986
rect 268016 685976 268068 685982
rect 268016 685918 268068 685924
rect 260196 685908 260248 685914
rect 260196 685850 260248 685856
rect 259840 673426 260144 673454
rect 239772 665304 239824 665310
rect 239772 665246 239824 665252
rect 239784 664714 239812 665246
rect 259840 664714 259868 673426
rect 239784 664686 240074 664714
rect 259394 664686 259868 664714
rect 249536 664142 249734 664170
rect 249536 663794 249564 664142
rect 249536 663766 249656 663794
rect 249628 662318 249656 663766
rect 260208 662318 260236 685850
rect 268028 683876 268056 685918
rect 277688 683876 277716 685986
rect 287336 685908 287388 685914
rect 287336 685850 287388 685856
rect 287348 683876 287376 685850
rect 266266 674248 266322 674257
rect 266266 674183 266322 674192
rect 262218 673568 262274 673577
rect 262218 673503 262274 673512
rect 262232 665174 262260 673503
rect 266280 665174 266308 674183
rect 262220 665168 262272 665174
rect 262220 665110 262272 665116
rect 266268 665168 266320 665174
rect 266268 665110 266320 665116
rect 287532 664714 287560 685986
rect 287704 685976 287756 685982
rect 287704 685918 287756 685924
rect 287716 665514 287744 685918
rect 289084 685908 289136 685914
rect 289084 685850 289136 685856
rect 287704 665508 287756 665514
rect 287704 665450 287756 665456
rect 287362 664686 287560 664714
rect 249616 662312 249668 662318
rect 249616 662254 249668 662260
rect 260196 662312 260248 662318
rect 260196 662254 260248 662260
rect 268028 662250 268056 664020
rect 277688 662386 277716 664020
rect 289096 662386 289124 685850
rect 296364 683890 296392 686054
rect 305368 686044 305420 686050
rect 305368 685986 305420 685992
rect 296056 683862 296392 683890
rect 305380 683890 305408 685986
rect 315488 685976 315540 685982
rect 315488 685918 315540 685924
rect 315028 685908 315080 685914
rect 315028 685850 315080 685856
rect 315040 683890 315068 685850
rect 305380 683862 305716 683890
rect 315040 683862 315376 683890
rect 289820 683188 289872 683194
rect 289820 683130 289872 683136
rect 293868 683188 293920 683194
rect 293868 683130 293920 683136
rect 289832 673577 289860 683130
rect 293880 674257 293908 683130
rect 293866 674248 293922 674257
rect 293866 674183 293922 674192
rect 289818 673568 289874 673577
rect 289818 673503 289874 673512
rect 295708 665508 295760 665514
rect 295708 665450 295760 665456
rect 295720 664714 295748 665450
rect 315500 664714 315528 685918
rect 316684 685908 316736 685914
rect 316684 685850 316736 685856
rect 295720 664686 296056 664714
rect 315376 664686 315528 664714
rect 305716 664006 306052 664034
rect 306024 662386 306052 664006
rect 316696 662386 316724 685850
rect 316788 665514 316816 686054
rect 317418 673568 317474 673577
rect 317418 673503 317474 673512
rect 316776 665508 316828 665514
rect 316776 665450 316828 665456
rect 317432 665174 317460 673503
rect 317420 665168 317472 665174
rect 317420 665110 317472 665116
rect 277676 662380 277728 662386
rect 277676 662322 277728 662328
rect 289084 662380 289136 662386
rect 289084 662322 289136 662328
rect 306012 662380 306064 662386
rect 306012 662322 306064 662328
rect 316684 662380 316736 662386
rect 316684 662322 316736 662328
rect 238852 662244 238904 662250
rect 238852 662186 238904 662192
rect 268016 662244 268068 662250
rect 268016 662186 268068 662192
rect 267832 658504 267884 658510
rect 267832 658446 267884 658452
rect 267004 658436 267056 658442
rect 267004 658378 267056 658384
rect 240600 658300 240652 658306
rect 240600 658242 240652 658248
rect 250260 658300 250312 658306
rect 250260 658242 250312 658248
rect 261484 658300 261536 658306
rect 261484 658242 261536 658248
rect 240612 656948 240640 658242
rect 250272 656948 250300 658242
rect 259946 656254 260144 656282
rect 238668 655648 238720 655654
rect 238668 655590 238720 655596
rect 238680 647465 238708 655590
rect 238666 647456 238722 647465
rect 238666 647391 238722 647400
rect 240612 634710 240640 637092
rect 240600 634704 240652 634710
rect 240600 634646 240652 634652
rect 250272 634642 250300 637092
rect 259932 634778 259960 637092
rect 260116 634778 260144 656254
rect 259920 634772 259972 634778
rect 259920 634714 259972 634720
rect 260104 634772 260156 634778
rect 260104 634714 260156 634720
rect 261496 634642 261524 658242
rect 262220 655580 262272 655586
rect 262220 655522 262272 655528
rect 266268 655580 266320 655586
rect 266268 655522 266320 655528
rect 262232 646785 262260 655522
rect 266280 647465 266308 655522
rect 266266 647456 266322 647465
rect 266266 647391 266322 647400
rect 262218 646776 262274 646785
rect 262218 646711 262274 646720
rect 267016 634710 267044 658378
rect 267844 654134 267872 658446
rect 295432 658436 295484 658442
rect 295432 658378 295484 658384
rect 268292 658300 268344 658306
rect 268292 658242 268344 658248
rect 277952 658300 278004 658306
rect 277952 658242 278004 658248
rect 289084 658300 289136 658306
rect 289084 658242 289136 658248
rect 268304 656962 268332 658242
rect 277964 656962 277992 658242
rect 268304 656934 268640 656962
rect 277964 656934 278300 656962
rect 287960 656254 288112 656282
rect 267844 654106 268240 654134
rect 268212 637786 268240 654106
rect 268212 637758 268640 637786
rect 278300 637078 278636 637106
rect 278608 634710 278636 637078
rect 287624 637078 287960 637106
rect 287624 634778 287652 637078
rect 288084 634778 288112 656254
rect 287612 634772 287664 634778
rect 287612 634714 287664 634720
rect 288072 634772 288124 634778
rect 288072 634714 288124 634720
rect 289096 634710 289124 658242
rect 289820 655648 289872 655654
rect 289820 655590 289872 655596
rect 293868 655648 293920 655654
rect 293868 655590 293920 655596
rect 289832 646785 289860 655590
rect 293880 647465 293908 655590
rect 295444 654134 295472 658378
rect 306288 658368 306340 658374
rect 306288 658310 306340 658316
rect 296628 658300 296680 658306
rect 296628 658242 296680 658248
rect 296640 656948 296668 658242
rect 306300 656948 306328 658310
rect 318064 658300 318116 658306
rect 318064 658242 318116 658248
rect 315974 656934 316172 656962
rect 316144 654134 316172 656934
rect 317420 655580 317472 655586
rect 317420 655522 317472 655528
rect 295444 654106 296208 654134
rect 316144 654106 316724 654134
rect 293866 647456 293922 647465
rect 293866 647391 293922 647400
rect 289818 646776 289874 646785
rect 289818 646711 289874 646720
rect 296180 637786 296208 654106
rect 296180 637758 296654 637786
rect 306300 634710 306328 637092
rect 315960 634778 315988 637092
rect 316696 634778 316724 654106
rect 317432 646785 317460 655522
rect 317418 646776 317474 646785
rect 317418 646711 317474 646720
rect 315948 634772 316000 634778
rect 315948 634714 316000 634720
rect 316684 634772 316736 634778
rect 316684 634714 316736 634720
rect 318076 634710 318104 658242
rect 267004 634704 267056 634710
rect 267004 634646 267056 634652
rect 278596 634704 278648 634710
rect 278596 634646 278648 634652
rect 289084 634704 289136 634710
rect 289084 634646 289136 634652
rect 306288 634704 306340 634710
rect 306288 634646 306340 634652
rect 318064 634704 318116 634710
rect 318064 634646 318116 634652
rect 250260 634636 250312 634642
rect 250260 634578 250312 634584
rect 261484 634636 261536 634642
rect 261484 634578 261536 634584
rect 296352 632324 296404 632330
rect 296352 632266 296404 632272
rect 316776 632324 316828 632330
rect 316776 632266 316828 632272
rect 260104 632256 260156 632262
rect 260104 632198 260156 632204
rect 277676 632256 277728 632262
rect 277676 632198 277728 632204
rect 287520 632256 287572 632262
rect 287520 632198 287572 632204
rect 249708 632188 249760 632194
rect 249708 632130 249760 632136
rect 249720 629884 249748 632130
rect 259368 632120 259420 632126
rect 259368 632062 259420 632068
rect 259380 629884 259408 632062
rect 238864 629326 240074 629354
rect 238666 620256 238722 620265
rect 238666 620191 238722 620200
rect 238680 611250 238708 620191
rect 238668 611244 238720 611250
rect 238668 611186 238720 611192
rect 238864 608462 238892 629326
rect 260116 615494 260144 632198
rect 268016 632188 268068 632194
rect 268016 632130 268068 632136
rect 260196 632120 260248 632126
rect 260196 632062 260248 632068
rect 259840 615466 260144 615494
rect 239772 611992 239824 611998
rect 239772 611934 239824 611940
rect 239784 610722 239812 611934
rect 259840 610722 259868 615466
rect 239784 610694 240074 610722
rect 259394 610694 259868 610722
rect 249720 608530 249748 610028
rect 260208 608530 260236 632062
rect 268028 629884 268056 632130
rect 277688 629884 277716 632198
rect 287336 632120 287388 632126
rect 287336 632062 287388 632068
rect 287348 629884 287376 632062
rect 266266 620256 266322 620265
rect 266266 620191 266322 620200
rect 262218 619576 262274 619585
rect 262218 619511 262274 619520
rect 262232 611318 262260 619511
rect 266280 611318 266308 620191
rect 262220 611312 262272 611318
rect 262220 611254 262272 611260
rect 266268 611312 266320 611318
rect 266268 611254 266320 611260
rect 287532 610722 287560 632198
rect 287704 632188 287756 632194
rect 287704 632130 287756 632136
rect 287716 611930 287744 632130
rect 289084 632120 289136 632126
rect 289084 632062 289136 632068
rect 287704 611924 287756 611930
rect 287704 611866 287756 611872
rect 287362 610694 287560 610722
rect 249708 608524 249760 608530
rect 249708 608466 249760 608472
rect 260196 608524 260248 608530
rect 260196 608466 260248 608472
rect 268028 608462 268056 610028
rect 277688 608598 277716 610028
rect 289096 608598 289124 632062
rect 296364 629898 296392 632266
rect 305368 632256 305420 632262
rect 305368 632198 305420 632204
rect 296056 629870 296392 629898
rect 305380 629898 305408 632198
rect 315488 632188 315540 632194
rect 315488 632130 315540 632136
rect 315028 632120 315080 632126
rect 315028 632062 315080 632068
rect 315040 629898 315068 632062
rect 305380 629870 305716 629898
rect 315040 629870 315376 629898
rect 293866 620256 293922 620265
rect 293866 620191 293922 620200
rect 289818 619576 289874 619585
rect 289818 619511 289874 619520
rect 289832 611250 289860 619511
rect 293880 611250 293908 620191
rect 295708 611924 295760 611930
rect 295708 611866 295760 611872
rect 289820 611244 289872 611250
rect 289820 611186 289872 611192
rect 293868 611244 293920 611250
rect 293868 611186 293920 611192
rect 295720 610722 295748 611866
rect 315500 610722 315528 632130
rect 316684 632120 316736 632126
rect 316684 632062 316736 632068
rect 295720 610694 296056 610722
rect 315376 610694 315528 610722
rect 305716 610014 306052 610042
rect 306024 608598 306052 610014
rect 316696 608598 316724 632062
rect 316788 611930 316816 632266
rect 317418 619576 317474 619585
rect 317418 619511 317474 619520
rect 316776 611924 316828 611930
rect 316776 611866 316828 611872
rect 317432 611318 317460 619511
rect 317420 611312 317472 611318
rect 317420 611254 317472 611260
rect 277676 608592 277728 608598
rect 277676 608534 277728 608540
rect 289084 608592 289136 608598
rect 289084 608534 289136 608540
rect 306012 608592 306064 608598
rect 306012 608534 306064 608540
rect 316684 608592 316736 608598
rect 316684 608534 316736 608540
rect 238852 608456 238904 608462
rect 238852 608398 238904 608404
rect 268016 608456 268068 608462
rect 268016 608398 268068 608404
rect 267004 604648 267056 604654
rect 267004 604590 267056 604596
rect 277952 604648 278004 604654
rect 277952 604590 278004 604596
rect 295432 604648 295484 604654
rect 295432 604590 295484 604596
rect 240600 604512 240652 604518
rect 240600 604454 240652 604460
rect 250260 604512 250312 604518
rect 250260 604454 250312 604460
rect 261484 604512 261536 604518
rect 261484 604454 261536 604460
rect 240612 602956 240640 604454
rect 250272 602956 250300 604454
rect 259946 602262 260144 602290
rect 238668 601792 238720 601798
rect 238668 601734 238720 601740
rect 238680 593473 238708 601734
rect 238666 593464 238722 593473
rect 238666 593399 238722 593408
rect 240612 580922 240640 583100
rect 240600 580916 240652 580922
rect 240600 580858 240652 580864
rect 250272 580854 250300 583100
rect 259932 580990 259960 583100
rect 260116 580990 260144 602262
rect 259920 580984 259972 580990
rect 259920 580926 259972 580932
rect 260104 580984 260156 580990
rect 260104 580926 260156 580932
rect 261496 580854 261524 604454
rect 262220 601724 262272 601730
rect 262220 601666 262272 601672
rect 266268 601724 266320 601730
rect 266268 601666 266320 601672
rect 262232 592793 262260 601666
rect 266280 593473 266308 601666
rect 266266 593464 266322 593473
rect 266266 593399 266322 593408
rect 262218 592784 262274 592793
rect 262218 592719 262274 592728
rect 267016 580922 267044 604590
rect 267832 604580 267884 604586
rect 267832 604522 267884 604528
rect 267844 596174 267872 604522
rect 268292 604512 268344 604518
rect 268292 604454 268344 604460
rect 268304 602970 268332 604454
rect 277964 602970 277992 604590
rect 289084 604512 289136 604518
rect 289084 604454 289136 604460
rect 268304 602942 268640 602970
rect 277964 602942 278300 602970
rect 287960 602262 288112 602290
rect 267844 596146 268240 596174
rect 268212 583794 268240 596146
rect 268212 583766 268640 583794
rect 278300 583086 278636 583114
rect 278608 580922 278636 583086
rect 287624 583086 287960 583114
rect 287624 580990 287652 583086
rect 288084 580990 288112 602262
rect 287612 580984 287664 580990
rect 287612 580926 287664 580932
rect 288072 580984 288124 580990
rect 288072 580926 288124 580932
rect 289096 580922 289124 604454
rect 289820 601792 289872 601798
rect 289820 601734 289872 601740
rect 293868 601792 293920 601798
rect 293868 601734 293920 601740
rect 289832 592793 289860 601734
rect 293880 593473 293908 601734
rect 295444 596174 295472 604590
rect 306288 604580 306340 604586
rect 306288 604522 306340 604528
rect 296628 604512 296680 604518
rect 296628 604454 296680 604460
rect 296640 602956 296668 604454
rect 306300 602956 306328 604522
rect 318064 604512 318116 604518
rect 318064 604454 318116 604460
rect 315974 602262 316080 602290
rect 316052 596174 316080 602262
rect 317420 601724 317472 601730
rect 317420 601666 317472 601672
rect 295444 596146 296208 596174
rect 316052 596146 316724 596174
rect 293866 593464 293922 593473
rect 293866 593399 293922 593408
rect 289818 592784 289874 592793
rect 289818 592719 289874 592728
rect 296180 583794 296208 596146
rect 296180 583766 296654 583794
rect 306300 580922 306328 583100
rect 315960 580990 315988 583100
rect 316696 580990 316724 596146
rect 317432 592793 317460 601666
rect 317418 592784 317474 592793
rect 317418 592719 317474 592728
rect 315948 580984 316000 580990
rect 315948 580926 316000 580932
rect 316684 580984 316736 580990
rect 316684 580926 316736 580932
rect 318076 580922 318104 604454
rect 267004 580916 267056 580922
rect 267004 580858 267056 580864
rect 278596 580916 278648 580922
rect 278596 580858 278648 580864
rect 289084 580916 289136 580922
rect 289084 580858 289136 580864
rect 306288 580916 306340 580922
rect 306288 580858 306340 580864
rect 318064 580916 318116 580922
rect 318064 580858 318116 580864
rect 250260 580848 250312 580854
rect 250260 580790 250312 580796
rect 261484 580848 261536 580854
rect 261484 580790 261536 580796
rect 296352 578468 296404 578474
rect 296352 578410 296404 578416
rect 316776 578468 316828 578474
rect 316776 578410 316828 578416
rect 260196 578400 260248 578406
rect 260196 578342 260248 578348
rect 277676 578400 277728 578406
rect 277676 578342 277728 578348
rect 287520 578400 287572 578406
rect 287520 578342 287572 578348
rect 249708 578332 249760 578338
rect 249708 578274 249760 578280
rect 249720 575892 249748 578274
rect 259368 578264 259420 578270
rect 259368 578206 259420 578212
rect 260104 578264 260156 578270
rect 260104 578206 260156 578212
rect 259380 575892 259408 578206
rect 238864 575334 240074 575362
rect 238666 566264 238722 566273
rect 238666 566199 238722 566208
rect 238680 557462 238708 566199
rect 238668 557456 238720 557462
rect 238668 557398 238720 557404
rect 238864 554606 238892 575334
rect 259736 562352 259788 562358
rect 259736 562294 259788 562300
rect 239772 558204 239824 558210
rect 239772 558146 239824 558152
rect 239784 556730 239812 558146
rect 259748 556730 259776 562294
rect 239784 556702 240074 556730
rect 259394 556702 259776 556730
rect 249720 554674 249748 556036
rect 260116 554674 260144 578206
rect 260208 562358 260236 578342
rect 268016 578332 268068 578338
rect 268016 578274 268068 578280
rect 268028 575892 268056 578274
rect 277688 575892 277716 578342
rect 287336 578264 287388 578270
rect 287336 578206 287388 578212
rect 287348 575892 287376 578206
rect 266266 566264 266322 566273
rect 266266 566199 266322 566208
rect 262218 565584 262274 565593
rect 262218 565519 262274 565528
rect 260196 562352 260248 562358
rect 260196 562294 260248 562300
rect 262232 557530 262260 565519
rect 266280 557530 266308 566199
rect 262220 557524 262272 557530
rect 262220 557466 262272 557472
rect 266268 557524 266320 557530
rect 266268 557466 266320 557472
rect 287532 556730 287560 578342
rect 287704 578332 287756 578338
rect 287704 578274 287756 578280
rect 287716 558890 287744 578274
rect 289084 578264 289136 578270
rect 289084 578206 289136 578212
rect 287704 558884 287756 558890
rect 287704 558826 287756 558832
rect 287362 556702 287560 556730
rect 249708 554668 249760 554674
rect 249708 554610 249760 554616
rect 260104 554668 260156 554674
rect 260104 554610 260156 554616
rect 268028 554606 268056 556036
rect 277688 554742 277716 556036
rect 289096 554742 289124 578206
rect 296364 575906 296392 578410
rect 305368 578400 305420 578406
rect 305368 578342 305420 578348
rect 296056 575878 296392 575906
rect 305380 575906 305408 578342
rect 315488 578332 315540 578338
rect 315488 578274 315540 578280
rect 315028 578264 315080 578270
rect 315028 578206 315080 578212
rect 315040 575906 315068 578206
rect 305380 575878 305716 575906
rect 315040 575878 315376 575906
rect 293866 566264 293922 566273
rect 293866 566199 293922 566208
rect 289818 565584 289874 565593
rect 289818 565519 289874 565528
rect 289832 557462 289860 565519
rect 293880 557462 293908 566199
rect 295708 558884 295760 558890
rect 295708 558826 295760 558832
rect 289820 557456 289872 557462
rect 289820 557398 289872 557404
rect 293868 557456 293920 557462
rect 293868 557398 293920 557404
rect 295720 556730 295748 558826
rect 315500 556730 315528 578274
rect 316684 578264 316736 578270
rect 316684 578206 316736 578212
rect 295720 556702 296056 556730
rect 315376 556702 315528 556730
rect 305716 556022 306052 556050
rect 306024 554742 306052 556022
rect 316696 554742 316724 578206
rect 316788 558890 316816 578410
rect 317418 565584 317474 565593
rect 317418 565519 317474 565528
rect 316776 558884 316828 558890
rect 316776 558826 316828 558832
rect 317432 557530 317460 565519
rect 317420 557524 317472 557530
rect 317420 557466 317472 557472
rect 277676 554736 277728 554742
rect 277676 554678 277728 554684
rect 289084 554736 289136 554742
rect 289084 554678 289136 554684
rect 306012 554736 306064 554742
rect 306012 554678 306064 554684
rect 316684 554736 316736 554742
rect 316684 554678 316736 554684
rect 238852 554600 238904 554606
rect 238852 554542 238904 554548
rect 268016 554600 268068 554606
rect 268016 554542 268068 554548
rect 267832 550792 267884 550798
rect 267832 550734 267884 550740
rect 295432 550792 295484 550798
rect 295432 550734 295484 550740
rect 267004 550724 267056 550730
rect 267004 550666 267056 550672
rect 240600 550656 240652 550662
rect 240600 550598 240652 550604
rect 250260 550656 250312 550662
rect 250260 550598 250312 550604
rect 261484 550656 261536 550662
rect 261484 550598 261536 550604
rect 240612 548964 240640 550598
rect 250272 548964 250300 550598
rect 259946 548270 260144 548298
rect 238666 539472 238722 539481
rect 238666 539407 238722 539416
rect 238680 529854 238708 539407
rect 238668 529848 238720 529854
rect 238668 529790 238720 529796
rect 240612 527066 240640 529108
rect 240600 527060 240652 527066
rect 240600 527002 240652 527008
rect 250272 526998 250300 529108
rect 259932 527134 259960 529108
rect 260116 527134 260144 548270
rect 259920 527128 259972 527134
rect 259920 527070 259972 527076
rect 260104 527128 260156 527134
rect 260104 527070 260156 527076
rect 261496 526998 261524 550598
rect 266266 539472 266322 539481
rect 266266 539407 266322 539416
rect 262218 538792 262274 538801
rect 262218 538727 262274 538736
rect 262232 529922 262260 538727
rect 266280 529922 266308 539407
rect 262220 529916 262272 529922
rect 262220 529858 262272 529864
rect 266268 529916 266320 529922
rect 266268 529858 266320 529864
rect 267016 527066 267044 550666
rect 267844 538214 267872 550734
rect 268292 550656 268344 550662
rect 268292 550598 268344 550604
rect 277952 550656 278004 550662
rect 277952 550598 278004 550604
rect 289084 550656 289136 550662
rect 289084 550598 289136 550604
rect 268304 548978 268332 550598
rect 277964 548978 277992 550598
rect 268304 548950 268640 548978
rect 277964 548950 278300 548978
rect 287960 548270 288112 548298
rect 267844 538186 268240 538214
rect 268212 529666 268240 538186
rect 268212 529638 268640 529666
rect 278300 529094 278636 529122
rect 278608 527066 278636 529094
rect 287624 529094 287960 529122
rect 287624 527134 287652 529094
rect 288084 527134 288112 548270
rect 287612 527128 287664 527134
rect 287612 527070 287664 527076
rect 288072 527128 288124 527134
rect 288072 527070 288124 527076
rect 289096 527066 289124 550598
rect 293866 539472 293922 539481
rect 293866 539407 293922 539416
rect 289818 538792 289874 538801
rect 289818 538727 289874 538736
rect 289832 529854 289860 538727
rect 293880 529854 293908 539407
rect 295444 538214 295472 550734
rect 306288 550724 306340 550730
rect 306288 550666 306340 550672
rect 296628 550656 296680 550662
rect 296628 550598 296680 550604
rect 296640 548964 296668 550598
rect 306300 548964 306328 550666
rect 318064 550656 318116 550662
rect 318064 550598 318116 550604
rect 315974 548270 316080 548298
rect 316052 547874 316080 548270
rect 316052 547846 316724 547874
rect 295444 538186 296208 538214
rect 289820 529848 289872 529854
rect 289820 529790 289872 529796
rect 293868 529848 293920 529854
rect 293868 529790 293920 529796
rect 296180 529666 296208 538186
rect 296180 529638 296654 529666
rect 306300 527066 306328 529108
rect 315960 527134 315988 529108
rect 316696 527134 316724 547846
rect 317418 538792 317474 538801
rect 317418 538727 317474 538736
rect 317432 529922 317460 538727
rect 317420 529916 317472 529922
rect 317420 529858 317472 529864
rect 315948 527128 316000 527134
rect 315948 527070 316000 527076
rect 316684 527128 316736 527134
rect 316684 527070 316736 527076
rect 318076 527066 318104 550598
rect 267004 527060 267056 527066
rect 267004 527002 267056 527008
rect 278596 527060 278648 527066
rect 278596 527002 278648 527008
rect 289084 527060 289136 527066
rect 289084 527002 289136 527008
rect 306288 527060 306340 527066
rect 306288 527002 306340 527008
rect 318064 527060 318116 527066
rect 318064 527002 318116 527008
rect 250260 526992 250312 526998
rect 250260 526934 250312 526940
rect 261484 526992 261536 526998
rect 261484 526934 261536 526940
rect 296352 523252 296404 523258
rect 296352 523194 296404 523200
rect 316776 523252 316828 523258
rect 316776 523194 316828 523200
rect 260196 523184 260248 523190
rect 260196 523126 260248 523132
rect 277676 523184 277728 523190
rect 277676 523126 277728 523132
rect 287520 523184 287572 523190
rect 287520 523126 287572 523132
rect 249708 523116 249760 523122
rect 249708 523058 249760 523064
rect 249720 521900 249748 523058
rect 259368 523048 259420 523054
rect 259368 522990 259420 522996
rect 260104 523048 260156 523054
rect 260104 522990 260156 522996
rect 259380 521900 259408 522990
rect 238864 521206 240074 521234
rect 238666 512272 238722 512281
rect 238666 512207 238722 512216
rect 238680 503674 238708 512207
rect 238668 503668 238720 503674
rect 238668 503610 238720 503616
rect 238864 500818 238892 521206
rect 259736 505640 259788 505646
rect 259736 505582 259788 505588
rect 239772 504280 239824 504286
rect 239772 504222 239824 504228
rect 239784 502738 239812 504222
rect 259748 502738 259776 505582
rect 239784 502710 240074 502738
rect 259394 502710 259776 502738
rect 249720 500886 249748 502044
rect 260116 500886 260144 522990
rect 260208 505646 260236 523126
rect 268016 523116 268068 523122
rect 268016 523058 268068 523064
rect 268028 521900 268056 523058
rect 277688 521900 277716 523126
rect 287336 523048 287388 523054
rect 287336 522990 287388 522996
rect 287348 521900 287376 522990
rect 262220 520328 262272 520334
rect 262220 520270 262272 520276
rect 266268 520328 266320 520334
rect 266268 520270 266320 520276
rect 262232 511601 262260 520270
rect 266280 512281 266308 520270
rect 266266 512272 266322 512281
rect 266266 512207 266322 512216
rect 262218 511592 262274 511601
rect 262218 511527 262274 511536
rect 260196 505640 260248 505646
rect 260196 505582 260248 505588
rect 287532 502738 287560 523126
rect 287704 523116 287756 523122
rect 287704 523058 287756 523064
rect 287716 504626 287744 523058
rect 289084 523048 289136 523054
rect 289084 522990 289136 522996
rect 287704 504620 287756 504626
rect 287704 504562 287756 504568
rect 287362 502710 287560 502738
rect 249708 500880 249760 500886
rect 249708 500822 249760 500828
rect 260104 500880 260156 500886
rect 260104 500822 260156 500828
rect 268028 500818 268056 502044
rect 277688 500954 277716 502044
rect 289096 500954 289124 522990
rect 296364 521914 296392 523194
rect 305368 523184 305420 523190
rect 305368 523126 305420 523132
rect 296056 521886 296392 521914
rect 305380 521914 305408 523126
rect 315488 523116 315540 523122
rect 315488 523058 315540 523064
rect 315028 523048 315080 523054
rect 315028 522990 315080 522996
rect 315040 521914 315068 522990
rect 305380 521886 305716 521914
rect 315040 521886 315376 521914
rect 293866 512272 293922 512281
rect 293866 512207 293922 512216
rect 289818 511592 289874 511601
rect 289818 511527 289874 511536
rect 289832 503674 289860 511527
rect 293880 503674 293908 512207
rect 295708 504620 295760 504626
rect 295708 504562 295760 504568
rect 289820 503668 289872 503674
rect 289820 503610 289872 503616
rect 293868 503668 293920 503674
rect 293868 503610 293920 503616
rect 295720 502738 295748 504562
rect 315500 502738 315528 523058
rect 316684 523048 316736 523054
rect 316684 522990 316736 522996
rect 295720 502710 296056 502738
rect 315376 502710 315528 502738
rect 305716 502030 306052 502058
rect 306024 500954 306052 502030
rect 316696 500954 316724 522990
rect 316788 503810 316816 523194
rect 317420 520328 317472 520334
rect 317420 520270 317472 520276
rect 317432 511601 317460 520270
rect 317418 511592 317474 511601
rect 317418 511527 317474 511536
rect 316776 503804 316828 503810
rect 316776 503746 316828 503752
rect 277676 500948 277728 500954
rect 277676 500890 277728 500896
rect 289084 500948 289136 500954
rect 289084 500890 289136 500896
rect 306012 500948 306064 500954
rect 306012 500890 306064 500896
rect 316684 500948 316736 500954
rect 316684 500890 316736 500896
rect 238852 500812 238904 500818
rect 238852 500754 238904 500760
rect 268016 500812 268068 500818
rect 268016 500754 268068 500760
rect 267004 497004 267056 497010
rect 267004 496946 267056 496952
rect 277952 497004 278004 497010
rect 277952 496946 278004 496952
rect 296168 497004 296220 497010
rect 296168 496946 296220 496952
rect 240600 496868 240652 496874
rect 240600 496810 240652 496816
rect 250260 496868 250312 496874
rect 250260 496810 250312 496816
rect 261484 496868 261536 496874
rect 261484 496810 261536 496816
rect 240612 494972 240640 496810
rect 250272 494972 250300 496810
rect 259946 494278 260144 494306
rect 238666 485480 238722 485489
rect 238666 485415 238722 485424
rect 238680 475998 238708 485415
rect 238668 475992 238720 475998
rect 238668 475934 238720 475940
rect 240612 473278 240640 475116
rect 240600 473272 240652 473278
rect 240600 473214 240652 473220
rect 250272 473210 250300 475116
rect 259932 473346 259960 475116
rect 260116 473346 260144 494278
rect 259920 473340 259972 473346
rect 259920 473282 259972 473288
rect 260104 473340 260156 473346
rect 260104 473282 260156 473288
rect 261496 473210 261524 496810
rect 266266 485480 266322 485489
rect 266266 485415 266322 485424
rect 262218 484800 262274 484809
rect 262218 484735 262274 484744
rect 262232 476066 262260 484735
rect 266280 476066 266308 485415
rect 262220 476060 262272 476066
rect 262220 476002 262272 476008
rect 266268 476060 266320 476066
rect 266268 476002 266320 476008
rect 267016 473278 267044 496946
rect 268200 496936 268252 496942
rect 268200 496878 268252 496884
rect 268212 475674 268240 496878
rect 268292 496868 268344 496874
rect 268292 496810 268344 496816
rect 268304 494986 268332 496810
rect 277964 494986 277992 496946
rect 289084 496868 289136 496874
rect 289084 496810 289136 496816
rect 268304 494958 268640 494986
rect 277964 494958 278300 494986
rect 287960 494278 288112 494306
rect 268212 475646 268640 475674
rect 278300 475102 278636 475130
rect 278608 473278 278636 475102
rect 287624 475102 287960 475130
rect 287624 473346 287652 475102
rect 288084 473346 288112 494278
rect 287612 473340 287664 473346
rect 287612 473282 287664 473288
rect 288072 473340 288124 473346
rect 288072 473282 288124 473288
rect 289096 473278 289124 496810
rect 293866 485480 293922 485489
rect 293866 485415 293922 485424
rect 289818 484800 289874 484809
rect 289818 484735 289874 484744
rect 289832 475998 289860 484735
rect 293880 475998 293908 485415
rect 289820 475992 289872 475998
rect 289820 475934 289872 475940
rect 293868 475992 293920 475998
rect 293868 475934 293920 475940
rect 296180 475674 296208 496946
rect 306288 496936 306340 496942
rect 306288 496878 306340 496884
rect 296628 496868 296680 496874
rect 296628 496810 296680 496816
rect 296640 494972 296668 496810
rect 306300 494972 306328 496878
rect 318064 496868 318116 496874
rect 318064 496810 318116 496816
rect 315974 494278 316172 494306
rect 316144 489914 316172 494278
rect 316144 489886 316724 489914
rect 296180 475646 296654 475674
rect 306300 473278 306328 475116
rect 315960 473346 315988 475116
rect 316696 473346 316724 489886
rect 317418 484800 317474 484809
rect 317418 484735 317474 484744
rect 317432 476066 317460 484735
rect 317420 476060 317472 476066
rect 317420 476002 317472 476008
rect 315948 473340 316000 473346
rect 315948 473282 316000 473288
rect 316684 473340 316736 473346
rect 316684 473282 316736 473288
rect 318076 473278 318104 496810
rect 267004 473272 267056 473278
rect 267004 473214 267056 473220
rect 278596 473272 278648 473278
rect 278596 473214 278648 473220
rect 289084 473272 289136 473278
rect 289084 473214 289136 473220
rect 306288 473272 306340 473278
rect 306288 473214 306340 473220
rect 318064 473272 318116 473278
rect 318064 473214 318116 473220
rect 250260 473204 250312 473210
rect 250260 473146 250312 473152
rect 261484 473204 261536 473210
rect 261484 473146 261536 473152
rect 296352 469464 296404 469470
rect 296352 469406 296404 469412
rect 316776 469464 316828 469470
rect 316776 469406 316828 469412
rect 260104 469396 260156 469402
rect 260104 469338 260156 469344
rect 277676 469396 277728 469402
rect 277676 469338 277728 469344
rect 287520 469396 287572 469402
rect 287520 469338 287572 469344
rect 249708 469328 249760 469334
rect 249708 469270 249760 469276
rect 249720 467908 249748 469270
rect 259368 469260 259420 469266
rect 259368 469202 259420 469208
rect 259380 467908 259408 469202
rect 238864 467214 240074 467242
rect 238668 466540 238720 466546
rect 238668 466482 238720 466488
rect 238680 458289 238708 466482
rect 238666 458280 238722 458289
rect 238666 458215 238722 458224
rect 238864 445602 238892 467214
rect 260116 451274 260144 469338
rect 268016 469328 268068 469334
rect 268016 469270 268068 469276
rect 260196 469260 260248 469266
rect 260196 469202 260248 469208
rect 259840 451246 260144 451274
rect 239772 449948 239824 449954
rect 239772 449890 239824 449896
rect 239784 448746 239812 449890
rect 259840 448746 259868 451246
rect 239784 448718 240074 448746
rect 259394 448718 259868 448746
rect 249720 445670 249748 448052
rect 260208 445670 260236 469202
rect 268028 467908 268056 469270
rect 277688 467908 277716 469338
rect 287336 469260 287388 469266
rect 287336 469202 287388 469208
rect 287348 467908 287376 469202
rect 262220 466472 262272 466478
rect 262220 466414 262272 466420
rect 266268 466472 266320 466478
rect 266268 466414 266320 466420
rect 262232 457609 262260 466414
rect 266280 458289 266308 466414
rect 266266 458280 266322 458289
rect 266266 458215 266322 458224
rect 262218 457600 262274 457609
rect 262218 457535 262274 457544
rect 287532 448746 287560 469338
rect 287704 469328 287756 469334
rect 287704 469270 287756 469276
rect 287716 449954 287744 469270
rect 289084 469260 289136 469266
rect 289084 469202 289136 469208
rect 287704 449948 287756 449954
rect 287704 449890 287756 449896
rect 287362 448718 287560 448746
rect 249708 445664 249760 445670
rect 249708 445606 249760 445612
rect 260196 445664 260248 445670
rect 260196 445606 260248 445612
rect 268028 445602 268056 448052
rect 277688 445738 277716 448052
rect 289096 445738 289124 469202
rect 296364 467922 296392 469406
rect 305368 469396 305420 469402
rect 305368 469338 305420 469344
rect 296056 467894 296392 467922
rect 305380 467922 305408 469338
rect 315488 469328 315540 469334
rect 315488 469270 315540 469276
rect 315028 469260 315080 469266
rect 315028 469202 315080 469208
rect 315040 467922 315068 469202
rect 305380 467894 305716 467922
rect 315040 467894 315376 467922
rect 289820 466540 289872 466546
rect 289820 466482 289872 466488
rect 293868 466540 293920 466546
rect 293868 466482 293920 466488
rect 289832 457609 289860 466482
rect 293880 458289 293908 466482
rect 293866 458280 293922 458289
rect 293866 458215 293922 458224
rect 289818 457600 289874 457609
rect 289818 457535 289874 457544
rect 295708 449948 295760 449954
rect 295708 449890 295760 449896
rect 295720 448746 295748 449890
rect 315500 448746 315528 469270
rect 316684 469260 316736 469266
rect 316684 469202 316736 469208
rect 295720 448718 296056 448746
rect 315376 448718 315528 448746
rect 305716 448038 306052 448066
rect 306024 445738 306052 448038
rect 316696 445738 316724 469202
rect 316788 449954 316816 469406
rect 317420 466472 317472 466478
rect 317420 466414 317472 466420
rect 317432 457609 317460 466414
rect 317418 457600 317474 457609
rect 317418 457535 317474 457544
rect 316776 449948 316828 449954
rect 316776 449890 316828 449896
rect 277676 445732 277728 445738
rect 277676 445674 277728 445680
rect 289084 445732 289136 445738
rect 289084 445674 289136 445680
rect 306012 445732 306064 445738
rect 306012 445674 306064 445680
rect 316684 445732 316736 445738
rect 316684 445674 316736 445680
rect 238852 445596 238904 445602
rect 238852 445538 238904 445544
rect 268016 445596 268068 445602
rect 268016 445538 268068 445544
rect 267004 443148 267056 443154
rect 267004 443090 267056 443096
rect 277952 443148 278004 443154
rect 277952 443090 278004 443096
rect 295432 443148 295484 443154
rect 295432 443090 295484 443096
rect 240600 443012 240652 443018
rect 240600 442954 240652 442960
rect 250260 443012 250312 443018
rect 250260 442954 250312 442960
rect 261484 443012 261536 443018
rect 261484 442954 261536 442960
rect 240612 440980 240640 442954
rect 250272 440980 250300 442954
rect 259946 440286 260144 440314
rect 238666 431488 238722 431497
rect 238666 431423 238722 431432
rect 238680 422278 238708 431423
rect 238668 422272 238720 422278
rect 238668 422214 238720 422220
rect 240612 419422 240640 421124
rect 240600 419416 240652 419422
rect 240600 419358 240652 419364
rect 250272 419354 250300 421124
rect 259932 419490 259960 421124
rect 260116 419490 260144 440286
rect 259920 419484 259972 419490
rect 259920 419426 259972 419432
rect 260104 419484 260156 419490
rect 260104 419426 260156 419432
rect 261496 419354 261524 442954
rect 262220 440292 262272 440298
rect 262220 440234 262272 440240
rect 266268 440292 266320 440298
rect 266268 440234 266320 440240
rect 262232 430817 262260 440234
rect 266280 431497 266308 440234
rect 266266 431488 266322 431497
rect 266266 431423 266322 431432
rect 262218 430808 262274 430817
rect 262218 430743 262274 430752
rect 267016 419422 267044 443090
rect 267832 443080 267884 443086
rect 267832 443022 267884 443028
rect 267844 441614 267872 443022
rect 268292 443012 268344 443018
rect 268292 442954 268344 442960
rect 267844 441586 268240 441614
rect 268212 421682 268240 441586
rect 268304 440994 268332 442954
rect 277964 440994 277992 443090
rect 289084 443012 289136 443018
rect 289084 442954 289136 442960
rect 268304 440966 268640 440994
rect 277964 440966 278300 440994
rect 287960 440286 288112 440314
rect 268212 421654 268640 421682
rect 278300 421110 278636 421138
rect 278608 419422 278636 421110
rect 287624 421110 287960 421138
rect 287624 419490 287652 421110
rect 288084 419490 288112 440286
rect 287612 419484 287664 419490
rect 287612 419426 287664 419432
rect 288072 419484 288124 419490
rect 288072 419426 288124 419432
rect 289096 419422 289124 442954
rect 295444 441614 295472 443090
rect 306288 443080 306340 443086
rect 306288 443022 306340 443028
rect 296628 443012 296680 443018
rect 296628 442954 296680 442960
rect 295444 441586 296208 441614
rect 293866 431488 293922 431497
rect 293866 431423 293922 431432
rect 289818 430808 289874 430817
rect 289818 430743 289874 430752
rect 289832 422278 289860 430743
rect 293880 422278 293908 431423
rect 289820 422272 289872 422278
rect 289820 422214 289872 422220
rect 293868 422272 293920 422278
rect 293868 422214 293920 422220
rect 296180 421682 296208 441586
rect 296640 440980 296668 442954
rect 306300 440980 306328 443022
rect 318064 443012 318116 443018
rect 318064 442954 318116 442960
rect 315974 440286 316172 440314
rect 316144 431954 316172 440286
rect 317420 440292 317472 440298
rect 317420 440234 317472 440240
rect 316144 431926 316724 431954
rect 296180 421654 296654 421682
rect 306300 419422 306328 421124
rect 315960 419490 315988 421124
rect 316696 419490 316724 431926
rect 317432 430817 317460 440234
rect 317418 430808 317474 430817
rect 317418 430743 317474 430752
rect 315948 419484 316000 419490
rect 315948 419426 316000 419432
rect 316684 419484 316736 419490
rect 316684 419426 316736 419432
rect 318076 419422 318104 442954
rect 267004 419416 267056 419422
rect 267004 419358 267056 419364
rect 278596 419416 278648 419422
rect 278596 419358 278648 419364
rect 289084 419416 289136 419422
rect 289084 419358 289136 419364
rect 306288 419416 306340 419422
rect 306288 419358 306340 419364
rect 318064 419416 318116 419422
rect 318064 419358 318116 419364
rect 250260 419348 250312 419354
rect 250260 419290 250312 419296
rect 261484 419348 261536 419354
rect 261484 419290 261536 419296
rect 296352 415676 296404 415682
rect 296352 415618 296404 415624
rect 316776 415676 316828 415682
rect 316776 415618 316828 415624
rect 260104 415608 260156 415614
rect 260104 415550 260156 415556
rect 277676 415608 277728 415614
rect 277676 415550 277728 415556
rect 287520 415608 287572 415614
rect 287520 415550 287572 415556
rect 249708 415540 249760 415546
rect 249708 415482 249760 415488
rect 249720 413916 249748 415482
rect 259368 415472 259420 415478
rect 259368 415414 259420 415420
rect 259380 413916 259408 415414
rect 238864 413222 240074 413250
rect 238666 404288 238722 404297
rect 238666 404223 238722 404232
rect 238680 394602 238708 404223
rect 238668 394596 238720 394602
rect 238668 394538 238720 394544
rect 238864 391814 238892 413222
rect 260116 402974 260144 415550
rect 268016 415540 268068 415546
rect 268016 415482 268068 415488
rect 260196 415472 260248 415478
rect 260196 415414 260248 415420
rect 259840 402946 260144 402974
rect 239772 395072 239824 395078
rect 239772 395014 239824 395020
rect 239784 394754 239812 395014
rect 259840 394754 259868 402946
rect 239784 394726 240074 394754
rect 259394 394726 259868 394754
rect 249720 391882 249748 394060
rect 260208 391882 260236 415414
rect 268028 413916 268056 415482
rect 277688 413916 277716 415550
rect 287336 415472 287388 415478
rect 287336 415414 287388 415420
rect 287348 413916 287376 415414
rect 266266 404288 266322 404297
rect 266266 404223 266322 404232
rect 262218 403608 262274 403617
rect 262218 403543 262274 403552
rect 262232 394670 262260 403543
rect 266280 394670 266308 404223
rect 287532 394754 287560 415550
rect 287704 415540 287756 415546
rect 287704 415482 287756 415488
rect 287716 395146 287744 415482
rect 289084 415472 289136 415478
rect 289084 415414 289136 415420
rect 287704 395140 287756 395146
rect 287704 395082 287756 395088
rect 287362 394726 287560 394754
rect 262220 394664 262272 394670
rect 262220 394606 262272 394612
rect 266268 394664 266320 394670
rect 266268 394606 266320 394612
rect 249708 391876 249760 391882
rect 249708 391818 249760 391824
rect 260196 391876 260248 391882
rect 260196 391818 260248 391824
rect 268028 391814 268056 394060
rect 277688 391950 277716 394060
rect 289096 391950 289124 415414
rect 296364 413930 296392 415618
rect 305368 415608 305420 415614
rect 305368 415550 305420 415556
rect 296056 413902 296392 413930
rect 305380 413930 305408 415550
rect 315488 415540 315540 415546
rect 315488 415482 315540 415488
rect 315028 415472 315080 415478
rect 315028 415414 315080 415420
rect 315040 413930 315068 415414
rect 305380 413902 305716 413930
rect 315040 413902 315376 413930
rect 293866 404288 293922 404297
rect 293866 404223 293922 404232
rect 289818 403608 289874 403617
rect 289818 403543 289874 403552
rect 289832 394602 289860 403543
rect 293880 394602 293908 404223
rect 295800 395140 295852 395146
rect 295800 395082 295852 395088
rect 295812 394754 295840 395082
rect 315500 394754 315528 415482
rect 316684 415472 316736 415478
rect 316684 415414 316736 415420
rect 295812 394726 296056 394754
rect 315376 394726 315528 394754
rect 289820 394596 289872 394602
rect 289820 394538 289872 394544
rect 293868 394596 293920 394602
rect 293868 394538 293920 394544
rect 305716 394046 306052 394074
rect 306024 391950 306052 394046
rect 316696 391950 316724 415414
rect 316788 395146 316816 415618
rect 317418 403608 317474 403617
rect 317418 403543 317474 403552
rect 316776 395140 316828 395146
rect 316776 395082 316828 395088
rect 317432 394670 317460 403543
rect 317420 394664 317472 394670
rect 317420 394606 317472 394612
rect 277676 391944 277728 391950
rect 277676 391886 277728 391892
rect 289084 391944 289136 391950
rect 289084 391886 289136 391892
rect 306012 391944 306064 391950
rect 306012 391886 306064 391892
rect 316684 391944 316736 391950
rect 316684 391886 316736 391892
rect 238852 391808 238904 391814
rect 238852 391750 238904 391756
rect 268016 391808 268068 391814
rect 268016 391750 268068 391756
rect 267004 389360 267056 389366
rect 267004 389302 267056 389308
rect 277952 389360 278004 389366
rect 277952 389302 278004 389308
rect 295432 389360 295484 389366
rect 295432 389302 295484 389308
rect 240600 389224 240652 389230
rect 240600 389166 240652 389172
rect 250260 389224 250312 389230
rect 250260 389166 250312 389172
rect 261484 389224 261536 389230
rect 261484 389166 261536 389172
rect 240612 386852 240640 389166
rect 250272 386852 250300 389166
rect 238668 386504 238720 386510
rect 238668 386446 238720 386452
rect 238680 377505 238708 386446
rect 259946 386294 260144 386322
rect 238666 377496 238722 377505
rect 238666 377431 238722 377440
rect 240612 365634 240640 367132
rect 240600 365628 240652 365634
rect 240600 365570 240652 365576
rect 250272 365566 250300 367132
rect 259932 365702 259960 367132
rect 260116 365702 260144 386294
rect 259920 365696 259972 365702
rect 259920 365638 259972 365644
rect 260104 365696 260156 365702
rect 260104 365638 260156 365644
rect 261496 365566 261524 389166
rect 262220 386436 262272 386442
rect 262220 386378 262272 386384
rect 266268 386436 266320 386442
rect 266268 386378 266320 386384
rect 262232 376825 262260 386378
rect 266280 377505 266308 386378
rect 266266 377496 266322 377505
rect 266266 377431 266322 377440
rect 262218 376816 262274 376825
rect 262218 376751 262274 376760
rect 267016 365634 267044 389302
rect 267832 389292 267884 389298
rect 267832 389234 267884 389240
rect 267844 383654 267872 389234
rect 268292 389224 268344 389230
rect 268292 389166 268344 389172
rect 268304 386866 268332 389166
rect 277964 386866 277992 389302
rect 289084 389224 289136 389230
rect 289084 389166 289136 389172
rect 268304 386838 268640 386866
rect 277964 386838 278300 386866
rect 287960 386294 288112 386322
rect 267844 383626 268240 383654
rect 268212 367690 268240 383626
rect 268212 367662 268640 367690
rect 278300 367118 278636 367146
rect 278608 365634 278636 367118
rect 287624 367118 287960 367146
rect 287624 365702 287652 367118
rect 288084 365702 288112 386294
rect 287612 365696 287664 365702
rect 287612 365638 287664 365644
rect 288072 365696 288124 365702
rect 288072 365638 288124 365644
rect 289096 365634 289124 389166
rect 289820 386504 289872 386510
rect 289820 386446 289872 386452
rect 293868 386504 293920 386510
rect 293868 386446 293920 386452
rect 289832 376825 289860 386446
rect 293880 377505 293908 386446
rect 295444 383654 295472 389302
rect 306288 389292 306340 389298
rect 306288 389234 306340 389240
rect 296628 389224 296680 389230
rect 296628 389166 296680 389172
rect 296640 386852 296668 389166
rect 306300 386852 306328 389234
rect 318064 389224 318116 389230
rect 318064 389166 318116 389172
rect 315974 386430 316080 386458
rect 316052 383654 316080 386430
rect 317420 386436 317472 386442
rect 317420 386378 317472 386384
rect 295444 383626 296208 383654
rect 316052 383626 316724 383654
rect 293866 377496 293922 377505
rect 293866 377431 293922 377440
rect 289818 376816 289874 376825
rect 289818 376751 289874 376760
rect 296180 367690 296208 383626
rect 296180 367662 296654 367690
rect 306300 365634 306328 367132
rect 315960 365702 315988 367132
rect 316696 365702 316724 383626
rect 317432 376825 317460 386378
rect 317418 376816 317474 376825
rect 317418 376751 317474 376760
rect 315948 365696 316000 365702
rect 315948 365638 316000 365644
rect 316684 365696 316736 365702
rect 316684 365638 316736 365644
rect 318076 365634 318104 389166
rect 267004 365628 267056 365634
rect 267004 365570 267056 365576
rect 278596 365628 278648 365634
rect 278596 365570 278648 365576
rect 289084 365628 289136 365634
rect 289084 365570 289136 365576
rect 306288 365628 306340 365634
rect 306288 365570 306340 365576
rect 318064 365628 318116 365634
rect 318064 365570 318116 365576
rect 250260 365560 250312 365566
rect 250260 365502 250312 365508
rect 261484 365560 261536 365566
rect 261484 365502 261536 365508
rect 249708 361752 249760 361758
rect 249708 361694 249760 361700
rect 260104 361752 260156 361758
rect 260104 361694 260156 361700
rect 277676 361752 277728 361758
rect 277676 361694 277728 361700
rect 296352 361752 296404 361758
rect 296352 361694 296404 361700
rect 316776 361752 316828 361758
rect 316776 361694 316828 361700
rect 249720 359924 249748 361694
rect 259368 361616 259420 361622
rect 259368 361558 259420 361564
rect 259380 359924 259408 361558
rect 238864 359230 240074 359258
rect 238666 350296 238722 350305
rect 238666 350231 238722 350240
rect 238680 340814 238708 350231
rect 238668 340808 238720 340814
rect 238668 340750 238720 340756
rect 238864 337958 238892 359230
rect 260116 345014 260144 361694
rect 268016 361684 268068 361690
rect 268016 361626 268068 361632
rect 260196 361616 260248 361622
rect 260196 361558 260248 361564
rect 259840 344986 260144 345014
rect 239772 341420 239824 341426
rect 239772 341362 239824 341368
rect 239784 340762 239812 341362
rect 259840 340762 259868 344986
rect 239784 340734 240074 340762
rect 259394 340734 259868 340762
rect 249720 338026 249748 340068
rect 260208 338026 260236 361558
rect 268028 359924 268056 361626
rect 277688 359924 277716 361694
rect 287704 361684 287756 361690
rect 287704 361626 287756 361632
rect 287336 361616 287388 361622
rect 287336 361558 287388 361564
rect 287348 359924 287376 361558
rect 287520 358828 287572 358834
rect 287520 358770 287572 358776
rect 266266 350296 266322 350305
rect 266266 350231 266322 350240
rect 262218 349616 262274 349625
rect 262218 349551 262274 349560
rect 262232 340882 262260 349551
rect 266280 340882 266308 350231
rect 262220 340876 262272 340882
rect 262220 340818 262272 340824
rect 266268 340876 266320 340882
rect 266268 340818 266320 340824
rect 287532 340762 287560 358770
rect 287716 341562 287744 361626
rect 289084 361616 289136 361622
rect 289084 361558 289136 361564
rect 287704 341556 287756 341562
rect 287704 341498 287756 341504
rect 287362 340734 287560 340762
rect 249708 338020 249760 338026
rect 249708 337962 249760 337968
rect 260196 338020 260248 338026
rect 260196 337962 260248 337968
rect 268028 337958 268056 340068
rect 277688 338094 277716 340068
rect 289096 338094 289124 361558
rect 296364 359938 296392 361694
rect 315488 361684 315540 361690
rect 315488 361626 315540 361632
rect 315028 361616 315080 361622
rect 315028 361558 315080 361564
rect 296056 359910 296392 359938
rect 315040 359938 315068 361558
rect 315040 359910 315376 359938
rect 305368 359304 305420 359310
rect 305420 359252 305716 359258
rect 305368 359246 305716 359252
rect 305380 359230 305716 359246
rect 293866 350296 293922 350305
rect 293866 350231 293922 350240
rect 289818 349616 289874 349625
rect 289818 349551 289874 349560
rect 289832 340814 289860 349551
rect 293880 340814 293908 350231
rect 295708 341556 295760 341562
rect 295708 341498 295760 341504
rect 289820 340808 289872 340814
rect 289820 340750 289872 340756
rect 293868 340808 293920 340814
rect 293868 340750 293920 340756
rect 295720 340762 295748 341498
rect 315500 340762 315528 361626
rect 316684 361616 316736 361622
rect 316684 361558 316736 361564
rect 295720 340734 296056 340762
rect 315376 340734 315528 340762
rect 305716 340054 306052 340082
rect 306024 338094 306052 340054
rect 316696 338094 316724 361558
rect 316788 341290 316816 361694
rect 317418 349616 317474 349625
rect 317418 349551 317474 349560
rect 316776 341284 316828 341290
rect 316776 341226 316828 341232
rect 317432 340882 317460 349551
rect 317420 340876 317472 340882
rect 317420 340818 317472 340824
rect 277676 338088 277728 338094
rect 277676 338030 277728 338036
rect 289084 338088 289136 338094
rect 289084 338030 289136 338036
rect 306012 338088 306064 338094
rect 306012 338030 306064 338036
rect 316684 338088 316736 338094
rect 316684 338030 316736 338036
rect 238852 337952 238904 337958
rect 238852 337894 238904 337900
rect 268016 337952 268068 337958
rect 268016 337894 268068 337900
rect 261484 335504 261536 335510
rect 261484 335446 261536 335452
rect 268292 335504 268344 335510
rect 268292 335446 268344 335452
rect 295432 335504 295484 335510
rect 295432 335446 295484 335452
rect 240600 335368 240652 335374
rect 240600 335310 240652 335316
rect 250260 335368 250312 335374
rect 250260 335310 250312 335316
rect 240612 332860 240640 335310
rect 250272 332860 250300 335310
rect 259946 332302 260144 332330
rect 238666 322960 238722 322969
rect 238666 322895 238722 322904
rect 238680 314634 238708 322895
rect 238668 314628 238720 314634
rect 238668 314570 238720 314576
rect 240612 311778 240640 313140
rect 240600 311772 240652 311778
rect 240600 311714 240652 311720
rect 250272 311710 250300 313140
rect 259932 311846 259960 313140
rect 260116 311846 260144 332302
rect 259920 311840 259972 311846
rect 259920 311782 259972 311788
rect 260104 311840 260156 311846
rect 260104 311782 260156 311788
rect 261496 311710 261524 335446
rect 267832 335436 267884 335442
rect 267832 335378 267884 335384
rect 267004 335368 267056 335374
rect 267004 335310 267056 335316
rect 262220 331356 262272 331362
rect 262220 331298 262272 331304
rect 262232 322833 262260 331298
rect 266266 322960 266322 322969
rect 266266 322895 266322 322904
rect 262218 322824 262274 322833
rect 262218 322759 262274 322768
rect 266280 314566 266308 322895
rect 266268 314560 266320 314566
rect 266268 314502 266320 314508
rect 267016 311778 267044 335310
rect 267844 325694 267872 335378
rect 268304 332874 268332 335446
rect 277952 335368 278004 335374
rect 277952 335310 278004 335316
rect 289084 335368 289136 335374
rect 289084 335310 289136 335316
rect 277964 332874 277992 335310
rect 268304 332846 268640 332874
rect 277964 332846 278300 332874
rect 287960 332302 288112 332330
rect 267844 325666 268240 325694
rect 268212 313698 268240 325666
rect 268212 313670 268640 313698
rect 278300 313126 278636 313154
rect 278608 311778 278636 313126
rect 287624 313126 287960 313154
rect 287624 311846 287652 313126
rect 288084 311846 288112 332302
rect 287612 311840 287664 311846
rect 287612 311782 287664 311788
rect 288072 311840 288124 311846
rect 288072 311782 288124 311788
rect 289096 311778 289124 335310
rect 293868 331288 293920 331294
rect 293868 331230 293920 331236
rect 293880 324057 293908 331230
rect 295444 325694 295472 335446
rect 306288 335436 306340 335442
rect 306288 335378 306340 335384
rect 296536 335368 296588 335374
rect 296536 335310 296588 335316
rect 296548 332874 296576 335310
rect 296548 332846 296654 332874
rect 306300 332860 306328 335378
rect 318064 335368 318116 335374
rect 318064 335310 318116 335316
rect 315974 332302 316172 332330
rect 316144 325694 316172 332302
rect 295444 325666 296208 325694
rect 316144 325666 316724 325694
rect 293866 324048 293922 324057
rect 293866 323983 293922 323992
rect 289818 322144 289874 322153
rect 289818 322079 289874 322088
rect 289832 314634 289860 322079
rect 289820 314628 289872 314634
rect 289820 314570 289872 314576
rect 296180 313698 296208 325666
rect 296180 313670 296654 313698
rect 306300 311778 306328 313140
rect 315960 311846 315988 313140
rect 316696 311846 316724 325666
rect 317418 322144 317474 322153
rect 317418 322079 317474 322088
rect 317432 314566 317460 322079
rect 317420 314560 317472 314566
rect 317420 314502 317472 314508
rect 315948 311840 316000 311846
rect 315948 311782 316000 311788
rect 316684 311840 316736 311846
rect 316684 311782 316736 311788
rect 318076 311778 318104 335310
rect 267004 311772 267056 311778
rect 267004 311714 267056 311720
rect 278596 311772 278648 311778
rect 278596 311714 278648 311720
rect 289084 311772 289136 311778
rect 289084 311714 289136 311720
rect 306288 311772 306340 311778
rect 306288 311714 306340 311720
rect 318064 311772 318116 311778
rect 318064 311714 318116 311720
rect 250260 311704 250312 311710
rect 250260 311646 250312 311652
rect 261484 311704 261536 311710
rect 261484 311646 261536 311652
rect 296352 308032 296404 308038
rect 296352 307974 296404 307980
rect 316776 308032 316828 308038
rect 316776 307974 316828 307980
rect 260196 307964 260248 307970
rect 260196 307906 260248 307912
rect 277676 307964 277728 307970
rect 277676 307906 277728 307912
rect 287520 307964 287572 307970
rect 287520 307906 287572 307912
rect 249708 307896 249760 307902
rect 249708 307838 249760 307844
rect 249720 305932 249748 307838
rect 259368 307828 259420 307834
rect 259368 307770 259420 307776
rect 260104 307828 260156 307834
rect 260104 307770 260156 307776
rect 259380 305932 259408 307770
rect 238864 305238 240074 305266
rect 238666 296304 238722 296313
rect 238666 296239 238722 296248
rect 238680 286958 238708 296239
rect 238668 286952 238720 286958
rect 238668 286894 238720 286900
rect 238864 284170 238892 305238
rect 259736 291916 259788 291922
rect 259736 291858 259788 291864
rect 239772 287972 239824 287978
rect 239772 287914 239824 287920
rect 239784 286770 239812 287914
rect 259748 286770 259776 291858
rect 239784 286742 240074 286770
rect 259394 286742 259776 286770
rect 249720 284238 249748 286076
rect 260116 284238 260144 307770
rect 260208 291922 260236 307906
rect 268016 307896 268068 307902
rect 268016 307838 268068 307844
rect 268028 305932 268056 307838
rect 277688 305932 277716 307906
rect 287336 307828 287388 307834
rect 287336 307770 287388 307776
rect 287348 305932 287376 307770
rect 266266 296304 266322 296313
rect 266266 296239 266322 296248
rect 262218 295624 262274 295633
rect 262218 295559 262274 295568
rect 260196 291916 260248 291922
rect 260196 291858 260248 291864
rect 262232 287026 262260 295559
rect 266280 287026 266308 296239
rect 262220 287020 262272 287026
rect 262220 286962 262272 286968
rect 266268 287020 266320 287026
rect 266268 286962 266320 286968
rect 287532 286770 287560 307906
rect 287704 307896 287756 307902
rect 287704 307838 287756 307844
rect 287716 288386 287744 307838
rect 289084 307828 289136 307834
rect 289084 307770 289136 307776
rect 287704 288380 287756 288386
rect 287704 288322 287756 288328
rect 287362 286742 287560 286770
rect 249708 284232 249760 284238
rect 249708 284174 249760 284180
rect 260104 284232 260156 284238
rect 260104 284174 260156 284180
rect 268028 284170 268056 286076
rect 277688 284306 277716 286076
rect 289096 284306 289124 307770
rect 296364 305946 296392 307974
rect 305368 307964 305420 307970
rect 305368 307906 305420 307912
rect 296056 305918 296392 305946
rect 305380 305946 305408 307906
rect 315488 307896 315540 307902
rect 315488 307838 315540 307844
rect 315028 307828 315080 307834
rect 315028 307770 315080 307776
rect 315040 305946 315068 307770
rect 305380 305918 305716 305946
rect 315040 305918 315376 305946
rect 293866 296304 293922 296313
rect 293866 296239 293922 296248
rect 289818 295624 289874 295633
rect 289818 295559 289874 295568
rect 289832 286958 289860 295559
rect 293880 286958 293908 296239
rect 295708 288380 295760 288386
rect 295708 288322 295760 288328
rect 289820 286952 289872 286958
rect 289820 286894 289872 286900
rect 293868 286952 293920 286958
rect 293868 286894 293920 286900
rect 295720 286770 295748 288322
rect 315500 286770 315528 307838
rect 316684 307828 316736 307834
rect 316684 307770 316736 307776
rect 295720 286742 296056 286770
rect 315376 286742 315528 286770
rect 305716 286062 306052 286090
rect 306024 284306 306052 286062
rect 316696 284306 316724 307770
rect 316788 288386 316816 307974
rect 317418 295624 317474 295633
rect 317418 295559 317474 295568
rect 316776 288380 316828 288386
rect 316776 288322 316828 288328
rect 317432 287026 317460 295559
rect 317420 287020 317472 287026
rect 317420 286962 317472 286968
rect 277676 284300 277728 284306
rect 277676 284242 277728 284248
rect 289084 284300 289136 284306
rect 289084 284242 289136 284248
rect 306012 284300 306064 284306
rect 306012 284242 306064 284248
rect 316684 284300 316736 284306
rect 316684 284242 316736 284248
rect 238852 284164 238904 284170
rect 238852 284106 238904 284112
rect 268016 284164 268068 284170
rect 268016 284106 268068 284112
rect 267004 280356 267056 280362
rect 267004 280298 267056 280304
rect 277952 280356 278004 280362
rect 277952 280298 278004 280304
rect 295432 280356 295484 280362
rect 295432 280298 295484 280304
rect 240600 280220 240652 280226
rect 240600 280162 240652 280168
rect 250260 280220 250312 280226
rect 250260 280162 250312 280168
rect 261484 280220 261536 280226
rect 261484 280162 261536 280168
rect 240612 278868 240640 280162
rect 250272 278868 250300 280162
rect 259946 278310 260144 278338
rect 238668 277432 238720 277438
rect 238668 277374 238720 277380
rect 238680 269929 238708 277374
rect 238666 269920 238722 269929
rect 238666 269855 238722 269864
rect 240612 256630 240640 259148
rect 240600 256624 240652 256630
rect 240600 256566 240652 256572
rect 250272 256562 250300 259148
rect 259932 256698 259960 259148
rect 260116 256698 260144 278310
rect 259920 256692 259972 256698
rect 259920 256634 259972 256640
rect 260104 256692 260156 256698
rect 260104 256634 260156 256640
rect 261496 256562 261524 280162
rect 262220 277500 262272 277506
rect 262220 277442 262272 277448
rect 266268 277500 266320 277506
rect 266268 277442 266320 277448
rect 262232 269113 262260 277442
rect 266280 269929 266308 277442
rect 266266 269920 266322 269929
rect 266266 269855 266322 269864
rect 262218 269104 262274 269113
rect 262218 269039 262274 269048
rect 267016 256630 267044 280298
rect 267832 280288 267884 280294
rect 267832 280230 267884 280236
rect 267844 267734 267872 280230
rect 268292 280220 268344 280226
rect 268292 280162 268344 280168
rect 268304 278882 268332 280162
rect 277964 278882 277992 280298
rect 289084 280220 289136 280226
rect 289084 280162 289136 280168
rect 268304 278854 268640 278882
rect 277964 278854 278300 278882
rect 287960 278310 288112 278338
rect 267844 267706 268240 267734
rect 268212 259706 268240 267706
rect 268212 259678 268640 259706
rect 278300 259134 278636 259162
rect 278608 256630 278636 259134
rect 287624 259134 287960 259162
rect 287624 256698 287652 259134
rect 288084 256698 288112 278310
rect 287612 256692 287664 256698
rect 287612 256634 287664 256640
rect 288072 256692 288124 256698
rect 288072 256634 288124 256640
rect 289096 256630 289124 280162
rect 289820 277432 289872 277438
rect 289820 277374 289872 277380
rect 293868 277432 293920 277438
rect 293868 277374 293920 277380
rect 289832 269113 289860 277374
rect 293880 270065 293908 277374
rect 293866 270056 293922 270065
rect 293866 269991 293922 270000
rect 289818 269104 289874 269113
rect 289818 269039 289874 269048
rect 295444 267734 295472 280298
rect 306288 280288 306340 280294
rect 306288 280230 306340 280236
rect 296628 280220 296680 280226
rect 296628 280162 296680 280168
rect 296640 278868 296668 280162
rect 306300 278868 306328 280230
rect 318064 280220 318116 280226
rect 318064 280162 318116 280168
rect 315974 278310 316172 278338
rect 316144 277394 316172 278310
rect 317420 277500 317472 277506
rect 317420 277442 317472 277448
rect 316144 277366 316724 277394
rect 295444 267706 296208 267734
rect 296180 259706 296208 267706
rect 296180 259678 296654 259706
rect 306300 256630 306328 259148
rect 315960 256698 315988 259148
rect 316696 256698 316724 277366
rect 317432 269113 317460 277442
rect 317418 269104 317474 269113
rect 317418 269039 317474 269048
rect 315948 256692 316000 256698
rect 315948 256634 316000 256640
rect 316684 256692 316736 256698
rect 316684 256634 316736 256640
rect 318076 256630 318104 280162
rect 267004 256624 267056 256630
rect 267004 256566 267056 256572
rect 278596 256624 278648 256630
rect 278596 256566 278648 256572
rect 289084 256624 289136 256630
rect 289084 256566 289136 256572
rect 306288 256624 306340 256630
rect 306288 256566 306340 256572
rect 318064 256624 318116 256630
rect 318064 256566 318116 256572
rect 250260 256556 250312 256562
rect 250260 256498 250312 256504
rect 261484 256556 261536 256562
rect 261484 256498 261536 256504
rect 296352 254176 296404 254182
rect 296352 254118 296404 254124
rect 316776 254176 316828 254182
rect 316776 254118 316828 254124
rect 260104 254108 260156 254114
rect 260104 254050 260156 254056
rect 277676 254108 277728 254114
rect 277676 254050 277728 254056
rect 287520 254108 287572 254114
rect 287520 254050 287572 254056
rect 249708 254040 249760 254046
rect 249708 253982 249760 253988
rect 249720 251940 249748 253982
rect 259368 253972 259420 253978
rect 259368 253914 259420 253920
rect 259380 251940 259408 253914
rect 238668 251320 238720 251326
rect 238668 251262 238720 251268
rect 238680 242321 238708 251262
rect 238864 251246 240074 251274
rect 238666 242312 238722 242321
rect 238666 242247 238722 242256
rect 238864 230314 238892 251246
rect 260116 238754 260144 254050
rect 268016 254040 268068 254046
rect 268016 253982 268068 253988
rect 260196 253972 260248 253978
rect 260196 253914 260248 253920
rect 259840 238726 260144 238754
rect 239772 233572 239824 233578
rect 239772 233514 239824 233520
rect 239784 232778 239812 233514
rect 259840 232778 259868 238726
rect 239784 232750 240074 232778
rect 259394 232750 259868 232778
rect 249720 230382 249748 232084
rect 260208 230382 260236 253914
rect 268028 251940 268056 253982
rect 277688 251940 277716 254050
rect 287336 253972 287388 253978
rect 287336 253914 287388 253920
rect 287348 251940 287376 253914
rect 262220 251252 262272 251258
rect 262220 251194 262272 251200
rect 266268 251252 266320 251258
rect 266268 251194 266320 251200
rect 262232 241641 262260 251194
rect 266280 242321 266308 251194
rect 266266 242312 266322 242321
rect 266266 242247 266322 242256
rect 262218 241632 262274 241641
rect 262218 241567 262274 241576
rect 287532 232778 287560 254050
rect 287704 254040 287756 254046
rect 287704 253982 287756 253988
rect 287716 233578 287744 253982
rect 289084 253972 289136 253978
rect 289084 253914 289136 253920
rect 287704 233572 287756 233578
rect 287704 233514 287756 233520
rect 287362 232750 287560 232778
rect 249708 230376 249760 230382
rect 249708 230318 249760 230324
rect 260196 230376 260248 230382
rect 260196 230318 260248 230324
rect 268028 230314 268056 232084
rect 277688 230450 277716 232084
rect 289096 230450 289124 253914
rect 296364 251954 296392 254118
rect 305368 254108 305420 254114
rect 305368 254050 305420 254056
rect 296056 251926 296392 251954
rect 305380 251954 305408 254050
rect 315488 254040 315540 254046
rect 315488 253982 315540 253988
rect 315028 253972 315080 253978
rect 315028 253914 315080 253920
rect 315040 251954 315068 253914
rect 305380 251926 305716 251954
rect 315040 251926 315376 251954
rect 289820 251320 289872 251326
rect 289820 251262 289872 251268
rect 293868 251320 293920 251326
rect 293868 251262 293920 251268
rect 289832 241641 289860 251262
rect 293880 242321 293908 251262
rect 293866 242312 293922 242321
rect 293866 242247 293922 242256
rect 289818 241632 289874 241641
rect 289818 241567 289874 241576
rect 295708 233572 295760 233578
rect 295708 233514 295760 233520
rect 295720 232778 295748 233514
rect 315500 232778 315528 253982
rect 316684 253972 316736 253978
rect 316684 253914 316736 253920
rect 295720 232750 296056 232778
rect 315376 232750 315528 232778
rect 305716 232070 306052 232098
rect 306024 230450 306052 232070
rect 316696 230450 316724 253914
rect 316788 233442 316816 254118
rect 317420 251252 317472 251258
rect 317420 251194 317472 251200
rect 317432 241641 317460 251194
rect 317418 241632 317474 241641
rect 317418 241567 317474 241576
rect 316776 233436 316828 233442
rect 316776 233378 316828 233384
rect 277676 230444 277728 230450
rect 277676 230386 277728 230392
rect 289084 230444 289136 230450
rect 289084 230386 289136 230392
rect 306012 230444 306064 230450
rect 306012 230386 306064 230392
rect 316684 230444 316736 230450
rect 316684 230386 316736 230392
rect 238852 230308 238904 230314
rect 238852 230250 238904 230256
rect 268016 230308 268068 230314
rect 268016 230250 268068 230256
rect 261484 226500 261536 226506
rect 261484 226442 261536 226448
rect 268292 226500 268344 226506
rect 268292 226442 268344 226448
rect 296168 226500 296220 226506
rect 296168 226442 296220 226448
rect 240600 226364 240652 226370
rect 240600 226306 240652 226312
rect 250260 226364 250312 226370
rect 250260 226306 250312 226312
rect 240612 224876 240640 226306
rect 250272 224876 250300 226306
rect 259946 224318 260144 224346
rect 238668 223712 238720 223718
rect 238668 223654 238720 223660
rect 238680 215393 238708 223654
rect 238666 215384 238722 215393
rect 238666 215319 238722 215328
rect 240612 202774 240640 205020
rect 240600 202768 240652 202774
rect 240600 202710 240652 202716
rect 250272 202706 250300 205020
rect 259932 202842 259960 205020
rect 260116 202842 260144 224318
rect 259920 202836 259972 202842
rect 259920 202778 259972 202784
rect 260104 202836 260156 202842
rect 260104 202778 260156 202784
rect 261496 202706 261524 226442
rect 268200 226432 268252 226438
rect 268200 226374 268252 226380
rect 267004 226364 267056 226370
rect 267004 226306 267056 226312
rect 262220 223644 262272 223650
rect 262220 223586 262272 223592
rect 266268 223644 266320 223650
rect 266268 223586 266320 223592
rect 262232 214713 262260 223586
rect 266280 215393 266308 223586
rect 266266 215384 266322 215393
rect 266266 215319 266322 215328
rect 262218 214704 262274 214713
rect 262218 214639 262274 214648
rect 267016 202774 267044 226306
rect 268212 205714 268240 226374
rect 268304 224890 268332 226442
rect 277952 226364 278004 226370
rect 277952 226306 278004 226312
rect 289084 226364 289136 226370
rect 289084 226306 289136 226312
rect 277964 224890 277992 226306
rect 268304 224862 268640 224890
rect 277964 224862 278300 224890
rect 287960 224318 288112 224346
rect 268212 205686 268640 205714
rect 278300 205006 278636 205034
rect 278608 202774 278636 205006
rect 287624 205006 287960 205034
rect 287624 202842 287652 205006
rect 288084 202842 288112 224318
rect 287612 202836 287664 202842
rect 287612 202778 287664 202784
rect 288072 202836 288124 202842
rect 288072 202778 288124 202784
rect 289096 202774 289124 226306
rect 289820 223712 289872 223718
rect 289820 223654 289872 223660
rect 293868 223712 293920 223718
rect 293868 223654 293920 223660
rect 289832 214713 289860 223654
rect 293880 215393 293908 223654
rect 293866 215384 293922 215393
rect 293866 215319 293922 215328
rect 289818 214704 289874 214713
rect 289818 214639 289874 214648
rect 296180 205714 296208 226442
rect 306288 226432 306340 226438
rect 306288 226374 306340 226380
rect 296628 226364 296680 226370
rect 296628 226306 296680 226312
rect 296640 224876 296668 226306
rect 306300 224876 306328 226374
rect 318064 226364 318116 226370
rect 318064 226306 318116 226312
rect 315974 224318 316172 224346
rect 316144 219434 316172 224318
rect 317420 223644 317472 223650
rect 317420 223586 317472 223592
rect 316144 219406 316724 219434
rect 296180 205686 296654 205714
rect 306300 202774 306328 205020
rect 315960 202842 315988 205020
rect 316696 202842 316724 219406
rect 317432 214713 317460 223586
rect 317418 214704 317474 214713
rect 317418 214639 317474 214648
rect 315948 202836 316000 202842
rect 315948 202778 316000 202784
rect 316684 202836 316736 202842
rect 316684 202778 316736 202784
rect 318076 202774 318104 226306
rect 267004 202768 267056 202774
rect 267004 202710 267056 202716
rect 278596 202768 278648 202774
rect 278596 202710 278648 202716
rect 289084 202768 289136 202774
rect 289084 202710 289136 202716
rect 306288 202768 306340 202774
rect 306288 202710 306340 202716
rect 318064 202768 318116 202774
rect 318064 202710 318116 202716
rect 250260 202700 250312 202706
rect 250260 202642 250312 202648
rect 261484 202700 261536 202706
rect 261484 202642 261536 202648
rect 296352 200388 296404 200394
rect 296352 200330 296404 200336
rect 316776 200388 316828 200394
rect 316776 200330 316828 200336
rect 249708 200320 249760 200326
rect 249708 200262 249760 200268
rect 260196 200320 260248 200326
rect 260196 200262 260248 200268
rect 277676 200320 277728 200326
rect 277676 200262 277728 200268
rect 287520 200320 287572 200326
rect 287520 200262 287572 200268
rect 249720 197948 249748 200262
rect 259368 200184 259420 200190
rect 259368 200126 259420 200132
rect 260104 200184 260156 200190
rect 260104 200126 260156 200132
rect 259380 197948 259408 200126
rect 238864 197254 240074 197282
rect 238666 188320 238722 188329
rect 238666 188255 238722 188264
rect 238680 179314 238708 188255
rect 238668 179308 238720 179314
rect 238668 179250 238720 179256
rect 238864 176526 238892 197254
rect 259736 185632 259788 185638
rect 259736 185574 259788 185580
rect 239772 179920 239824 179926
rect 239772 179862 239824 179868
rect 239784 178786 239812 179862
rect 259748 178786 259776 185574
rect 239784 178758 240074 178786
rect 259394 178758 259776 178786
rect 249720 176594 249748 178092
rect 260116 176594 260144 200126
rect 260208 185638 260236 200262
rect 268016 200252 268068 200258
rect 268016 200194 268068 200200
rect 268028 197948 268056 200194
rect 277688 197948 277716 200262
rect 287336 200184 287388 200190
rect 287336 200126 287388 200132
rect 287348 197948 287376 200126
rect 266266 188320 266322 188329
rect 266266 188255 266322 188264
rect 262218 187640 262274 187649
rect 262218 187575 262274 187584
rect 260196 185632 260248 185638
rect 260196 185574 260248 185580
rect 262232 179382 262260 187575
rect 266280 179382 266308 188255
rect 262220 179376 262272 179382
rect 262220 179318 262272 179324
rect 266268 179376 266320 179382
rect 266268 179318 266320 179324
rect 287532 178786 287560 200262
rect 287704 200252 287756 200258
rect 287704 200194 287756 200200
rect 287716 179450 287744 200194
rect 289084 200184 289136 200190
rect 289084 200126 289136 200132
rect 287704 179444 287756 179450
rect 287704 179386 287756 179392
rect 287362 178758 287560 178786
rect 249708 176588 249760 176594
rect 249708 176530 249760 176536
rect 260104 176588 260156 176594
rect 260104 176530 260156 176536
rect 268028 176526 268056 178092
rect 277688 176662 277716 178092
rect 289096 176662 289124 200126
rect 296364 197962 296392 200330
rect 305368 200320 305420 200326
rect 305368 200262 305420 200268
rect 296056 197934 296392 197962
rect 305380 197962 305408 200262
rect 315488 200252 315540 200258
rect 315488 200194 315540 200200
rect 315028 200184 315080 200190
rect 315028 200126 315080 200132
rect 315040 197962 315068 200126
rect 305380 197934 305716 197962
rect 315040 197934 315376 197962
rect 293866 188320 293922 188329
rect 293866 188255 293922 188264
rect 289818 187640 289874 187649
rect 289818 187575 289874 187584
rect 289832 179314 289860 187575
rect 293880 179314 293908 188255
rect 295708 179444 295760 179450
rect 295708 179386 295760 179392
rect 289820 179308 289872 179314
rect 289820 179250 289872 179256
rect 293868 179308 293920 179314
rect 293868 179250 293920 179256
rect 295720 178786 295748 179386
rect 315500 178786 315528 200194
rect 316684 200184 316736 200190
rect 316684 200126 316736 200132
rect 295720 178758 296056 178786
rect 315376 178758 315528 178786
rect 305716 178078 306052 178106
rect 306024 176662 306052 178078
rect 316696 176662 316724 200126
rect 316788 179518 316816 200330
rect 317418 187640 317474 187649
rect 317418 187575 317474 187584
rect 316776 179512 316828 179518
rect 316776 179454 316828 179460
rect 317432 179382 317460 187575
rect 317420 179376 317472 179382
rect 317420 179318 317472 179324
rect 277676 176656 277728 176662
rect 277676 176598 277728 176604
rect 289084 176656 289136 176662
rect 289084 176598 289136 176604
rect 306012 176656 306064 176662
rect 306012 176598 306064 176604
rect 316684 176656 316736 176662
rect 316684 176598 316736 176604
rect 238852 176520 238904 176526
rect 238852 176462 238904 176468
rect 268016 176520 268068 176526
rect 268016 176462 268068 176468
rect 261484 172712 261536 172718
rect 261484 172654 261536 172660
rect 268292 172712 268344 172718
rect 268292 172654 268344 172660
rect 295432 172712 295484 172718
rect 295432 172654 295484 172660
rect 240600 172576 240652 172582
rect 240600 172518 240652 172524
rect 250260 172576 250312 172582
rect 250260 172518 250312 172524
rect 240612 170884 240640 172518
rect 250272 170884 250300 172518
rect 259946 170326 260144 170354
rect 238666 161392 238722 161401
rect 238666 161327 238722 161336
rect 238680 151706 238708 161327
rect 238668 151700 238720 151706
rect 238668 151642 238720 151648
rect 240612 148986 240640 151028
rect 240600 148980 240652 148986
rect 240600 148922 240652 148928
rect 250272 148918 250300 151028
rect 259932 149054 259960 151028
rect 260116 149054 260144 170326
rect 259920 149048 259972 149054
rect 259920 148990 259972 148996
rect 260104 149048 260156 149054
rect 260104 148990 260156 148996
rect 261496 148918 261524 172654
rect 267832 172644 267884 172650
rect 267832 172586 267884 172592
rect 267004 172576 267056 172582
rect 267004 172518 267056 172524
rect 266266 161392 266322 161401
rect 266266 161327 266322 161336
rect 262218 160712 262274 160721
rect 262218 160647 262274 160656
rect 262232 151774 262260 160647
rect 266280 151774 266308 161327
rect 262220 151768 262272 151774
rect 262220 151710 262272 151716
rect 266268 151768 266320 151774
rect 266268 151710 266320 151716
rect 267016 148986 267044 172518
rect 267844 171134 267872 172586
rect 267844 171106 268240 171134
rect 268212 151722 268240 171106
rect 268304 170898 268332 172654
rect 277952 172576 278004 172582
rect 277952 172518 278004 172524
rect 289084 172576 289136 172582
rect 289084 172518 289136 172524
rect 277964 170898 277992 172518
rect 268304 170870 268640 170898
rect 277964 170870 278300 170898
rect 287960 170326 288112 170354
rect 268212 151694 268640 151722
rect 278300 151014 278636 151042
rect 278608 148986 278636 151014
rect 287624 151014 287960 151042
rect 287624 149054 287652 151014
rect 288084 149054 288112 170326
rect 287612 149048 287664 149054
rect 287612 148990 287664 148996
rect 288072 149048 288124 149054
rect 288072 148990 288124 148996
rect 289096 148986 289124 172518
rect 295444 171134 295472 172654
rect 306288 172644 306340 172650
rect 306288 172586 306340 172592
rect 296628 172576 296680 172582
rect 296628 172518 296680 172524
rect 295444 171106 296208 171134
rect 293866 161392 293922 161401
rect 293866 161327 293922 161336
rect 289818 160712 289874 160721
rect 289818 160647 289874 160656
rect 289832 151706 289860 160647
rect 293880 151706 293908 161327
rect 296180 151722 296208 171106
rect 296640 170884 296668 172518
rect 306300 170884 306328 172586
rect 318064 172576 318116 172582
rect 318064 172518 318116 172524
rect 315974 170326 316080 170354
rect 316052 161474 316080 170326
rect 316052 161446 316724 161474
rect 289820 151700 289872 151706
rect 289820 151642 289872 151648
rect 293868 151700 293920 151706
rect 296180 151694 296654 151722
rect 293868 151642 293920 151648
rect 306300 148986 306328 151028
rect 315960 149054 315988 151028
rect 316696 149054 316724 161446
rect 317418 160712 317474 160721
rect 317418 160647 317474 160656
rect 317432 151774 317460 160647
rect 317420 151768 317472 151774
rect 317420 151710 317472 151716
rect 315948 149048 316000 149054
rect 315948 148990 316000 148996
rect 316684 149048 316736 149054
rect 316684 148990 316736 148996
rect 318076 148986 318104 172518
rect 267004 148980 267056 148986
rect 267004 148922 267056 148928
rect 278596 148980 278648 148986
rect 278596 148922 278648 148928
rect 289084 148980 289136 148986
rect 289084 148922 289136 148928
rect 306288 148980 306340 148986
rect 306288 148922 306340 148928
rect 318064 148980 318116 148986
rect 318064 148922 318116 148928
rect 250260 148912 250312 148918
rect 250260 148854 250312 148860
rect 261484 148912 261536 148918
rect 261484 148854 261536 148860
rect 296352 146532 296404 146538
rect 296352 146474 296404 146480
rect 316776 146532 316828 146538
rect 316776 146474 316828 146480
rect 260196 146464 260248 146470
rect 260196 146406 260248 146412
rect 277676 146464 277728 146470
rect 277676 146406 277728 146412
rect 287520 146464 287572 146470
rect 287520 146406 287572 146412
rect 249708 146396 249760 146402
rect 249708 146338 249760 146344
rect 249720 143956 249748 146338
rect 259368 146328 259420 146334
rect 259368 146270 259420 146276
rect 260104 146328 260156 146334
rect 260104 146270 260156 146276
rect 259380 143956 259408 146270
rect 238864 143262 240074 143290
rect 238666 134328 238722 134337
rect 238666 134263 238722 134272
rect 238680 125526 238708 134263
rect 238668 125520 238720 125526
rect 238668 125462 238720 125468
rect 238864 122670 238892 143262
rect 259736 128308 259788 128314
rect 259736 128250 259788 128256
rect 239772 126948 239824 126954
rect 239772 126890 239824 126896
rect 239784 124794 239812 126890
rect 259748 124794 259776 128250
rect 239784 124766 240074 124794
rect 259394 124766 259776 124794
rect 249720 122738 249748 124100
rect 260116 122738 260144 146270
rect 260208 128314 260236 146406
rect 268016 146396 268068 146402
rect 268016 146338 268068 146344
rect 268028 143956 268056 146338
rect 277688 143956 277716 146406
rect 287336 146328 287388 146334
rect 287336 146270 287388 146276
rect 287348 143956 287376 146270
rect 266266 134328 266322 134337
rect 266266 134263 266322 134272
rect 262218 133648 262274 133657
rect 262218 133583 262274 133592
rect 260196 128308 260248 128314
rect 260196 128250 260248 128256
rect 262232 125594 262260 133583
rect 266280 125594 266308 134263
rect 262220 125588 262272 125594
rect 262220 125530 262272 125536
rect 266268 125588 266320 125594
rect 266268 125530 266320 125536
rect 287532 124794 287560 146406
rect 287704 146396 287756 146402
rect 287704 146338 287756 146344
rect 287716 126138 287744 146338
rect 289084 146328 289136 146334
rect 289084 146270 289136 146276
rect 287704 126132 287756 126138
rect 287704 126074 287756 126080
rect 287362 124766 287560 124794
rect 249708 122732 249760 122738
rect 249708 122674 249760 122680
rect 260104 122732 260156 122738
rect 260104 122674 260156 122680
rect 268028 122670 268056 124100
rect 277688 122806 277716 124100
rect 289096 122806 289124 146270
rect 296364 143970 296392 146474
rect 305368 146464 305420 146470
rect 305368 146406 305420 146412
rect 296056 143942 296392 143970
rect 305380 143970 305408 146406
rect 315488 146396 315540 146402
rect 315488 146338 315540 146344
rect 315028 146328 315080 146334
rect 315028 146270 315080 146276
rect 315040 143970 315068 146270
rect 305380 143942 305716 143970
rect 315040 143942 315376 143970
rect 293866 134328 293922 134337
rect 293866 134263 293922 134272
rect 289818 133648 289874 133657
rect 289818 133583 289874 133592
rect 289832 125526 289860 133583
rect 293880 125526 293908 134263
rect 295708 126132 295760 126138
rect 295708 126074 295760 126080
rect 289820 125520 289872 125526
rect 289820 125462 289872 125468
rect 293868 125520 293920 125526
rect 293868 125462 293920 125468
rect 295720 124794 295748 126074
rect 315500 124794 315528 146338
rect 316684 146328 316736 146334
rect 316684 146270 316736 146276
rect 295720 124766 296056 124794
rect 315376 124766 315528 124794
rect 305716 124086 306052 124114
rect 306024 122806 306052 124086
rect 316696 122806 316724 146270
rect 316788 126138 316816 146474
rect 317418 133648 317474 133657
rect 317418 133583 317474 133592
rect 316776 126132 316828 126138
rect 316776 126074 316828 126080
rect 317432 125594 317460 133583
rect 317420 125588 317472 125594
rect 317420 125530 317472 125536
rect 277676 122800 277728 122806
rect 277676 122742 277728 122748
rect 289084 122800 289136 122806
rect 289084 122742 289136 122748
rect 306012 122800 306064 122806
rect 306012 122742 306064 122748
rect 316684 122800 316736 122806
rect 316684 122742 316736 122748
rect 238852 122664 238904 122670
rect 238852 122606 238904 122612
rect 268016 122664 268068 122670
rect 268016 122606 268068 122612
rect 267004 118856 267056 118862
rect 267004 118798 267056 118804
rect 277952 118856 278004 118862
rect 277952 118798 278004 118804
rect 295432 118856 295484 118862
rect 295432 118798 295484 118804
rect 240600 118720 240652 118726
rect 240600 118662 240652 118668
rect 250260 118720 250312 118726
rect 250260 118662 250312 118668
rect 261484 118720 261536 118726
rect 261484 118662 261536 118668
rect 240612 116892 240640 118662
rect 250272 116892 250300 118662
rect 259946 116334 260144 116362
rect 238666 107400 238722 107409
rect 238666 107335 238722 107344
rect 238680 97918 238708 107335
rect 238668 97912 238720 97918
rect 238668 97854 238720 97860
rect 240612 95130 240640 97036
rect 240600 95124 240652 95130
rect 240600 95066 240652 95072
rect 250272 95062 250300 97036
rect 259932 95198 259960 97036
rect 260116 95198 260144 116334
rect 259920 95192 259972 95198
rect 259920 95134 259972 95140
rect 260104 95192 260156 95198
rect 260104 95134 260156 95140
rect 261496 95062 261524 118662
rect 266266 107400 266322 107409
rect 266266 107335 266322 107344
rect 262218 106720 262274 106729
rect 262218 106655 262274 106664
rect 262232 97986 262260 106655
rect 266280 97986 266308 107335
rect 262220 97980 262272 97986
rect 262220 97922 262272 97928
rect 266268 97980 266320 97986
rect 266268 97922 266320 97928
rect 267016 95130 267044 118798
rect 267832 118788 267884 118794
rect 267832 118730 267884 118736
rect 267844 113174 267872 118730
rect 268292 118720 268344 118726
rect 268292 118662 268344 118668
rect 268304 116906 268332 118662
rect 277964 116906 277992 118798
rect 289084 118720 289136 118726
rect 289084 118662 289136 118668
rect 268304 116878 268640 116906
rect 277964 116878 278300 116906
rect 287960 116334 288112 116362
rect 267844 113146 268240 113174
rect 268212 97730 268240 113146
rect 268212 97702 268640 97730
rect 278300 97022 278636 97050
rect 278608 95130 278636 97022
rect 287624 97022 287960 97050
rect 287624 95198 287652 97022
rect 288084 95198 288112 116334
rect 287612 95192 287664 95198
rect 287612 95134 287664 95140
rect 288072 95192 288124 95198
rect 288072 95134 288124 95140
rect 289096 95130 289124 118662
rect 295444 113174 295472 118798
rect 306288 118788 306340 118794
rect 306288 118730 306340 118736
rect 296628 118720 296680 118726
rect 296628 118662 296680 118668
rect 296640 116892 296668 118662
rect 306300 116892 306328 118730
rect 318064 118720 318116 118726
rect 318064 118662 318116 118668
rect 315974 116334 316080 116362
rect 316052 113174 316080 116334
rect 295444 113146 296208 113174
rect 316052 113146 316724 113174
rect 293866 107400 293922 107409
rect 293866 107335 293922 107344
rect 289818 106720 289874 106729
rect 289818 106655 289874 106664
rect 289832 97918 289860 106655
rect 293880 97918 293908 107335
rect 289820 97912 289872 97918
rect 289820 97854 289872 97860
rect 293868 97912 293920 97918
rect 293868 97854 293920 97860
rect 296180 97730 296208 113146
rect 296180 97702 296654 97730
rect 306300 95130 306328 97036
rect 315960 95198 315988 97036
rect 316696 95198 316724 113146
rect 317418 106720 317474 106729
rect 317418 106655 317474 106664
rect 317432 97986 317460 106655
rect 317420 97980 317472 97986
rect 317420 97922 317472 97928
rect 315948 95192 316000 95198
rect 315948 95134 316000 95140
rect 316684 95192 316736 95198
rect 316684 95134 316736 95140
rect 318076 95130 318104 118662
rect 267004 95124 267056 95130
rect 267004 95066 267056 95072
rect 278596 95124 278648 95130
rect 278596 95066 278648 95072
rect 289084 95124 289136 95130
rect 289084 95066 289136 95072
rect 306288 95124 306340 95130
rect 306288 95066 306340 95072
rect 318064 95124 318116 95130
rect 318064 95066 318116 95072
rect 250260 95056 250312 95062
rect 250260 94998 250312 95004
rect 261484 95056 261536 95062
rect 261484 94998 261536 95004
rect 249708 91248 249760 91254
rect 249708 91190 249760 91196
rect 260196 91248 260248 91254
rect 260196 91190 260248 91196
rect 277676 91248 277728 91254
rect 277676 91190 277728 91196
rect 287520 91248 287572 91254
rect 287520 91190 287572 91196
rect 305368 91248 305420 91254
rect 305368 91190 305420 91196
rect 315488 91248 315540 91254
rect 315488 91190 315540 91196
rect 249720 89964 249748 91190
rect 259368 91112 259420 91118
rect 259368 91054 259420 91060
rect 260104 91112 260156 91118
rect 260104 91054 260156 91060
rect 259380 89964 259408 91054
rect 238864 89270 240074 89298
rect 238666 80336 238722 80345
rect 238666 80271 238722 80280
rect 238680 71738 238708 80271
rect 238668 71732 238720 71738
rect 238668 71674 238720 71680
rect 238864 68882 238892 89270
rect 239772 72344 239824 72350
rect 239772 72286 239824 72292
rect 259736 72344 259788 72350
rect 259736 72286 259788 72292
rect 239784 70666 239812 72286
rect 259748 70666 259776 72286
rect 239784 70638 240074 70666
rect 259394 70638 259776 70666
rect 249720 68950 249748 70108
rect 260116 68950 260144 91054
rect 260208 72350 260236 91190
rect 268016 91180 268068 91186
rect 268016 91122 268068 91128
rect 268028 89964 268056 91122
rect 277688 89964 277716 91190
rect 287336 91112 287388 91118
rect 287336 91054 287388 91060
rect 287348 89964 287376 91054
rect 262220 88392 262272 88398
rect 262220 88334 262272 88340
rect 266268 88392 266320 88398
rect 266268 88334 266320 88340
rect 262232 79665 262260 88334
rect 266280 80345 266308 88334
rect 266266 80336 266322 80345
rect 266266 80271 266322 80280
rect 262218 79656 262274 79665
rect 262218 79591 262274 79600
rect 260196 72344 260248 72350
rect 260196 72286 260248 72292
rect 287532 70666 287560 91190
rect 287704 91180 287756 91186
rect 287704 91122 287756 91128
rect 296352 91180 296404 91186
rect 296352 91122 296404 91128
rect 287716 72146 287744 91122
rect 289084 91112 289136 91118
rect 289084 91054 289136 91060
rect 287704 72140 287756 72146
rect 287704 72082 287756 72088
rect 287362 70638 287560 70666
rect 249708 68944 249760 68950
rect 249708 68886 249760 68892
rect 260104 68944 260156 68950
rect 260104 68886 260156 68892
rect 268028 68882 268056 70108
rect 277688 69018 277716 70108
rect 289096 69018 289124 91054
rect 296364 89978 296392 91122
rect 296056 89950 296392 89978
rect 305380 89978 305408 91190
rect 315028 91112 315080 91118
rect 315028 91054 315080 91060
rect 315040 89978 315068 91054
rect 305380 89950 305716 89978
rect 315040 89950 315376 89978
rect 293866 80336 293922 80345
rect 293866 80271 293922 80280
rect 289818 79656 289874 79665
rect 289818 79591 289874 79600
rect 289832 71738 289860 79591
rect 293880 71738 293908 80271
rect 295708 72140 295760 72146
rect 295708 72082 295760 72088
rect 289820 71732 289872 71738
rect 289820 71674 289872 71680
rect 293868 71732 293920 71738
rect 293868 71674 293920 71680
rect 295720 70666 295748 72082
rect 315500 70666 315528 91190
rect 316776 91180 316828 91186
rect 316776 91122 316828 91128
rect 316684 91112 316736 91118
rect 316684 91054 316736 91060
rect 295720 70638 296056 70666
rect 315376 70638 315528 70666
rect 305716 70094 306052 70122
rect 306024 69018 306052 70094
rect 316696 69018 316724 91054
rect 316788 72350 316816 91122
rect 317420 88392 317472 88398
rect 317420 88334 317472 88340
rect 317432 79665 317460 88334
rect 317418 79656 317474 79665
rect 317418 79591 317474 79600
rect 316776 72344 316828 72350
rect 316776 72286 316828 72292
rect 277676 69012 277728 69018
rect 277676 68954 277728 68960
rect 289084 69012 289136 69018
rect 289084 68954 289136 68960
rect 306012 69012 306064 69018
rect 306012 68954 306064 68960
rect 316684 69012 316736 69018
rect 316684 68954 316736 68960
rect 238852 68876 238904 68882
rect 238852 68818 238904 68824
rect 268016 68876 268068 68882
rect 268016 68818 268068 68824
rect 261484 65068 261536 65074
rect 261484 65010 261536 65016
rect 268292 65068 268344 65074
rect 268292 65010 268344 65016
rect 295432 65068 295484 65074
rect 295432 65010 295484 65016
rect 240600 64932 240652 64938
rect 240600 64874 240652 64880
rect 250260 64932 250312 64938
rect 250260 64874 250312 64880
rect 240612 62900 240640 64874
rect 250272 62900 250300 64874
rect 259946 62206 260144 62234
rect 238666 53408 238722 53417
rect 238666 53343 238722 53352
rect 238680 44130 238708 53343
rect 238668 44124 238720 44130
rect 238668 44066 238720 44072
rect 240612 41342 240640 43044
rect 240600 41336 240652 41342
rect 240600 41278 240652 41284
rect 250272 41274 250300 43044
rect 259932 41410 259960 43044
rect 260116 41410 260144 62206
rect 259920 41404 259972 41410
rect 259920 41346 259972 41352
rect 260104 41404 260156 41410
rect 260104 41346 260156 41352
rect 261496 41274 261524 65010
rect 267832 65000 267884 65006
rect 267832 64942 267884 64948
rect 267004 64932 267056 64938
rect 267004 64874 267056 64880
rect 262220 62144 262272 62150
rect 262220 62086 262272 62092
rect 266268 62144 266320 62150
rect 266268 62086 266320 62092
rect 262232 52737 262260 62086
rect 266280 53417 266308 62086
rect 266266 53408 266322 53417
rect 266266 53343 266322 53352
rect 262218 52728 262274 52737
rect 262218 52663 262274 52672
rect 267016 41342 267044 64874
rect 267844 55214 267872 64942
rect 268304 62914 268332 65010
rect 277952 64932 278004 64938
rect 277952 64874 278004 64880
rect 289084 64932 289136 64938
rect 289084 64874 289136 64880
rect 277964 62914 277992 64874
rect 268304 62886 268640 62914
rect 277964 62886 278300 62914
rect 287960 62206 288112 62234
rect 267844 55186 268240 55214
rect 268212 43738 268240 55186
rect 268212 43710 268640 43738
rect 278300 43030 278636 43058
rect 278608 41342 278636 43030
rect 287624 43030 287960 43058
rect 287624 41410 287652 43030
rect 288084 41410 288112 62206
rect 287612 41404 287664 41410
rect 287612 41346 287664 41352
rect 288072 41404 288124 41410
rect 288072 41346 288124 41352
rect 289096 41342 289124 64874
rect 295444 55214 295472 65010
rect 306288 65000 306340 65006
rect 306288 64942 306340 64948
rect 296628 64932 296680 64938
rect 296628 64874 296680 64880
rect 296640 62900 296668 64874
rect 306300 62900 306328 64942
rect 318064 64932 318116 64938
rect 318064 64874 318116 64880
rect 315974 62206 316080 62234
rect 316052 55214 316080 62206
rect 317420 62144 317472 62150
rect 317420 62086 317472 62092
rect 295444 55186 296208 55214
rect 316052 55186 316724 55214
rect 293866 53408 293922 53417
rect 293866 53343 293922 53352
rect 289818 52728 289874 52737
rect 289818 52663 289874 52672
rect 289832 44130 289860 52663
rect 293880 44130 293908 53343
rect 289820 44124 289872 44130
rect 289820 44066 289872 44072
rect 293868 44124 293920 44130
rect 293868 44066 293920 44072
rect 296180 43738 296208 55186
rect 296180 43710 296654 43738
rect 306300 41342 306328 43044
rect 315960 41410 315988 43044
rect 316696 41410 316724 55186
rect 317432 52737 317460 62086
rect 317418 52728 317474 52737
rect 317418 52663 317474 52672
rect 315948 41404 316000 41410
rect 315948 41346 316000 41352
rect 316684 41404 316736 41410
rect 316684 41346 316736 41352
rect 318076 41342 318104 64874
rect 267004 41336 267056 41342
rect 267004 41278 267056 41284
rect 278596 41336 278648 41342
rect 278596 41278 278648 41284
rect 289084 41336 289136 41342
rect 289084 41278 289136 41284
rect 306288 41336 306340 41342
rect 306288 41278 306340 41284
rect 318064 41336 318116 41342
rect 318064 41278 318116 41284
rect 250260 41268 250312 41274
rect 250260 41210 250312 41216
rect 261484 41268 261536 41274
rect 261484 41210 261536 41216
rect 234620 39364 234672 39370
rect 234620 39306 234672 39312
rect 322216 38350 322244 700470
rect 364996 700398 365024 703520
rect 397472 700398 397500 703520
rect 364984 700392 365036 700398
rect 364984 700334 365036 700340
rect 378784 700392 378836 700398
rect 378784 700334 378836 700340
rect 397460 700392 397512 700398
rect 397460 700334 397512 700340
rect 345664 686044 345716 686050
rect 345664 685986 345716 685992
rect 361672 686044 361724 686050
rect 361672 685986 361724 685992
rect 371516 686044 371568 686050
rect 371516 685986 371568 685992
rect 333704 685976 333756 685982
rect 333704 685918 333756 685924
rect 333716 683876 333744 685918
rect 343364 685908 343416 685914
rect 343364 685850 343416 685856
rect 344284 685908 344336 685914
rect 344284 685850 344336 685856
rect 343376 683876 343404 685850
rect 323044 683318 324070 683346
rect 322846 674248 322902 674257
rect 322846 674183 322902 674192
rect 322860 665174 322888 674183
rect 322848 665168 322900 665174
rect 322848 665110 322900 665116
rect 323044 662250 323072 683318
rect 323676 665508 323728 665514
rect 323676 665450 323728 665456
rect 323688 664714 323716 665450
rect 343548 665100 343600 665106
rect 343548 665042 343600 665048
rect 343560 664714 343588 665042
rect 323688 664686 324070 664714
rect 343390 664686 343588 664714
rect 333730 664006 333928 664034
rect 333900 662318 333928 664006
rect 344296 662318 344324 685850
rect 345020 683188 345072 683194
rect 345020 683130 345072 683136
rect 345032 673577 345060 683130
rect 345018 673568 345074 673577
rect 345018 673503 345074 673512
rect 345676 665106 345704 685986
rect 352012 685976 352064 685982
rect 352012 685918 352064 685924
rect 352024 683876 352052 685918
rect 361684 683876 361712 685986
rect 371332 685908 371384 685914
rect 371332 685850 371384 685856
rect 371344 683876 371372 685850
rect 350448 683256 350500 683262
rect 350448 683198 350500 683204
rect 350460 674257 350488 683198
rect 350446 674248 350502 674257
rect 350446 674183 350502 674192
rect 345664 665100 345716 665106
rect 345664 665042 345716 665048
rect 371528 664714 371556 685986
rect 374644 685976 374696 685982
rect 374644 685918 374696 685924
rect 373264 685908 373316 685914
rect 373264 685850 373316 685856
rect 371358 664686 371556 664714
rect 333888 662312 333940 662318
rect 333888 662254 333940 662260
rect 344284 662312 344336 662318
rect 344284 662254 344336 662260
rect 352024 662250 352052 664020
rect 361684 662386 361712 664020
rect 373276 662386 373304 685850
rect 373998 673568 374054 673577
rect 373998 673503 374054 673512
rect 374012 665174 374040 673503
rect 374000 665168 374052 665174
rect 374000 665110 374052 665116
rect 361672 662380 361724 662386
rect 361672 662322 361724 662328
rect 373264 662380 373316 662386
rect 373264 662322 373316 662328
rect 374656 662318 374684 685918
rect 378048 683188 378100 683194
rect 378048 683130 378100 683136
rect 378060 674257 378088 683130
rect 378046 674248 378102 674257
rect 378046 674183 378102 674192
rect 374644 662312 374696 662318
rect 374644 662254 374696 662260
rect 323032 662244 323084 662250
rect 323032 662186 323084 662192
rect 352012 662244 352064 662250
rect 352012 662186 352064 662192
rect 334256 658436 334308 658442
rect 334256 658378 334308 658384
rect 352012 658436 352064 658442
rect 352012 658378 352064 658384
rect 324596 658300 324648 658306
rect 324596 658242 324648 658248
rect 324608 656948 324636 658242
rect 334268 656948 334296 658378
rect 347044 658368 347096 658374
rect 347044 658310 347096 658316
rect 343942 656254 344140 656282
rect 322848 655580 322900 655586
rect 322848 655522 322900 655528
rect 322860 647465 322888 655522
rect 322846 647456 322902 647465
rect 322846 647391 322902 647400
rect 324608 634710 324636 637092
rect 324596 634704 324648 634710
rect 324596 634646 324648 634652
rect 334268 634642 334296 637092
rect 343928 634778 343956 637092
rect 344112 634778 344140 656254
rect 345020 655648 345072 655654
rect 345020 655590 345072 655596
rect 345032 646785 345060 655590
rect 345018 646776 345074 646785
rect 345018 646711 345074 646720
rect 343916 634772 343968 634778
rect 343916 634714 343968 634720
rect 344100 634772 344152 634778
rect 344100 634714 344152 634720
rect 347056 634710 347084 658310
rect 348424 658300 348476 658306
rect 348424 658242 348476 658248
rect 347044 634704 347096 634710
rect 347044 634646 347096 634652
rect 348436 634642 348464 658242
rect 350448 655716 350500 655722
rect 350448 655658 350500 655664
rect 350460 647465 350488 655658
rect 352024 654134 352052 658378
rect 361948 658368 362000 658374
rect 361948 658310 362000 658316
rect 352288 658300 352340 658306
rect 352288 658242 352340 658248
rect 352300 656962 352328 658242
rect 361960 656962 361988 658310
rect 373264 658300 373316 658306
rect 373264 658242 373316 658248
rect 352300 656934 352636 656962
rect 361960 656934 362296 656962
rect 371956 656254 372108 656282
rect 352024 654106 352236 654134
rect 350446 647456 350502 647465
rect 350446 647391 350502 647400
rect 352208 637786 352236 654106
rect 352208 637758 352636 637786
rect 362296 637078 362632 637106
rect 362604 634710 362632 637078
rect 371620 637078 371956 637106
rect 371620 634778 371648 637078
rect 372080 634778 372108 656254
rect 371608 634772 371660 634778
rect 371608 634714 371660 634720
rect 372068 634772 372120 634778
rect 372068 634714 372120 634720
rect 373276 634710 373304 658242
rect 378048 655648 378100 655654
rect 378048 655590 378100 655596
rect 374000 655580 374052 655586
rect 374000 655522 374052 655528
rect 374012 646785 374040 655522
rect 378060 647465 378088 655590
rect 378046 647456 378102 647465
rect 378046 647391 378102 647400
rect 373998 646776 374054 646785
rect 373998 646711 374054 646720
rect 362592 634704 362644 634710
rect 362592 634646 362644 634652
rect 373264 634704 373316 634710
rect 373264 634646 373316 634652
rect 334256 634636 334308 634642
rect 334256 634578 334308 634584
rect 348424 634636 348476 634642
rect 348424 634578 348476 634584
rect 345664 632256 345716 632262
rect 345664 632198 345716 632204
rect 361672 632256 361724 632262
rect 361672 632198 361724 632204
rect 371516 632256 371568 632262
rect 371516 632198 371568 632204
rect 333704 632188 333756 632194
rect 333704 632130 333756 632136
rect 333716 629884 333744 632130
rect 343364 632120 343416 632126
rect 343364 632062 343416 632068
rect 344284 632120 344336 632126
rect 344284 632062 344336 632068
rect 343376 629884 343404 632062
rect 323044 629326 324070 629354
rect 322846 620256 322902 620265
rect 322846 620191 322902 620200
rect 322860 611318 322888 620191
rect 322848 611312 322900 611318
rect 322848 611254 322900 611260
rect 323044 608462 323072 629326
rect 323676 611924 323728 611930
rect 323676 611866 323728 611872
rect 323688 610722 323716 611866
rect 323688 610694 324070 610722
rect 333716 608530 333744 610028
rect 343376 608598 343404 610028
rect 343364 608592 343416 608598
rect 343364 608534 343416 608540
rect 344296 608530 344324 632062
rect 345018 619576 345074 619585
rect 345018 619511 345074 619520
rect 345032 611250 345060 619511
rect 345020 611244 345072 611250
rect 345020 611186 345072 611192
rect 345676 608598 345704 632198
rect 352012 632188 352064 632194
rect 352012 632130 352064 632136
rect 352024 629884 352052 632130
rect 361684 629884 361712 632198
rect 371332 632120 371384 632126
rect 371332 632062 371384 632068
rect 371344 629884 371372 632062
rect 350446 620256 350502 620265
rect 350446 620191 350502 620200
rect 350460 611182 350488 620191
rect 350448 611176 350500 611182
rect 350448 611118 350500 611124
rect 371528 610722 371556 632198
rect 374644 632188 374696 632194
rect 374644 632130 374696 632136
rect 373264 632120 373316 632126
rect 373264 632062 373316 632068
rect 371358 610694 371556 610722
rect 345664 608592 345716 608598
rect 345664 608534 345716 608540
rect 333704 608524 333756 608530
rect 333704 608466 333756 608472
rect 344284 608524 344336 608530
rect 344284 608466 344336 608472
rect 352024 608462 352052 610028
rect 361684 608598 361712 610028
rect 373276 608598 373304 632062
rect 373998 619576 374054 619585
rect 373998 619511 374054 619520
rect 374012 611318 374040 619511
rect 374000 611312 374052 611318
rect 374000 611254 374052 611260
rect 361672 608592 361724 608598
rect 361672 608534 361724 608540
rect 373264 608592 373316 608598
rect 373264 608534 373316 608540
rect 374656 608530 374684 632130
rect 378046 620256 378102 620265
rect 378046 620191 378102 620200
rect 378060 611250 378088 620191
rect 378048 611244 378100 611250
rect 378048 611186 378100 611192
rect 374644 608524 374696 608530
rect 374644 608466 374696 608472
rect 323032 608456 323084 608462
rect 323032 608398 323084 608404
rect 352012 608456 352064 608462
rect 352012 608398 352064 608404
rect 334256 604648 334308 604654
rect 334256 604590 334308 604596
rect 352012 604648 352064 604654
rect 352012 604590 352064 604596
rect 324596 604512 324648 604518
rect 324596 604454 324648 604460
rect 324608 602956 324636 604454
rect 334268 602956 334296 604590
rect 347044 604580 347096 604586
rect 347044 604522 347096 604528
rect 343942 602262 344140 602290
rect 322848 601724 322900 601730
rect 322848 601666 322900 601672
rect 322860 593473 322888 601666
rect 322846 593464 322902 593473
rect 322846 593399 322902 593408
rect 324608 580922 324636 583100
rect 324596 580916 324648 580922
rect 324596 580858 324648 580864
rect 334268 580854 334296 583100
rect 343928 580990 343956 583100
rect 344112 580990 344140 602262
rect 345020 601792 345072 601798
rect 345020 601734 345072 601740
rect 345032 592793 345060 601734
rect 345018 592784 345074 592793
rect 345018 592719 345074 592728
rect 343916 580984 343968 580990
rect 343916 580926 343968 580932
rect 344100 580984 344152 580990
rect 344100 580926 344152 580932
rect 347056 580922 347084 604522
rect 348424 604512 348476 604518
rect 348424 604454 348476 604460
rect 347044 580916 347096 580922
rect 347044 580858 347096 580864
rect 348436 580854 348464 604454
rect 350448 601860 350500 601866
rect 350448 601802 350500 601808
rect 350460 593473 350488 601802
rect 352024 596174 352052 604590
rect 361948 604580 362000 604586
rect 361948 604522 362000 604528
rect 352288 604512 352340 604518
rect 352288 604454 352340 604460
rect 352300 602970 352328 604454
rect 361960 602970 361988 604522
rect 373264 604512 373316 604518
rect 373264 604454 373316 604460
rect 352300 602942 352636 602970
rect 361960 602942 362296 602970
rect 371956 602262 372108 602290
rect 352024 596146 352236 596174
rect 350446 593464 350502 593473
rect 350446 593399 350502 593408
rect 352208 583794 352236 596146
rect 352208 583766 352636 583794
rect 362296 583086 362632 583114
rect 362604 580922 362632 583086
rect 371620 583086 371956 583114
rect 371620 580990 371648 583086
rect 372080 580990 372108 602262
rect 371608 580984 371660 580990
rect 371608 580926 371660 580932
rect 372068 580984 372120 580990
rect 372068 580926 372120 580932
rect 373276 580922 373304 604454
rect 378048 601792 378100 601798
rect 378048 601734 378100 601740
rect 374000 601724 374052 601730
rect 374000 601666 374052 601672
rect 374012 592793 374040 601666
rect 378060 593473 378088 601734
rect 378046 593464 378102 593473
rect 378046 593399 378102 593408
rect 373998 592784 374054 592793
rect 373998 592719 374054 592728
rect 362592 580916 362644 580922
rect 362592 580858 362644 580864
rect 373264 580916 373316 580922
rect 373264 580858 373316 580864
rect 334256 580848 334308 580854
rect 334256 580790 334308 580796
rect 348424 580848 348476 580854
rect 348424 580790 348476 580796
rect 345664 578400 345716 578406
rect 345664 578342 345716 578348
rect 361672 578400 361724 578406
rect 361672 578342 361724 578348
rect 371516 578400 371568 578406
rect 371516 578342 371568 578348
rect 333704 578332 333756 578338
rect 333704 578274 333756 578280
rect 333716 575892 333744 578274
rect 343364 578264 343416 578270
rect 343364 578206 343416 578212
rect 344284 578264 344336 578270
rect 344284 578206 344336 578212
rect 343376 575892 343404 578206
rect 323044 575334 324070 575362
rect 322846 566264 322902 566273
rect 322846 566199 322902 566208
rect 322860 557530 322888 566199
rect 322848 557524 322900 557530
rect 322848 557466 322900 557472
rect 323044 554606 323072 575334
rect 323676 558884 323728 558890
rect 323676 558826 323728 558832
rect 323688 556730 323716 558826
rect 343548 557456 343600 557462
rect 343548 557398 343600 557404
rect 343560 556730 343588 557398
rect 323688 556702 324070 556730
rect 343390 556702 343588 556730
rect 333716 554674 333744 556036
rect 344296 554674 344324 578206
rect 345018 565584 345074 565593
rect 345018 565519 345074 565528
rect 345032 557394 345060 565519
rect 345676 557462 345704 578342
rect 352012 578332 352064 578338
rect 352012 578274 352064 578280
rect 352024 575892 352052 578274
rect 361684 575892 361712 578342
rect 371332 578264 371384 578270
rect 371332 578206 371384 578212
rect 371344 575892 371372 578206
rect 350446 566264 350502 566273
rect 350446 566199 350502 566208
rect 345664 557456 345716 557462
rect 345664 557398 345716 557404
rect 350460 557394 350488 566199
rect 345020 557388 345072 557394
rect 345020 557330 345072 557336
rect 350448 557388 350500 557394
rect 350448 557330 350500 557336
rect 371528 556730 371556 578342
rect 374644 578332 374696 578338
rect 374644 578274 374696 578280
rect 373264 578264 373316 578270
rect 373264 578206 373316 578212
rect 371358 556702 371556 556730
rect 333704 554668 333756 554674
rect 333704 554610 333756 554616
rect 344284 554668 344336 554674
rect 344284 554610 344336 554616
rect 352024 554606 352052 556036
rect 361684 554742 361712 556036
rect 373276 554742 373304 578206
rect 373998 565584 374054 565593
rect 373998 565519 374054 565528
rect 374012 557530 374040 565519
rect 374000 557524 374052 557530
rect 374000 557466 374052 557472
rect 374656 554742 374684 578274
rect 378046 566264 378102 566273
rect 378046 566199 378102 566208
rect 378060 557462 378088 566199
rect 378048 557456 378100 557462
rect 378048 557398 378100 557404
rect 361672 554736 361724 554742
rect 361672 554678 361724 554684
rect 373264 554736 373316 554742
rect 373264 554678 373316 554684
rect 374644 554736 374696 554742
rect 374644 554678 374696 554684
rect 323032 554600 323084 554606
rect 323032 554542 323084 554548
rect 352012 554600 352064 554606
rect 352012 554542 352064 554548
rect 352012 550860 352064 550866
rect 352012 550802 352064 550808
rect 334256 550792 334308 550798
rect 334256 550734 334308 550740
rect 345664 550792 345716 550798
rect 345664 550734 345716 550740
rect 324596 550656 324648 550662
rect 324596 550598 324648 550604
rect 324608 548964 324636 550598
rect 334268 548964 334296 550734
rect 343942 548270 344140 548298
rect 322846 539472 322902 539481
rect 322846 539407 322902 539416
rect 322860 529922 322888 539407
rect 322848 529916 322900 529922
rect 322848 529858 322900 529864
rect 324608 527066 324636 529108
rect 324596 527060 324648 527066
rect 324596 527002 324648 527008
rect 334268 526998 334296 529108
rect 343928 527134 343956 529108
rect 344112 527134 344140 548270
rect 345018 538792 345074 538801
rect 345018 538727 345074 538736
rect 345032 529854 345060 538727
rect 345020 529848 345072 529854
rect 345020 529790 345072 529796
rect 343916 527128 343968 527134
rect 343916 527070 343968 527076
rect 344100 527128 344152 527134
rect 344100 527070 344152 527076
rect 345676 527066 345704 550734
rect 347044 550656 347096 550662
rect 347044 550598 347096 550604
rect 345664 527060 345716 527066
rect 345664 527002 345716 527008
rect 347056 526998 347084 550598
rect 350446 539472 350502 539481
rect 350446 539407 350502 539416
rect 350460 529786 350488 539407
rect 352024 538214 352052 550802
rect 352288 550656 352340 550662
rect 352288 550598 352340 550604
rect 361948 550656 362000 550662
rect 361948 550598 362000 550604
rect 373264 550656 373316 550662
rect 373264 550598 373316 550604
rect 352300 548978 352328 550598
rect 361960 548978 361988 550598
rect 352300 548950 352636 548978
rect 361960 548950 362296 548978
rect 371956 548270 372108 548298
rect 352024 538186 352236 538214
rect 350448 529780 350500 529786
rect 350448 529722 350500 529728
rect 352208 529666 352236 538186
rect 352208 529638 352636 529666
rect 362296 529094 362632 529122
rect 362604 527066 362632 529094
rect 371620 529094 371956 529122
rect 371620 527134 371648 529094
rect 372080 527134 372108 548270
rect 371608 527128 371660 527134
rect 371608 527070 371660 527076
rect 372068 527128 372120 527134
rect 372068 527070 372120 527076
rect 373276 527066 373304 550598
rect 378046 539472 378102 539481
rect 378046 539407 378102 539416
rect 373998 538792 374054 538801
rect 373998 538727 374054 538736
rect 374012 529922 374040 538727
rect 374000 529916 374052 529922
rect 374000 529858 374052 529864
rect 378060 529854 378088 539407
rect 378048 529848 378100 529854
rect 378048 529790 378100 529796
rect 362592 527060 362644 527066
rect 362592 527002 362644 527008
rect 373264 527060 373316 527066
rect 373264 527002 373316 527008
rect 334256 526992 334308 526998
rect 334256 526934 334308 526940
rect 347044 526992 347096 526998
rect 347044 526934 347096 526940
rect 345664 523184 345716 523190
rect 345664 523126 345716 523132
rect 361672 523184 361724 523190
rect 361672 523126 361724 523132
rect 371516 523184 371568 523190
rect 371516 523126 371568 523132
rect 333704 523116 333756 523122
rect 333704 523058 333756 523064
rect 333716 521900 333744 523058
rect 343364 523048 343416 523054
rect 343364 522990 343416 522996
rect 344284 523048 344336 523054
rect 344284 522990 344336 522996
rect 343376 521900 343404 522990
rect 323044 521206 324070 521234
rect 322848 520328 322900 520334
rect 322848 520270 322900 520276
rect 322860 512281 322888 520270
rect 322846 512272 322902 512281
rect 322846 512207 322902 512216
rect 323044 500818 323072 521206
rect 323676 503804 323728 503810
rect 323676 503746 323728 503752
rect 323688 502738 323716 503746
rect 323688 502710 324070 502738
rect 333716 500886 333744 502044
rect 343376 500954 343404 502044
rect 343364 500948 343416 500954
rect 343364 500890 343416 500896
rect 344296 500886 344324 522990
rect 345018 511592 345074 511601
rect 345018 511527 345074 511536
rect 345032 503674 345060 511527
rect 345020 503668 345072 503674
rect 345020 503610 345072 503616
rect 345676 500954 345704 523126
rect 352012 523116 352064 523122
rect 352012 523058 352064 523064
rect 352024 521900 352052 523058
rect 361684 521900 361712 523126
rect 371332 523048 371384 523054
rect 371332 522990 371384 522996
rect 371344 521900 371372 522990
rect 350446 512272 350502 512281
rect 350446 512207 350502 512216
rect 350460 503674 350488 512207
rect 350448 503668 350500 503674
rect 350448 503610 350500 503616
rect 371528 502738 371556 523126
rect 374644 523116 374696 523122
rect 374644 523058 374696 523064
rect 373264 523048 373316 523054
rect 373264 522990 373316 522996
rect 371358 502710 371556 502738
rect 345664 500948 345716 500954
rect 345664 500890 345716 500896
rect 333704 500880 333756 500886
rect 333704 500822 333756 500828
rect 344284 500880 344336 500886
rect 344284 500822 344336 500828
rect 352024 500818 352052 502044
rect 361684 500954 361712 502044
rect 373276 500954 373304 522990
rect 374000 520328 374052 520334
rect 374000 520270 374052 520276
rect 374012 511601 374040 520270
rect 373998 511592 374054 511601
rect 373998 511527 374054 511536
rect 361672 500948 361724 500954
rect 361672 500890 361724 500896
rect 373264 500948 373316 500954
rect 373264 500890 373316 500896
rect 374656 500886 374684 523058
rect 378048 520328 378100 520334
rect 378048 520270 378100 520276
rect 378060 512281 378088 520270
rect 378046 512272 378102 512281
rect 378046 512207 378102 512216
rect 374644 500880 374696 500886
rect 374644 500822 374696 500828
rect 323032 500812 323084 500818
rect 323032 500754 323084 500760
rect 352012 500812 352064 500818
rect 352012 500754 352064 500760
rect 334256 497004 334308 497010
rect 334256 496946 334308 496952
rect 352196 497004 352248 497010
rect 352196 496946 352248 496952
rect 324596 496868 324648 496874
rect 324596 496810 324648 496816
rect 324608 494972 324636 496810
rect 334268 494972 334296 496946
rect 345664 496936 345716 496942
rect 345664 496878 345716 496884
rect 343942 494278 344140 494306
rect 322846 485480 322902 485489
rect 322846 485415 322902 485424
rect 322860 476066 322888 485415
rect 322848 476060 322900 476066
rect 322848 476002 322900 476008
rect 324608 473278 324636 475116
rect 324596 473272 324648 473278
rect 324596 473214 324648 473220
rect 334268 473210 334296 475116
rect 343928 473346 343956 475116
rect 344112 473346 344140 494278
rect 345018 484800 345074 484809
rect 345018 484735 345074 484744
rect 345032 475998 345060 484735
rect 345020 475992 345072 475998
rect 345020 475934 345072 475940
rect 343916 473340 343968 473346
rect 343916 473282 343968 473288
rect 344100 473340 344152 473346
rect 344100 473282 344152 473288
rect 345676 473278 345704 496878
rect 347044 496868 347096 496874
rect 347044 496810 347096 496816
rect 345664 473272 345716 473278
rect 345664 473214 345716 473220
rect 347056 473210 347084 496810
rect 350446 485480 350502 485489
rect 350446 485415 350502 485424
rect 350460 475930 350488 485415
rect 350448 475924 350500 475930
rect 350448 475866 350500 475872
rect 352208 475674 352236 496946
rect 361948 496936 362000 496942
rect 361948 496878 362000 496884
rect 352288 496868 352340 496874
rect 352288 496810 352340 496816
rect 352300 494986 352328 496810
rect 361960 494986 361988 496878
rect 373264 496868 373316 496874
rect 373264 496810 373316 496816
rect 352300 494958 352636 494986
rect 361960 494958 362296 494986
rect 371956 494278 372108 494306
rect 352208 475646 352636 475674
rect 362296 475102 362632 475130
rect 362604 473278 362632 475102
rect 371620 475102 371956 475130
rect 371620 473346 371648 475102
rect 372080 473346 372108 494278
rect 371608 473340 371660 473346
rect 371608 473282 371660 473288
rect 372068 473340 372120 473346
rect 372068 473282 372120 473288
rect 373276 473278 373304 496810
rect 378046 485480 378102 485489
rect 378046 485415 378102 485424
rect 373998 484800 374054 484809
rect 373998 484735 374054 484744
rect 374012 476066 374040 484735
rect 374000 476060 374052 476066
rect 374000 476002 374052 476008
rect 378060 475998 378088 485415
rect 378048 475992 378100 475998
rect 378048 475934 378100 475940
rect 362592 473272 362644 473278
rect 362592 473214 362644 473220
rect 373264 473272 373316 473278
rect 373264 473214 373316 473220
rect 334256 473204 334308 473210
rect 334256 473146 334308 473152
rect 347044 473204 347096 473210
rect 347044 473146 347096 473152
rect 345664 469396 345716 469402
rect 345664 469338 345716 469344
rect 361672 469396 361724 469402
rect 361672 469338 361724 469344
rect 371516 469396 371568 469402
rect 371516 469338 371568 469344
rect 333704 469328 333756 469334
rect 333704 469270 333756 469276
rect 333716 467908 333744 469270
rect 343364 469260 343416 469266
rect 343364 469202 343416 469208
rect 344284 469260 344336 469266
rect 344284 469202 344336 469208
rect 343376 467908 343404 469202
rect 323044 467214 324070 467242
rect 322848 466472 322900 466478
rect 322848 466414 322900 466420
rect 322860 458289 322888 466414
rect 322846 458280 322902 458289
rect 322846 458215 322902 458224
rect 323044 445602 323072 467214
rect 323676 449948 323728 449954
rect 323676 449890 323728 449896
rect 323688 448746 323716 449890
rect 323688 448718 324070 448746
rect 343640 448520 343692 448526
rect 343390 448468 343640 448474
rect 343390 448462 343692 448468
rect 343390 448446 343680 448462
rect 333716 445670 333744 448052
rect 344296 445670 344324 469202
rect 345020 466540 345072 466546
rect 345020 466482 345072 466488
rect 345032 457609 345060 466482
rect 345018 457600 345074 457609
rect 345018 457535 345074 457544
rect 345676 448526 345704 469338
rect 352012 469328 352064 469334
rect 352012 469270 352064 469276
rect 352024 467908 352052 469270
rect 361684 467908 361712 469338
rect 371332 469260 371384 469266
rect 371332 469202 371384 469208
rect 371344 467908 371372 469202
rect 350448 466608 350500 466614
rect 350448 466550 350500 466556
rect 350460 458289 350488 466550
rect 350446 458280 350502 458289
rect 350446 458215 350502 458224
rect 371528 448746 371556 469338
rect 374644 469328 374696 469334
rect 374644 469270 374696 469276
rect 373264 469260 373316 469266
rect 373264 469202 373316 469208
rect 371358 448718 371556 448746
rect 345664 448520 345716 448526
rect 345664 448462 345716 448468
rect 333704 445664 333756 445670
rect 333704 445606 333756 445612
rect 344284 445664 344336 445670
rect 344284 445606 344336 445612
rect 352024 445602 352052 448052
rect 361684 445738 361712 448052
rect 373276 445738 373304 469202
rect 374000 466472 374052 466478
rect 374000 466414 374052 466420
rect 374012 457609 374040 466414
rect 373998 457600 374054 457609
rect 373998 457535 374054 457544
rect 361672 445732 361724 445738
rect 361672 445674 361724 445680
rect 373264 445732 373316 445738
rect 373264 445674 373316 445680
rect 374656 445670 374684 469270
rect 378048 466540 378100 466546
rect 378048 466482 378100 466488
rect 378060 458289 378088 466482
rect 378046 458280 378102 458289
rect 378046 458215 378102 458224
rect 374644 445664 374696 445670
rect 374644 445606 374696 445612
rect 323032 445596 323084 445602
rect 323032 445538 323084 445544
rect 352012 445596 352064 445602
rect 352012 445538 352064 445544
rect 334256 443148 334308 443154
rect 334256 443090 334308 443096
rect 352012 443148 352064 443154
rect 352012 443090 352064 443096
rect 324596 443012 324648 443018
rect 324596 442954 324648 442960
rect 324608 440980 324636 442954
rect 334268 440980 334296 443090
rect 345664 443080 345716 443086
rect 345664 443022 345716 443028
rect 322848 440292 322900 440298
rect 343942 440286 344140 440314
rect 322848 440234 322900 440240
rect 322860 431497 322888 440234
rect 322846 431488 322902 431497
rect 322846 431423 322902 431432
rect 324608 419422 324636 421124
rect 324596 419416 324648 419422
rect 324596 419358 324648 419364
rect 334268 419354 334296 421124
rect 343928 419490 343956 421124
rect 344112 419490 344140 440286
rect 345018 430808 345074 430817
rect 345018 430743 345074 430752
rect 345032 422278 345060 430743
rect 345020 422272 345072 422278
rect 345020 422214 345072 422220
rect 343916 419484 343968 419490
rect 343916 419426 343968 419432
rect 344100 419484 344152 419490
rect 344100 419426 344152 419432
rect 345676 419422 345704 443022
rect 347044 443012 347096 443018
rect 347044 442954 347096 442960
rect 345664 419416 345716 419422
rect 345664 419358 345716 419364
rect 347056 419354 347084 442954
rect 352024 441614 352052 443090
rect 361948 443080 362000 443086
rect 361948 443022 362000 443028
rect 352288 443012 352340 443018
rect 352288 442954 352340 442960
rect 352024 441586 352236 441614
rect 350446 431488 350502 431497
rect 350446 431423 350502 431432
rect 350460 422278 350488 431423
rect 350448 422272 350500 422278
rect 350448 422214 350500 422220
rect 352208 421682 352236 441586
rect 352300 440994 352328 442954
rect 361960 440994 361988 443022
rect 373264 443012 373316 443018
rect 373264 442954 373316 442960
rect 352300 440966 352636 440994
rect 361960 440966 362296 440994
rect 371956 440286 372108 440314
rect 352208 421654 352636 421682
rect 362296 421110 362632 421138
rect 362604 419422 362632 421110
rect 371620 421110 371956 421138
rect 371620 419490 371648 421110
rect 372080 419490 372108 440286
rect 371608 419484 371660 419490
rect 371608 419426 371660 419432
rect 372068 419484 372120 419490
rect 372068 419426 372120 419432
rect 373276 419422 373304 442954
rect 374000 440292 374052 440298
rect 374000 440234 374052 440240
rect 378048 440292 378100 440298
rect 378048 440234 378100 440240
rect 374012 430817 374040 440234
rect 378060 431497 378088 440234
rect 378046 431488 378102 431497
rect 378046 431423 378102 431432
rect 373998 430808 374054 430817
rect 373998 430743 374054 430752
rect 362592 419416 362644 419422
rect 362592 419358 362644 419364
rect 373264 419416 373316 419422
rect 373264 419358 373316 419364
rect 334256 419348 334308 419354
rect 334256 419290 334308 419296
rect 347044 419348 347096 419354
rect 347044 419290 347096 419296
rect 345664 415608 345716 415614
rect 345664 415550 345716 415556
rect 361672 415608 361724 415614
rect 361672 415550 361724 415556
rect 371516 415608 371568 415614
rect 371516 415550 371568 415556
rect 333704 415540 333756 415546
rect 333704 415482 333756 415488
rect 333716 413916 333744 415482
rect 343364 415472 343416 415478
rect 343364 415414 343416 415420
rect 344284 415472 344336 415478
rect 344284 415414 344336 415420
rect 343376 413916 343404 415414
rect 323044 413222 324070 413250
rect 322846 404288 322902 404297
rect 322846 404223 322902 404232
rect 322860 394670 322888 404223
rect 322848 394664 322900 394670
rect 322848 394606 322900 394612
rect 323044 391814 323072 413222
rect 323676 395140 323728 395146
rect 323676 395082 323728 395088
rect 323688 394754 323716 395082
rect 323688 394726 324070 394754
rect 343390 394602 343680 394618
rect 343390 394596 343692 394602
rect 343390 394590 343640 394596
rect 343640 394538 343692 394544
rect 333716 391882 333744 394060
rect 344296 391882 344324 415414
rect 345018 403608 345074 403617
rect 345018 403543 345074 403552
rect 345032 394534 345060 403543
rect 345676 394602 345704 415550
rect 352012 415540 352064 415546
rect 352012 415482 352064 415488
rect 352024 413916 352052 415482
rect 361684 413916 361712 415550
rect 371332 415472 371384 415478
rect 371332 415414 371384 415420
rect 371344 413916 371372 415414
rect 350446 404288 350502 404297
rect 350446 404223 350502 404232
rect 345664 394596 345716 394602
rect 345664 394538 345716 394544
rect 350460 394534 350488 404223
rect 371528 394754 371556 415550
rect 374644 415540 374696 415546
rect 374644 415482 374696 415488
rect 373264 415472 373316 415478
rect 373264 415414 373316 415420
rect 371358 394726 371556 394754
rect 345020 394528 345072 394534
rect 345020 394470 345072 394476
rect 350448 394528 350500 394534
rect 350448 394470 350500 394476
rect 333704 391876 333756 391882
rect 333704 391818 333756 391824
rect 344284 391876 344336 391882
rect 344284 391818 344336 391824
rect 352024 391814 352052 394060
rect 361684 391950 361712 394060
rect 373276 391950 373304 415414
rect 373998 403608 374054 403617
rect 373998 403543 374054 403552
rect 374012 394670 374040 403543
rect 374000 394664 374052 394670
rect 374000 394606 374052 394612
rect 361672 391944 361724 391950
rect 361672 391886 361724 391892
rect 373264 391944 373316 391950
rect 373264 391886 373316 391892
rect 374656 391882 374684 415482
rect 378046 404288 378102 404297
rect 378046 404223 378102 404232
rect 378060 394602 378088 404223
rect 378048 394596 378100 394602
rect 378048 394538 378100 394544
rect 374644 391876 374696 391882
rect 374644 391818 374696 391824
rect 323032 391808 323084 391814
rect 323032 391750 323084 391756
rect 352012 391808 352064 391814
rect 352012 391750 352064 391756
rect 334256 389360 334308 389366
rect 334256 389302 334308 389308
rect 352012 389360 352064 389366
rect 352012 389302 352064 389308
rect 324596 389224 324648 389230
rect 324596 389166 324648 389172
rect 324608 386852 324636 389166
rect 334268 386852 334296 389302
rect 345664 389292 345716 389298
rect 345664 389234 345716 389240
rect 345020 386504 345072 386510
rect 345020 386446 345072 386452
rect 322848 386436 322900 386442
rect 322848 386378 322900 386384
rect 322860 377505 322888 386378
rect 343942 386294 344140 386322
rect 322846 377496 322902 377505
rect 322846 377431 322902 377440
rect 324608 365634 324636 367132
rect 324596 365628 324648 365634
rect 324596 365570 324648 365576
rect 334268 365566 334296 367132
rect 343928 365702 343956 367132
rect 344112 365702 344140 386294
rect 345032 376825 345060 386446
rect 345018 376816 345074 376825
rect 345018 376751 345074 376760
rect 343916 365696 343968 365702
rect 343916 365638 343968 365644
rect 344100 365696 344152 365702
rect 344100 365638 344152 365644
rect 345676 365634 345704 389234
rect 347044 389224 347096 389230
rect 347044 389166 347096 389172
rect 345664 365628 345716 365634
rect 345664 365570 345716 365576
rect 347056 365566 347084 389166
rect 350448 386572 350500 386578
rect 350448 386514 350500 386520
rect 350460 377505 350488 386514
rect 352024 383654 352052 389302
rect 361948 389292 362000 389298
rect 361948 389234 362000 389240
rect 352288 389224 352340 389230
rect 352288 389166 352340 389172
rect 352300 386866 352328 389166
rect 361960 386866 361988 389234
rect 373264 389224 373316 389230
rect 373264 389166 373316 389172
rect 352300 386838 352636 386866
rect 361960 386838 362296 386866
rect 371956 386294 372108 386322
rect 352024 383626 352236 383654
rect 350446 377496 350502 377505
rect 350446 377431 350502 377440
rect 352208 367690 352236 383626
rect 352208 367662 352636 367690
rect 362296 367118 362632 367146
rect 362604 365634 362632 367118
rect 371620 367118 371956 367146
rect 371620 365702 371648 367118
rect 372080 365702 372108 386294
rect 371608 365696 371660 365702
rect 371608 365638 371660 365644
rect 372068 365696 372120 365702
rect 372068 365638 372120 365644
rect 373276 365634 373304 389166
rect 378048 386504 378100 386510
rect 378048 386446 378100 386452
rect 374000 386436 374052 386442
rect 374000 386378 374052 386384
rect 374012 377369 374040 386378
rect 378060 377505 378088 386446
rect 378046 377496 378102 377505
rect 378046 377431 378102 377440
rect 373998 377360 374054 377369
rect 373998 377295 374054 377304
rect 362592 365628 362644 365634
rect 362592 365570 362644 365576
rect 373264 365628 373316 365634
rect 373264 365570 373316 365576
rect 334256 365560 334308 365566
rect 334256 365502 334308 365508
rect 347044 365560 347096 365566
rect 347044 365502 347096 365508
rect 345664 361752 345716 361758
rect 345664 361694 345716 361700
rect 361672 361752 361724 361758
rect 361672 361694 361724 361700
rect 371516 361752 371568 361758
rect 371516 361694 371568 361700
rect 333704 361684 333756 361690
rect 333704 361626 333756 361632
rect 333716 359924 333744 361626
rect 343364 361616 343416 361622
rect 343364 361558 343416 361564
rect 344284 361616 344336 361622
rect 344284 361558 344336 361564
rect 343376 359924 343404 361558
rect 323044 359230 324070 359258
rect 322846 350296 322902 350305
rect 322846 350231 322902 350240
rect 322860 340882 322888 350231
rect 322848 340876 322900 340882
rect 322848 340818 322900 340824
rect 323044 337958 323072 359230
rect 323676 341284 323728 341290
rect 323676 341226 323728 341232
rect 323688 340762 323716 341226
rect 323688 340734 324070 340762
rect 343390 340746 343680 340762
rect 343390 340740 343692 340746
rect 343390 340734 343640 340740
rect 343640 340682 343692 340688
rect 333716 338026 333744 340068
rect 344296 338026 344324 361558
rect 345018 349616 345074 349625
rect 345018 349551 345074 349560
rect 345032 340814 345060 349551
rect 345020 340808 345072 340814
rect 345020 340750 345072 340756
rect 345676 340746 345704 361694
rect 352012 361684 352064 361690
rect 352012 361626 352064 361632
rect 352024 359924 352052 361626
rect 361684 359924 361712 361694
rect 371332 361616 371384 361622
rect 371332 361558 371384 361564
rect 371344 359924 371372 361558
rect 350446 350296 350502 350305
rect 350446 350231 350502 350240
rect 350460 340746 350488 350231
rect 371528 340762 371556 361694
rect 374644 361684 374696 361690
rect 374644 361626 374696 361632
rect 373264 361616 373316 361622
rect 373264 361558 373316 361564
rect 345664 340740 345716 340746
rect 345664 340682 345716 340688
rect 350448 340740 350500 340746
rect 371358 340734 371556 340762
rect 350448 340682 350500 340688
rect 333704 338020 333756 338026
rect 333704 337962 333756 337968
rect 344284 338020 344336 338026
rect 344284 337962 344336 337968
rect 352024 337958 352052 340068
rect 361684 338094 361712 340068
rect 373276 338094 373304 361558
rect 373998 349616 374054 349625
rect 373998 349551 374054 349560
rect 374012 340882 374040 349551
rect 374000 340876 374052 340882
rect 374000 340818 374052 340824
rect 374656 338094 374684 361626
rect 378046 350296 378102 350305
rect 378046 350231 378102 350240
rect 378060 340814 378088 350231
rect 378048 340808 378100 340814
rect 378048 340750 378100 340756
rect 361672 338088 361724 338094
rect 361672 338030 361724 338036
rect 373264 338088 373316 338094
rect 373264 338030 373316 338036
rect 374644 338088 374696 338094
rect 374644 338030 374696 338036
rect 323032 337952 323084 337958
rect 323032 337894 323084 337900
rect 352012 337952 352064 337958
rect 352012 337894 352064 337900
rect 334256 335504 334308 335510
rect 334256 335446 334308 335452
rect 324596 335368 324648 335374
rect 324596 335310 324648 335316
rect 324608 332860 324636 335310
rect 334268 332860 334296 335446
rect 352012 335436 352064 335442
rect 352012 335378 352064 335384
rect 347044 335368 347096 335374
rect 347044 335310 347096 335316
rect 343942 332302 344140 332330
rect 322846 322960 322902 322969
rect 322846 322895 322902 322904
rect 322860 314634 322888 322895
rect 322848 314628 322900 314634
rect 322848 314570 322900 314576
rect 324608 311778 324636 313140
rect 324596 311772 324648 311778
rect 324596 311714 324648 311720
rect 334268 311710 334296 313140
rect 343928 311846 343956 313140
rect 344112 311846 344140 332302
rect 345020 331288 345072 331294
rect 345020 331230 345072 331236
rect 345032 322833 345060 331230
rect 345018 322824 345074 322833
rect 345018 322759 345074 322768
rect 343916 311840 343968 311846
rect 343916 311782 343968 311788
rect 344100 311840 344152 311846
rect 344100 311782 344152 311788
rect 347056 311778 347084 335310
rect 348424 332580 348476 332586
rect 348424 332522 348476 332528
rect 347044 311772 347096 311778
rect 347044 311714 347096 311720
rect 348436 311710 348464 332522
rect 352024 325694 352052 335378
rect 361948 335368 362000 335374
rect 361948 335310 362000 335316
rect 373264 335368 373316 335374
rect 373264 335310 373316 335316
rect 361960 332874 361988 335310
rect 361960 332846 362296 332874
rect 352300 332586 352636 332602
rect 352288 332580 352636 332586
rect 352340 332574 352636 332580
rect 352288 332522 352340 332528
rect 371956 332302 372108 332330
rect 352024 325666 352236 325694
rect 350446 322960 350502 322969
rect 350446 322895 350502 322904
rect 350460 314566 350488 322895
rect 350448 314560 350500 314566
rect 350448 314502 350500 314508
rect 352208 313698 352236 325666
rect 352208 313670 352636 313698
rect 362296 313126 362632 313154
rect 362604 311778 362632 313126
rect 371620 313126 371956 313154
rect 371620 311846 371648 313126
rect 372080 311846 372108 332302
rect 371608 311840 371660 311846
rect 371608 311782 371660 311788
rect 372068 311840 372120 311846
rect 372068 311782 372120 311788
rect 373276 311778 373304 335310
rect 378046 322960 378102 322969
rect 378046 322895 378102 322904
rect 373998 322144 374054 322153
rect 373998 322079 374054 322088
rect 374012 314634 374040 322079
rect 378060 314634 378088 322895
rect 374000 314628 374052 314634
rect 374000 314570 374052 314576
rect 378048 314628 378100 314634
rect 378048 314570 378100 314576
rect 362592 311772 362644 311778
rect 362592 311714 362644 311720
rect 373264 311772 373316 311778
rect 373264 311714 373316 311720
rect 334256 311704 334308 311710
rect 334256 311646 334308 311652
rect 348424 311704 348476 311710
rect 348424 311646 348476 311652
rect 345664 307964 345716 307970
rect 345664 307906 345716 307912
rect 361672 307964 361724 307970
rect 361672 307906 361724 307912
rect 371516 307964 371568 307970
rect 371516 307906 371568 307912
rect 333704 307896 333756 307902
rect 333704 307838 333756 307844
rect 333716 305932 333744 307838
rect 343364 307828 343416 307834
rect 343364 307770 343416 307776
rect 344284 307828 344336 307834
rect 344284 307770 344336 307776
rect 343376 305932 343404 307770
rect 323044 305238 324070 305266
rect 322846 296304 322902 296313
rect 322846 296239 322902 296248
rect 322860 287026 322888 296239
rect 322848 287020 322900 287026
rect 322848 286962 322900 286968
rect 323044 284170 323072 305238
rect 323676 288380 323728 288386
rect 323676 288322 323728 288328
rect 323688 286770 323716 288322
rect 343548 286952 343600 286958
rect 343548 286894 343600 286900
rect 343560 286770 343588 286894
rect 323688 286742 324070 286770
rect 343390 286742 343588 286770
rect 333716 284238 333744 286076
rect 344296 284238 344324 307770
rect 345018 295624 345074 295633
rect 345018 295559 345074 295568
rect 345032 286890 345060 295559
rect 345676 286958 345704 307906
rect 352012 307896 352064 307902
rect 352012 307838 352064 307844
rect 352024 305932 352052 307838
rect 361684 305932 361712 307906
rect 371332 307828 371384 307834
rect 371332 307770 371384 307776
rect 371344 305932 371372 307770
rect 350446 296304 350502 296313
rect 350446 296239 350502 296248
rect 345664 286952 345716 286958
rect 345664 286894 345716 286900
rect 350460 286890 350488 296239
rect 345020 286884 345072 286890
rect 345020 286826 345072 286832
rect 350448 286884 350500 286890
rect 350448 286826 350500 286832
rect 371528 286770 371556 307906
rect 374644 307896 374696 307902
rect 374644 307838 374696 307844
rect 373264 307828 373316 307834
rect 373264 307770 373316 307776
rect 371358 286742 371556 286770
rect 333704 284232 333756 284238
rect 333704 284174 333756 284180
rect 344284 284232 344336 284238
rect 344284 284174 344336 284180
rect 352024 284170 352052 286076
rect 361684 284306 361712 286076
rect 373276 284306 373304 307770
rect 373998 295624 374054 295633
rect 373998 295559 374054 295568
rect 374012 287026 374040 295559
rect 374000 287020 374052 287026
rect 374000 286962 374052 286968
rect 374656 284306 374684 307838
rect 378046 296304 378102 296313
rect 378046 296239 378102 296248
rect 378060 286958 378088 296239
rect 378048 286952 378100 286958
rect 378048 286894 378100 286900
rect 361672 284300 361724 284306
rect 361672 284242 361724 284248
rect 373264 284300 373316 284306
rect 373264 284242 373316 284248
rect 374644 284300 374696 284306
rect 374644 284242 374696 284248
rect 323032 284164 323084 284170
rect 323032 284106 323084 284112
rect 352012 284164 352064 284170
rect 352012 284106 352064 284112
rect 352012 280424 352064 280430
rect 352012 280366 352064 280372
rect 334256 280356 334308 280362
rect 334256 280298 334308 280304
rect 347044 280356 347096 280362
rect 347044 280298 347096 280304
rect 324596 280220 324648 280226
rect 324596 280162 324648 280168
rect 324608 278868 324636 280162
rect 334268 278868 334296 280298
rect 343942 278310 344140 278338
rect 322848 277500 322900 277506
rect 322848 277442 322900 277448
rect 322860 270065 322888 277442
rect 322846 270056 322902 270065
rect 322846 269991 322902 270000
rect 324608 256630 324636 259148
rect 324596 256624 324648 256630
rect 324596 256566 324648 256572
rect 334268 256562 334296 259148
rect 343928 256698 343956 259148
rect 344112 256698 344140 278310
rect 345020 277432 345072 277438
rect 345020 277374 345072 277380
rect 345032 269113 345060 277374
rect 345018 269104 345074 269113
rect 345018 269039 345074 269048
rect 343916 256692 343968 256698
rect 343916 256634 343968 256640
rect 344100 256692 344152 256698
rect 344100 256634 344152 256640
rect 347056 256630 347084 280298
rect 348424 280220 348476 280226
rect 348424 280162 348476 280168
rect 347044 256624 347096 256630
rect 347044 256566 347096 256572
rect 348436 256562 348464 280162
rect 350448 277432 350500 277438
rect 350448 277374 350500 277380
rect 350460 270065 350488 277374
rect 350446 270056 350502 270065
rect 350446 269991 350502 270000
rect 352024 267734 352052 280366
rect 352288 280220 352340 280226
rect 352288 280162 352340 280168
rect 361948 280220 362000 280226
rect 361948 280162 362000 280168
rect 373264 280220 373316 280226
rect 373264 280162 373316 280168
rect 352300 278882 352328 280162
rect 361960 278882 361988 280162
rect 352300 278854 352636 278882
rect 361960 278854 362296 278882
rect 371956 278310 372108 278338
rect 352024 267706 352236 267734
rect 352208 259706 352236 267706
rect 352208 259678 352636 259706
rect 362296 259134 362632 259162
rect 362604 256630 362632 259134
rect 371620 259134 371956 259162
rect 371620 256698 371648 259134
rect 372080 256698 372108 278310
rect 371608 256692 371660 256698
rect 371608 256634 371660 256640
rect 372068 256692 372120 256698
rect 372068 256634 372120 256640
rect 373276 256630 373304 280162
rect 374000 277500 374052 277506
rect 374000 277442 374052 277448
rect 378048 277500 378100 277506
rect 378048 277442 378100 277448
rect 374012 269113 374040 277442
rect 378060 270065 378088 277442
rect 378046 270056 378102 270065
rect 378046 269991 378102 270000
rect 373998 269104 374054 269113
rect 373998 269039 374054 269048
rect 362592 256624 362644 256630
rect 362592 256566 362644 256572
rect 373264 256624 373316 256630
rect 373264 256566 373316 256572
rect 334256 256556 334308 256562
rect 334256 256498 334308 256504
rect 348424 256556 348476 256562
rect 348424 256498 348476 256504
rect 345664 254108 345716 254114
rect 345664 254050 345716 254056
rect 361672 254108 361724 254114
rect 361672 254050 361724 254056
rect 371516 254108 371568 254114
rect 371516 254050 371568 254056
rect 333704 254040 333756 254046
rect 333704 253982 333756 253988
rect 333716 251940 333744 253982
rect 343364 253972 343416 253978
rect 343364 253914 343416 253920
rect 344284 253972 344336 253978
rect 344284 253914 344336 253920
rect 343376 251940 343404 253914
rect 322848 251252 322900 251258
rect 322848 251194 322900 251200
rect 323044 251246 324070 251274
rect 322860 242321 322888 251194
rect 322846 242312 322902 242321
rect 322846 242247 322902 242256
rect 323044 230314 323072 251246
rect 323676 233436 323728 233442
rect 323676 233378 323728 233384
rect 323688 232778 323716 233378
rect 323688 232750 324070 232778
rect 343390 232762 343680 232778
rect 343390 232756 343692 232762
rect 343390 232750 343640 232756
rect 343640 232698 343692 232704
rect 333716 230382 333744 232084
rect 344296 230382 344324 253914
rect 345020 251320 345072 251326
rect 345020 251262 345072 251268
rect 345032 241641 345060 251262
rect 345018 241632 345074 241641
rect 345018 241567 345074 241576
rect 345676 232762 345704 254050
rect 352012 254040 352064 254046
rect 352012 253982 352064 253988
rect 352024 251940 352052 253982
rect 361684 251940 361712 254050
rect 371332 253972 371384 253978
rect 371332 253914 371384 253920
rect 371344 251940 371372 253914
rect 350448 251388 350500 251394
rect 350448 251330 350500 251336
rect 350460 242321 350488 251330
rect 350446 242312 350502 242321
rect 350446 242247 350502 242256
rect 371528 232778 371556 254050
rect 374644 254040 374696 254046
rect 374644 253982 374696 253988
rect 373264 253972 373316 253978
rect 373264 253914 373316 253920
rect 345664 232756 345716 232762
rect 371358 232750 371556 232778
rect 345664 232698 345716 232704
rect 333704 230376 333756 230382
rect 333704 230318 333756 230324
rect 344284 230376 344336 230382
rect 344284 230318 344336 230324
rect 352024 230314 352052 232084
rect 361684 230450 361712 232084
rect 373276 230450 373304 253914
rect 374000 251252 374052 251258
rect 374000 251194 374052 251200
rect 374012 241641 374040 251194
rect 373998 241632 374054 241641
rect 373998 241567 374054 241576
rect 361672 230444 361724 230450
rect 361672 230386 361724 230392
rect 373264 230444 373316 230450
rect 373264 230386 373316 230392
rect 374656 230382 374684 253982
rect 378048 251320 378100 251326
rect 378048 251262 378100 251268
rect 378060 242321 378088 251262
rect 378046 242312 378102 242321
rect 378046 242247 378102 242256
rect 374644 230376 374696 230382
rect 374644 230318 374696 230324
rect 323032 230308 323084 230314
rect 323032 230250 323084 230256
rect 352012 230308 352064 230314
rect 352012 230250 352064 230256
rect 334256 226500 334308 226506
rect 334256 226442 334308 226448
rect 352196 226500 352248 226506
rect 352196 226442 352248 226448
rect 324596 226364 324648 226370
rect 324596 226306 324648 226312
rect 324608 224876 324636 226306
rect 334268 224876 334296 226442
rect 347044 226432 347096 226438
rect 347044 226374 347096 226380
rect 343942 224318 344140 224346
rect 322848 223644 322900 223650
rect 322848 223586 322900 223592
rect 322860 215393 322888 223586
rect 322846 215384 322902 215393
rect 322846 215319 322902 215328
rect 324608 202774 324636 205020
rect 324596 202768 324648 202774
rect 324596 202710 324648 202716
rect 334268 202706 334296 205020
rect 343928 202842 343956 205020
rect 344112 202842 344140 224318
rect 345020 223712 345072 223718
rect 345020 223654 345072 223660
rect 345032 214713 345060 223654
rect 345018 214704 345074 214713
rect 345018 214639 345074 214648
rect 343916 202836 343968 202842
rect 343916 202778 343968 202784
rect 344100 202836 344152 202842
rect 344100 202778 344152 202784
rect 347056 202774 347084 226374
rect 348424 226364 348476 226370
rect 348424 226306 348476 226312
rect 347044 202768 347096 202774
rect 347044 202710 347096 202716
rect 348436 202706 348464 226306
rect 350448 223780 350500 223786
rect 350448 223722 350500 223728
rect 350460 215393 350488 223722
rect 350446 215384 350502 215393
rect 350446 215319 350502 215328
rect 352208 205714 352236 226442
rect 361948 226432 362000 226438
rect 361948 226374 362000 226380
rect 352288 226364 352340 226370
rect 352288 226306 352340 226312
rect 352300 224890 352328 226306
rect 361960 224890 361988 226374
rect 373264 226364 373316 226370
rect 373264 226306 373316 226312
rect 352300 224862 352636 224890
rect 361960 224862 362296 224890
rect 371956 224318 372108 224346
rect 352208 205686 352636 205714
rect 362296 205006 362632 205034
rect 362604 202774 362632 205006
rect 371620 205006 371956 205034
rect 371620 202842 371648 205006
rect 372080 202842 372108 224318
rect 371608 202836 371660 202842
rect 371608 202778 371660 202784
rect 372068 202836 372120 202842
rect 372068 202778 372120 202784
rect 373276 202774 373304 226306
rect 378048 223712 378100 223718
rect 378048 223654 378100 223660
rect 374000 223644 374052 223650
rect 374000 223586 374052 223592
rect 374012 215257 374040 223586
rect 378060 215393 378088 223654
rect 378046 215384 378102 215393
rect 378046 215319 378102 215328
rect 373998 215248 374054 215257
rect 373998 215183 374054 215192
rect 362592 202768 362644 202774
rect 362592 202710 362644 202716
rect 373264 202768 373316 202774
rect 373264 202710 373316 202716
rect 334256 202700 334308 202706
rect 334256 202642 334308 202648
rect 348424 202700 348476 202706
rect 348424 202642 348476 202648
rect 345664 200320 345716 200326
rect 345664 200262 345716 200268
rect 361672 200320 361724 200326
rect 361672 200262 361724 200268
rect 371516 200320 371568 200326
rect 371516 200262 371568 200268
rect 333704 200252 333756 200258
rect 333704 200194 333756 200200
rect 333716 197948 333744 200194
rect 343364 200184 343416 200190
rect 343364 200126 343416 200132
rect 344284 200184 344336 200190
rect 344284 200126 344336 200132
rect 343376 197948 343404 200126
rect 323044 197254 324070 197282
rect 322846 188320 322902 188329
rect 322846 188255 322902 188264
rect 322860 179382 322888 188255
rect 322848 179376 322900 179382
rect 322848 179318 322900 179324
rect 323044 176526 323072 197254
rect 323676 179512 323728 179518
rect 323676 179454 323728 179460
rect 323688 178786 323716 179454
rect 343548 179308 343600 179314
rect 343548 179250 343600 179256
rect 343560 178786 343588 179250
rect 323688 178758 324070 178786
rect 343390 178758 343588 178786
rect 333716 176594 333744 178092
rect 344296 176594 344324 200126
rect 345018 187640 345074 187649
rect 345018 187575 345074 187584
rect 345032 179246 345060 187575
rect 345676 179314 345704 200262
rect 352012 200252 352064 200258
rect 352012 200194 352064 200200
rect 352024 197948 352052 200194
rect 361684 197948 361712 200262
rect 371332 200184 371384 200190
rect 371332 200126 371384 200132
rect 371344 197948 371372 200126
rect 350446 188320 350502 188329
rect 350446 188255 350502 188264
rect 345664 179308 345716 179314
rect 345664 179250 345716 179256
rect 350460 179246 350488 188255
rect 345020 179240 345072 179246
rect 345020 179182 345072 179188
rect 350448 179240 350500 179246
rect 350448 179182 350500 179188
rect 371528 178786 371556 200262
rect 374644 200252 374696 200258
rect 374644 200194 374696 200200
rect 373264 200184 373316 200190
rect 373264 200126 373316 200132
rect 371358 178758 371556 178786
rect 333704 176588 333756 176594
rect 333704 176530 333756 176536
rect 344284 176588 344336 176594
rect 344284 176530 344336 176536
rect 352024 176526 352052 178092
rect 361684 176662 361712 178092
rect 373276 176662 373304 200126
rect 373998 187640 374054 187649
rect 373998 187575 374054 187584
rect 374012 179382 374040 187575
rect 374000 179376 374052 179382
rect 374000 179318 374052 179324
rect 374656 176662 374684 200194
rect 378046 188320 378102 188329
rect 378046 188255 378102 188264
rect 378060 179314 378088 188255
rect 378048 179308 378100 179314
rect 378048 179250 378100 179256
rect 361672 176656 361724 176662
rect 361672 176598 361724 176604
rect 373264 176656 373316 176662
rect 373264 176598 373316 176604
rect 374644 176656 374696 176662
rect 374644 176598 374696 176604
rect 323032 176520 323084 176526
rect 323032 176462 323084 176468
rect 352012 176520 352064 176526
rect 352012 176462 352064 176468
rect 334256 172712 334308 172718
rect 334256 172654 334308 172660
rect 352012 172712 352064 172718
rect 352012 172654 352064 172660
rect 324596 172576 324648 172582
rect 324596 172518 324648 172524
rect 324608 170884 324636 172518
rect 334268 170884 334296 172654
rect 345664 172644 345716 172650
rect 345664 172586 345716 172592
rect 343942 170326 344140 170354
rect 322846 161392 322902 161401
rect 322846 161327 322902 161336
rect 322860 151774 322888 161327
rect 322848 151768 322900 151774
rect 322848 151710 322900 151716
rect 324608 148986 324636 151028
rect 324596 148980 324648 148986
rect 324596 148922 324648 148928
rect 334268 148918 334296 151028
rect 343928 149054 343956 151028
rect 344112 149054 344140 170326
rect 345018 160712 345074 160721
rect 345018 160647 345074 160656
rect 345032 151706 345060 160647
rect 345020 151700 345072 151706
rect 345020 151642 345072 151648
rect 343916 149048 343968 149054
rect 343916 148990 343968 148996
rect 344100 149048 344152 149054
rect 344100 148990 344152 148996
rect 345676 148986 345704 172586
rect 347044 172576 347096 172582
rect 347044 172518 347096 172524
rect 345664 148980 345716 148986
rect 345664 148922 345716 148928
rect 347056 148918 347084 172518
rect 352024 171134 352052 172654
rect 361948 172644 362000 172650
rect 361948 172586 362000 172592
rect 352288 172576 352340 172582
rect 352288 172518 352340 172524
rect 352024 171106 352236 171134
rect 350446 161392 350502 161401
rect 350446 161327 350502 161336
rect 350460 151638 350488 161327
rect 352208 151722 352236 171106
rect 352300 170898 352328 172518
rect 361960 170898 361988 172586
rect 373264 172576 373316 172582
rect 373264 172518 373316 172524
rect 352300 170870 352636 170898
rect 361960 170870 362296 170898
rect 371956 170326 372108 170354
rect 352208 151694 352636 151722
rect 350448 151632 350500 151638
rect 350448 151574 350500 151580
rect 362296 151014 362632 151042
rect 362604 148986 362632 151014
rect 371620 151014 371956 151042
rect 371620 149054 371648 151014
rect 372080 149054 372108 170326
rect 371608 149048 371660 149054
rect 371608 148990 371660 148996
rect 372068 149048 372120 149054
rect 372068 148990 372120 148996
rect 373276 148986 373304 172518
rect 378046 161392 378102 161401
rect 378046 161327 378102 161336
rect 373998 160712 374054 160721
rect 373998 160647 374054 160656
rect 374012 151774 374040 160647
rect 374000 151768 374052 151774
rect 374000 151710 374052 151716
rect 378060 151706 378088 161327
rect 378048 151700 378100 151706
rect 378048 151642 378100 151648
rect 362592 148980 362644 148986
rect 362592 148922 362644 148928
rect 373264 148980 373316 148986
rect 373264 148922 373316 148928
rect 334256 148912 334308 148918
rect 334256 148854 334308 148860
rect 347044 148912 347096 148918
rect 347044 148854 347096 148860
rect 345664 146464 345716 146470
rect 345664 146406 345716 146412
rect 361672 146464 361724 146470
rect 361672 146406 361724 146412
rect 371516 146464 371568 146470
rect 371516 146406 371568 146412
rect 333704 146396 333756 146402
rect 333704 146338 333756 146344
rect 333716 143956 333744 146338
rect 343364 146328 343416 146334
rect 343364 146270 343416 146276
rect 344284 146328 344336 146334
rect 344284 146270 344336 146276
rect 343376 143956 343404 146270
rect 323044 143262 324070 143290
rect 322846 134328 322902 134337
rect 322846 134263 322902 134272
rect 322860 125594 322888 134263
rect 322848 125588 322900 125594
rect 322848 125530 322900 125536
rect 323044 122670 323072 143262
rect 323676 126132 323728 126138
rect 323676 126074 323728 126080
rect 323688 124794 323716 126074
rect 343548 124840 343600 124846
rect 323688 124766 324070 124794
rect 343390 124788 343548 124794
rect 343390 124782 343600 124788
rect 343390 124766 343588 124782
rect 333716 122738 333744 124100
rect 344296 122738 344324 146270
rect 345018 133648 345074 133657
rect 345018 133583 345074 133592
rect 345032 125526 345060 133583
rect 345020 125520 345072 125526
rect 345020 125462 345072 125468
rect 345676 124846 345704 146406
rect 352012 146396 352064 146402
rect 352012 146338 352064 146344
rect 352024 143956 352052 146338
rect 361684 143956 361712 146406
rect 371332 146328 371384 146334
rect 371332 146270 371384 146276
rect 371344 143956 371372 146270
rect 350446 134328 350502 134337
rect 350446 134263 350502 134272
rect 350460 125458 350488 134263
rect 350448 125452 350500 125458
rect 350448 125394 350500 125400
rect 345664 124840 345716 124846
rect 371528 124794 371556 146406
rect 374644 146396 374696 146402
rect 374644 146338 374696 146344
rect 373264 146328 373316 146334
rect 373264 146270 373316 146276
rect 345664 124782 345716 124788
rect 371358 124766 371556 124794
rect 333704 122732 333756 122738
rect 333704 122674 333756 122680
rect 344284 122732 344336 122738
rect 344284 122674 344336 122680
rect 352024 122670 352052 124100
rect 361684 122806 361712 124100
rect 373276 122806 373304 146270
rect 373998 133648 374054 133657
rect 373998 133583 374054 133592
rect 374012 125594 374040 133583
rect 374000 125588 374052 125594
rect 374000 125530 374052 125536
rect 361672 122800 361724 122806
rect 361672 122742 361724 122748
rect 373264 122800 373316 122806
rect 373264 122742 373316 122748
rect 374656 122738 374684 146338
rect 378046 134328 378102 134337
rect 378046 134263 378102 134272
rect 378060 125526 378088 134263
rect 378048 125520 378100 125526
rect 378048 125462 378100 125468
rect 374644 122732 374696 122738
rect 374644 122674 374696 122680
rect 323032 122664 323084 122670
rect 323032 122606 323084 122612
rect 352012 122664 352064 122670
rect 352012 122606 352064 122612
rect 334256 118856 334308 118862
rect 334256 118798 334308 118804
rect 352012 118856 352064 118862
rect 352012 118798 352064 118804
rect 324596 118720 324648 118726
rect 324596 118662 324648 118668
rect 324608 116892 324636 118662
rect 334268 116892 334296 118798
rect 345664 118788 345716 118794
rect 345664 118730 345716 118736
rect 343942 116334 344140 116362
rect 322846 107400 322902 107409
rect 322846 107335 322902 107344
rect 322860 97986 322888 107335
rect 322848 97980 322900 97986
rect 322848 97922 322900 97928
rect 324608 95130 324636 97036
rect 324596 95124 324648 95130
rect 324596 95066 324648 95072
rect 334268 95062 334296 97036
rect 343928 95198 343956 97036
rect 344112 95198 344140 116334
rect 345018 106720 345074 106729
rect 345018 106655 345074 106664
rect 345032 97918 345060 106655
rect 345020 97912 345072 97918
rect 345020 97854 345072 97860
rect 343916 95192 343968 95198
rect 343916 95134 343968 95140
rect 344100 95192 344152 95198
rect 344100 95134 344152 95140
rect 345676 95130 345704 118730
rect 347044 118720 347096 118726
rect 347044 118662 347096 118668
rect 345664 95124 345716 95130
rect 345664 95066 345716 95072
rect 347056 95062 347084 118662
rect 352024 113174 352052 118798
rect 361948 118788 362000 118794
rect 361948 118730 362000 118736
rect 352288 118720 352340 118726
rect 352288 118662 352340 118668
rect 352300 116906 352328 118662
rect 361960 116906 361988 118730
rect 373264 118720 373316 118726
rect 373264 118662 373316 118668
rect 352300 116878 352636 116906
rect 361960 116878 362296 116906
rect 371956 116334 372108 116362
rect 352024 113146 352236 113174
rect 350446 107400 350502 107409
rect 350446 107335 350502 107344
rect 350460 97850 350488 107335
rect 350448 97844 350500 97850
rect 350448 97786 350500 97792
rect 352208 97730 352236 113146
rect 352208 97702 352636 97730
rect 362296 97022 362632 97050
rect 362604 95130 362632 97022
rect 371620 97022 371956 97050
rect 371620 95198 371648 97022
rect 372080 95198 372108 116334
rect 371608 95192 371660 95198
rect 371608 95134 371660 95140
rect 372068 95192 372120 95198
rect 372068 95134 372120 95140
rect 373276 95130 373304 118662
rect 378046 107400 378102 107409
rect 378046 107335 378102 107344
rect 373998 106720 374054 106729
rect 373998 106655 374054 106664
rect 374012 97986 374040 106655
rect 374000 97980 374052 97986
rect 374000 97922 374052 97928
rect 378060 97918 378088 107335
rect 378048 97912 378100 97918
rect 378048 97854 378100 97860
rect 362592 95124 362644 95130
rect 362592 95066 362644 95072
rect 373264 95124 373316 95130
rect 373264 95066 373316 95072
rect 334256 95056 334308 95062
rect 334256 94998 334308 95004
rect 347044 95056 347096 95062
rect 347044 94998 347096 95004
rect 333704 91248 333756 91254
rect 333704 91190 333756 91196
rect 345664 91248 345716 91254
rect 345664 91190 345716 91196
rect 361672 91248 361724 91254
rect 361672 91190 361724 91196
rect 371516 91248 371568 91254
rect 371516 91190 371568 91196
rect 333716 89964 333744 91190
rect 343364 91112 343416 91118
rect 343364 91054 343416 91060
rect 344284 91112 344336 91118
rect 344284 91054 344336 91060
rect 343376 89964 343404 91054
rect 323044 89270 324070 89298
rect 322848 88392 322900 88398
rect 322848 88334 322900 88340
rect 322860 80345 322888 88334
rect 322846 80336 322902 80345
rect 322846 80271 322902 80280
rect 323044 68882 323072 89270
rect 323676 72344 323728 72350
rect 323676 72286 323728 72292
rect 323688 70666 323716 72286
rect 343548 71664 343600 71670
rect 343548 71606 343600 71612
rect 343560 70666 343588 71606
rect 323688 70638 324070 70666
rect 343390 70638 343588 70666
rect 333716 68950 333744 70108
rect 344296 68950 344324 91054
rect 345018 79656 345074 79665
rect 345018 79591 345074 79600
rect 345032 71738 345060 79591
rect 345020 71732 345072 71738
rect 345020 71674 345072 71680
rect 345676 71670 345704 91190
rect 352012 91180 352064 91186
rect 352012 91122 352064 91128
rect 352024 89964 352052 91122
rect 361684 89964 361712 91190
rect 371332 91112 371384 91118
rect 371332 91054 371384 91060
rect 371344 89964 371372 91054
rect 350446 80336 350502 80345
rect 350446 80271 350502 80280
rect 350460 71738 350488 80271
rect 350448 71732 350500 71738
rect 350448 71674 350500 71680
rect 345664 71664 345716 71670
rect 345664 71606 345716 71612
rect 371528 70666 371556 91190
rect 374644 91180 374696 91186
rect 374644 91122 374696 91128
rect 373264 91112 373316 91118
rect 373264 91054 373316 91060
rect 371358 70638 371556 70666
rect 333704 68944 333756 68950
rect 333704 68886 333756 68892
rect 344284 68944 344336 68950
rect 344284 68886 344336 68892
rect 352024 68882 352052 70108
rect 361684 69018 361712 70108
rect 373276 69018 373304 91054
rect 374000 88392 374052 88398
rect 374000 88334 374052 88340
rect 374012 79665 374040 88334
rect 373998 79656 374054 79665
rect 373998 79591 374054 79600
rect 361672 69012 361724 69018
rect 361672 68954 361724 68960
rect 373264 69012 373316 69018
rect 373264 68954 373316 68960
rect 374656 68950 374684 91122
rect 378048 88392 378100 88398
rect 378048 88334 378100 88340
rect 378060 80345 378088 88334
rect 378046 80336 378102 80345
rect 378046 80271 378102 80280
rect 374644 68944 374696 68950
rect 374644 68886 374696 68892
rect 323032 68876 323084 68882
rect 323032 68818 323084 68824
rect 352012 68876 352064 68882
rect 352012 68818 352064 68824
rect 334256 65068 334308 65074
rect 334256 65010 334308 65016
rect 352012 65068 352064 65074
rect 352012 65010 352064 65016
rect 324596 64932 324648 64938
rect 324596 64874 324648 64880
rect 324608 62900 324636 64874
rect 334268 62900 334296 65010
rect 345664 65000 345716 65006
rect 345664 64942 345716 64948
rect 343942 62206 344140 62234
rect 322848 62144 322900 62150
rect 322848 62086 322900 62092
rect 322860 53417 322888 62086
rect 322846 53408 322902 53417
rect 322846 53343 322902 53352
rect 324608 41342 324636 43044
rect 324596 41336 324648 41342
rect 324596 41278 324648 41284
rect 334268 41274 334296 43044
rect 343928 41410 343956 43044
rect 344112 41410 344140 62206
rect 345018 52728 345074 52737
rect 345018 52663 345074 52672
rect 345032 44130 345060 52663
rect 345020 44124 345072 44130
rect 345020 44066 345072 44072
rect 343916 41404 343968 41410
rect 343916 41346 343968 41352
rect 344100 41404 344152 41410
rect 344100 41346 344152 41352
rect 345676 41342 345704 64942
rect 347044 64932 347096 64938
rect 347044 64874 347096 64880
rect 345664 41336 345716 41342
rect 345664 41278 345716 41284
rect 347056 41274 347084 64874
rect 352024 55214 352052 65010
rect 361948 65000 362000 65006
rect 361948 64942 362000 64948
rect 352288 64932 352340 64938
rect 352288 64874 352340 64880
rect 352300 62914 352328 64874
rect 361960 62914 361988 64942
rect 373264 64932 373316 64938
rect 373264 64874 373316 64880
rect 352300 62886 352636 62914
rect 361960 62886 362296 62914
rect 371956 62206 372108 62234
rect 352024 55186 352236 55214
rect 350446 53408 350502 53417
rect 350446 53343 350502 53352
rect 350460 44130 350488 53343
rect 350448 44124 350500 44130
rect 350448 44066 350500 44072
rect 352208 43738 352236 55186
rect 352208 43710 352636 43738
rect 362296 43030 362632 43058
rect 362604 41342 362632 43030
rect 371620 43030 371956 43058
rect 371620 41410 371648 43030
rect 372080 41410 372108 62206
rect 371608 41404 371660 41410
rect 371608 41346 371660 41352
rect 372068 41404 372120 41410
rect 372068 41346 372120 41352
rect 373276 41342 373304 64874
rect 374000 62144 374052 62150
rect 374000 62086 374052 62092
rect 378048 62144 378100 62150
rect 378048 62086 378100 62092
rect 374012 52737 374040 62086
rect 378060 53417 378088 62086
rect 378046 53408 378102 53417
rect 378046 53343 378102 53352
rect 373998 52728 374054 52737
rect 373998 52663 374054 52672
rect 362592 41336 362644 41342
rect 362592 41278 362644 41284
rect 373264 41336 373316 41342
rect 373264 41278 373316 41284
rect 334256 41268 334308 41274
rect 334256 41210 334308 41216
rect 347044 41268 347096 41274
rect 347044 41210 347096 41216
rect 322204 38344 322256 38350
rect 322204 38286 322256 38292
rect 249708 37460 249760 37466
rect 249708 37402 249760 37408
rect 260196 37460 260248 37466
rect 260196 37402 260248 37408
rect 277676 37460 277728 37466
rect 277676 37402 277728 37408
rect 287520 37460 287572 37466
rect 287520 37402 287572 37408
rect 305368 37460 305420 37466
rect 305368 37402 305420 37408
rect 345664 37460 345716 37466
rect 345664 37402 345716 37408
rect 361672 37460 361724 37466
rect 361672 37402 361724 37408
rect 371516 37460 371568 37466
rect 371516 37402 371568 37408
rect 239404 37324 239456 37330
rect 239404 37266 239456 37272
rect 238668 34604 238720 34610
rect 238668 34546 238720 34552
rect 238680 26353 238708 34546
rect 238852 30796 238904 30802
rect 238852 30738 238904 30744
rect 238666 26344 238722 26353
rect 238666 26279 238722 26288
rect 233884 15088 233936 15094
rect 233884 15030 233936 15036
rect 156052 13388 156104 13394
rect 156052 13330 156104 13336
rect 183652 13388 183704 13394
rect 183652 13330 183704 13336
rect 211712 13388 211764 13394
rect 211712 13330 211764 13336
rect 222016 13388 222068 13394
rect 222016 13330 222068 13336
rect 99472 13320 99524 13326
rect 99472 13262 99524 13268
rect 109684 13320 109736 13326
rect 109684 13262 109736 13268
rect 120724 13320 120776 13326
rect 120724 13262 120776 13268
rect 127072 13320 127124 13326
rect 127072 13262 127124 13268
rect 137652 13320 137704 13326
rect 137652 13262 137704 13268
rect 148324 13320 148376 13326
rect 148324 13262 148376 13268
rect 238864 13258 238892 30738
rect 239416 13394 239444 37266
rect 249720 35972 249748 37402
rect 259368 37324 259420 37330
rect 259368 37266 259420 37272
rect 260104 37324 260156 37330
rect 260104 37266 260156 37272
rect 259380 35972 259408 37266
rect 239784 35278 240074 35306
rect 239784 30802 239812 35278
rect 239772 30796 239824 30802
rect 239772 30738 239824 30744
rect 259736 21480 259788 21486
rect 259736 21422 259788 21428
rect 239772 18012 239824 18018
rect 239772 17954 239824 17960
rect 239784 16674 239812 17954
rect 259748 16674 259776 21422
rect 239784 16646 240074 16674
rect 259394 16646 259776 16674
rect 249720 13802 249748 16116
rect 260116 13802 260144 37266
rect 260208 21486 260236 37402
rect 268016 37392 268068 37398
rect 268016 37334 268068 37340
rect 268028 35972 268056 37334
rect 277688 35972 277716 37402
rect 287336 37324 287388 37330
rect 287336 37266 287388 37272
rect 287348 35972 287376 37266
rect 266268 34672 266320 34678
rect 266268 34614 266320 34620
rect 262220 34536 262272 34542
rect 262220 34478 262272 34484
rect 262232 25673 262260 34478
rect 266280 26353 266308 34614
rect 266266 26344 266322 26353
rect 266266 26279 266322 26288
rect 262218 25664 262274 25673
rect 262218 25599 262274 25608
rect 260196 21480 260248 21486
rect 260196 21422 260248 21428
rect 287532 16674 287560 37402
rect 287704 37392 287756 37398
rect 287704 37334 287756 37340
rect 296168 37392 296220 37398
rect 296168 37334 296220 37340
rect 287716 18290 287744 37334
rect 289084 37324 289136 37330
rect 289084 37266 289136 37272
rect 287704 18284 287756 18290
rect 287704 18226 287756 18232
rect 287362 16646 287560 16674
rect 249708 13796 249760 13802
rect 249708 13738 249760 13744
rect 260104 13796 260156 13802
rect 260104 13738 260156 13744
rect 239404 13388 239456 13394
rect 239404 13330 239456 13336
rect 268028 13258 268056 16116
rect 277688 13802 277716 16116
rect 289096 13802 289124 37266
rect 296180 35986 296208 37334
rect 296056 35958 296208 35986
rect 305380 35986 305408 37402
rect 316776 37392 316828 37398
rect 316776 37334 316828 37340
rect 322296 37392 322348 37398
rect 322296 37334 322348 37340
rect 333704 37392 333756 37398
rect 333704 37334 333756 37340
rect 315028 37324 315080 37330
rect 315028 37266 315080 37272
rect 316684 37324 316736 37330
rect 316684 37266 316736 37272
rect 315040 35986 315068 37266
rect 305380 35958 305716 35986
rect 315040 35958 315376 35986
rect 289820 34604 289872 34610
rect 289820 34546 289872 34552
rect 289832 25673 289860 34546
rect 293868 34536 293920 34542
rect 293868 34478 293920 34484
rect 293880 26353 293908 34478
rect 293866 26344 293922 26353
rect 293866 26279 293922 26288
rect 289818 25664 289874 25673
rect 289818 25599 289874 25608
rect 295708 18284 295760 18290
rect 295708 18226 295760 18232
rect 295720 16674 295748 18226
rect 295720 16646 296056 16674
rect 305716 16102 306052 16130
rect 315376 16102 315712 16130
rect 306024 13802 306052 16102
rect 277676 13796 277728 13802
rect 277676 13738 277728 13744
rect 289084 13796 289136 13802
rect 289084 13738 289136 13744
rect 306012 13796 306064 13802
rect 306012 13738 306064 13744
rect 315684 13394 315712 16102
rect 316696 13802 316724 37266
rect 316788 18154 316816 37334
rect 317420 34672 317472 34678
rect 317420 34614 317472 34620
rect 317432 25673 317460 34614
rect 317418 25664 317474 25673
rect 317418 25599 317474 25608
rect 316776 18148 316828 18154
rect 316776 18090 316828 18096
rect 316684 13796 316736 13802
rect 316684 13738 316736 13744
rect 322308 13394 322336 37334
rect 333716 35972 333744 37334
rect 343364 37324 343416 37330
rect 343364 37266 343416 37272
rect 344284 37324 344336 37330
rect 344284 37266 344336 37272
rect 343376 35972 343404 37266
rect 323044 35278 324070 35306
rect 322848 34604 322900 34610
rect 322848 34546 322900 34552
rect 322860 26353 322888 34546
rect 322846 26344 322902 26353
rect 322846 26279 322902 26288
rect 323044 13394 323072 35278
rect 323676 18148 323728 18154
rect 323676 18090 323728 18096
rect 323688 16674 323716 18090
rect 323688 16646 324070 16674
rect 343548 16584 343600 16590
rect 343390 16532 343548 16538
rect 343390 16526 343600 16532
rect 343390 16510 343588 16526
rect 315672 13388 315724 13394
rect 315672 13330 315724 13336
rect 322296 13388 322348 13394
rect 322296 13330 322348 13336
rect 323032 13388 323084 13394
rect 323032 13330 323084 13336
rect 333716 13326 333744 16116
rect 344296 13326 344324 37266
rect 345020 34536 345072 34542
rect 345020 34478 345072 34484
rect 345032 25673 345060 34478
rect 345018 25664 345074 25673
rect 345018 25599 345074 25608
rect 345676 16590 345704 37402
rect 352012 37392 352064 37398
rect 352012 37334 352064 37340
rect 352024 35972 352052 37334
rect 361684 35972 361712 37402
rect 371332 37324 371384 37330
rect 371332 37266 371384 37272
rect 371344 35972 371372 37266
rect 350448 34536 350500 34542
rect 350448 34478 350500 34484
rect 350460 26353 350488 34478
rect 350446 26344 350502 26353
rect 350446 26279 350502 26288
rect 371528 16674 371556 37402
rect 374644 37392 374696 37398
rect 374644 37334 374696 37340
rect 373264 37324 373316 37330
rect 373264 37266 373316 37272
rect 371358 16646 371556 16674
rect 345664 16584 345716 16590
rect 345664 16526 345716 16532
rect 352024 13394 352052 16116
rect 361684 13802 361712 16116
rect 373276 13802 373304 37266
rect 374000 34604 374052 34610
rect 374000 34546 374052 34552
rect 374012 25673 374040 34546
rect 373998 25664 374054 25673
rect 373998 25599 374054 25608
rect 374656 13802 374684 37334
rect 378048 34604 378100 34610
rect 378048 34546 378100 34552
rect 378060 26353 378088 34546
rect 378046 26344 378102 26353
rect 378046 26279 378102 26288
rect 361672 13796 361724 13802
rect 361672 13738 361724 13744
rect 373264 13796 373316 13802
rect 373264 13738 373316 13744
rect 374644 13796 374696 13802
rect 374644 13738 374696 13744
rect 378796 13462 378824 700334
rect 408040 686112 408092 686118
rect 408040 686054 408092 686060
rect 428648 686112 428700 686118
rect 428648 686054 428700 686060
rect 389364 686044 389416 686050
rect 389364 685986 389416 685992
rect 399484 686044 399536 686050
rect 399484 685986 399536 685992
rect 389376 683890 389404 685986
rect 399024 685908 399076 685914
rect 399024 685850 399076 685856
rect 399036 683890 399064 685850
rect 389376 683862 389712 683890
rect 399036 683862 399372 683890
rect 379624 683318 380052 683346
rect 379624 662386 379652 683318
rect 399496 664714 399524 685986
rect 400864 685908 400916 685914
rect 400864 685850 400916 685856
rect 399372 664686 399524 664714
rect 379716 664006 380052 664034
rect 389712 664006 390048 664034
rect 379612 662380 379664 662386
rect 379612 662322 379664 662328
rect 379716 662318 379744 664006
rect 390020 662318 390048 664006
rect 400876 662318 400904 685850
rect 408052 683876 408080 686054
rect 417700 686044 417752 686050
rect 417700 685986 417752 685992
rect 417712 683876 417740 685986
rect 428556 685976 428608 685982
rect 428556 685918 428608 685924
rect 427360 685908 427412 685914
rect 427360 685850 427412 685856
rect 428464 685908 428516 685914
rect 428464 685850 428516 685856
rect 427372 683876 427400 685850
rect 401600 683256 401652 683262
rect 401600 683198 401652 683204
rect 401612 673577 401640 683198
rect 405646 674248 405702 674257
rect 405646 674183 405702 674192
rect 401598 673568 401654 673577
rect 401598 673503 401654 673512
rect 405660 665174 405688 674183
rect 405648 665168 405700 665174
rect 405648 665110 405700 665116
rect 427728 665100 427780 665106
rect 427728 665042 427780 665048
rect 427740 664714 427768 665042
rect 427386 664686 427768 664714
rect 408052 662386 408080 664020
rect 408040 662380 408092 662386
rect 408040 662322 408092 662328
rect 417712 662318 417740 664020
rect 428476 662318 428504 685850
rect 428568 665106 428596 685918
rect 428660 665854 428688 686054
rect 428648 665848 428700 665854
rect 428648 665790 428700 665796
rect 428556 665100 428608 665106
rect 428556 665042 428608 665048
rect 379704 662312 379756 662318
rect 379704 662254 379756 662260
rect 390008 662312 390060 662318
rect 390008 662254 390060 662260
rect 400864 662312 400916 662318
rect 400864 662254 400916 662260
rect 417700 662312 417752 662318
rect 417700 662254 417752 662260
rect 428464 662312 428516 662318
rect 428464 662254 428516 662260
rect 379612 658436 379664 658442
rect 379612 658378 379664 658384
rect 418252 658436 418304 658442
rect 418252 658378 418304 658384
rect 379624 654134 379652 658378
rect 390284 658368 390336 658374
rect 390284 658310 390336 658316
rect 400864 658368 400916 658374
rect 400864 658310 400916 658316
rect 408592 658368 408644 658374
rect 408592 658310 408644 658316
rect 380624 658300 380676 658306
rect 380624 658242 380676 658248
rect 380636 656948 380664 658242
rect 390296 656948 390324 658310
rect 399970 656254 400352 656282
rect 400324 655246 400352 656254
rect 400312 655240 400364 655246
rect 400312 655182 400364 655188
rect 379624 654106 380296 654134
rect 380268 637786 380296 654106
rect 380268 637758 380650 637786
rect 390296 634710 390324 637092
rect 399956 634778 399984 637092
rect 399944 634772 399996 634778
rect 399944 634714 399996 634720
rect 400876 634710 400904 658310
rect 408604 656948 408632 658310
rect 418264 656948 418292 658378
rect 428464 658300 428516 658306
rect 428464 658242 428516 658248
rect 427938 656254 428136 656282
rect 401600 655716 401652 655722
rect 401600 655658 401652 655664
rect 400956 655240 401008 655246
rect 400956 655182 401008 655188
rect 400968 634778 400996 655182
rect 401612 646785 401640 655658
rect 408408 655580 408460 655586
rect 408408 655522 408460 655528
rect 408420 648009 408448 655522
rect 408406 648000 408462 648009
rect 408406 647935 408462 647944
rect 401598 646776 401654 646785
rect 401598 646711 401654 646720
rect 400956 634772 401008 634778
rect 400956 634714 401008 634720
rect 408604 634710 408632 637092
rect 390284 634704 390336 634710
rect 390284 634646 390336 634652
rect 400864 634704 400916 634710
rect 400864 634646 400916 634652
rect 408592 634704 408644 634710
rect 408592 634646 408644 634652
rect 418264 634642 418292 637092
rect 427924 634778 427952 637092
rect 428108 634778 428136 656254
rect 427912 634772 427964 634778
rect 427912 634714 427964 634720
rect 428096 634772 428148 634778
rect 428096 634714 428148 634720
rect 428476 634710 428504 658242
rect 428464 634704 428516 634710
rect 428464 634646 428516 634652
rect 418252 634636 418304 634642
rect 418252 634578 418304 634584
rect 408040 632324 408092 632330
rect 408040 632266 408092 632272
rect 428648 632324 428700 632330
rect 428648 632266 428700 632272
rect 389364 632256 389416 632262
rect 389364 632198 389416 632204
rect 399484 632256 399536 632262
rect 399484 632198 399536 632204
rect 389376 629898 389404 632198
rect 399024 632120 399076 632126
rect 399024 632062 399076 632068
rect 399036 629898 399064 632062
rect 389376 629870 389712 629898
rect 399036 629870 399372 629898
rect 379624 629326 380052 629354
rect 379624 608598 379652 629326
rect 399496 610722 399524 632198
rect 400864 632120 400916 632126
rect 400864 632062 400916 632068
rect 399372 610694 399524 610722
rect 379716 610014 380052 610042
rect 389712 610014 390048 610042
rect 379612 608592 379664 608598
rect 379612 608534 379664 608540
rect 379716 608530 379744 610014
rect 390020 608530 390048 610014
rect 400876 608530 400904 632062
rect 408052 629884 408080 632266
rect 417700 632256 417752 632262
rect 417700 632198 417752 632204
rect 417712 629884 417740 632198
rect 428464 632188 428516 632194
rect 428464 632130 428516 632136
rect 427360 632120 427412 632126
rect 427360 632062 427412 632068
rect 427372 629884 427400 632062
rect 405646 620256 405702 620265
rect 405646 620191 405702 620200
rect 401598 619576 401654 619585
rect 401598 619511 401654 619520
rect 401612 611182 401640 619511
rect 405660 611318 405688 620191
rect 428476 615494 428504 632130
rect 428556 632120 428608 632126
rect 428556 632062 428608 632068
rect 427832 615466 428504 615494
rect 405648 611312 405700 611318
rect 405648 611254 405700 611260
rect 401600 611176 401652 611182
rect 401600 611118 401652 611124
rect 427832 610722 427860 615466
rect 427386 610694 427860 610722
rect 408052 608598 408080 610028
rect 408040 608592 408092 608598
rect 408040 608534 408092 608540
rect 417712 608530 417740 610028
rect 428568 608530 428596 632062
rect 428660 612066 428688 632266
rect 428648 612060 428700 612066
rect 428648 612002 428700 612008
rect 379704 608524 379756 608530
rect 379704 608466 379756 608472
rect 390008 608524 390060 608530
rect 390008 608466 390060 608472
rect 400864 608524 400916 608530
rect 400864 608466 400916 608472
rect 417700 608524 417752 608530
rect 417700 608466 417752 608472
rect 428556 608524 428608 608530
rect 428556 608466 428608 608472
rect 379612 604648 379664 604654
rect 379612 604590 379664 604596
rect 418252 604648 418304 604654
rect 418252 604590 418304 604596
rect 379624 596174 379652 604590
rect 390284 604580 390336 604586
rect 390284 604522 390336 604528
rect 400956 604580 401008 604586
rect 400956 604522 401008 604528
rect 408592 604580 408644 604586
rect 408592 604522 408644 604528
rect 380624 604512 380676 604518
rect 380624 604454 380676 604460
rect 380636 602956 380664 604454
rect 390296 602956 390324 604522
rect 399970 602262 400904 602290
rect 379624 596146 380296 596174
rect 380268 583794 380296 596146
rect 380268 583766 380650 583794
rect 390296 580922 390324 583100
rect 399956 580990 399984 583100
rect 400876 580990 400904 602262
rect 399944 580984 399996 580990
rect 399944 580926 399996 580932
rect 400864 580984 400916 580990
rect 400864 580926 400916 580932
rect 400968 580922 400996 604522
rect 408604 602956 408632 604522
rect 418264 602956 418292 604590
rect 428464 604512 428516 604518
rect 428464 604454 428516 604460
rect 427938 602262 428136 602290
rect 401600 601860 401652 601866
rect 401600 601802 401652 601808
rect 401612 592793 401640 601802
rect 405648 601724 405700 601730
rect 405648 601666 405700 601672
rect 405660 593473 405688 601666
rect 405646 593464 405702 593473
rect 405646 593399 405702 593408
rect 401598 592784 401654 592793
rect 401598 592719 401654 592728
rect 408604 580922 408632 583100
rect 390284 580916 390336 580922
rect 390284 580858 390336 580864
rect 400956 580916 401008 580922
rect 400956 580858 401008 580864
rect 408592 580916 408644 580922
rect 408592 580858 408644 580864
rect 418264 580854 418292 583100
rect 427924 580990 427952 583100
rect 428108 580990 428136 602262
rect 427912 580984 427964 580990
rect 427912 580926 427964 580932
rect 428096 580984 428148 580990
rect 428096 580926 428148 580932
rect 428476 580922 428504 604454
rect 428464 580916 428516 580922
rect 428464 580858 428516 580864
rect 418252 580848 418304 580854
rect 418252 580790 418304 580796
rect 408040 578468 408092 578474
rect 408040 578410 408092 578416
rect 428648 578468 428700 578474
rect 428648 578410 428700 578416
rect 389364 578400 389416 578406
rect 389364 578342 389416 578348
rect 399484 578400 399536 578406
rect 399484 578342 399536 578348
rect 389376 575906 389404 578342
rect 399024 578264 399076 578270
rect 399024 578206 399076 578212
rect 399036 575906 399064 578206
rect 389376 575878 389712 575906
rect 399036 575878 399372 575906
rect 379624 575334 380052 575362
rect 379624 554674 379652 575334
rect 399496 556730 399524 578342
rect 400864 578264 400916 578270
rect 400864 578206 400916 578212
rect 399372 556702 399524 556730
rect 379716 556022 380052 556050
rect 389712 556022 390048 556050
rect 379716 554742 379744 556022
rect 379704 554736 379756 554742
rect 379704 554678 379756 554684
rect 390020 554674 390048 556022
rect 400876 554674 400904 578206
rect 408052 575892 408080 578410
rect 417700 578400 417752 578406
rect 417700 578342 417752 578348
rect 417712 575892 417740 578342
rect 428464 578332 428516 578338
rect 428464 578274 428516 578280
rect 427360 578264 427412 578270
rect 427360 578206 427412 578212
rect 427372 575892 427400 578206
rect 405646 566264 405702 566273
rect 405646 566199 405702 566208
rect 401598 565584 401654 565593
rect 401598 565519 401654 565528
rect 401612 557394 401640 565519
rect 405660 557530 405688 566199
rect 428476 557534 428504 578274
rect 428556 578264 428608 578270
rect 428556 578206 428608 578212
rect 405648 557524 405700 557530
rect 405648 557466 405700 557472
rect 427832 557506 428504 557534
rect 401600 557388 401652 557394
rect 401600 557330 401652 557336
rect 427832 556730 427860 557506
rect 427386 556702 427860 556730
rect 408052 554742 408080 556036
rect 408040 554736 408092 554742
rect 408040 554678 408092 554684
rect 417712 554674 417740 556036
rect 428568 554674 428596 578206
rect 428660 558210 428688 578410
rect 428648 558204 428700 558210
rect 428648 558146 428700 558152
rect 379612 554668 379664 554674
rect 379612 554610 379664 554616
rect 390008 554668 390060 554674
rect 390008 554610 390060 554616
rect 400864 554668 400916 554674
rect 400864 554610 400916 554616
rect 417700 554668 417752 554674
rect 417700 554610 417752 554616
rect 428556 554668 428608 554674
rect 428556 554610 428608 554616
rect 379612 550792 379664 550798
rect 379612 550734 379664 550740
rect 418252 550792 418304 550798
rect 418252 550734 418304 550740
rect 379624 538214 379652 550734
rect 390284 550724 390336 550730
rect 390284 550666 390336 550672
rect 400956 550724 401008 550730
rect 400956 550666 401008 550672
rect 408592 550724 408644 550730
rect 408592 550666 408644 550672
rect 380624 550656 380676 550662
rect 380624 550598 380676 550604
rect 380636 548964 380664 550598
rect 390296 548964 390324 550666
rect 399970 548270 400904 548298
rect 379624 538186 380296 538214
rect 380268 529666 380296 538186
rect 380268 529638 380650 529666
rect 390296 527066 390324 529108
rect 399956 527134 399984 529108
rect 400876 527134 400904 548270
rect 399944 527128 399996 527134
rect 399944 527070 399996 527076
rect 400864 527128 400916 527134
rect 400864 527070 400916 527076
rect 400968 527066 400996 550666
rect 408604 548964 408632 550666
rect 418264 548964 418292 550734
rect 428464 550656 428516 550662
rect 428464 550598 428516 550604
rect 427938 548270 428136 548298
rect 405646 539472 405702 539481
rect 405646 539407 405702 539416
rect 401598 538792 401654 538801
rect 401598 538727 401654 538736
rect 401612 529786 401640 538727
rect 405660 529922 405688 539407
rect 405648 529916 405700 529922
rect 405648 529858 405700 529864
rect 401600 529780 401652 529786
rect 401600 529722 401652 529728
rect 408604 527066 408632 529108
rect 390284 527060 390336 527066
rect 390284 527002 390336 527008
rect 400956 527060 401008 527066
rect 400956 527002 401008 527008
rect 408592 527060 408644 527066
rect 408592 527002 408644 527008
rect 418264 526998 418292 529108
rect 427924 527134 427952 529108
rect 428108 527134 428136 548270
rect 427912 527128 427964 527134
rect 427912 527070 427964 527076
rect 428096 527128 428148 527134
rect 428096 527070 428148 527076
rect 428476 527066 428504 550598
rect 428464 527060 428516 527066
rect 428464 527002 428516 527008
rect 418252 526992 418304 526998
rect 418252 526934 418304 526940
rect 408040 523252 408092 523258
rect 408040 523194 408092 523200
rect 428648 523252 428700 523258
rect 428648 523194 428700 523200
rect 389364 523184 389416 523190
rect 389364 523126 389416 523132
rect 399484 523184 399536 523190
rect 399484 523126 399536 523132
rect 389376 521914 389404 523126
rect 399024 523048 399076 523054
rect 399024 522990 399076 522996
rect 399036 521914 399064 522990
rect 389376 521886 389712 521914
rect 399036 521886 399372 521914
rect 379624 521206 380052 521234
rect 379624 500954 379652 521206
rect 399496 502738 399524 523126
rect 400864 523048 400916 523054
rect 400864 522990 400916 522996
rect 399372 502710 399524 502738
rect 379716 502030 380052 502058
rect 389712 502030 390048 502058
rect 379612 500948 379664 500954
rect 379612 500890 379664 500896
rect 379716 500886 379744 502030
rect 390020 500886 390048 502030
rect 400876 500886 400904 522990
rect 408052 521900 408080 523194
rect 417700 523184 417752 523190
rect 417700 523126 417752 523132
rect 417712 521900 417740 523126
rect 428464 523116 428516 523122
rect 428464 523058 428516 523064
rect 427360 523048 427412 523054
rect 427360 522990 427412 522996
rect 427372 521900 427400 522990
rect 405646 512272 405702 512281
rect 405646 512207 405702 512216
rect 401598 511592 401654 511601
rect 401598 511527 401654 511536
rect 401612 503674 401640 511527
rect 405660 503674 405688 512207
rect 428476 509234 428504 523058
rect 428556 523048 428608 523054
rect 428556 522990 428608 522996
rect 427832 509206 428504 509234
rect 401600 503668 401652 503674
rect 401600 503610 401652 503616
rect 405648 503668 405700 503674
rect 405648 503610 405700 503616
rect 427832 502738 427860 509206
rect 427386 502710 427860 502738
rect 408052 500954 408080 502044
rect 408040 500948 408092 500954
rect 408040 500890 408092 500896
rect 417712 500886 417740 502044
rect 428568 500886 428596 522990
rect 428660 504422 428688 523194
rect 428648 504416 428700 504422
rect 428648 504358 428700 504364
rect 379704 500880 379756 500886
rect 379704 500822 379756 500828
rect 390008 500880 390060 500886
rect 390008 500822 390060 500828
rect 400864 500880 400916 500886
rect 400864 500822 400916 500828
rect 417700 500880 417752 500886
rect 417700 500822 417752 500828
rect 428556 500880 428608 500886
rect 428556 500822 428608 500828
rect 380256 497004 380308 497010
rect 380256 496946 380308 496952
rect 418252 497004 418304 497010
rect 418252 496946 418304 496952
rect 380268 475674 380296 496946
rect 390284 496936 390336 496942
rect 390284 496878 390336 496884
rect 400956 496936 401008 496942
rect 400956 496878 401008 496884
rect 408592 496936 408644 496942
rect 408592 496878 408644 496884
rect 380624 496868 380676 496874
rect 380624 496810 380676 496816
rect 380636 494972 380664 496810
rect 390296 494972 390324 496878
rect 399970 494278 400904 494306
rect 380268 475646 380650 475674
rect 390296 473278 390324 475116
rect 399956 473346 399984 475116
rect 400876 473346 400904 494278
rect 399944 473340 399996 473346
rect 399944 473282 399996 473288
rect 400864 473340 400916 473346
rect 400864 473282 400916 473288
rect 400968 473278 400996 496878
rect 408604 494972 408632 496878
rect 418264 494972 418292 496946
rect 428464 496868 428516 496874
rect 428464 496810 428516 496816
rect 427938 494278 428136 494306
rect 405646 485480 405702 485489
rect 405646 485415 405702 485424
rect 401598 484800 401654 484809
rect 401598 484735 401654 484744
rect 401612 475930 401640 484735
rect 405660 476066 405688 485415
rect 405648 476060 405700 476066
rect 405648 476002 405700 476008
rect 401600 475924 401652 475930
rect 401600 475866 401652 475872
rect 408604 473278 408632 475116
rect 390284 473272 390336 473278
rect 390284 473214 390336 473220
rect 400956 473272 401008 473278
rect 400956 473214 401008 473220
rect 408592 473272 408644 473278
rect 408592 473214 408644 473220
rect 418264 473210 418292 475116
rect 427924 473346 427952 475116
rect 428108 473346 428136 494278
rect 427912 473340 427964 473346
rect 427912 473282 427964 473288
rect 428096 473340 428148 473346
rect 428096 473282 428148 473288
rect 428476 473278 428504 496810
rect 428464 473272 428516 473278
rect 428464 473214 428516 473220
rect 418252 473204 418304 473210
rect 418252 473146 418304 473152
rect 408040 469464 408092 469470
rect 408040 469406 408092 469412
rect 428648 469464 428700 469470
rect 428648 469406 428700 469412
rect 389364 469396 389416 469402
rect 389364 469338 389416 469344
rect 399484 469396 399536 469402
rect 399484 469338 399536 469344
rect 389376 467922 389404 469338
rect 399024 469260 399076 469266
rect 399024 469202 399076 469208
rect 399036 467922 399064 469202
rect 389376 467894 389712 467922
rect 399036 467894 399372 467922
rect 379624 467214 380052 467242
rect 379624 445738 379652 467214
rect 399496 448746 399524 469338
rect 400864 469260 400916 469266
rect 400864 469202 400916 469208
rect 399372 448718 399524 448746
rect 379716 448038 380052 448066
rect 389712 448038 390048 448066
rect 379612 445732 379664 445738
rect 379612 445674 379664 445680
rect 379716 445670 379744 448038
rect 390020 445670 390048 448038
rect 400876 445670 400904 469202
rect 408052 467908 408080 469406
rect 417700 469396 417752 469402
rect 417700 469338 417752 469344
rect 417712 467908 417740 469338
rect 428464 469328 428516 469334
rect 428464 469270 428516 469276
rect 427360 469260 427412 469266
rect 427360 469202 427412 469208
rect 427372 467908 427400 469202
rect 401600 466608 401652 466614
rect 401600 466550 401652 466556
rect 401612 457609 401640 466550
rect 405648 466472 405700 466478
rect 405648 466414 405700 466420
rect 405660 458289 405688 466414
rect 405646 458280 405702 458289
rect 405646 458215 405702 458224
rect 401598 457600 401654 457609
rect 401598 457535 401654 457544
rect 428476 451274 428504 469270
rect 428556 469260 428608 469266
rect 428556 469202 428608 469208
rect 427832 451246 428504 451274
rect 427832 448474 427860 451246
rect 427386 448446 427860 448474
rect 408052 445738 408080 448052
rect 408040 445732 408092 445738
rect 408040 445674 408092 445680
rect 417712 445670 417740 448052
rect 428568 445670 428596 469202
rect 428660 450566 428688 469406
rect 428648 450560 428700 450566
rect 428648 450502 428700 450508
rect 379704 445664 379756 445670
rect 379704 445606 379756 445612
rect 390008 445664 390060 445670
rect 390008 445606 390060 445612
rect 400864 445664 400916 445670
rect 400864 445606 400916 445612
rect 417700 445664 417752 445670
rect 417700 445606 417752 445612
rect 428556 445664 428608 445670
rect 428556 445606 428608 445612
rect 379612 443148 379664 443154
rect 379612 443090 379664 443096
rect 418252 443148 418304 443154
rect 418252 443090 418304 443096
rect 379624 441614 379652 443090
rect 390284 443080 390336 443086
rect 390284 443022 390336 443028
rect 400864 443080 400916 443086
rect 400864 443022 400916 443028
rect 408592 443080 408644 443086
rect 408592 443022 408644 443028
rect 380624 443012 380676 443018
rect 380624 442954 380676 442960
rect 379624 441586 380296 441614
rect 380268 421682 380296 441586
rect 380636 440980 380664 442954
rect 390296 440980 390324 443022
rect 399970 440286 400352 440314
rect 400324 436150 400352 440286
rect 400312 436144 400364 436150
rect 400312 436086 400364 436092
rect 380268 421654 380650 421682
rect 390296 419422 390324 421124
rect 399956 419490 399984 421124
rect 399944 419484 399996 419490
rect 399944 419426 399996 419432
rect 400876 419422 400904 443022
rect 408604 440980 408632 443022
rect 418264 440980 418292 443090
rect 428464 443012 428516 443018
rect 428464 442954 428516 442960
rect 427938 440286 428136 440314
rect 400956 436144 401008 436150
rect 400956 436086 401008 436092
rect 400968 419490 400996 436086
rect 405646 431488 405702 431497
rect 405646 431423 405702 431432
rect 401598 430808 401654 430817
rect 401598 430743 401654 430752
rect 401612 422278 401640 430743
rect 405660 422278 405688 431423
rect 401600 422272 401652 422278
rect 401600 422214 401652 422220
rect 405648 422272 405700 422278
rect 405648 422214 405700 422220
rect 400956 419484 401008 419490
rect 400956 419426 401008 419432
rect 408604 419422 408632 421124
rect 390284 419416 390336 419422
rect 390284 419358 390336 419364
rect 400864 419416 400916 419422
rect 400864 419358 400916 419364
rect 408592 419416 408644 419422
rect 408592 419358 408644 419364
rect 418264 419354 418292 421124
rect 427924 419490 427952 421124
rect 428108 419490 428136 440286
rect 427912 419484 427964 419490
rect 427912 419426 427964 419432
rect 428096 419484 428148 419490
rect 428096 419426 428148 419432
rect 428476 419422 428504 442954
rect 428464 419416 428516 419422
rect 428464 419358 428516 419364
rect 418252 419348 418304 419354
rect 418252 419290 418304 419296
rect 408040 415676 408092 415682
rect 408040 415618 408092 415624
rect 428648 415676 428700 415682
rect 428648 415618 428700 415624
rect 389364 415608 389416 415614
rect 389364 415550 389416 415556
rect 399484 415608 399536 415614
rect 399484 415550 399536 415556
rect 389376 413930 389404 415550
rect 399024 415472 399076 415478
rect 399024 415414 399076 415420
rect 399036 413930 399064 415414
rect 389376 413902 389712 413930
rect 399036 413902 399372 413930
rect 379624 413222 380052 413250
rect 379624 391950 379652 413222
rect 399496 394754 399524 415550
rect 400864 415472 400916 415478
rect 400864 415414 400916 415420
rect 399372 394726 399524 394754
rect 379716 394046 380052 394074
rect 389712 394046 390048 394074
rect 379612 391944 379664 391950
rect 379612 391886 379664 391892
rect 379716 391882 379744 394046
rect 390020 391882 390048 394046
rect 400876 391882 400904 415414
rect 408052 413916 408080 415618
rect 417700 415608 417752 415614
rect 417700 415550 417752 415556
rect 417712 413916 417740 415550
rect 428464 415540 428516 415546
rect 428464 415482 428516 415488
rect 427360 415472 427412 415478
rect 427360 415414 427412 415420
rect 427372 413916 427400 415414
rect 405646 404288 405702 404297
rect 405646 404223 405702 404232
rect 401598 403608 401654 403617
rect 401598 403543 401654 403552
rect 401612 394534 401640 403543
rect 405660 394670 405688 404223
rect 428476 402974 428504 415482
rect 428556 415472 428608 415478
rect 428556 415414 428608 415420
rect 427832 402946 428504 402974
rect 405648 394664 405700 394670
rect 427832 394618 427860 402946
rect 405648 394606 405700 394612
rect 427386 394590 427860 394618
rect 401600 394528 401652 394534
rect 401600 394470 401652 394476
rect 408052 391950 408080 394060
rect 408040 391944 408092 391950
rect 408040 391886 408092 391892
rect 417712 391882 417740 394060
rect 428568 391882 428596 415414
rect 428660 395350 428688 415618
rect 428648 395344 428700 395350
rect 428648 395286 428700 395292
rect 379704 391876 379756 391882
rect 379704 391818 379756 391824
rect 390008 391876 390060 391882
rect 390008 391818 390060 391824
rect 400864 391876 400916 391882
rect 400864 391818 400916 391824
rect 417700 391876 417752 391882
rect 417700 391818 417752 391824
rect 428556 391876 428608 391882
rect 428556 391818 428608 391824
rect 379612 389360 379664 389366
rect 379612 389302 379664 389308
rect 418252 389360 418304 389366
rect 418252 389302 418304 389308
rect 379624 383654 379652 389302
rect 390284 389292 390336 389298
rect 390284 389234 390336 389240
rect 400956 389292 401008 389298
rect 400956 389234 401008 389240
rect 408592 389292 408644 389298
rect 408592 389234 408644 389240
rect 380624 389224 380676 389230
rect 380624 389166 380676 389172
rect 380636 386852 380664 389166
rect 390296 386852 390324 389234
rect 399970 386430 400904 386458
rect 379624 383626 380296 383654
rect 380268 367690 380296 383626
rect 380268 367662 380650 367690
rect 390296 365634 390324 367132
rect 399956 365702 399984 367132
rect 400876 365702 400904 386430
rect 399944 365696 399996 365702
rect 399944 365638 399996 365644
rect 400864 365696 400916 365702
rect 400864 365638 400916 365644
rect 400968 365634 400996 389234
rect 408604 386852 408632 389234
rect 418264 386852 418292 389302
rect 428464 389224 428516 389230
rect 428464 389166 428516 389172
rect 401600 386572 401652 386578
rect 401600 386514 401652 386520
rect 401612 376825 401640 386514
rect 405648 386436 405700 386442
rect 405648 386378 405700 386384
rect 405660 377505 405688 386378
rect 427938 386294 428136 386322
rect 405646 377496 405702 377505
rect 405646 377431 405702 377440
rect 401598 376816 401654 376825
rect 401598 376751 401654 376760
rect 408604 365634 408632 367132
rect 390284 365628 390336 365634
rect 390284 365570 390336 365576
rect 400956 365628 401008 365634
rect 400956 365570 401008 365576
rect 408592 365628 408644 365634
rect 408592 365570 408644 365576
rect 418264 365566 418292 367132
rect 427924 365702 427952 367132
rect 428108 365702 428136 386294
rect 427912 365696 427964 365702
rect 427912 365638 427964 365644
rect 428096 365696 428148 365702
rect 428096 365638 428148 365644
rect 428476 365634 428504 389166
rect 428464 365628 428516 365634
rect 428464 365570 428516 365576
rect 418252 365560 418304 365566
rect 418252 365502 418304 365508
rect 389364 361752 389416 361758
rect 389364 361694 389416 361700
rect 399484 361752 399536 361758
rect 399484 361694 399536 361700
rect 417700 361752 417752 361758
rect 417700 361694 417752 361700
rect 428464 361752 428516 361758
rect 428464 361694 428516 361700
rect 389376 359938 389404 361694
rect 399024 361616 399076 361622
rect 399024 361558 399076 361564
rect 399036 359938 399064 361558
rect 389376 359910 389712 359938
rect 399036 359910 399372 359938
rect 379624 359230 380052 359258
rect 379624 338026 379652 359230
rect 399496 340762 399524 361694
rect 408040 361684 408092 361690
rect 408040 361626 408092 361632
rect 400864 361616 400916 361622
rect 400864 361558 400916 361564
rect 399372 340734 399524 340762
rect 379716 340054 380052 340082
rect 389712 340054 390048 340082
rect 379716 338094 379744 340054
rect 379704 338088 379756 338094
rect 379704 338030 379756 338036
rect 390020 338026 390048 340054
rect 400876 338026 400904 361558
rect 408052 359924 408080 361626
rect 417712 359924 417740 361694
rect 427360 361616 427412 361622
rect 427360 361558 427412 361564
rect 427372 359924 427400 361558
rect 405646 350296 405702 350305
rect 405646 350231 405702 350240
rect 401598 349616 401654 349625
rect 401598 349551 401654 349560
rect 401612 340746 401640 349551
rect 405660 340882 405688 350231
rect 428476 345014 428504 361694
rect 428648 361684 428700 361690
rect 428648 361626 428700 361632
rect 428556 361616 428608 361622
rect 428556 361558 428608 361564
rect 427832 344986 428504 345014
rect 405648 340876 405700 340882
rect 405648 340818 405700 340824
rect 427832 340762 427860 344986
rect 401600 340740 401652 340746
rect 427386 340734 427860 340762
rect 401600 340682 401652 340688
rect 408052 338094 408080 340068
rect 408040 338088 408092 338094
rect 408040 338030 408092 338036
rect 417712 338026 417740 340068
rect 428568 338026 428596 361558
rect 428660 341562 428688 361626
rect 428648 341556 428700 341562
rect 428648 341498 428700 341504
rect 379612 338020 379664 338026
rect 379612 337962 379664 337968
rect 390008 338020 390060 338026
rect 390008 337962 390060 337968
rect 400864 338020 400916 338026
rect 400864 337962 400916 337968
rect 417700 338020 417752 338026
rect 417700 337962 417752 337968
rect 428556 338020 428608 338026
rect 428556 337962 428608 337968
rect 379612 335504 379664 335510
rect 379612 335446 379664 335452
rect 418252 335504 418304 335510
rect 418252 335446 418304 335452
rect 379624 325694 379652 335446
rect 390284 335436 390336 335442
rect 390284 335378 390336 335384
rect 400864 335436 400916 335442
rect 400864 335378 400916 335384
rect 408592 335436 408644 335442
rect 408592 335378 408644 335384
rect 380624 335368 380676 335374
rect 380624 335310 380676 335316
rect 380636 332860 380664 335310
rect 390296 332860 390324 335378
rect 399970 332302 400352 332330
rect 400324 329050 400352 332302
rect 400312 329044 400364 329050
rect 400312 328986 400364 328992
rect 379624 325666 380296 325694
rect 380268 313698 380296 325666
rect 380268 313670 380650 313698
rect 390296 311778 390324 313140
rect 399956 311846 399984 313140
rect 399944 311840 399996 311846
rect 399944 311782 399996 311788
rect 400876 311778 400904 335378
rect 408604 332860 408632 335378
rect 418264 332860 418292 335446
rect 428464 335368 428516 335374
rect 428464 335310 428516 335316
rect 427938 332302 428136 332330
rect 405648 331288 405700 331294
rect 405648 331230 405700 331236
rect 400956 329044 401008 329050
rect 400956 328986 401008 328992
rect 400968 311846 400996 328986
rect 405660 324057 405688 331230
rect 405646 324048 405702 324057
rect 405646 323983 405702 323992
rect 401598 322144 401654 322153
rect 401598 322079 401654 322088
rect 401612 314566 401640 322079
rect 401600 314560 401652 314566
rect 401600 314502 401652 314508
rect 400956 311840 401008 311846
rect 400956 311782 401008 311788
rect 408604 311778 408632 313140
rect 390284 311772 390336 311778
rect 390284 311714 390336 311720
rect 400864 311772 400916 311778
rect 400864 311714 400916 311720
rect 408592 311772 408644 311778
rect 408592 311714 408644 311720
rect 418264 311710 418292 313140
rect 427924 311846 427952 313140
rect 428108 311846 428136 332302
rect 427912 311840 427964 311846
rect 427912 311782 427964 311788
rect 428096 311840 428148 311846
rect 428096 311782 428148 311788
rect 428476 311778 428504 335310
rect 428464 311772 428516 311778
rect 428464 311714 428516 311720
rect 418252 311704 418304 311710
rect 418252 311646 418304 311652
rect 408040 308032 408092 308038
rect 408040 307974 408092 307980
rect 428648 308032 428700 308038
rect 428648 307974 428700 307980
rect 389364 307964 389416 307970
rect 389364 307906 389416 307912
rect 399484 307964 399536 307970
rect 399484 307906 399536 307912
rect 389376 305946 389404 307906
rect 399024 307828 399076 307834
rect 399024 307770 399076 307776
rect 399036 305946 399064 307770
rect 389376 305918 389712 305946
rect 399036 305918 399372 305946
rect 379624 305238 380052 305266
rect 379624 284238 379652 305238
rect 399496 286770 399524 307906
rect 400864 307828 400916 307834
rect 400864 307770 400916 307776
rect 399372 286742 399524 286770
rect 379716 286062 380052 286090
rect 389712 286062 390048 286090
rect 379716 284306 379744 286062
rect 379704 284300 379756 284306
rect 379704 284242 379756 284248
rect 390020 284238 390048 286062
rect 400876 284238 400904 307770
rect 408052 305932 408080 307974
rect 417700 307964 417752 307970
rect 417700 307906 417752 307912
rect 417712 305932 417740 307906
rect 428556 307896 428608 307902
rect 428556 307838 428608 307844
rect 427360 307828 427412 307834
rect 427360 307770 427412 307776
rect 428464 307828 428516 307834
rect 428464 307770 428516 307776
rect 427372 305932 427400 307770
rect 405646 296304 405702 296313
rect 405646 296239 405702 296248
rect 401598 295624 401654 295633
rect 401598 295559 401654 295568
rect 401612 286890 401640 295559
rect 405660 287026 405688 296239
rect 405648 287020 405700 287026
rect 405648 286962 405700 286968
rect 401600 286884 401652 286890
rect 401600 286826 401652 286832
rect 427728 286816 427780 286822
rect 427386 286764 427728 286770
rect 427386 286758 427780 286764
rect 427386 286742 427768 286758
rect 408052 284306 408080 286076
rect 408040 284300 408092 284306
rect 408040 284242 408092 284248
rect 417712 284238 417740 286076
rect 428476 284238 428504 307770
rect 428568 286822 428596 307838
rect 428660 287706 428688 307974
rect 428648 287700 428700 287706
rect 428648 287642 428700 287648
rect 428556 286816 428608 286822
rect 428556 286758 428608 286764
rect 379612 284232 379664 284238
rect 379612 284174 379664 284180
rect 390008 284232 390060 284238
rect 390008 284174 390060 284180
rect 400864 284232 400916 284238
rect 400864 284174 400916 284180
rect 417700 284232 417752 284238
rect 417700 284174 417752 284180
rect 428464 284232 428516 284238
rect 428464 284174 428516 284180
rect 379612 280356 379664 280362
rect 379612 280298 379664 280304
rect 418252 280356 418304 280362
rect 418252 280298 418304 280304
rect 379624 267734 379652 280298
rect 390284 280288 390336 280294
rect 390284 280230 390336 280236
rect 400864 280288 400916 280294
rect 400864 280230 400916 280236
rect 408592 280288 408644 280294
rect 408592 280230 408644 280236
rect 380624 280220 380676 280226
rect 380624 280162 380676 280168
rect 380636 278868 380664 280162
rect 390296 278868 390324 280230
rect 399970 278310 400352 278338
rect 400324 272610 400352 278310
rect 400312 272604 400364 272610
rect 400312 272546 400364 272552
rect 379624 267706 380296 267734
rect 380268 259706 380296 267706
rect 380268 259678 380650 259706
rect 390296 256630 390324 259148
rect 399956 256698 399984 259148
rect 399944 256692 399996 256698
rect 399944 256634 399996 256640
rect 400876 256630 400904 280230
rect 408604 278868 408632 280230
rect 418264 278868 418292 280298
rect 428464 280220 428516 280226
rect 428464 280162 428516 280168
rect 427938 278310 428136 278338
rect 401600 277432 401652 277438
rect 401600 277374 401652 277380
rect 405648 277432 405700 277438
rect 405648 277374 405700 277380
rect 400956 272604 401008 272610
rect 400956 272546 401008 272552
rect 400968 256698 400996 272546
rect 401612 269113 401640 277374
rect 405660 270065 405688 277374
rect 405646 270056 405702 270065
rect 405646 269991 405702 270000
rect 401598 269104 401654 269113
rect 401598 269039 401654 269048
rect 400956 256692 401008 256698
rect 400956 256634 401008 256640
rect 408604 256630 408632 259148
rect 390284 256624 390336 256630
rect 390284 256566 390336 256572
rect 400864 256624 400916 256630
rect 400864 256566 400916 256572
rect 408592 256624 408644 256630
rect 408592 256566 408644 256572
rect 418264 256562 418292 259148
rect 427924 256698 427952 259148
rect 428108 256698 428136 278310
rect 427912 256692 427964 256698
rect 427912 256634 427964 256640
rect 428096 256692 428148 256698
rect 428096 256634 428148 256640
rect 428476 256630 428504 280162
rect 428464 256624 428516 256630
rect 428464 256566 428516 256572
rect 418252 256556 418304 256562
rect 418252 256498 418304 256504
rect 408040 254176 408092 254182
rect 408040 254118 408092 254124
rect 428648 254176 428700 254182
rect 428648 254118 428700 254124
rect 389364 254108 389416 254114
rect 389364 254050 389416 254056
rect 399484 254108 399536 254114
rect 399484 254050 399536 254056
rect 389376 251954 389404 254050
rect 399024 253972 399076 253978
rect 399024 253914 399076 253920
rect 399036 251954 399064 253914
rect 389376 251926 389712 251954
rect 399036 251926 399372 251954
rect 379624 251246 380052 251274
rect 379624 230450 379652 251246
rect 399496 232778 399524 254050
rect 400864 253972 400916 253978
rect 400864 253914 400916 253920
rect 399372 232750 399524 232778
rect 379716 232070 380052 232098
rect 389712 232070 390048 232098
rect 379612 230444 379664 230450
rect 379612 230386 379664 230392
rect 379716 230382 379744 232070
rect 390020 230382 390048 232070
rect 400876 230382 400904 253914
rect 408052 251940 408080 254118
rect 417700 254108 417752 254114
rect 417700 254050 417752 254056
rect 417712 251940 417740 254050
rect 428556 254040 428608 254046
rect 428556 253982 428608 253988
rect 427360 253972 427412 253978
rect 427360 253914 427412 253920
rect 428464 253972 428516 253978
rect 428464 253914 428516 253920
rect 427372 251940 427400 253914
rect 401600 251388 401652 251394
rect 401600 251330 401652 251336
rect 401612 241641 401640 251330
rect 405648 251252 405700 251258
rect 405648 251194 405700 251200
rect 405660 242321 405688 251194
rect 405646 242312 405702 242321
rect 405646 242247 405702 242256
rect 401598 241632 401654 241641
rect 401598 241567 401654 241576
rect 427728 233232 427780 233238
rect 427728 233174 427780 233180
rect 427740 232778 427768 233174
rect 427386 232750 427768 232778
rect 408052 230450 408080 232084
rect 408040 230444 408092 230450
rect 408040 230386 408092 230392
rect 417712 230382 417740 232084
rect 428476 230382 428504 253914
rect 428568 233238 428596 253982
rect 428660 233918 428688 254118
rect 428648 233912 428700 233918
rect 428648 233854 428700 233860
rect 428556 233232 428608 233238
rect 428556 233174 428608 233180
rect 379704 230376 379756 230382
rect 379704 230318 379756 230324
rect 390008 230376 390060 230382
rect 390008 230318 390060 230324
rect 400864 230376 400916 230382
rect 400864 230318 400916 230324
rect 417700 230376 417752 230382
rect 417700 230318 417752 230324
rect 428464 230376 428516 230382
rect 428464 230318 428516 230324
rect 380256 226500 380308 226506
rect 380256 226442 380308 226448
rect 418252 226500 418304 226506
rect 418252 226442 418304 226448
rect 380268 205714 380296 226442
rect 390284 226432 390336 226438
rect 390284 226374 390336 226380
rect 400956 226432 401008 226438
rect 400956 226374 401008 226380
rect 408592 226432 408644 226438
rect 408592 226374 408644 226380
rect 380624 226364 380676 226370
rect 380624 226306 380676 226312
rect 380636 224876 380664 226306
rect 390296 224876 390324 226374
rect 399970 224318 400904 224346
rect 380268 205686 380650 205714
rect 390296 202774 390324 205020
rect 399956 202842 399984 205020
rect 400876 202842 400904 224318
rect 399944 202836 399996 202842
rect 399944 202778 399996 202784
rect 400864 202836 400916 202842
rect 400864 202778 400916 202784
rect 400968 202774 400996 226374
rect 408604 224876 408632 226374
rect 418264 224876 418292 226442
rect 428464 226364 428516 226370
rect 428464 226306 428516 226312
rect 427938 224318 428136 224346
rect 401600 223780 401652 223786
rect 401600 223722 401652 223728
rect 401612 214713 401640 223722
rect 405648 223644 405700 223650
rect 405648 223586 405700 223592
rect 405660 215393 405688 223586
rect 405646 215384 405702 215393
rect 405646 215319 405702 215328
rect 401598 214704 401654 214713
rect 401598 214639 401654 214648
rect 408604 202774 408632 205020
rect 390284 202768 390336 202774
rect 390284 202710 390336 202716
rect 400956 202768 401008 202774
rect 400956 202710 401008 202716
rect 408592 202768 408644 202774
rect 408592 202710 408644 202716
rect 418264 202706 418292 205020
rect 427924 202842 427952 205020
rect 428108 202842 428136 224318
rect 427912 202836 427964 202842
rect 427912 202778 427964 202784
rect 428096 202836 428148 202842
rect 428096 202778 428148 202784
rect 428476 202774 428504 226306
rect 428464 202768 428516 202774
rect 428464 202710 428516 202716
rect 418252 202700 418304 202706
rect 418252 202642 418304 202648
rect 408040 200388 408092 200394
rect 408040 200330 408092 200336
rect 428648 200388 428700 200394
rect 428648 200330 428700 200336
rect 389364 200320 389416 200326
rect 389364 200262 389416 200268
rect 399484 200320 399536 200326
rect 399484 200262 399536 200268
rect 389376 197962 389404 200262
rect 399024 200184 399076 200190
rect 399024 200126 399076 200132
rect 399036 197962 399064 200126
rect 389376 197934 389712 197962
rect 399036 197934 399372 197962
rect 379624 197254 380052 197282
rect 379624 176594 379652 197254
rect 399496 178786 399524 200262
rect 400864 200184 400916 200190
rect 400864 200126 400916 200132
rect 399372 178758 399524 178786
rect 379716 178078 380052 178106
rect 389712 178078 390048 178106
rect 379716 176662 379744 178078
rect 379704 176656 379756 176662
rect 379704 176598 379756 176604
rect 390020 176594 390048 178078
rect 400876 176594 400904 200126
rect 408052 197948 408080 200330
rect 417700 200320 417752 200326
rect 417700 200262 417752 200268
rect 417712 197948 417740 200262
rect 428464 200252 428516 200258
rect 428464 200194 428516 200200
rect 427360 200184 427412 200190
rect 427360 200126 427412 200132
rect 427372 197948 427400 200126
rect 405646 188320 405702 188329
rect 405646 188255 405702 188264
rect 401598 187640 401654 187649
rect 401598 187575 401654 187584
rect 401612 179246 401640 187575
rect 405660 179382 405688 188255
rect 428476 180794 428504 200194
rect 428556 200184 428608 200190
rect 428556 200126 428608 200132
rect 427832 180766 428504 180794
rect 405648 179376 405700 179382
rect 405648 179318 405700 179324
rect 401600 179240 401652 179246
rect 401600 179182 401652 179188
rect 427832 178786 427860 180766
rect 427386 178758 427860 178786
rect 408052 176662 408080 178092
rect 408040 176656 408092 176662
rect 408040 176598 408092 176604
rect 417712 176594 417740 178092
rect 428568 176594 428596 200126
rect 428660 180130 428688 200330
rect 428648 180124 428700 180130
rect 428648 180066 428700 180072
rect 379612 176588 379664 176594
rect 379612 176530 379664 176536
rect 390008 176588 390060 176594
rect 390008 176530 390060 176536
rect 400864 176588 400916 176594
rect 400864 176530 400916 176536
rect 417700 176588 417752 176594
rect 417700 176530 417752 176536
rect 428556 176588 428608 176594
rect 428556 176530 428608 176536
rect 379612 172712 379664 172718
rect 379612 172654 379664 172660
rect 418252 172712 418304 172718
rect 418252 172654 418304 172660
rect 379624 171134 379652 172654
rect 390284 172644 390336 172650
rect 390284 172586 390336 172592
rect 400956 172644 401008 172650
rect 400956 172586 401008 172592
rect 408592 172644 408644 172650
rect 408592 172586 408644 172592
rect 380624 172576 380676 172582
rect 380624 172518 380676 172524
rect 379624 171106 380296 171134
rect 380268 151722 380296 171106
rect 380636 170884 380664 172518
rect 390296 170884 390324 172586
rect 399970 170326 400904 170354
rect 380268 151694 380650 151722
rect 390296 148986 390324 151028
rect 399956 149054 399984 151028
rect 400876 149054 400904 170326
rect 399944 149048 399996 149054
rect 399944 148990 399996 148996
rect 400864 149048 400916 149054
rect 400864 148990 400916 148996
rect 400968 148986 400996 172586
rect 408604 170884 408632 172586
rect 418264 170884 418292 172654
rect 428464 172576 428516 172582
rect 428464 172518 428516 172524
rect 427938 170326 428136 170354
rect 405646 161392 405702 161401
rect 405646 161327 405702 161336
rect 401598 160712 401654 160721
rect 401598 160647 401654 160656
rect 401612 151638 401640 160647
rect 405660 151774 405688 161327
rect 405648 151768 405700 151774
rect 405648 151710 405700 151716
rect 401600 151632 401652 151638
rect 401600 151574 401652 151580
rect 408604 148986 408632 151028
rect 390284 148980 390336 148986
rect 390284 148922 390336 148928
rect 400956 148980 401008 148986
rect 400956 148922 401008 148928
rect 408592 148980 408644 148986
rect 408592 148922 408644 148928
rect 418264 148918 418292 151028
rect 427924 149054 427952 151028
rect 428108 149054 428136 170326
rect 427912 149048 427964 149054
rect 427912 148990 427964 148996
rect 428096 149048 428148 149054
rect 428096 148990 428148 148996
rect 428476 148986 428504 172518
rect 428464 148980 428516 148986
rect 428464 148922 428516 148928
rect 418252 148912 418304 148918
rect 418252 148854 418304 148860
rect 408040 146532 408092 146538
rect 408040 146474 408092 146480
rect 428648 146532 428700 146538
rect 428648 146474 428700 146480
rect 389364 146464 389416 146470
rect 389364 146406 389416 146412
rect 399484 146464 399536 146470
rect 399484 146406 399536 146412
rect 389376 143970 389404 146406
rect 399024 146328 399076 146334
rect 399024 146270 399076 146276
rect 399036 143970 399064 146270
rect 389376 143942 389712 143970
rect 399036 143942 399372 143970
rect 379624 143262 380052 143290
rect 379624 122806 379652 143262
rect 399496 124794 399524 146406
rect 400864 146328 400916 146334
rect 400864 146270 400916 146276
rect 399372 124766 399524 124794
rect 379716 124086 380052 124114
rect 389712 124086 390048 124114
rect 379612 122800 379664 122806
rect 379612 122742 379664 122748
rect 379716 122738 379744 124086
rect 390020 122738 390048 124086
rect 400876 122738 400904 146270
rect 408052 143956 408080 146474
rect 417700 146464 417752 146470
rect 417700 146406 417752 146412
rect 417712 143956 417740 146406
rect 428464 146396 428516 146402
rect 428464 146338 428516 146344
rect 427360 146328 427412 146334
rect 427360 146270 427412 146276
rect 427372 143956 427400 146270
rect 405646 134328 405702 134337
rect 405646 134263 405702 134272
rect 401598 133648 401654 133657
rect 401598 133583 401654 133592
rect 401612 125458 401640 133583
rect 405660 125594 405688 134263
rect 428476 132494 428504 146338
rect 428556 146328 428608 146334
rect 428556 146270 428608 146276
rect 427832 132466 428504 132494
rect 405648 125588 405700 125594
rect 405648 125530 405700 125536
rect 401600 125452 401652 125458
rect 401600 125394 401652 125400
rect 427832 124794 427860 132466
rect 427386 124766 427860 124794
rect 408052 122806 408080 124100
rect 408040 122800 408092 122806
rect 408040 122742 408092 122748
rect 417712 122738 417740 124100
rect 428568 122738 428596 146270
rect 428660 126274 428688 146474
rect 428648 126268 428700 126274
rect 428648 126210 428700 126216
rect 379704 122732 379756 122738
rect 379704 122674 379756 122680
rect 390008 122732 390060 122738
rect 390008 122674 390060 122680
rect 400864 122732 400916 122738
rect 400864 122674 400916 122680
rect 417700 122732 417752 122738
rect 417700 122674 417752 122680
rect 428556 122732 428608 122738
rect 428556 122674 428608 122680
rect 379612 118856 379664 118862
rect 379612 118798 379664 118804
rect 418252 118856 418304 118862
rect 418252 118798 418304 118804
rect 379624 113174 379652 118798
rect 390284 118788 390336 118794
rect 390284 118730 390336 118736
rect 400956 118788 401008 118794
rect 400956 118730 401008 118736
rect 408592 118788 408644 118794
rect 408592 118730 408644 118736
rect 380624 118720 380676 118726
rect 380624 118662 380676 118668
rect 380636 116892 380664 118662
rect 390296 116892 390324 118730
rect 399970 116334 400904 116362
rect 379624 113146 380296 113174
rect 380268 97730 380296 113146
rect 380268 97702 380650 97730
rect 390296 95130 390324 97036
rect 399956 95198 399984 97036
rect 400876 95198 400904 116334
rect 399944 95192 399996 95198
rect 399944 95134 399996 95140
rect 400864 95192 400916 95198
rect 400864 95134 400916 95140
rect 400968 95130 400996 118730
rect 408604 116892 408632 118730
rect 418264 116892 418292 118798
rect 428464 118720 428516 118726
rect 428464 118662 428516 118668
rect 427938 116334 428136 116362
rect 405646 107400 405702 107409
rect 405646 107335 405702 107344
rect 401598 106720 401654 106729
rect 401598 106655 401654 106664
rect 401612 97850 401640 106655
rect 405660 97986 405688 107335
rect 405648 97980 405700 97986
rect 405648 97922 405700 97928
rect 401600 97844 401652 97850
rect 401600 97786 401652 97792
rect 408604 95130 408632 97036
rect 390284 95124 390336 95130
rect 390284 95066 390336 95072
rect 400956 95124 401008 95130
rect 400956 95066 401008 95072
rect 408592 95124 408644 95130
rect 408592 95066 408644 95072
rect 418264 95062 418292 97036
rect 427924 95198 427952 97036
rect 428108 95198 428136 116334
rect 427912 95192 427964 95198
rect 427912 95134 427964 95140
rect 428096 95192 428148 95198
rect 428096 95134 428148 95140
rect 428476 95130 428504 118662
rect 428464 95124 428516 95130
rect 428464 95066 428516 95072
rect 418252 95056 418304 95062
rect 418252 94998 418304 95004
rect 408040 91316 408092 91322
rect 408040 91258 408092 91264
rect 428648 91316 428700 91322
rect 428648 91258 428700 91264
rect 389364 91248 389416 91254
rect 389364 91190 389416 91196
rect 399484 91248 399536 91254
rect 399484 91190 399536 91196
rect 389376 89978 389404 91190
rect 399024 91112 399076 91118
rect 399024 91054 399076 91060
rect 399036 89978 399064 91054
rect 389376 89950 389712 89978
rect 399036 89950 399372 89978
rect 379624 89270 380052 89298
rect 379624 69018 379652 89270
rect 399496 70666 399524 91190
rect 400864 91112 400916 91118
rect 400864 91054 400916 91060
rect 399372 70638 399524 70666
rect 379716 70094 380052 70122
rect 389712 70094 390048 70122
rect 379612 69012 379664 69018
rect 379612 68954 379664 68960
rect 379716 68950 379744 70094
rect 390020 68950 390048 70094
rect 400876 68950 400904 91054
rect 408052 89964 408080 91258
rect 417700 91248 417752 91254
rect 417700 91190 417752 91196
rect 417712 89964 417740 91190
rect 428464 91180 428516 91186
rect 428464 91122 428516 91128
rect 427360 91112 427412 91118
rect 427360 91054 427412 91060
rect 427372 89964 427400 91054
rect 405648 88800 405700 88806
rect 405648 88742 405700 88748
rect 405660 80345 405688 88742
rect 405646 80336 405702 80345
rect 405646 80271 405702 80280
rect 401598 79656 401654 79665
rect 401598 79591 401654 79600
rect 401612 71738 401640 79591
rect 428476 74534 428504 91122
rect 428556 91112 428608 91118
rect 428556 91054 428608 91060
rect 427832 74506 428504 74534
rect 401600 71732 401652 71738
rect 401600 71674 401652 71680
rect 427832 70666 427860 74506
rect 427386 70638 427860 70666
rect 408052 69018 408080 70108
rect 408040 69012 408092 69018
rect 408040 68954 408092 68960
rect 417712 68950 417740 70108
rect 428568 68950 428596 91054
rect 428660 72486 428688 91258
rect 428648 72480 428700 72486
rect 428648 72422 428700 72428
rect 379704 68944 379756 68950
rect 379704 68886 379756 68892
rect 390008 68944 390060 68950
rect 390008 68886 390060 68892
rect 400864 68944 400916 68950
rect 400864 68886 400916 68892
rect 417700 68944 417752 68950
rect 417700 68886 417752 68892
rect 428556 68944 428608 68950
rect 428556 68886 428608 68892
rect 379612 65068 379664 65074
rect 379612 65010 379664 65016
rect 418252 65068 418304 65074
rect 418252 65010 418304 65016
rect 379624 55214 379652 65010
rect 390284 65000 390336 65006
rect 390284 64942 390336 64948
rect 400864 65000 400916 65006
rect 400864 64942 400916 64948
rect 408592 65000 408644 65006
rect 408592 64942 408644 64948
rect 380624 64932 380676 64938
rect 380624 64874 380676 64880
rect 380636 62900 380664 64874
rect 390296 62900 390324 64942
rect 399970 62206 400352 62234
rect 400324 58750 400352 62206
rect 400312 58744 400364 58750
rect 400312 58686 400364 58692
rect 379624 55186 380296 55214
rect 380268 43738 380296 55186
rect 380268 43710 380650 43738
rect 390296 41342 390324 43044
rect 399956 41410 399984 43044
rect 399944 41404 399996 41410
rect 399944 41346 399996 41352
rect 400876 41342 400904 64942
rect 408604 62900 408632 64942
rect 418264 62900 418292 65010
rect 428464 64932 428516 64938
rect 428464 64874 428516 64880
rect 427938 62206 428136 62234
rect 400956 58744 401008 58750
rect 400956 58686 401008 58692
rect 400968 41410 400996 58686
rect 405646 53408 405702 53417
rect 405646 53343 405702 53352
rect 401598 52728 401654 52737
rect 401598 52663 401654 52672
rect 401612 44130 401640 52663
rect 405660 44130 405688 53343
rect 401600 44124 401652 44130
rect 401600 44066 401652 44072
rect 405648 44124 405700 44130
rect 405648 44066 405700 44072
rect 400956 41404 401008 41410
rect 400956 41346 401008 41352
rect 408604 41342 408632 43044
rect 390284 41336 390336 41342
rect 390284 41278 390336 41284
rect 400864 41336 400916 41342
rect 400864 41278 400916 41284
rect 408592 41336 408644 41342
rect 408592 41278 408644 41284
rect 418264 41274 418292 43044
rect 427924 41410 427952 43044
rect 428108 41410 428136 62206
rect 427912 41404 427964 41410
rect 427912 41346 427964 41352
rect 428096 41404 428148 41410
rect 428096 41346 428148 41352
rect 428476 41342 428504 64874
rect 428464 41336 428516 41342
rect 428464 41278 428516 41284
rect 418252 41268 418304 41274
rect 418252 41210 418304 41216
rect 389364 37460 389416 37466
rect 389364 37402 389416 37408
rect 399484 37460 399536 37466
rect 399484 37402 399536 37408
rect 417700 37460 417752 37466
rect 417700 37402 417752 37408
rect 389376 35986 389404 37402
rect 399024 37324 399076 37330
rect 399024 37266 399076 37272
rect 399036 35986 399064 37266
rect 389376 35958 389712 35986
rect 399036 35958 399372 35986
rect 379624 35278 380052 35306
rect 379624 13462 379652 35278
rect 399496 16674 399524 37402
rect 408040 37392 408092 37398
rect 408040 37334 408092 37340
rect 400864 37324 400916 37330
rect 400864 37266 400916 37272
rect 399372 16646 399524 16674
rect 379716 16102 380052 16130
rect 389712 16102 390048 16130
rect 379716 13802 379744 16102
rect 390020 13802 390048 16102
rect 400876 13802 400904 37266
rect 408052 35972 408080 37334
rect 417712 35972 417740 37402
rect 428556 37392 428608 37398
rect 428556 37334 428608 37340
rect 427360 37324 427412 37330
rect 427360 37266 427412 37272
rect 428464 37324 428516 37330
rect 428464 37266 428516 37272
rect 427372 35972 427400 37266
rect 401600 34536 401652 34542
rect 401600 34478 401652 34484
rect 405648 34536 405700 34542
rect 405648 34478 405700 34484
rect 401612 25673 401640 34478
rect 405660 26353 405688 34478
rect 405646 26344 405702 26353
rect 405646 26279 405702 26288
rect 401598 25664 401654 25673
rect 401598 25599 401654 25608
rect 427728 16584 427780 16590
rect 427386 16532 427728 16538
rect 427386 16526 427780 16532
rect 427386 16510 427768 16526
rect 379704 13796 379756 13802
rect 379704 13738 379756 13744
rect 390008 13796 390060 13802
rect 390008 13738 390060 13744
rect 400864 13796 400916 13802
rect 400864 13738 400916 13744
rect 408052 13462 408080 16116
rect 417712 13462 417740 16116
rect 428476 13462 428504 37266
rect 428568 18630 428596 37334
rect 428556 18624 428608 18630
rect 428556 18566 428608 18572
rect 429212 15162 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 456064 686044 456116 686050
rect 456064 685986 456116 685992
rect 445668 685976 445720 685982
rect 445668 685918 445720 685924
rect 445680 683876 445708 685918
rect 455328 685908 455380 685914
rect 455328 685850 455380 685856
rect 455340 683876 455368 685850
rect 434824 683318 436034 683346
rect 429292 683188 429344 683194
rect 429292 683130 429344 683136
rect 434628 683188 434680 683194
rect 434628 683130 434680 683136
rect 429304 673577 429332 683130
rect 434640 674257 434668 683130
rect 434626 674248 434682 674257
rect 434626 674183 434682 674192
rect 429290 673568 429346 673577
rect 429290 673503 429346 673512
rect 434824 662250 434852 683318
rect 456076 673454 456104 685986
rect 456156 685908 456208 685914
rect 456156 685850 456208 685856
rect 455800 673426 456104 673454
rect 435732 665848 435784 665854
rect 435732 665790 435784 665796
rect 435744 664714 435772 665790
rect 455800 664714 455828 673426
rect 435744 664686 436034 664714
rect 455354 664686 455828 664714
rect 445680 662318 445708 664020
rect 456168 662318 456196 685850
rect 462226 674248 462282 674257
rect 462226 674183 462282 674192
rect 458178 673568 458234 673577
rect 458178 673503 458234 673512
rect 458192 665174 458220 673503
rect 462240 665174 462268 674183
rect 458180 665168 458232 665174
rect 458180 665110 458232 665116
rect 462228 665168 462280 665174
rect 462228 665110 462280 665116
rect 445668 662312 445720 662318
rect 445668 662254 445720 662260
rect 456156 662312 456208 662318
rect 456156 662254 456208 662260
rect 434812 662244 434864 662250
rect 434812 662186 434864 662192
rect 429844 658368 429896 658374
rect 429844 658310 429896 658316
rect 436284 658368 436336 658374
rect 436284 658310 436336 658316
rect 457444 658368 457496 658374
rect 457444 658310 457496 658316
rect 429292 655648 429344 655654
rect 429292 655590 429344 655596
rect 429304 646785 429332 655590
rect 429290 646776 429346 646785
rect 429290 646711 429346 646720
rect 429856 634642 429884 658310
rect 436296 656962 436324 658310
rect 445944 658300 445996 658306
rect 445944 658242 445996 658248
rect 445956 656962 445984 658242
rect 436296 656934 436632 656962
rect 445956 656934 446292 656962
rect 455952 656254 456104 656282
rect 436468 655648 436520 655654
rect 436468 655590 436520 655596
rect 436480 654090 436508 655590
rect 434628 654084 434680 654090
rect 434628 654026 434680 654032
rect 436468 654084 436520 654090
rect 436468 654026 436520 654032
rect 434640 647465 434668 654026
rect 434626 647456 434682 647465
rect 434626 647391 434682 647400
rect 436632 637078 436968 637106
rect 446292 637078 446628 637106
rect 436940 634710 436968 637078
rect 436928 634704 436980 634710
rect 436928 634646 436980 634652
rect 446600 634642 446628 637078
rect 455616 637078 455952 637106
rect 455616 634778 455644 637078
rect 456076 634778 456104 656254
rect 455604 634772 455656 634778
rect 455604 634714 455656 634720
rect 456064 634772 456116 634778
rect 456064 634714 456116 634720
rect 457456 634642 457484 658310
rect 458180 655580 458232 655586
rect 458180 655522 458232 655528
rect 458192 646785 458220 655522
rect 458178 646776 458234 646785
rect 458178 646711 458234 646720
rect 429844 634636 429896 634642
rect 429844 634578 429896 634584
rect 446588 634636 446640 634642
rect 446588 634578 446640 634584
rect 457444 634636 457496 634642
rect 457444 634578 457496 634584
rect 456156 632256 456208 632262
rect 456156 632198 456208 632204
rect 445668 632188 445720 632194
rect 445668 632130 445720 632136
rect 445680 629884 445708 632130
rect 455328 632120 455380 632126
rect 455328 632062 455380 632068
rect 456064 632120 456116 632126
rect 456064 632062 456116 632068
rect 455340 629884 455368 632062
rect 434824 629326 436034 629354
rect 434626 620256 434682 620265
rect 434626 620191 434682 620200
rect 429290 619576 429346 619585
rect 429290 619511 429346 619520
rect 429304 611250 429332 619511
rect 434640 611250 434668 620191
rect 429292 611244 429344 611250
rect 429292 611186 429344 611192
rect 434628 611244 434680 611250
rect 434628 611186 434680 611192
rect 434824 608462 434852 629326
rect 455696 612808 455748 612814
rect 455696 612750 455748 612756
rect 435732 612060 435784 612066
rect 435732 612002 435784 612008
rect 435744 610722 435772 612002
rect 455708 610722 455736 612750
rect 435744 610694 436034 610722
rect 455354 610694 455736 610722
rect 445680 608530 445708 610028
rect 456076 608530 456104 632062
rect 456168 612814 456196 632198
rect 462226 620256 462282 620265
rect 462226 620191 462282 620200
rect 458178 619576 458234 619585
rect 458178 619511 458234 619520
rect 456156 612808 456208 612814
rect 456156 612750 456208 612756
rect 458192 611318 458220 619511
rect 458180 611312 458232 611318
rect 458180 611254 458232 611260
rect 462240 611182 462268 620191
rect 462228 611176 462280 611182
rect 462228 611118 462280 611124
rect 445668 608524 445720 608530
rect 445668 608466 445720 608472
rect 456064 608524 456116 608530
rect 456064 608466 456116 608472
rect 434812 608456 434864 608462
rect 434812 608398 434864 608404
rect 429844 604580 429896 604586
rect 429844 604522 429896 604528
rect 436284 604580 436336 604586
rect 436284 604522 436336 604528
rect 429292 601792 429344 601798
rect 429292 601734 429344 601740
rect 429304 592793 429332 601734
rect 429290 592784 429346 592793
rect 429290 592719 429346 592728
rect 429856 580854 429884 604522
rect 436296 602970 436324 604522
rect 445944 604512 445996 604518
rect 445944 604454 445996 604460
rect 457444 604512 457496 604518
rect 457444 604454 457496 604460
rect 445956 602970 445984 604454
rect 436296 602942 436632 602970
rect 445956 602942 446292 602970
rect 455952 602262 456104 602290
rect 434628 601792 434680 601798
rect 434628 601734 434680 601740
rect 434640 593473 434668 601734
rect 434626 593464 434682 593473
rect 434626 593399 434682 593408
rect 436632 583086 436968 583114
rect 446292 583086 446628 583114
rect 436940 580922 436968 583086
rect 436928 580916 436980 580922
rect 436928 580858 436980 580864
rect 446600 580854 446628 583086
rect 455616 583086 455952 583114
rect 455616 580990 455644 583086
rect 456076 580990 456104 602262
rect 455604 580984 455656 580990
rect 455604 580926 455656 580932
rect 456064 580984 456116 580990
rect 456064 580926 456116 580932
rect 457456 580854 457484 604454
rect 462228 601860 462280 601866
rect 462228 601802 462280 601808
rect 458180 601724 458232 601730
rect 458180 601666 458232 601672
rect 458192 592793 458220 601666
rect 462240 593473 462268 601802
rect 462226 593464 462282 593473
rect 462226 593399 462282 593408
rect 458178 592784 458234 592793
rect 458178 592719 458234 592728
rect 429844 580848 429896 580854
rect 429844 580790 429896 580796
rect 446588 580848 446640 580854
rect 446588 580790 446640 580796
rect 457444 580848 457496 580854
rect 457444 580790 457496 580796
rect 456156 578400 456208 578406
rect 456156 578342 456208 578348
rect 445668 578332 445720 578338
rect 445668 578274 445720 578280
rect 445680 575892 445708 578274
rect 455328 578264 455380 578270
rect 455328 578206 455380 578212
rect 456064 578264 456116 578270
rect 456064 578206 456116 578212
rect 455340 575892 455368 578206
rect 434824 575334 436034 575362
rect 434626 566264 434682 566273
rect 434626 566199 434682 566208
rect 429290 565584 429346 565593
rect 429290 565519 429346 565528
rect 429304 557462 429332 565519
rect 434640 557462 434668 566199
rect 429292 557456 429344 557462
rect 429292 557398 429344 557404
rect 434628 557456 434680 557462
rect 434628 557398 434680 557404
rect 434824 554606 434852 575334
rect 455696 562352 455748 562358
rect 455696 562294 455748 562300
rect 435732 558204 435784 558210
rect 435732 558146 435784 558152
rect 435744 556730 435772 558146
rect 455708 556730 455736 562294
rect 435744 556702 436034 556730
rect 455354 556702 455736 556730
rect 445680 554674 445708 556036
rect 456076 554674 456104 578206
rect 456168 562358 456196 578342
rect 462226 566264 462282 566273
rect 462226 566199 462282 566208
rect 458178 565584 458234 565593
rect 458178 565519 458234 565528
rect 456156 562352 456208 562358
rect 456156 562294 456208 562300
rect 458192 557530 458220 565519
rect 458180 557524 458232 557530
rect 458180 557466 458232 557472
rect 462240 557394 462268 566199
rect 462228 557388 462280 557394
rect 462228 557330 462280 557336
rect 445668 554668 445720 554674
rect 445668 554610 445720 554616
rect 456064 554668 456116 554674
rect 456064 554610 456116 554616
rect 434812 554600 434864 554606
rect 434812 554542 434864 554548
rect 429844 550724 429896 550730
rect 429844 550666 429896 550672
rect 436284 550724 436336 550730
rect 436284 550666 436336 550672
rect 457444 550724 457496 550730
rect 457444 550666 457496 550672
rect 429290 538792 429346 538801
rect 429290 538727 429346 538736
rect 429304 529854 429332 538727
rect 429292 529848 429344 529854
rect 429292 529790 429344 529796
rect 429856 526998 429884 550666
rect 436296 548978 436324 550666
rect 445944 550656 445996 550662
rect 445944 550598 445996 550604
rect 445956 548978 445984 550598
rect 436296 548950 436632 548978
rect 445956 548950 446292 548978
rect 455952 548270 456104 548298
rect 434626 539472 434682 539481
rect 434626 539407 434682 539416
rect 434640 529854 434668 539407
rect 434628 529848 434680 529854
rect 434628 529790 434680 529796
rect 436632 529094 436968 529122
rect 446292 529094 446628 529122
rect 436940 527066 436968 529094
rect 436928 527060 436980 527066
rect 436928 527002 436980 527008
rect 446600 526998 446628 529094
rect 455616 529094 455952 529122
rect 455616 527134 455644 529094
rect 456076 527134 456104 548270
rect 455604 527128 455656 527134
rect 455604 527070 455656 527076
rect 456064 527128 456116 527134
rect 456064 527070 456116 527076
rect 457456 526998 457484 550666
rect 462226 539472 462282 539481
rect 462226 539407 462282 539416
rect 458178 538792 458234 538801
rect 458178 538727 458234 538736
rect 458192 529922 458220 538727
rect 458180 529916 458232 529922
rect 458180 529858 458232 529864
rect 462240 529786 462268 539407
rect 462228 529780 462280 529786
rect 462228 529722 462280 529728
rect 429844 526992 429896 526998
rect 429844 526934 429896 526940
rect 446588 526992 446640 526998
rect 446588 526934 446640 526940
rect 457444 526992 457496 526998
rect 457444 526934 457496 526940
rect 456156 523184 456208 523190
rect 456156 523126 456208 523132
rect 445668 523116 445720 523122
rect 445668 523058 445720 523064
rect 445680 521900 445708 523058
rect 455328 523048 455380 523054
rect 455328 522990 455380 522996
rect 456064 523048 456116 523054
rect 456064 522990 456116 522996
rect 455340 521900 455368 522990
rect 434824 521206 436034 521234
rect 429292 520328 429344 520334
rect 429292 520270 429344 520276
rect 434628 520328 434680 520334
rect 434628 520270 434680 520276
rect 429304 511601 429332 520270
rect 434640 512281 434668 520270
rect 434626 512272 434682 512281
rect 434626 512207 434682 512216
rect 429290 511592 429346 511601
rect 429290 511527 429346 511536
rect 434824 500818 434852 521206
rect 455696 505640 455748 505646
rect 455696 505582 455748 505588
rect 435732 504416 435784 504422
rect 435732 504358 435784 504364
rect 435744 502738 435772 504358
rect 455708 502738 455736 505582
rect 435744 502710 436034 502738
rect 455354 502710 455736 502738
rect 445680 500886 445708 502044
rect 456076 500886 456104 522990
rect 456168 505646 456196 523126
rect 462226 512272 462282 512281
rect 462226 512207 462282 512216
rect 458178 511592 458234 511601
rect 458178 511527 458234 511536
rect 456156 505640 456208 505646
rect 456156 505582 456208 505588
rect 458192 503674 458220 511527
rect 462240 503674 462268 512207
rect 458180 503668 458232 503674
rect 458180 503610 458232 503616
rect 462228 503668 462280 503674
rect 462228 503610 462280 503616
rect 445668 500880 445720 500886
rect 445668 500822 445720 500828
rect 456064 500880 456116 500886
rect 456064 500822 456116 500828
rect 434812 500812 434864 500818
rect 434812 500754 434864 500760
rect 429844 496936 429896 496942
rect 429844 496878 429896 496884
rect 436284 496936 436336 496942
rect 436284 496878 436336 496884
rect 457444 496936 457496 496942
rect 457444 496878 457496 496884
rect 429290 484800 429346 484809
rect 429290 484735 429346 484744
rect 429304 475998 429332 484735
rect 429292 475992 429344 475998
rect 429292 475934 429344 475940
rect 429856 473210 429884 496878
rect 436296 494986 436324 496878
rect 445944 496868 445996 496874
rect 445944 496810 445996 496816
rect 445956 494986 445984 496810
rect 436296 494958 436632 494986
rect 445956 494958 446292 494986
rect 455952 494278 456104 494306
rect 434626 485480 434682 485489
rect 434626 485415 434682 485424
rect 434640 475930 434668 485415
rect 434628 475924 434680 475930
rect 434628 475866 434680 475872
rect 436632 475102 436968 475130
rect 446292 475102 446628 475130
rect 436940 473278 436968 475102
rect 436928 473272 436980 473278
rect 436928 473214 436980 473220
rect 446600 473210 446628 475102
rect 455616 475102 455952 475130
rect 455616 473346 455644 475102
rect 456076 473346 456104 494278
rect 455604 473340 455656 473346
rect 455604 473282 455656 473288
rect 456064 473340 456116 473346
rect 456064 473282 456116 473288
rect 457456 473210 457484 496878
rect 462226 485480 462282 485489
rect 462226 485415 462282 485424
rect 458178 484800 458234 484809
rect 458178 484735 458234 484744
rect 458192 476066 458220 484735
rect 458180 476060 458232 476066
rect 458180 476002 458232 476008
rect 462240 475998 462268 485415
rect 462228 475992 462280 475998
rect 462228 475934 462280 475940
rect 429844 473204 429896 473210
rect 429844 473146 429896 473152
rect 446588 473204 446640 473210
rect 446588 473146 446640 473152
rect 457444 473204 457496 473210
rect 457444 473146 457496 473152
rect 456156 469396 456208 469402
rect 456156 469338 456208 469344
rect 445668 469328 445720 469334
rect 445668 469270 445720 469276
rect 445680 467908 445708 469270
rect 455328 469260 455380 469266
rect 455328 469202 455380 469208
rect 456064 469260 456116 469266
rect 456064 469202 456116 469208
rect 455340 467908 455368 469202
rect 434824 467214 436034 467242
rect 429292 466540 429344 466546
rect 429292 466482 429344 466488
rect 434628 466540 434680 466546
rect 434628 466482 434680 466488
rect 429304 457609 429332 466482
rect 434640 458289 434668 466482
rect 434626 458280 434682 458289
rect 434626 458215 434682 458224
rect 429290 457600 429346 457609
rect 429290 457535 429346 457544
rect 434824 445602 434852 467214
rect 435732 450560 435784 450566
rect 435732 450502 435784 450508
rect 435744 448746 435772 450502
rect 455696 449676 455748 449682
rect 455696 449618 455748 449624
rect 455708 448746 455736 449618
rect 435744 448718 436034 448746
rect 455354 448718 455736 448746
rect 445680 445670 445708 448052
rect 456076 445670 456104 469202
rect 456168 449682 456196 469338
rect 462228 466608 462280 466614
rect 462228 466550 462280 466556
rect 458180 466472 458232 466478
rect 458180 466414 458232 466420
rect 458192 457609 458220 466414
rect 462240 458289 462268 466550
rect 462226 458280 462282 458289
rect 462226 458215 462282 458224
rect 458178 457600 458234 457609
rect 458178 457535 458234 457544
rect 456156 449676 456208 449682
rect 456156 449618 456208 449624
rect 445668 445664 445720 445670
rect 445668 445606 445720 445612
rect 456064 445664 456116 445670
rect 456064 445606 456116 445612
rect 434812 445596 434864 445602
rect 434812 445538 434864 445544
rect 429844 443080 429896 443086
rect 429844 443022 429896 443028
rect 436284 443080 436336 443086
rect 436284 443022 436336 443028
rect 429292 440292 429344 440298
rect 429292 440234 429344 440240
rect 429304 430817 429332 440234
rect 429290 430808 429346 430817
rect 429290 430743 429346 430752
rect 429856 419354 429884 443022
rect 436296 440994 436324 443022
rect 445944 443012 445996 443018
rect 445944 442954 445996 442960
rect 457444 443012 457496 443018
rect 457444 442954 457496 442960
rect 445956 440994 445984 442954
rect 436296 440966 436632 440994
rect 445956 440966 446292 440994
rect 434628 440292 434680 440298
rect 455952 440286 456104 440314
rect 434628 440234 434680 440240
rect 434640 431497 434668 440234
rect 434626 431488 434682 431497
rect 434626 431423 434682 431432
rect 436632 421110 436968 421138
rect 446292 421110 446628 421138
rect 436940 419422 436968 421110
rect 436928 419416 436980 419422
rect 436928 419358 436980 419364
rect 446600 419354 446628 421110
rect 455616 421110 455952 421138
rect 455616 419490 455644 421110
rect 456076 419490 456104 440286
rect 455604 419484 455656 419490
rect 455604 419426 455656 419432
rect 456064 419484 456116 419490
rect 456064 419426 456116 419432
rect 457456 419354 457484 442954
rect 462226 431488 462282 431497
rect 462226 431423 462282 431432
rect 458178 430808 458234 430817
rect 458178 430743 458234 430752
rect 458192 422278 458220 430743
rect 462240 422278 462268 431423
rect 458180 422272 458232 422278
rect 458180 422214 458232 422220
rect 462228 422272 462280 422278
rect 462228 422214 462280 422220
rect 429844 419348 429896 419354
rect 429844 419290 429896 419296
rect 446588 419348 446640 419354
rect 446588 419290 446640 419296
rect 457444 419348 457496 419354
rect 457444 419290 457496 419296
rect 456064 415608 456116 415614
rect 456064 415550 456116 415556
rect 445668 415540 445720 415546
rect 445668 415482 445720 415488
rect 445680 413916 445708 415482
rect 455328 415472 455380 415478
rect 455328 415414 455380 415420
rect 455340 413916 455368 415414
rect 434824 413222 436034 413250
rect 434626 404288 434682 404297
rect 434626 404223 434682 404232
rect 429290 403608 429346 403617
rect 429290 403543 429346 403552
rect 429304 394602 429332 403543
rect 429292 394596 429344 394602
rect 429292 394538 429344 394544
rect 434640 394534 434668 404223
rect 434628 394528 434680 394534
rect 434628 394470 434680 394476
rect 434824 391814 434852 413222
rect 456076 402974 456104 415550
rect 456156 415472 456208 415478
rect 456156 415414 456208 415420
rect 455800 402946 456104 402974
rect 435732 395344 435784 395350
rect 435732 395286 435784 395292
rect 435744 394754 435772 395286
rect 455800 394754 455828 402946
rect 435744 394726 436034 394754
rect 455354 394726 455828 394754
rect 445680 391882 445708 394060
rect 456168 391882 456196 415414
rect 462226 404288 462282 404297
rect 462226 404223 462282 404232
rect 458178 403608 458234 403617
rect 458178 403543 458234 403552
rect 458192 394670 458220 403543
rect 458180 394664 458232 394670
rect 458180 394606 458232 394612
rect 462240 394602 462268 404223
rect 462228 394596 462280 394602
rect 462228 394538 462280 394544
rect 445668 391876 445720 391882
rect 445668 391818 445720 391824
rect 456156 391876 456208 391882
rect 456156 391818 456208 391824
rect 434812 391808 434864 391814
rect 434812 391750 434864 391756
rect 429844 389292 429896 389298
rect 429844 389234 429896 389240
rect 436284 389292 436336 389298
rect 436284 389234 436336 389240
rect 457444 389292 457496 389298
rect 457444 389234 457496 389240
rect 429292 386504 429344 386510
rect 429292 386446 429344 386452
rect 429304 376825 429332 386446
rect 429290 376816 429346 376825
rect 429290 376751 429346 376760
rect 429856 365566 429884 389234
rect 436296 386866 436324 389234
rect 445944 389224 445996 389230
rect 445944 389166 445996 389172
rect 445956 386866 445984 389166
rect 436296 386838 436632 386866
rect 445956 386838 446292 386866
rect 434628 386504 434680 386510
rect 434628 386446 434680 386452
rect 434640 377505 434668 386446
rect 455952 386294 456104 386322
rect 434626 377496 434682 377505
rect 434626 377431 434682 377440
rect 436632 367118 436968 367146
rect 446292 367118 446628 367146
rect 436940 365634 436968 367118
rect 436928 365628 436980 365634
rect 436928 365570 436980 365576
rect 446600 365566 446628 367118
rect 455616 367118 455952 367146
rect 455616 365702 455644 367118
rect 456076 365702 456104 386294
rect 455604 365696 455656 365702
rect 455604 365638 455656 365644
rect 456064 365696 456116 365702
rect 456064 365638 456116 365644
rect 457456 365566 457484 389234
rect 462228 386572 462280 386578
rect 462228 386514 462280 386520
rect 458180 386436 458232 386442
rect 458180 386378 458232 386384
rect 458192 376825 458220 386378
rect 462240 377505 462268 386514
rect 462226 377496 462282 377505
rect 462226 377431 462282 377440
rect 458178 376816 458234 376825
rect 458178 376751 458234 376760
rect 429844 365560 429896 365566
rect 429844 365502 429896 365508
rect 446588 365560 446640 365566
rect 446588 365502 446640 365508
rect 457444 365560 457496 365566
rect 457444 365502 457496 365508
rect 445668 361752 445720 361758
rect 445668 361694 445720 361700
rect 456064 361752 456116 361758
rect 456064 361694 456116 361700
rect 445680 359924 445708 361694
rect 455328 361616 455380 361622
rect 455328 361558 455380 361564
rect 455340 359924 455368 361558
rect 434824 359230 436034 359258
rect 434626 350296 434682 350305
rect 434626 350231 434682 350240
rect 429290 349616 429346 349625
rect 429290 349551 429346 349560
rect 429304 340814 429332 349551
rect 434640 340814 434668 350231
rect 429292 340808 429344 340814
rect 429292 340750 429344 340756
rect 434628 340808 434680 340814
rect 434628 340750 434680 340756
rect 434824 337958 434852 359230
rect 456076 345014 456104 361694
rect 456156 361616 456208 361622
rect 456156 361558 456208 361564
rect 455800 344986 456104 345014
rect 435732 341556 435784 341562
rect 435732 341498 435784 341504
rect 435744 340762 435772 341498
rect 455800 340762 455828 344986
rect 435744 340734 436034 340762
rect 455354 340734 455828 340762
rect 445680 338026 445708 340068
rect 456168 338026 456196 361558
rect 462226 350296 462282 350305
rect 462226 350231 462282 350240
rect 458178 349616 458234 349625
rect 458178 349551 458234 349560
rect 458192 340882 458220 349551
rect 458180 340876 458232 340882
rect 458180 340818 458232 340824
rect 462240 340746 462268 350231
rect 462228 340740 462280 340746
rect 462228 340682 462280 340688
rect 445668 338020 445720 338026
rect 445668 337962 445720 337968
rect 456156 338020 456208 338026
rect 456156 337962 456208 337968
rect 434812 337952 434864 337958
rect 434812 337894 434864 337900
rect 429844 335436 429896 335442
rect 429844 335378 429896 335384
rect 436284 335436 436336 335442
rect 436284 335378 436336 335384
rect 457444 335436 457496 335442
rect 457444 335378 457496 335384
rect 429290 322144 429346 322153
rect 429290 322079 429346 322088
rect 429304 314634 429332 322079
rect 429292 314628 429344 314634
rect 429292 314570 429344 314576
rect 429856 311710 429884 335378
rect 436296 332874 436324 335378
rect 445944 335368 445996 335374
rect 445944 335310 445996 335316
rect 445956 332874 445984 335310
rect 436296 332846 436632 332874
rect 445956 332846 446292 332874
rect 455952 332302 456104 332330
rect 434626 322960 434682 322969
rect 434626 322895 434682 322904
rect 434640 314634 434668 322895
rect 434628 314628 434680 314634
rect 434628 314570 434680 314576
rect 436632 313126 436968 313154
rect 446292 313126 446628 313154
rect 436940 311778 436968 313126
rect 436928 311772 436980 311778
rect 436928 311714 436980 311720
rect 446600 311710 446628 313126
rect 455616 313126 455952 313154
rect 455616 311846 455644 313126
rect 456076 311846 456104 332302
rect 455604 311840 455656 311846
rect 455604 311782 455656 311788
rect 456064 311840 456116 311846
rect 456064 311782 456116 311788
rect 457456 311710 457484 335378
rect 458180 331288 458232 331294
rect 458180 331230 458232 331236
rect 458192 322833 458220 331230
rect 462226 322960 462282 322969
rect 462226 322895 462282 322904
rect 458178 322824 458234 322833
rect 458178 322759 458234 322768
rect 462240 314566 462268 322895
rect 462228 314560 462280 314566
rect 462228 314502 462280 314508
rect 429844 311704 429896 311710
rect 429844 311646 429896 311652
rect 446588 311704 446640 311710
rect 446588 311646 446640 311652
rect 457444 311704 457496 311710
rect 457444 311646 457496 311652
rect 456156 307964 456208 307970
rect 456156 307906 456208 307912
rect 445668 307896 445720 307902
rect 445668 307838 445720 307844
rect 445680 305932 445708 307838
rect 455328 307828 455380 307834
rect 455328 307770 455380 307776
rect 456064 307828 456116 307834
rect 456064 307770 456116 307776
rect 455340 305932 455368 307770
rect 434824 305238 436034 305266
rect 434626 296304 434682 296313
rect 434626 296239 434682 296248
rect 429290 295624 429346 295633
rect 429290 295559 429346 295568
rect 429304 286958 429332 295559
rect 434640 286958 434668 296239
rect 429292 286952 429344 286958
rect 429292 286894 429344 286900
rect 434628 286952 434680 286958
rect 434628 286894 434680 286900
rect 434824 284170 434852 305238
rect 455696 291916 455748 291922
rect 455696 291858 455748 291864
rect 435732 287700 435784 287706
rect 435732 287642 435784 287648
rect 435744 286770 435772 287642
rect 455708 286770 455736 291858
rect 435744 286742 436034 286770
rect 455354 286742 455736 286770
rect 445680 284238 445708 286076
rect 456076 284238 456104 307770
rect 456168 291922 456196 307906
rect 462226 296304 462282 296313
rect 462226 296239 462282 296248
rect 458178 295624 458234 295633
rect 458178 295559 458234 295568
rect 456156 291916 456208 291922
rect 456156 291858 456208 291864
rect 458192 287026 458220 295559
rect 458180 287020 458232 287026
rect 458180 286962 458232 286968
rect 462240 286890 462268 296239
rect 462228 286884 462280 286890
rect 462228 286826 462280 286832
rect 445668 284232 445720 284238
rect 445668 284174 445720 284180
rect 456064 284232 456116 284238
rect 456064 284174 456116 284180
rect 434812 284164 434864 284170
rect 434812 284106 434864 284112
rect 429844 280288 429896 280294
rect 429844 280230 429896 280236
rect 436284 280288 436336 280294
rect 436284 280230 436336 280236
rect 457444 280288 457496 280294
rect 457444 280230 457496 280236
rect 429292 277500 429344 277506
rect 429292 277442 429344 277448
rect 429304 269113 429332 277442
rect 429290 269104 429346 269113
rect 429290 269039 429346 269048
rect 429856 256562 429884 280230
rect 436296 278882 436324 280230
rect 445944 280220 445996 280226
rect 445944 280162 445996 280168
rect 445956 278882 445984 280162
rect 436296 278854 436632 278882
rect 445956 278854 446292 278882
rect 455952 278310 456104 278338
rect 434628 277500 434680 277506
rect 434628 277442 434680 277448
rect 434640 270065 434668 277442
rect 434626 270056 434682 270065
rect 434626 269991 434682 270000
rect 436632 259134 436968 259162
rect 446292 259134 446628 259162
rect 436940 256630 436968 259134
rect 436928 256624 436980 256630
rect 436928 256566 436980 256572
rect 446600 256562 446628 259134
rect 455616 259134 455952 259162
rect 455616 256698 455644 259134
rect 456076 256698 456104 278310
rect 455604 256692 455656 256698
rect 455604 256634 455656 256640
rect 456064 256692 456116 256698
rect 456064 256634 456116 256640
rect 457456 256562 457484 280230
rect 462228 277568 462280 277574
rect 462228 277510 462280 277516
rect 458180 277432 458232 277438
rect 458180 277374 458232 277380
rect 458192 269113 458220 277374
rect 462240 270065 462268 277510
rect 462226 270056 462282 270065
rect 462226 269991 462282 270000
rect 458178 269104 458234 269113
rect 458178 269039 458234 269048
rect 429844 256556 429896 256562
rect 429844 256498 429896 256504
rect 446588 256556 446640 256562
rect 446588 256498 446640 256504
rect 457444 256556 457496 256562
rect 457444 256498 457496 256504
rect 456064 254108 456116 254114
rect 456064 254050 456116 254056
rect 445668 254040 445720 254046
rect 445668 253982 445720 253988
rect 445680 251940 445708 253982
rect 455328 253972 455380 253978
rect 455328 253914 455380 253920
rect 455340 251940 455368 253914
rect 429292 251320 429344 251326
rect 429292 251262 429344 251268
rect 434628 251320 434680 251326
rect 434628 251262 434680 251268
rect 429304 241641 429332 251262
rect 434640 242321 434668 251262
rect 434824 251246 436034 251274
rect 434626 242312 434682 242321
rect 434626 242247 434682 242256
rect 429290 241632 429346 241641
rect 429290 241567 429346 241576
rect 434824 230314 434852 251246
rect 456076 238754 456104 254050
rect 456156 253972 456208 253978
rect 456156 253914 456208 253920
rect 455800 238726 456104 238754
rect 435732 233912 435784 233918
rect 435732 233854 435784 233860
rect 435744 232778 435772 233854
rect 455800 232778 455828 238726
rect 435744 232750 436034 232778
rect 455354 232750 455828 232778
rect 445680 230382 445708 232084
rect 456168 230382 456196 253914
rect 462228 251388 462280 251394
rect 462228 251330 462280 251336
rect 458180 251252 458232 251258
rect 458180 251194 458232 251200
rect 458192 241641 458220 251194
rect 462240 242321 462268 251330
rect 462226 242312 462282 242321
rect 462226 242247 462282 242256
rect 458178 241632 458234 241641
rect 458178 241567 458234 241576
rect 445668 230376 445720 230382
rect 445668 230318 445720 230324
rect 456156 230376 456208 230382
rect 456156 230318 456208 230324
rect 434812 230308 434864 230314
rect 434812 230250 434864 230256
rect 429844 226432 429896 226438
rect 429844 226374 429896 226380
rect 436284 226432 436336 226438
rect 436284 226374 436336 226380
rect 429292 223712 429344 223718
rect 429292 223654 429344 223660
rect 429304 214713 429332 223654
rect 429290 214704 429346 214713
rect 429290 214639 429346 214648
rect 429856 202706 429884 226374
rect 436296 224890 436324 226374
rect 445944 226364 445996 226370
rect 445944 226306 445996 226312
rect 457444 226364 457496 226370
rect 457444 226306 457496 226312
rect 445956 224890 445984 226306
rect 436296 224862 436632 224890
rect 445956 224862 446292 224890
rect 455952 224318 456104 224346
rect 434628 223712 434680 223718
rect 434628 223654 434680 223660
rect 434640 215393 434668 223654
rect 434626 215384 434682 215393
rect 434626 215319 434682 215328
rect 436632 205006 436968 205034
rect 446292 205006 446628 205034
rect 436940 202774 436968 205006
rect 436928 202768 436980 202774
rect 436928 202710 436980 202716
rect 446600 202706 446628 205006
rect 455616 205006 455952 205034
rect 455616 202842 455644 205006
rect 456076 202842 456104 224318
rect 455604 202836 455656 202842
rect 455604 202778 455656 202784
rect 456064 202836 456116 202842
rect 456064 202778 456116 202784
rect 457456 202706 457484 226306
rect 462228 223780 462280 223786
rect 462228 223722 462280 223728
rect 458180 223644 458232 223650
rect 458180 223586 458232 223592
rect 458192 214713 458220 223586
rect 462240 215393 462268 223722
rect 462226 215384 462282 215393
rect 462226 215319 462282 215328
rect 458178 214704 458234 214713
rect 458178 214639 458234 214648
rect 429844 202700 429896 202706
rect 429844 202642 429896 202648
rect 446588 202700 446640 202706
rect 446588 202642 446640 202648
rect 457444 202700 457496 202706
rect 457444 202642 457496 202648
rect 456156 200320 456208 200326
rect 456156 200262 456208 200268
rect 445668 200252 445720 200258
rect 445668 200194 445720 200200
rect 445680 197948 445708 200194
rect 455328 200184 455380 200190
rect 455328 200126 455380 200132
rect 456064 200184 456116 200190
rect 456064 200126 456116 200132
rect 455340 197948 455368 200126
rect 434824 197254 436034 197282
rect 434626 188320 434682 188329
rect 434626 188255 434682 188264
rect 429290 187640 429346 187649
rect 429290 187575 429346 187584
rect 429304 179314 429332 187575
rect 434640 179314 434668 188255
rect 429292 179308 429344 179314
rect 429292 179250 429344 179256
rect 434628 179308 434680 179314
rect 434628 179250 434680 179256
rect 434824 176526 434852 197254
rect 455696 185632 455748 185638
rect 455696 185574 455748 185580
rect 435732 180124 435784 180130
rect 435732 180066 435784 180072
rect 435744 178786 435772 180066
rect 455708 178786 455736 185574
rect 435744 178758 436034 178786
rect 455354 178758 455736 178786
rect 445680 176594 445708 178092
rect 456076 176594 456104 200126
rect 456168 185638 456196 200262
rect 462226 188320 462282 188329
rect 462226 188255 462282 188264
rect 458178 187640 458234 187649
rect 458178 187575 458234 187584
rect 456156 185632 456208 185638
rect 456156 185574 456208 185580
rect 458192 179382 458220 187575
rect 458180 179376 458232 179382
rect 458180 179318 458232 179324
rect 462240 179246 462268 188255
rect 462228 179240 462280 179246
rect 462228 179182 462280 179188
rect 445668 176588 445720 176594
rect 445668 176530 445720 176536
rect 456064 176588 456116 176594
rect 456064 176530 456116 176536
rect 434812 176520 434864 176526
rect 434812 176462 434864 176468
rect 429844 172644 429896 172650
rect 429844 172586 429896 172592
rect 436284 172644 436336 172650
rect 436284 172586 436336 172592
rect 457444 172644 457496 172650
rect 457444 172586 457496 172592
rect 429290 160712 429346 160721
rect 429290 160647 429346 160656
rect 429304 151706 429332 160647
rect 429292 151700 429344 151706
rect 429292 151642 429344 151648
rect 429856 148918 429884 172586
rect 436296 170898 436324 172586
rect 445944 172576 445996 172582
rect 445944 172518 445996 172524
rect 445956 170898 445984 172518
rect 436296 170870 436632 170898
rect 445956 170870 446292 170898
rect 455952 170326 456104 170354
rect 434626 161392 434682 161401
rect 434626 161327 434682 161336
rect 434640 151706 434668 161327
rect 434628 151700 434680 151706
rect 434628 151642 434680 151648
rect 436632 151014 436968 151042
rect 446292 151014 446628 151042
rect 436940 148986 436968 151014
rect 436928 148980 436980 148986
rect 436928 148922 436980 148928
rect 446600 148918 446628 151014
rect 455616 151014 455952 151042
rect 455616 149054 455644 151014
rect 456076 149054 456104 170326
rect 455604 149048 455656 149054
rect 455604 148990 455656 148996
rect 456064 149048 456116 149054
rect 456064 148990 456116 148996
rect 457456 148918 457484 172586
rect 462226 161392 462282 161401
rect 462226 161327 462282 161336
rect 458178 160712 458234 160721
rect 458178 160647 458234 160656
rect 458192 151774 458220 160647
rect 458180 151768 458232 151774
rect 458180 151710 458232 151716
rect 462240 151638 462268 161327
rect 462228 151632 462280 151638
rect 462228 151574 462280 151580
rect 429844 148912 429896 148918
rect 429844 148854 429896 148860
rect 446588 148912 446640 148918
rect 446588 148854 446640 148860
rect 457444 148912 457496 148918
rect 457444 148854 457496 148860
rect 456156 146464 456208 146470
rect 456156 146406 456208 146412
rect 445668 146396 445720 146402
rect 445668 146338 445720 146344
rect 445680 143956 445708 146338
rect 455328 146328 455380 146334
rect 455328 146270 455380 146276
rect 456064 146328 456116 146334
rect 456064 146270 456116 146276
rect 455340 143956 455368 146270
rect 434824 143262 436034 143290
rect 434626 134328 434682 134337
rect 434626 134263 434682 134272
rect 429290 133648 429346 133657
rect 429290 133583 429346 133592
rect 429304 125526 429332 133583
rect 434640 125526 434668 134263
rect 429292 125520 429344 125526
rect 429292 125462 429344 125468
rect 434628 125520 434680 125526
rect 434628 125462 434680 125468
rect 434824 122670 434852 143262
rect 455696 128308 455748 128314
rect 455696 128250 455748 128256
rect 435732 126268 435784 126274
rect 435732 126210 435784 126216
rect 435744 124794 435772 126210
rect 455708 124794 455736 128250
rect 435744 124766 436034 124794
rect 455354 124766 455736 124794
rect 445680 122738 445708 124100
rect 456076 122738 456104 146270
rect 456168 128314 456196 146406
rect 462226 134328 462282 134337
rect 462226 134263 462282 134272
rect 458178 133648 458234 133657
rect 458178 133583 458234 133592
rect 456156 128308 456208 128314
rect 456156 128250 456208 128256
rect 458192 125594 458220 133583
rect 458180 125588 458232 125594
rect 458180 125530 458232 125536
rect 462240 125458 462268 134263
rect 462228 125452 462280 125458
rect 462228 125394 462280 125400
rect 445668 122732 445720 122738
rect 445668 122674 445720 122680
rect 456064 122732 456116 122738
rect 456064 122674 456116 122680
rect 434812 122664 434864 122670
rect 434812 122606 434864 122612
rect 429844 118788 429896 118794
rect 429844 118730 429896 118736
rect 436284 118788 436336 118794
rect 436284 118730 436336 118736
rect 457444 118788 457496 118794
rect 457444 118730 457496 118736
rect 429290 106720 429346 106729
rect 429290 106655 429346 106664
rect 429304 97918 429332 106655
rect 429292 97912 429344 97918
rect 429292 97854 429344 97860
rect 429856 95062 429884 118730
rect 436296 116906 436324 118730
rect 445944 118720 445996 118726
rect 445944 118662 445996 118668
rect 445956 116906 445984 118662
rect 436296 116878 436632 116906
rect 445956 116878 446292 116906
rect 455952 116334 456104 116362
rect 434626 107400 434682 107409
rect 434626 107335 434682 107344
rect 434640 97918 434668 107335
rect 434628 97912 434680 97918
rect 434628 97854 434680 97860
rect 436632 97022 436968 97050
rect 446292 97022 446628 97050
rect 436940 95130 436968 97022
rect 436928 95124 436980 95130
rect 436928 95066 436980 95072
rect 446600 95062 446628 97022
rect 455616 97022 455952 97050
rect 455616 95198 455644 97022
rect 456076 95198 456104 116334
rect 455604 95192 455656 95198
rect 455604 95134 455656 95140
rect 456064 95192 456116 95198
rect 456064 95134 456116 95140
rect 457456 95062 457484 118730
rect 462226 107400 462282 107409
rect 462226 107335 462282 107344
rect 458178 106720 458234 106729
rect 458178 106655 458234 106664
rect 458192 97986 458220 106655
rect 458180 97980 458232 97986
rect 458180 97922 458232 97928
rect 462240 97850 462268 107335
rect 462228 97844 462280 97850
rect 462228 97786 462280 97792
rect 429844 95056 429896 95062
rect 429844 94998 429896 95004
rect 446588 95056 446640 95062
rect 446588 94998 446640 95004
rect 457444 95056 457496 95062
rect 457444 94998 457496 95004
rect 456156 91248 456208 91254
rect 456156 91190 456208 91196
rect 445668 91180 445720 91186
rect 445668 91122 445720 91128
rect 445680 89964 445708 91122
rect 455328 91112 455380 91118
rect 455328 91054 455380 91060
rect 456064 91112 456116 91118
rect 456064 91054 456116 91060
rect 455340 89964 455368 91054
rect 434824 89270 436034 89298
rect 434628 88868 434680 88874
rect 434628 88810 434680 88816
rect 429292 88392 429344 88398
rect 429292 88334 429344 88340
rect 429304 79665 429332 88334
rect 434640 80345 434668 88810
rect 434626 80336 434682 80345
rect 434626 80271 434682 80280
rect 429290 79656 429346 79665
rect 429290 79591 429346 79600
rect 434824 68882 434852 89270
rect 435732 72480 435784 72486
rect 435732 72422 435784 72428
rect 435744 70666 435772 72422
rect 455696 72344 455748 72350
rect 455696 72286 455748 72292
rect 455708 70666 455736 72286
rect 435744 70638 436034 70666
rect 455354 70638 455736 70666
rect 445680 68950 445708 70108
rect 456076 68950 456104 91054
rect 456168 72350 456196 91190
rect 458180 88800 458232 88806
rect 458180 88742 458232 88748
rect 458192 79665 458220 88742
rect 462226 80336 462282 80345
rect 462226 80271 462282 80280
rect 458178 79656 458234 79665
rect 458178 79591 458234 79600
rect 456156 72344 456208 72350
rect 456156 72286 456208 72292
rect 462240 71738 462268 80271
rect 462228 71732 462280 71738
rect 462228 71674 462280 71680
rect 445668 68944 445720 68950
rect 445668 68886 445720 68892
rect 456064 68944 456116 68950
rect 456064 68886 456116 68892
rect 434812 68876 434864 68882
rect 434812 68818 434864 68824
rect 429844 65000 429896 65006
rect 429844 64942 429896 64948
rect 436284 65000 436336 65006
rect 436284 64942 436336 64948
rect 457444 65000 457496 65006
rect 457444 64942 457496 64948
rect 429292 62144 429344 62150
rect 429292 62086 429344 62092
rect 429304 52737 429332 62086
rect 429290 52728 429346 52737
rect 429290 52663 429346 52672
rect 429856 41274 429884 64942
rect 436296 62914 436324 64942
rect 445944 64932 445996 64938
rect 445944 64874 445996 64880
rect 445956 62914 445984 64874
rect 436296 62886 436632 62914
rect 445956 62886 446292 62914
rect 455952 62206 456104 62234
rect 434628 62144 434680 62150
rect 434628 62086 434680 62092
rect 434640 53417 434668 62086
rect 434626 53408 434682 53417
rect 434626 53343 434682 53352
rect 436632 43030 436968 43058
rect 446292 43030 446628 43058
rect 436940 41342 436968 43030
rect 436928 41336 436980 41342
rect 436928 41278 436980 41284
rect 446600 41274 446628 43030
rect 455616 43030 455952 43058
rect 455616 41410 455644 43030
rect 456076 41410 456104 62206
rect 455604 41404 455656 41410
rect 455604 41346 455656 41352
rect 456064 41404 456116 41410
rect 456064 41346 456116 41352
rect 457456 41274 457484 64942
rect 462226 53408 462282 53417
rect 462226 53343 462282 53352
rect 458178 52728 458234 52737
rect 458178 52663 458234 52672
rect 458192 44130 458220 52663
rect 462240 44130 462268 53343
rect 458180 44124 458232 44130
rect 458180 44066 458232 44072
rect 462228 44124 462280 44130
rect 462228 44066 462280 44072
rect 429844 41268 429896 41274
rect 429844 41210 429896 41216
rect 446588 41268 446640 41274
rect 446588 41210 446640 41216
rect 457444 41268 457496 41274
rect 457444 41210 457496 41216
rect 462332 38282 462360 703520
rect 494808 700466 494836 703520
rect 494796 700460 494848 700466
rect 494796 700402 494848 700408
rect 527192 700398 527220 703520
rect 518164 700392 518216 700398
rect 518164 700334 518216 700340
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 492036 686112 492088 686118
rect 492036 686054 492088 686060
rect 512736 686112 512788 686118
rect 512736 686054 512788 686060
rect 473360 686044 473412 686050
rect 473360 685986 473412 685992
rect 483480 686044 483532 686050
rect 483480 685986 483532 685992
rect 464344 685976 464396 685982
rect 464344 685918 464396 685924
rect 464356 683890 464384 685918
rect 464048 683862 464384 683890
rect 473372 683890 473400 685986
rect 483020 685908 483072 685914
rect 483020 685850 483072 685856
rect 483032 683890 483060 685850
rect 473372 683862 473708 683890
rect 483032 683862 483368 683890
rect 483492 664714 483520 685986
rect 483664 685976 483716 685982
rect 483664 685918 483716 685924
rect 483676 665310 483704 685918
rect 485044 685908 485096 685914
rect 485044 685850 485096 685856
rect 483664 665304 483716 665310
rect 483664 665246 483716 665252
rect 483368 664686 483520 664714
rect 463804 664006 464048 664034
rect 473708 664006 474044 664034
rect 463804 662250 463832 664006
rect 474016 662386 474044 664006
rect 485056 662386 485084 685850
rect 492048 683876 492076 686054
rect 501696 686044 501748 686050
rect 501696 685986 501748 685992
rect 501708 683876 501736 685986
rect 511448 685976 511500 685982
rect 511448 685918 511500 685924
rect 511356 685908 511408 685914
rect 511356 685850 511408 685856
rect 511368 683876 511396 685850
rect 485780 683188 485832 683194
rect 485780 683130 485832 683136
rect 489828 683188 489880 683194
rect 489828 683130 489880 683136
rect 485792 673577 485820 683130
rect 489840 674257 489868 683130
rect 489826 674248 489882 674257
rect 489826 674183 489882 674192
rect 485778 673568 485834 673577
rect 485778 673503 485834 673512
rect 491668 665304 491720 665310
rect 491668 665246 491720 665252
rect 491680 664714 491708 665246
rect 511460 664714 511488 685918
rect 512644 685908 512696 685914
rect 512644 685850 512696 685856
rect 491680 664686 492062 664714
rect 511382 664686 511488 664714
rect 501708 662386 501736 664020
rect 512656 662386 512684 685850
rect 512748 665310 512776 686054
rect 513378 673568 513434 673577
rect 513378 673503 513434 673512
rect 512736 665304 512788 665310
rect 512736 665246 512788 665252
rect 513392 665174 513420 673503
rect 513380 665168 513432 665174
rect 513380 665110 513432 665116
rect 474004 662380 474056 662386
rect 474004 662322 474056 662328
rect 485044 662380 485096 662386
rect 485044 662322 485096 662328
rect 501696 662380 501748 662386
rect 501696 662322 501748 662328
rect 512644 662380 512696 662386
rect 512644 662322 512696 662328
rect 463792 662244 463844 662250
rect 463792 662186 463844 662192
rect 463792 658436 463844 658442
rect 463792 658378 463844 658384
rect 491392 658436 491444 658442
rect 491392 658378 491444 658384
rect 462964 658300 463016 658306
rect 462964 658242 463016 658248
rect 462976 634710 463004 658242
rect 463804 654134 463832 658378
rect 464620 658368 464672 658374
rect 464620 658310 464672 658316
rect 464632 656948 464660 658310
rect 474280 658300 474332 658306
rect 474280 658242 474332 658248
rect 485044 658300 485096 658306
rect 485044 658242 485096 658248
rect 474292 656948 474320 658242
rect 483966 656254 484072 656282
rect 464436 655716 464488 655722
rect 464436 655658 464488 655664
rect 463804 654106 464200 654134
rect 464172 637786 464200 654106
rect 464448 648009 464476 655658
rect 464434 648000 464490 648009
rect 464434 647935 464490 647944
rect 464172 637758 464646 637786
rect 474292 634710 474320 637092
rect 483952 634778 483980 637092
rect 484044 634778 484072 656254
rect 483940 634772 483992 634778
rect 483940 634714 483992 634720
rect 484032 634772 484084 634778
rect 484032 634714 484084 634720
rect 485056 634710 485084 658242
rect 485780 655648 485832 655654
rect 485780 655590 485832 655596
rect 485792 646785 485820 655590
rect 489828 655580 489880 655586
rect 489828 655522 489880 655528
rect 489840 647465 489868 655522
rect 491404 654134 491432 658378
rect 502248 658368 502300 658374
rect 502248 658310 502300 658316
rect 512644 658368 512696 658374
rect 512644 658310 512696 658316
rect 492588 658300 492640 658306
rect 492588 658242 492640 658248
rect 492600 656948 492628 658242
rect 502260 656948 502288 658310
rect 511934 656266 512132 656282
rect 511934 656260 512144 656266
rect 511934 656254 512092 656260
rect 512092 656202 512144 656208
rect 491404 654106 492168 654134
rect 489826 647456 489882 647465
rect 489826 647391 489882 647400
rect 485778 646776 485834 646785
rect 485778 646711 485834 646720
rect 492140 637786 492168 654106
rect 492140 637758 492614 637786
rect 502260 634710 502288 637092
rect 511920 634778 511948 637092
rect 511908 634772 511960 634778
rect 511908 634714 511960 634720
rect 512656 634710 512684 658310
rect 514024 656260 514076 656266
rect 514024 656202 514076 656208
rect 513380 655716 513432 655722
rect 513380 655658 513432 655664
rect 513392 646785 513420 655658
rect 513378 646776 513434 646785
rect 513378 646711 513434 646720
rect 514036 634778 514064 656202
rect 514024 634772 514076 634778
rect 514024 634714 514076 634720
rect 462964 634704 463016 634710
rect 462964 634646 463016 634652
rect 474280 634704 474332 634710
rect 474280 634646 474332 634652
rect 485044 634704 485096 634710
rect 485044 634646 485096 634652
rect 502248 634704 502300 634710
rect 502248 634646 502300 634652
rect 512644 634704 512696 634710
rect 512644 634646 512696 634652
rect 492036 632324 492088 632330
rect 492036 632266 492088 632272
rect 512736 632324 512788 632330
rect 512736 632266 512788 632272
rect 473360 632256 473412 632262
rect 473360 632198 473412 632204
rect 483480 632256 483532 632262
rect 483480 632198 483532 632204
rect 464344 632188 464396 632194
rect 464344 632130 464396 632136
rect 464356 629898 464384 632130
rect 464048 629870 464384 629898
rect 473372 629898 473400 632198
rect 483020 632120 483072 632126
rect 483020 632062 483072 632068
rect 483032 629898 483060 632062
rect 473372 629870 473708 629898
rect 483032 629870 483368 629898
rect 483492 610722 483520 632198
rect 483664 632188 483716 632194
rect 483664 632130 483716 632136
rect 483676 611794 483704 632130
rect 485044 632120 485096 632126
rect 485044 632062 485096 632068
rect 483664 611788 483716 611794
rect 483664 611730 483716 611736
rect 483368 610694 483520 610722
rect 463712 610014 464048 610042
rect 473708 610014 474044 610042
rect 463712 608462 463740 610014
rect 474016 608598 474044 610014
rect 485056 608598 485084 632062
rect 492048 629884 492076 632266
rect 501696 632256 501748 632262
rect 501696 632198 501748 632204
rect 501708 629884 501736 632198
rect 511448 632188 511500 632194
rect 511448 632130 511500 632136
rect 511356 632120 511408 632126
rect 511356 632062 511408 632068
rect 511368 629884 511396 632062
rect 489826 620256 489882 620265
rect 489826 620191 489882 620200
rect 485778 619576 485834 619585
rect 485778 619511 485834 619520
rect 485792 611250 485820 619511
rect 489840 611318 489868 620191
rect 491668 611788 491720 611794
rect 491668 611730 491720 611736
rect 489828 611312 489880 611318
rect 489828 611254 489880 611260
rect 485780 611244 485832 611250
rect 485780 611186 485832 611192
rect 491680 610722 491708 611730
rect 511460 610722 511488 632130
rect 512644 632120 512696 632126
rect 512644 632062 512696 632068
rect 491680 610694 492062 610722
rect 511382 610694 511488 610722
rect 501708 608598 501736 610028
rect 512656 608598 512684 632062
rect 512748 611794 512776 632266
rect 513378 619576 513434 619585
rect 513378 619511 513434 619520
rect 512736 611788 512788 611794
rect 512736 611730 512788 611736
rect 513392 611182 513420 619511
rect 513380 611176 513432 611182
rect 513380 611118 513432 611124
rect 474004 608592 474056 608598
rect 474004 608534 474056 608540
rect 485044 608592 485096 608598
rect 485044 608534 485096 608540
rect 501696 608592 501748 608598
rect 501696 608534 501748 608540
rect 512644 608592 512696 608598
rect 512644 608534 512696 608540
rect 463700 608456 463752 608462
rect 463700 608398 463752 608404
rect 462964 604648 463016 604654
rect 462964 604590 463016 604596
rect 474280 604648 474332 604654
rect 474280 604590 474332 604596
rect 491392 604648 491444 604654
rect 491392 604590 491444 604596
rect 462976 580922 463004 604590
rect 463792 604580 463844 604586
rect 463792 604522 463844 604528
rect 463804 596174 463832 604522
rect 464620 604512 464672 604518
rect 464620 604454 464672 604460
rect 464632 602956 464660 604454
rect 474292 602956 474320 604590
rect 485044 604512 485096 604518
rect 485044 604454 485096 604460
rect 483966 602262 484072 602290
rect 463804 596146 464200 596174
rect 464172 583794 464200 596146
rect 464172 583766 464646 583794
rect 474292 580922 474320 583100
rect 483952 580990 483980 583100
rect 484044 580990 484072 602262
rect 483940 580984 483992 580990
rect 483940 580926 483992 580932
rect 484032 580984 484084 580990
rect 484032 580926 484084 580932
rect 485056 580922 485084 604454
rect 485780 601792 485832 601798
rect 485780 601734 485832 601740
rect 485792 592793 485820 601734
rect 489828 601724 489880 601730
rect 489828 601666 489880 601672
rect 489840 593473 489868 601666
rect 491404 596174 491432 604590
rect 502248 604580 502300 604586
rect 502248 604522 502300 604528
rect 512644 604580 512696 604586
rect 512644 604522 512696 604528
rect 492588 604512 492640 604518
rect 492588 604454 492640 604460
rect 492600 602956 492628 604454
rect 502260 602956 502288 604522
rect 511934 602274 512132 602290
rect 511934 602268 512144 602274
rect 511934 602262 512092 602268
rect 512092 602210 512144 602216
rect 491404 596146 492168 596174
rect 489826 593464 489882 593473
rect 489826 593399 489882 593408
rect 485778 592784 485834 592793
rect 485778 592719 485834 592728
rect 492140 583794 492168 596146
rect 492140 583766 492614 583794
rect 502260 580922 502288 583100
rect 511920 580990 511948 583100
rect 511908 580984 511960 580990
rect 511908 580926 511960 580932
rect 512656 580922 512684 604522
rect 514024 602268 514076 602274
rect 514024 602210 514076 602216
rect 513380 601860 513432 601866
rect 513380 601802 513432 601808
rect 513392 592793 513420 601802
rect 513378 592784 513434 592793
rect 513378 592719 513434 592728
rect 514036 580990 514064 602210
rect 514024 580984 514076 580990
rect 514024 580926 514076 580932
rect 462964 580916 463016 580922
rect 462964 580858 463016 580864
rect 474280 580916 474332 580922
rect 474280 580858 474332 580864
rect 485044 580916 485096 580922
rect 485044 580858 485096 580864
rect 502248 580916 502300 580922
rect 502248 580858 502300 580864
rect 512644 580916 512696 580922
rect 512644 580858 512696 580864
rect 492036 578468 492088 578474
rect 492036 578410 492088 578416
rect 512736 578468 512788 578474
rect 512736 578410 512788 578416
rect 473544 578400 473596 578406
rect 473544 578342 473596 578348
rect 483480 578400 483532 578406
rect 483480 578342 483532 578348
rect 464344 578332 464396 578338
rect 464344 578274 464396 578280
rect 464356 575906 464384 578274
rect 464048 575878 464384 575906
rect 473556 575906 473584 578342
rect 483204 578264 483256 578270
rect 483204 578206 483256 578212
rect 483216 575906 483244 578206
rect 473556 575878 473708 575906
rect 483216 575878 483368 575906
rect 483492 556730 483520 578342
rect 483664 578332 483716 578338
rect 483664 578274 483716 578280
rect 483676 558210 483704 578274
rect 485044 578264 485096 578270
rect 485044 578206 485096 578212
rect 483664 558204 483716 558210
rect 483664 558146 483716 558152
rect 483368 556702 483520 556730
rect 463712 556022 464048 556050
rect 473708 556022 474044 556050
rect 463712 554606 463740 556022
rect 474016 554742 474044 556022
rect 485056 554742 485084 578206
rect 492048 575892 492076 578410
rect 501696 578400 501748 578406
rect 501696 578342 501748 578348
rect 501708 575892 501736 578342
rect 511448 578332 511500 578338
rect 511448 578274 511500 578280
rect 511356 578264 511408 578270
rect 511356 578206 511408 578212
rect 511368 575892 511396 578206
rect 489826 566264 489882 566273
rect 489826 566199 489882 566208
rect 485778 565584 485834 565593
rect 485778 565519 485834 565528
rect 485792 557462 485820 565519
rect 489840 557530 489868 566199
rect 491668 558204 491720 558210
rect 491668 558146 491720 558152
rect 489828 557524 489880 557530
rect 489828 557466 489880 557472
rect 485780 557456 485832 557462
rect 485780 557398 485832 557404
rect 491680 556730 491708 558146
rect 511460 556730 511488 578274
rect 512644 578264 512696 578270
rect 512644 578206 512696 578212
rect 491680 556702 492062 556730
rect 511382 556702 511488 556730
rect 501708 554742 501736 556036
rect 512656 554742 512684 578206
rect 512748 558210 512776 578410
rect 513378 565584 513434 565593
rect 513378 565519 513434 565528
rect 512736 558204 512788 558210
rect 512736 558146 512788 558152
rect 513392 557394 513420 565519
rect 513380 557388 513432 557394
rect 513380 557330 513432 557336
rect 474004 554736 474056 554742
rect 474004 554678 474056 554684
rect 485044 554736 485096 554742
rect 485044 554678 485096 554684
rect 501696 554736 501748 554742
rect 501696 554678 501748 554684
rect 512644 554736 512696 554742
rect 512644 554678 512696 554684
rect 463700 554600 463752 554606
rect 463700 554542 463752 554548
rect 463792 550860 463844 550866
rect 463792 550802 463844 550808
rect 462964 550656 463016 550662
rect 462964 550598 463016 550604
rect 462976 527066 463004 550598
rect 463804 538214 463832 550802
rect 491392 550792 491444 550798
rect 491392 550734 491444 550740
rect 464620 550724 464672 550730
rect 464620 550666 464672 550672
rect 464632 548964 464660 550666
rect 474280 550656 474332 550662
rect 474280 550598 474332 550604
rect 485044 550656 485096 550662
rect 485044 550598 485096 550604
rect 474292 548964 474320 550598
rect 483966 548270 484072 548298
rect 463804 538186 464200 538214
rect 464172 529666 464200 538186
rect 464172 529638 464646 529666
rect 474292 527066 474320 529108
rect 483952 527134 483980 529108
rect 484044 527134 484072 548270
rect 483940 527128 483992 527134
rect 483940 527070 483992 527076
rect 484032 527128 484084 527134
rect 484032 527070 484084 527076
rect 485056 527066 485084 550598
rect 489826 539472 489882 539481
rect 489826 539407 489882 539416
rect 485778 538792 485834 538801
rect 485778 538727 485834 538736
rect 485792 529854 485820 538727
rect 489840 529922 489868 539407
rect 491404 538214 491432 550734
rect 502248 550724 502300 550730
rect 502248 550666 502300 550672
rect 492588 550656 492640 550662
rect 492588 550598 492640 550604
rect 492600 548964 492628 550598
rect 502260 548964 502288 550666
rect 514024 550656 514076 550662
rect 514024 550598 514076 550604
rect 511934 548270 512132 548298
rect 491404 538186 492168 538214
rect 489828 529916 489880 529922
rect 489828 529858 489880 529864
rect 485780 529848 485832 529854
rect 485780 529790 485832 529796
rect 492140 529666 492168 538186
rect 492140 529638 492614 529666
rect 502260 527066 502288 529108
rect 511920 527134 511948 529108
rect 512104 527134 512132 548270
rect 513378 538792 513434 538801
rect 513378 538727 513434 538736
rect 513392 529786 513420 538727
rect 513380 529780 513432 529786
rect 513380 529722 513432 529728
rect 511908 527128 511960 527134
rect 511908 527070 511960 527076
rect 512092 527128 512144 527134
rect 512092 527070 512144 527076
rect 514036 527066 514064 550598
rect 462964 527060 463016 527066
rect 462964 527002 463016 527008
rect 474280 527060 474332 527066
rect 474280 527002 474332 527008
rect 485044 527060 485096 527066
rect 485044 527002 485096 527008
rect 502248 527060 502300 527066
rect 502248 527002 502300 527008
rect 514024 527060 514076 527066
rect 514024 527002 514076 527008
rect 492036 523252 492088 523258
rect 492036 523194 492088 523200
rect 512736 523252 512788 523258
rect 512736 523194 512788 523200
rect 473360 523184 473412 523190
rect 473360 523126 473412 523132
rect 483480 523184 483532 523190
rect 483480 523126 483532 523132
rect 464344 523116 464396 523122
rect 464344 523058 464396 523064
rect 464356 521914 464384 523058
rect 464048 521886 464384 521914
rect 473372 521914 473400 523126
rect 483020 523048 483072 523054
rect 483020 522990 483072 522996
rect 483032 521914 483060 522990
rect 473372 521886 473708 521914
rect 483032 521886 483368 521914
rect 483492 502738 483520 523126
rect 483664 523116 483716 523122
rect 483664 523058 483716 523064
rect 483676 504354 483704 523058
rect 485044 523048 485096 523054
rect 485044 522990 485096 522996
rect 483664 504348 483716 504354
rect 483664 504290 483716 504296
rect 483368 502710 483520 502738
rect 463712 502030 464048 502058
rect 473708 502030 474044 502058
rect 463712 500818 463740 502030
rect 474016 500954 474044 502030
rect 485056 500954 485084 522990
rect 492048 521900 492076 523194
rect 501696 523184 501748 523190
rect 501696 523126 501748 523132
rect 501708 521900 501736 523126
rect 511448 523116 511500 523122
rect 511448 523058 511500 523064
rect 511356 523048 511408 523054
rect 511356 522990 511408 522996
rect 511368 521900 511396 522990
rect 485780 520328 485832 520334
rect 485780 520270 485832 520276
rect 489828 520328 489880 520334
rect 489828 520270 489880 520276
rect 485792 511601 485820 520270
rect 489840 512281 489868 520270
rect 489826 512272 489882 512281
rect 489826 512207 489882 512216
rect 485778 511592 485834 511601
rect 485778 511527 485834 511536
rect 491668 504348 491720 504354
rect 491668 504290 491720 504296
rect 491680 502738 491708 504290
rect 511460 502738 511488 523058
rect 512644 523048 512696 523054
rect 512644 522990 512696 522996
rect 491680 502710 492062 502738
rect 511382 502710 511488 502738
rect 501708 500954 501736 502044
rect 512656 500954 512684 522990
rect 512748 504354 512776 523194
rect 513378 511592 513434 511601
rect 513378 511527 513434 511536
rect 512736 504348 512788 504354
rect 512736 504290 512788 504296
rect 513392 503674 513420 511527
rect 513380 503668 513432 503674
rect 513380 503610 513432 503616
rect 474004 500948 474056 500954
rect 474004 500890 474056 500896
rect 485044 500948 485096 500954
rect 485044 500890 485096 500896
rect 501696 500948 501748 500954
rect 501696 500890 501748 500896
rect 512644 500948 512696 500954
rect 512644 500890 512696 500896
rect 463700 500812 463752 500818
rect 463700 500754 463752 500760
rect 464160 497004 464212 497010
rect 464160 496946 464212 496952
rect 485044 497004 485096 497010
rect 485044 496946 485096 496952
rect 492588 497004 492640 497010
rect 492588 496946 492640 496952
rect 462964 496868 463016 496874
rect 462964 496810 463016 496816
rect 462976 473278 463004 496810
rect 464172 475674 464200 496946
rect 464620 496936 464672 496942
rect 464620 496878 464672 496884
rect 464632 494972 464660 496878
rect 474280 496868 474332 496874
rect 474280 496810 474332 496816
rect 474292 494972 474320 496810
rect 483966 494278 484072 494306
rect 464172 475646 464646 475674
rect 474292 473278 474320 475116
rect 483952 473346 483980 475116
rect 484044 473346 484072 494278
rect 483940 473340 483992 473346
rect 483940 473282 483992 473288
rect 484032 473340 484084 473346
rect 484032 473282 484084 473288
rect 485056 473278 485084 496946
rect 492128 496868 492180 496874
rect 492128 496810 492180 496816
rect 489826 485480 489882 485489
rect 489826 485415 489882 485424
rect 485778 484800 485834 484809
rect 485778 484735 485834 484744
rect 485792 475930 485820 484735
rect 489840 476066 489868 485415
rect 489828 476060 489880 476066
rect 489828 476002 489880 476008
rect 485780 475924 485832 475930
rect 485780 475866 485832 475872
rect 492140 475674 492168 496810
rect 492600 494972 492628 496946
rect 502248 496936 502300 496942
rect 502248 496878 502300 496884
rect 514024 496936 514076 496942
rect 514024 496878 514076 496884
rect 502260 494972 502288 496878
rect 511934 494278 512132 494306
rect 492140 475646 492614 475674
rect 502260 473278 502288 475116
rect 511920 473346 511948 475116
rect 512104 473346 512132 494278
rect 513378 484800 513434 484809
rect 513378 484735 513434 484744
rect 513392 475998 513420 484735
rect 513380 475992 513432 475998
rect 513380 475934 513432 475940
rect 511908 473340 511960 473346
rect 511908 473282 511960 473288
rect 512092 473340 512144 473346
rect 512092 473282 512144 473288
rect 514036 473278 514064 496878
rect 462964 473272 463016 473278
rect 462964 473214 463016 473220
rect 474280 473272 474332 473278
rect 474280 473214 474332 473220
rect 485044 473272 485096 473278
rect 485044 473214 485096 473220
rect 502248 473272 502300 473278
rect 502248 473214 502300 473220
rect 514024 473272 514076 473278
rect 514024 473214 514076 473220
rect 473360 469396 473412 469402
rect 473360 469338 473412 469344
rect 483480 469396 483532 469402
rect 483480 469338 483532 469344
rect 501696 469396 501748 469402
rect 501696 469338 501748 469344
rect 511448 469396 511500 469402
rect 511448 469338 511500 469344
rect 464344 469328 464396 469334
rect 464344 469270 464396 469276
rect 464356 467922 464384 469270
rect 464048 467894 464384 467922
rect 473372 467922 473400 469338
rect 483020 469260 483072 469266
rect 483020 469202 483072 469208
rect 483032 467922 483060 469202
rect 473372 467894 473708 467922
rect 483032 467894 483368 467922
rect 483492 448746 483520 469338
rect 483664 469328 483716 469334
rect 483664 469270 483716 469276
rect 492036 469328 492088 469334
rect 492036 469270 492088 469276
rect 483676 450362 483704 469270
rect 485044 469260 485096 469266
rect 485044 469202 485096 469208
rect 483664 450356 483716 450362
rect 483664 450298 483716 450304
rect 483368 448718 483520 448746
rect 463712 448038 464048 448066
rect 473708 448038 474044 448066
rect 463712 445602 463740 448038
rect 474016 445738 474044 448038
rect 485056 445738 485084 469202
rect 492048 467908 492076 469270
rect 501708 467908 501736 469338
rect 511356 469260 511408 469266
rect 511356 469202 511408 469208
rect 511368 467908 511396 469202
rect 485780 466540 485832 466546
rect 485780 466482 485832 466488
rect 485792 457609 485820 466482
rect 489828 466472 489880 466478
rect 489828 466414 489880 466420
rect 489840 458289 489868 466414
rect 489826 458280 489882 458289
rect 489826 458215 489882 458224
rect 485778 457600 485834 457609
rect 485778 457535 485834 457544
rect 491668 450356 491720 450362
rect 491668 450298 491720 450304
rect 491680 448746 491708 450298
rect 511460 448746 511488 469338
rect 512736 469328 512788 469334
rect 512736 469270 512788 469276
rect 512644 469260 512696 469266
rect 512644 469202 512696 469208
rect 491680 448718 492062 448746
rect 511382 448718 511488 448746
rect 501708 445738 501736 448052
rect 512656 445738 512684 469202
rect 512748 450498 512776 469270
rect 513380 466608 513432 466614
rect 513380 466550 513432 466556
rect 513392 457609 513420 466550
rect 513378 457600 513434 457609
rect 513378 457535 513434 457544
rect 512736 450492 512788 450498
rect 512736 450434 512788 450440
rect 474004 445732 474056 445738
rect 474004 445674 474056 445680
rect 485044 445732 485096 445738
rect 485044 445674 485096 445680
rect 501696 445732 501748 445738
rect 501696 445674 501748 445680
rect 512644 445732 512696 445738
rect 512644 445674 512696 445680
rect 463700 445596 463752 445602
rect 463700 445538 463752 445544
rect 462964 443148 463016 443154
rect 462964 443090 463016 443096
rect 474280 443148 474332 443154
rect 474280 443090 474332 443096
rect 485044 443148 485096 443154
rect 485044 443090 485096 443096
rect 492588 443148 492640 443154
rect 492588 443090 492640 443096
rect 462976 419422 463004 443090
rect 463792 443080 463844 443086
rect 463792 443022 463844 443028
rect 463804 441614 463832 443022
rect 464620 443012 464672 443018
rect 464620 442954 464672 442960
rect 463804 441586 464200 441614
rect 464172 421682 464200 441586
rect 464632 440980 464660 442954
rect 474292 440980 474320 443090
rect 483966 440286 484072 440314
rect 464172 421654 464646 421682
rect 474292 419422 474320 421124
rect 483952 419490 483980 421124
rect 484044 419490 484072 440286
rect 483940 419484 483992 419490
rect 483940 419426 483992 419432
rect 484032 419484 484084 419490
rect 484032 419426 484084 419432
rect 485056 419422 485084 443090
rect 491392 443012 491444 443018
rect 491392 442954 491444 442960
rect 491404 441614 491432 442954
rect 491404 441586 492168 441614
rect 485780 440292 485832 440298
rect 485780 440234 485832 440240
rect 489828 440292 489880 440298
rect 489828 440234 489880 440240
rect 485792 430817 485820 440234
rect 489840 431497 489868 440234
rect 489826 431488 489882 431497
rect 489826 431423 489882 431432
rect 485778 430808 485834 430817
rect 485778 430743 485834 430752
rect 492140 421682 492168 441586
rect 492600 440980 492628 443090
rect 502248 443080 502300 443086
rect 502248 443022 502300 443028
rect 514024 443080 514076 443086
rect 514024 443022 514076 443028
rect 502260 440980 502288 443022
rect 511934 440286 512132 440314
rect 492140 421654 492614 421682
rect 502260 419422 502288 421124
rect 511920 419490 511948 421124
rect 512104 419490 512132 440286
rect 513378 430808 513434 430817
rect 513378 430743 513434 430752
rect 513392 422278 513420 430743
rect 513380 422272 513432 422278
rect 513380 422214 513432 422220
rect 511908 419484 511960 419490
rect 511908 419426 511960 419432
rect 512092 419484 512144 419490
rect 512092 419426 512144 419432
rect 514036 419422 514064 443022
rect 462964 419416 463016 419422
rect 462964 419358 463016 419364
rect 474280 419416 474332 419422
rect 474280 419358 474332 419364
rect 485044 419416 485096 419422
rect 485044 419358 485096 419364
rect 502248 419416 502300 419422
rect 502248 419358 502300 419364
rect 514024 419416 514076 419422
rect 514024 419358 514076 419364
rect 473360 415608 473412 415614
rect 473360 415550 473412 415556
rect 483480 415608 483532 415614
rect 483480 415550 483532 415556
rect 501696 415608 501748 415614
rect 501696 415550 501748 415556
rect 511448 415608 511500 415614
rect 511448 415550 511500 415556
rect 464344 415540 464396 415546
rect 464344 415482 464396 415488
rect 464356 413930 464384 415482
rect 464048 413902 464384 413930
rect 473372 413930 473400 415550
rect 483020 415472 483072 415478
rect 483020 415414 483072 415420
rect 483032 413930 483060 415414
rect 473372 413902 473708 413930
rect 483032 413902 483368 413930
rect 483492 394754 483520 415550
rect 483664 415540 483716 415546
rect 483664 415482 483716 415488
rect 492036 415540 492088 415546
rect 492036 415482 492088 415488
rect 483676 395078 483704 415482
rect 485044 415472 485096 415478
rect 485044 415414 485096 415420
rect 483664 395072 483716 395078
rect 483664 395014 483716 395020
rect 483368 394726 483520 394754
rect 463804 394046 464048 394074
rect 473708 394046 474044 394074
rect 463804 391814 463832 394046
rect 474016 391950 474044 394046
rect 485056 391950 485084 415414
rect 492048 413916 492076 415482
rect 501708 413916 501736 415550
rect 511356 415472 511408 415478
rect 511356 415414 511408 415420
rect 511368 413916 511396 415414
rect 489826 404288 489882 404297
rect 489826 404223 489882 404232
rect 485778 403608 485834 403617
rect 485778 403543 485834 403552
rect 485792 394534 485820 403543
rect 489840 394670 489868 404223
rect 491668 395072 491720 395078
rect 491668 395014 491720 395020
rect 491680 394754 491708 395014
rect 511460 394754 511488 415550
rect 512736 415540 512788 415546
rect 512736 415482 512788 415488
rect 512644 415472 512696 415478
rect 512644 415414 512696 415420
rect 491680 394726 492062 394754
rect 511382 394726 511488 394754
rect 489828 394664 489880 394670
rect 489828 394606 489880 394612
rect 485780 394528 485832 394534
rect 485780 394470 485832 394476
rect 501708 391950 501736 394060
rect 512656 391950 512684 415414
rect 512748 395078 512776 415482
rect 513378 403608 513434 403617
rect 513378 403543 513434 403552
rect 512736 395072 512788 395078
rect 512736 395014 512788 395020
rect 513392 394602 513420 403543
rect 513380 394596 513432 394602
rect 513380 394538 513432 394544
rect 474004 391944 474056 391950
rect 474004 391886 474056 391892
rect 485044 391944 485096 391950
rect 485044 391886 485096 391892
rect 501696 391944 501748 391950
rect 501696 391886 501748 391892
rect 512644 391944 512696 391950
rect 512644 391886 512696 391892
rect 463792 391808 463844 391814
rect 463792 391750 463844 391756
rect 463792 389360 463844 389366
rect 463792 389302 463844 389308
rect 491392 389360 491444 389366
rect 491392 389302 491444 389308
rect 462964 389224 463016 389230
rect 462964 389166 463016 389172
rect 462976 365634 463004 389166
rect 463804 383654 463832 389302
rect 464620 389292 464672 389298
rect 464620 389234 464672 389240
rect 464632 386852 464660 389234
rect 474280 389224 474332 389230
rect 474280 389166 474332 389172
rect 485044 389224 485096 389230
rect 485044 389166 485096 389172
rect 474292 386852 474320 389166
rect 483966 386294 484072 386322
rect 463804 383626 464200 383654
rect 464172 367690 464200 383626
rect 464172 367662 464646 367690
rect 474292 365634 474320 367132
rect 483952 365702 483980 367132
rect 484044 365702 484072 386294
rect 483940 365696 483992 365702
rect 483940 365638 483992 365644
rect 484032 365696 484084 365702
rect 484032 365638 484084 365644
rect 485056 365634 485084 389166
rect 485780 386504 485832 386510
rect 485780 386446 485832 386452
rect 485792 376825 485820 386446
rect 489828 386436 489880 386442
rect 489828 386378 489880 386384
rect 489840 377505 489868 386378
rect 491404 383654 491432 389302
rect 502248 389292 502300 389298
rect 502248 389234 502300 389240
rect 514024 389292 514076 389298
rect 514024 389234 514076 389240
rect 492588 389224 492640 389230
rect 492588 389166 492640 389172
rect 492600 386852 492628 389166
rect 502260 386852 502288 389234
rect 513380 386572 513432 386578
rect 513380 386514 513432 386520
rect 511934 386294 512132 386322
rect 491404 383626 492168 383654
rect 489826 377496 489882 377505
rect 489826 377431 489882 377440
rect 485778 376816 485834 376825
rect 485778 376751 485834 376760
rect 492140 367690 492168 383626
rect 492140 367662 492614 367690
rect 502260 365634 502288 367132
rect 511920 365702 511948 367132
rect 512104 365702 512132 386294
rect 513392 376825 513420 386514
rect 513378 376816 513434 376825
rect 513378 376751 513434 376760
rect 511908 365696 511960 365702
rect 511908 365638 511960 365644
rect 512092 365696 512144 365702
rect 512092 365638 512144 365644
rect 514036 365634 514064 389234
rect 462964 365628 463016 365634
rect 462964 365570 463016 365576
rect 474280 365628 474332 365634
rect 474280 365570 474332 365576
rect 485044 365628 485096 365634
rect 485044 365570 485096 365576
rect 502248 365628 502300 365634
rect 502248 365570 502300 365576
rect 514024 365628 514076 365634
rect 514024 365570 514076 365576
rect 473360 361752 473412 361758
rect 473360 361694 473412 361700
rect 483480 361752 483532 361758
rect 483480 361694 483532 361700
rect 501696 361752 501748 361758
rect 501696 361694 501748 361700
rect 511448 361752 511500 361758
rect 511448 361694 511500 361700
rect 464344 361684 464396 361690
rect 464344 361626 464396 361632
rect 464356 359938 464384 361626
rect 464048 359910 464384 359938
rect 473372 359938 473400 361694
rect 483020 361616 483072 361622
rect 483020 361558 483072 361564
rect 483032 359938 483060 361558
rect 473372 359910 473708 359938
rect 483032 359910 483368 359938
rect 483492 340762 483520 361694
rect 483664 361684 483716 361690
rect 483664 361626 483716 361632
rect 492036 361684 492088 361690
rect 492036 361626 492088 361632
rect 483676 341426 483704 361626
rect 485044 361616 485096 361622
rect 485044 361558 485096 361564
rect 483664 341420 483716 341426
rect 483664 341362 483716 341368
rect 483368 340734 483520 340762
rect 463712 340054 464048 340082
rect 473708 340054 474044 340082
rect 463712 337958 463740 340054
rect 474016 338094 474044 340054
rect 485056 338094 485084 361558
rect 492048 359924 492076 361626
rect 501708 359924 501736 361694
rect 511356 361616 511408 361622
rect 511356 361558 511408 361564
rect 511368 359924 511396 361558
rect 489826 350296 489882 350305
rect 489826 350231 489882 350240
rect 485778 349616 485834 349625
rect 485778 349551 485834 349560
rect 485792 340814 485820 349551
rect 489840 340882 489868 350231
rect 491668 341420 491720 341426
rect 491668 341362 491720 341368
rect 489828 340876 489880 340882
rect 489828 340818 489880 340824
rect 485780 340808 485832 340814
rect 485780 340750 485832 340756
rect 491680 340762 491708 341362
rect 511460 340762 511488 361694
rect 512736 361684 512788 361690
rect 512736 361626 512788 361632
rect 512644 361616 512696 361622
rect 512644 361558 512696 361564
rect 491680 340734 492062 340762
rect 511382 340734 511488 340762
rect 501708 338094 501736 340068
rect 512656 338094 512684 361558
rect 512748 341970 512776 361626
rect 513378 349616 513434 349625
rect 513378 349551 513434 349560
rect 512736 341964 512788 341970
rect 512736 341906 512788 341912
rect 513392 340746 513420 349551
rect 513380 340740 513432 340746
rect 513380 340682 513432 340688
rect 474004 338088 474056 338094
rect 474004 338030 474056 338036
rect 485044 338088 485096 338094
rect 485044 338030 485096 338036
rect 501696 338088 501748 338094
rect 501696 338030 501748 338036
rect 512644 338088 512696 338094
rect 512644 338030 512696 338036
rect 463700 337952 463752 337958
rect 463700 337894 463752 337900
rect 463792 335504 463844 335510
rect 463792 335446 463844 335452
rect 491392 335504 491444 335510
rect 491392 335446 491444 335452
rect 462964 335368 463016 335374
rect 462964 335310 463016 335316
rect 462976 311778 463004 335310
rect 463804 325694 463832 335446
rect 464620 335436 464672 335442
rect 464620 335378 464672 335384
rect 464632 332860 464660 335378
rect 474280 335368 474332 335374
rect 474280 335310 474332 335316
rect 485044 335368 485096 335374
rect 485044 335310 485096 335316
rect 474292 332860 474320 335310
rect 483966 332302 484072 332330
rect 463804 325666 464200 325694
rect 464172 313698 464200 325666
rect 464172 313670 464646 313698
rect 474292 311778 474320 313140
rect 483952 311846 483980 313140
rect 484044 311846 484072 332302
rect 483940 311840 483992 311846
rect 483940 311782 483992 311788
rect 484032 311840 484084 311846
rect 484032 311782 484084 311788
rect 485056 311778 485084 335310
rect 489828 331288 489880 331294
rect 489828 331230 489880 331236
rect 489840 324057 489868 331230
rect 491404 325694 491432 335446
rect 502248 335436 502300 335442
rect 502248 335378 502300 335384
rect 512644 335436 512696 335442
rect 512644 335378 512696 335384
rect 492588 335368 492640 335374
rect 492588 335310 492640 335316
rect 492600 332860 492628 335310
rect 502260 332860 502288 335378
rect 511816 335368 511868 335374
rect 511816 335310 511868 335316
rect 511828 332874 511856 335310
rect 511828 332846 511934 332874
rect 491404 325666 492168 325694
rect 489826 324048 489882 324057
rect 489826 323983 489882 323992
rect 485778 322144 485834 322153
rect 485778 322079 485834 322088
rect 485792 314634 485820 322079
rect 485780 314628 485832 314634
rect 485780 314570 485832 314576
rect 492140 313698 492168 325666
rect 492140 313670 492614 313698
rect 502260 311778 502288 313140
rect 511920 311846 511948 313140
rect 511908 311840 511960 311846
rect 511908 311782 511960 311788
rect 512656 311778 512684 335378
rect 514024 335368 514076 335374
rect 514024 335310 514076 335316
rect 513378 322144 513434 322153
rect 513378 322079 513434 322088
rect 513392 314566 513420 322079
rect 513380 314560 513432 314566
rect 513380 314502 513432 314508
rect 514036 311846 514064 335310
rect 514024 311840 514076 311846
rect 514024 311782 514076 311788
rect 462964 311772 463016 311778
rect 462964 311714 463016 311720
rect 474280 311772 474332 311778
rect 474280 311714 474332 311720
rect 485044 311772 485096 311778
rect 485044 311714 485096 311720
rect 502248 311772 502300 311778
rect 502248 311714 502300 311720
rect 512644 311772 512696 311778
rect 512644 311714 512696 311720
rect 473544 307964 473596 307970
rect 473544 307906 473596 307912
rect 483480 307964 483532 307970
rect 483480 307906 483532 307912
rect 501696 307964 501748 307970
rect 501696 307906 501748 307912
rect 511448 307964 511500 307970
rect 511448 307906 511500 307912
rect 464344 307896 464396 307902
rect 464344 307838 464396 307844
rect 464356 305946 464384 307838
rect 464048 305918 464384 305946
rect 473556 305946 473584 307906
rect 483204 307828 483256 307834
rect 483204 307770 483256 307776
rect 483216 305946 483244 307770
rect 473556 305918 473708 305946
rect 483216 305918 483368 305946
rect 483492 286770 483520 307906
rect 483664 307896 483716 307902
rect 483664 307838 483716 307844
rect 492036 307896 492088 307902
rect 492036 307838 492088 307844
rect 483676 287434 483704 307838
rect 485044 307828 485096 307834
rect 485044 307770 485096 307776
rect 483664 287428 483716 287434
rect 483664 287370 483716 287376
rect 483368 286742 483520 286770
rect 463712 286062 464048 286090
rect 473708 286062 474044 286090
rect 463712 284170 463740 286062
rect 474016 284306 474044 286062
rect 485056 284306 485084 307770
rect 492048 305932 492076 307838
rect 501708 305932 501736 307906
rect 511356 307828 511408 307834
rect 511356 307770 511408 307776
rect 511368 305932 511396 307770
rect 489826 296304 489882 296313
rect 489826 296239 489882 296248
rect 485778 295624 485834 295633
rect 485778 295559 485834 295568
rect 485792 286958 485820 295559
rect 489840 287026 489868 296239
rect 491668 287428 491720 287434
rect 491668 287370 491720 287376
rect 489828 287020 489880 287026
rect 489828 286962 489880 286968
rect 485780 286952 485832 286958
rect 485780 286894 485832 286900
rect 491680 286770 491708 287370
rect 511460 286770 511488 307906
rect 512736 307896 512788 307902
rect 512736 307838 512788 307844
rect 512644 307828 512696 307834
rect 512644 307770 512696 307776
rect 491680 286742 492062 286770
rect 511382 286742 511488 286770
rect 501708 284306 501736 286076
rect 512656 284306 512684 307770
rect 512748 287570 512776 307838
rect 513378 295624 513434 295633
rect 513378 295559 513434 295568
rect 512736 287564 512788 287570
rect 512736 287506 512788 287512
rect 513392 286890 513420 295559
rect 513380 286884 513432 286890
rect 513380 286826 513432 286832
rect 474004 284300 474056 284306
rect 474004 284242 474056 284248
rect 485044 284300 485096 284306
rect 485044 284242 485096 284248
rect 501696 284300 501748 284306
rect 501696 284242 501748 284248
rect 512644 284300 512696 284306
rect 512644 284242 512696 284248
rect 463700 284164 463752 284170
rect 463700 284106 463752 284112
rect 463792 280424 463844 280430
rect 463792 280366 463844 280372
rect 462964 280220 463016 280226
rect 462964 280162 463016 280168
rect 462976 256630 463004 280162
rect 463804 267734 463832 280366
rect 491392 280356 491444 280362
rect 491392 280298 491444 280304
rect 464620 280288 464672 280294
rect 464620 280230 464672 280236
rect 464632 278868 464660 280230
rect 474280 280220 474332 280226
rect 474280 280162 474332 280168
rect 485044 280220 485096 280226
rect 485044 280162 485096 280168
rect 474292 278868 474320 280162
rect 483966 278310 484072 278338
rect 463804 267706 464200 267734
rect 464172 259706 464200 267706
rect 464172 259678 464646 259706
rect 474292 256630 474320 259148
rect 483952 256698 483980 259148
rect 484044 256698 484072 278310
rect 483940 256692 483992 256698
rect 483940 256634 483992 256640
rect 484032 256692 484084 256698
rect 484032 256634 484084 256640
rect 485056 256630 485084 280162
rect 485780 277500 485832 277506
rect 485780 277442 485832 277448
rect 485792 269113 485820 277442
rect 489828 277432 489880 277438
rect 489828 277374 489880 277380
rect 489840 269929 489868 277374
rect 489826 269920 489882 269929
rect 489826 269855 489882 269864
rect 485778 269104 485834 269113
rect 485778 269039 485834 269048
rect 491404 267734 491432 280298
rect 502248 280288 502300 280294
rect 502248 280230 502300 280236
rect 492588 280220 492640 280226
rect 492588 280162 492640 280168
rect 492600 278868 492628 280162
rect 502260 278868 502288 280230
rect 512644 280220 512696 280226
rect 512644 280162 512696 280168
rect 511934 278322 512132 278338
rect 511934 278316 512144 278322
rect 511934 278310 512092 278316
rect 512092 278258 512144 278264
rect 491404 267706 492168 267734
rect 492140 259706 492168 267706
rect 492140 259678 492614 259706
rect 502260 256630 502288 259148
rect 511920 256698 511948 259148
rect 511908 256692 511960 256698
rect 511908 256634 511960 256640
rect 512656 256630 512684 280162
rect 514024 278316 514076 278322
rect 514024 278258 514076 278264
rect 513380 277568 513432 277574
rect 513380 277510 513432 277516
rect 513392 269113 513420 277510
rect 513378 269104 513434 269113
rect 513378 269039 513434 269048
rect 514036 256698 514064 278258
rect 514024 256692 514076 256698
rect 514024 256634 514076 256640
rect 462964 256624 463016 256630
rect 462964 256566 463016 256572
rect 474280 256624 474332 256630
rect 474280 256566 474332 256572
rect 485044 256624 485096 256630
rect 485044 256566 485096 256572
rect 502248 256624 502300 256630
rect 502248 256566 502300 256572
rect 512644 256624 512696 256630
rect 512644 256566 512696 256572
rect 492036 254176 492088 254182
rect 492036 254118 492088 254124
rect 512736 254176 512788 254182
rect 512736 254118 512788 254124
rect 473360 254108 473412 254114
rect 473360 254050 473412 254056
rect 483480 254108 483532 254114
rect 483480 254050 483532 254056
rect 464344 254040 464396 254046
rect 464344 253982 464396 253988
rect 464356 251954 464384 253982
rect 464048 251926 464384 251954
rect 473372 251954 473400 254050
rect 483020 253972 483072 253978
rect 483020 253914 483072 253920
rect 483032 251954 483060 253914
rect 473372 251926 473708 251954
rect 483032 251926 483368 251954
rect 483492 232778 483520 254050
rect 483664 254040 483716 254046
rect 483664 253982 483716 253988
rect 483676 233442 483704 253982
rect 485044 253972 485096 253978
rect 485044 253914 485096 253920
rect 483664 233436 483716 233442
rect 483664 233378 483716 233384
rect 483368 232750 483520 232778
rect 463712 232070 464048 232098
rect 473708 232070 474044 232098
rect 463712 230314 463740 232070
rect 474016 230450 474044 232070
rect 485056 230450 485084 253914
rect 492048 251940 492076 254118
rect 501696 254108 501748 254114
rect 501696 254050 501748 254056
rect 501708 251940 501736 254050
rect 511448 254040 511500 254046
rect 511448 253982 511500 253988
rect 511356 253972 511408 253978
rect 511356 253914 511408 253920
rect 511368 251940 511396 253914
rect 485780 251320 485832 251326
rect 485780 251262 485832 251268
rect 485792 241641 485820 251262
rect 489828 251252 489880 251258
rect 489828 251194 489880 251200
rect 489840 242321 489868 251194
rect 489826 242312 489882 242321
rect 489826 242247 489882 242256
rect 485778 241632 485834 241641
rect 485778 241567 485834 241576
rect 491668 233436 491720 233442
rect 491668 233378 491720 233384
rect 491680 232778 491708 233378
rect 511460 232778 511488 253982
rect 512644 253972 512696 253978
rect 512644 253914 512696 253920
rect 491680 232750 492062 232778
rect 511382 232750 511488 232778
rect 501708 230450 501736 232084
rect 512656 230450 512684 253914
rect 512748 234258 512776 254118
rect 513380 251388 513432 251394
rect 513380 251330 513432 251336
rect 513392 241641 513420 251330
rect 513378 241632 513434 241641
rect 513378 241567 513434 241576
rect 512736 234252 512788 234258
rect 512736 234194 512788 234200
rect 474004 230444 474056 230450
rect 474004 230386 474056 230392
rect 485044 230444 485096 230450
rect 485044 230386 485096 230392
rect 501696 230444 501748 230450
rect 501696 230386 501748 230392
rect 512644 230444 512696 230450
rect 512644 230386 512696 230392
rect 463700 230308 463752 230314
rect 463700 230250 463752 230256
rect 462964 226500 463016 226506
rect 462964 226442 463016 226448
rect 474280 226500 474332 226506
rect 474280 226442 474332 226448
rect 492128 226500 492180 226506
rect 492128 226442 492180 226448
rect 462976 202774 463004 226442
rect 464160 226432 464212 226438
rect 464160 226374 464212 226380
rect 464172 205714 464200 226374
rect 464620 226364 464672 226370
rect 464620 226306 464672 226312
rect 464632 224876 464660 226306
rect 474292 224876 474320 226442
rect 485044 226364 485096 226370
rect 485044 226306 485096 226312
rect 483966 224318 484072 224346
rect 464172 205686 464646 205714
rect 474292 202774 474320 205020
rect 483952 202842 483980 205020
rect 484044 202842 484072 224318
rect 483940 202836 483992 202842
rect 483940 202778 483992 202784
rect 484032 202836 484084 202842
rect 484032 202778 484084 202784
rect 485056 202774 485084 226306
rect 485780 223712 485832 223718
rect 485780 223654 485832 223660
rect 485792 214713 485820 223654
rect 489828 223644 489880 223650
rect 489828 223586 489880 223592
rect 489840 215393 489868 223586
rect 489826 215384 489882 215393
rect 489826 215319 489882 215328
rect 485778 214704 485834 214713
rect 485778 214639 485834 214648
rect 492140 205714 492168 226442
rect 502248 226432 502300 226438
rect 502248 226374 502300 226380
rect 512644 226432 512696 226438
rect 512644 226374 512696 226380
rect 492588 226364 492640 226370
rect 492588 226306 492640 226312
rect 492600 224876 492628 226306
rect 502260 224876 502288 226374
rect 511934 224330 512224 224346
rect 511934 224324 512236 224330
rect 511934 224318 512184 224324
rect 512184 224266 512236 224272
rect 492140 205686 492614 205714
rect 502260 202774 502288 205020
rect 511920 202842 511948 205020
rect 511908 202836 511960 202842
rect 511908 202778 511960 202784
rect 512656 202774 512684 226374
rect 514024 224324 514076 224330
rect 514024 224266 514076 224272
rect 513380 223780 513432 223786
rect 513380 223722 513432 223728
rect 513392 214713 513420 223722
rect 513378 214704 513434 214713
rect 513378 214639 513434 214648
rect 514036 202842 514064 224266
rect 514024 202836 514076 202842
rect 514024 202778 514076 202784
rect 462964 202768 463016 202774
rect 462964 202710 463016 202716
rect 474280 202768 474332 202774
rect 474280 202710 474332 202716
rect 485044 202768 485096 202774
rect 485044 202710 485096 202716
rect 502248 202768 502300 202774
rect 502248 202710 502300 202716
rect 512644 202768 512696 202774
rect 512644 202710 512696 202716
rect 492036 200388 492088 200394
rect 492036 200330 492088 200336
rect 512736 200388 512788 200394
rect 512736 200330 512788 200336
rect 473544 200320 473596 200326
rect 473544 200262 473596 200268
rect 483480 200320 483532 200326
rect 483480 200262 483532 200268
rect 464344 200252 464396 200258
rect 464344 200194 464396 200200
rect 464356 197962 464384 200194
rect 464048 197934 464384 197962
rect 473556 197962 473584 200262
rect 483204 200184 483256 200190
rect 483204 200126 483256 200132
rect 483216 197962 483244 200126
rect 473556 197934 473708 197962
rect 483216 197934 483368 197962
rect 483492 178786 483520 200262
rect 483664 200252 483716 200258
rect 483664 200194 483716 200200
rect 483676 179722 483704 200194
rect 485044 200184 485096 200190
rect 485044 200126 485096 200132
rect 483664 179716 483716 179722
rect 483664 179658 483716 179664
rect 483368 178758 483520 178786
rect 463712 178078 464048 178106
rect 473708 178078 474044 178106
rect 463712 176526 463740 178078
rect 474016 176662 474044 178078
rect 485056 176662 485084 200126
rect 492048 197948 492076 200330
rect 501696 200320 501748 200326
rect 501696 200262 501748 200268
rect 501708 197948 501736 200262
rect 511448 200252 511500 200258
rect 511448 200194 511500 200200
rect 511356 200184 511408 200190
rect 511356 200126 511408 200132
rect 511368 197948 511396 200126
rect 489826 188320 489882 188329
rect 489826 188255 489882 188264
rect 485778 187640 485834 187649
rect 485778 187575 485834 187584
rect 485792 179314 485820 187575
rect 489840 179382 489868 188255
rect 491668 179716 491720 179722
rect 491668 179658 491720 179664
rect 489828 179376 489880 179382
rect 489828 179318 489880 179324
rect 485780 179308 485832 179314
rect 485780 179250 485832 179256
rect 491680 178786 491708 179658
rect 511460 178786 511488 200194
rect 512644 200184 512696 200190
rect 512644 200126 512696 200132
rect 491680 178758 492062 178786
rect 511382 178758 511488 178786
rect 501708 176662 501736 178092
rect 512656 176662 512684 200126
rect 512748 180266 512776 200330
rect 513378 187640 513434 187649
rect 513378 187575 513434 187584
rect 512736 180260 512788 180266
rect 512736 180202 512788 180208
rect 513392 179246 513420 187575
rect 513380 179240 513432 179246
rect 513380 179182 513432 179188
rect 474004 176656 474056 176662
rect 474004 176598 474056 176604
rect 485044 176656 485096 176662
rect 485044 176598 485096 176604
rect 501696 176656 501748 176662
rect 501696 176598 501748 176604
rect 512644 176656 512696 176662
rect 512644 176598 512696 176604
rect 463700 176520 463752 176526
rect 463700 176462 463752 176468
rect 463792 172712 463844 172718
rect 463792 172654 463844 172660
rect 485044 172712 485096 172718
rect 485044 172654 485096 172660
rect 492588 172712 492640 172718
rect 492588 172654 492640 172660
rect 462964 172576 463016 172582
rect 462964 172518 463016 172524
rect 462976 148986 463004 172518
rect 463804 171134 463832 172654
rect 464620 172644 464672 172650
rect 464620 172586 464672 172592
rect 463804 171106 464200 171134
rect 464172 151722 464200 171106
rect 464632 170884 464660 172586
rect 474280 172576 474332 172582
rect 474280 172518 474332 172524
rect 474292 170884 474320 172518
rect 483966 170326 484072 170354
rect 464172 151694 464646 151722
rect 474292 148986 474320 151028
rect 483952 149054 483980 151028
rect 484044 149054 484072 170326
rect 483940 149048 483992 149054
rect 483940 148990 483992 148996
rect 484032 149048 484084 149054
rect 484032 148990 484084 148996
rect 485056 148986 485084 172654
rect 491392 172576 491444 172582
rect 491392 172518 491444 172524
rect 491404 171134 491432 172518
rect 491404 171106 492168 171134
rect 489826 161392 489882 161401
rect 489826 161327 489882 161336
rect 485778 160712 485834 160721
rect 485778 160647 485834 160656
rect 485792 151706 485820 160647
rect 489840 151774 489868 161327
rect 489828 151768 489880 151774
rect 489828 151710 489880 151716
rect 492140 151722 492168 171106
rect 492600 170884 492628 172654
rect 502248 172644 502300 172650
rect 502248 172586 502300 172592
rect 514024 172644 514076 172650
rect 514024 172586 514076 172592
rect 502260 170884 502288 172586
rect 511934 170326 512132 170354
rect 485780 151700 485832 151706
rect 492140 151694 492614 151722
rect 485780 151642 485832 151648
rect 502260 148986 502288 151028
rect 511920 149054 511948 151028
rect 512104 149054 512132 170326
rect 513378 160712 513434 160721
rect 513378 160647 513434 160656
rect 513392 151638 513420 160647
rect 513380 151632 513432 151638
rect 513380 151574 513432 151580
rect 511908 149048 511960 149054
rect 511908 148990 511960 148996
rect 512092 149048 512144 149054
rect 512092 148990 512144 148996
rect 514036 148986 514064 172586
rect 462964 148980 463016 148986
rect 462964 148922 463016 148928
rect 474280 148980 474332 148986
rect 474280 148922 474332 148928
rect 485044 148980 485096 148986
rect 485044 148922 485096 148928
rect 502248 148980 502300 148986
rect 502248 148922 502300 148928
rect 514024 148980 514076 148986
rect 514024 148922 514076 148928
rect 492036 146532 492088 146538
rect 492036 146474 492088 146480
rect 512736 146532 512788 146538
rect 512736 146474 512788 146480
rect 473360 146464 473412 146470
rect 473360 146406 473412 146412
rect 483480 146464 483532 146470
rect 483480 146406 483532 146412
rect 464344 146396 464396 146402
rect 464344 146338 464396 146344
rect 464356 143970 464384 146338
rect 464048 143942 464384 143970
rect 473372 143970 473400 146406
rect 483020 146328 483072 146334
rect 483020 146270 483072 146276
rect 483032 143970 483060 146270
rect 473372 143942 473708 143970
rect 483032 143942 483368 143970
rect 483492 124794 483520 146406
rect 483664 146396 483716 146402
rect 483664 146338 483716 146344
rect 483676 126954 483704 146338
rect 485044 146328 485096 146334
rect 485044 146270 485096 146276
rect 483664 126948 483716 126954
rect 483664 126890 483716 126896
rect 483368 124766 483520 124794
rect 463804 124086 464048 124114
rect 473708 124086 474044 124114
rect 463804 122670 463832 124086
rect 474016 122806 474044 124086
rect 485056 122806 485084 146270
rect 492048 143956 492076 146474
rect 501696 146464 501748 146470
rect 501696 146406 501748 146412
rect 501708 143956 501736 146406
rect 511448 146396 511500 146402
rect 511448 146338 511500 146344
rect 511356 146328 511408 146334
rect 511356 146270 511408 146276
rect 511368 143956 511396 146270
rect 489826 134328 489882 134337
rect 489826 134263 489882 134272
rect 485778 133648 485834 133657
rect 485778 133583 485834 133592
rect 485792 125526 485820 133583
rect 489840 125594 489868 134263
rect 491668 126948 491720 126954
rect 491668 126890 491720 126896
rect 489828 125588 489880 125594
rect 489828 125530 489880 125536
rect 485780 125520 485832 125526
rect 485780 125462 485832 125468
rect 491680 124794 491708 126890
rect 511460 124794 511488 146338
rect 512644 146328 512696 146334
rect 512644 146270 512696 146276
rect 491680 124766 492062 124794
rect 511382 124766 511488 124794
rect 501708 122806 501736 124100
rect 512656 122806 512684 146270
rect 512748 126954 512776 146474
rect 513378 133648 513434 133657
rect 513378 133583 513434 133592
rect 512736 126948 512788 126954
rect 512736 126890 512788 126896
rect 513392 125458 513420 133583
rect 513380 125452 513432 125458
rect 513380 125394 513432 125400
rect 474004 122800 474056 122806
rect 474004 122742 474056 122748
rect 485044 122800 485096 122806
rect 485044 122742 485096 122748
rect 501696 122800 501748 122806
rect 501696 122742 501748 122748
rect 512644 122800 512696 122806
rect 512644 122742 512696 122748
rect 463792 122664 463844 122670
rect 463792 122606 463844 122612
rect 463792 118856 463844 118862
rect 463792 118798 463844 118804
rect 491392 118856 491444 118862
rect 491392 118798 491444 118804
rect 462964 118720 463016 118726
rect 462964 118662 463016 118668
rect 462976 95130 463004 118662
rect 463804 113174 463832 118798
rect 464620 118788 464672 118794
rect 464620 118730 464672 118736
rect 464632 116892 464660 118730
rect 474280 118720 474332 118726
rect 474280 118662 474332 118668
rect 485044 118720 485096 118726
rect 485044 118662 485096 118668
rect 474292 116892 474320 118662
rect 483966 116334 484072 116362
rect 463804 113146 464200 113174
rect 464172 97730 464200 113146
rect 464172 97702 464646 97730
rect 474292 95130 474320 97036
rect 483952 95198 483980 97036
rect 484044 95198 484072 116334
rect 483940 95192 483992 95198
rect 483940 95134 483992 95140
rect 484032 95192 484084 95198
rect 484032 95134 484084 95140
rect 485056 95130 485084 118662
rect 491404 113174 491432 118798
rect 502248 118788 502300 118794
rect 502248 118730 502300 118736
rect 514024 118788 514076 118794
rect 514024 118730 514076 118736
rect 492588 118720 492640 118726
rect 492588 118662 492640 118668
rect 492600 116892 492628 118662
rect 502260 116892 502288 118730
rect 511934 116334 512132 116362
rect 491404 113146 492168 113174
rect 489826 107400 489882 107409
rect 489826 107335 489882 107344
rect 485778 106720 485834 106729
rect 485778 106655 485834 106664
rect 485792 97918 485820 106655
rect 489840 97986 489868 107335
rect 489828 97980 489880 97986
rect 489828 97922 489880 97928
rect 485780 97912 485832 97918
rect 485780 97854 485832 97860
rect 492140 97730 492168 113146
rect 492140 97702 492614 97730
rect 502260 95130 502288 97036
rect 511920 95198 511948 97036
rect 512104 95198 512132 116334
rect 513378 106720 513434 106729
rect 513378 106655 513434 106664
rect 513392 97850 513420 106655
rect 513380 97844 513432 97850
rect 513380 97786 513432 97792
rect 511908 95192 511960 95198
rect 511908 95134 511960 95140
rect 512092 95192 512144 95198
rect 512092 95134 512144 95140
rect 514036 95130 514064 118730
rect 462964 95124 463016 95130
rect 462964 95066 463016 95072
rect 474280 95124 474332 95130
rect 474280 95066 474332 95072
rect 485044 95124 485096 95130
rect 485044 95066 485096 95072
rect 502248 95124 502300 95130
rect 502248 95066 502300 95072
rect 514024 95124 514076 95130
rect 514024 95066 514076 95072
rect 473360 91248 473412 91254
rect 473360 91190 473412 91196
rect 483480 91248 483532 91254
rect 483480 91190 483532 91196
rect 501696 91248 501748 91254
rect 501696 91190 501748 91196
rect 511448 91248 511500 91254
rect 511448 91190 511500 91196
rect 464344 91180 464396 91186
rect 464344 91122 464396 91128
rect 464356 89978 464384 91122
rect 464048 89950 464384 89978
rect 473372 89978 473400 91190
rect 483020 91112 483072 91118
rect 483020 91054 483072 91060
rect 483032 89978 483060 91054
rect 473372 89950 473708 89978
rect 483032 89950 483368 89978
rect 483492 70666 483520 91190
rect 483664 91180 483716 91186
rect 483664 91122 483716 91128
rect 492036 91180 492088 91186
rect 492036 91122 492088 91128
rect 483676 72282 483704 91122
rect 485044 91112 485096 91118
rect 485044 91054 485096 91060
rect 483664 72276 483716 72282
rect 483664 72218 483716 72224
rect 483368 70638 483520 70666
rect 463712 70094 464048 70122
rect 473708 70094 474044 70122
rect 463712 68882 463740 70094
rect 474016 69018 474044 70094
rect 485056 69018 485084 91054
rect 492048 89964 492076 91122
rect 501708 89964 501736 91190
rect 511356 91112 511408 91118
rect 511356 91054 511408 91060
rect 511368 89964 511396 91054
rect 485780 88868 485832 88874
rect 485780 88810 485832 88816
rect 485792 79665 485820 88810
rect 489828 88392 489880 88398
rect 489828 88334 489880 88340
rect 489840 80345 489868 88334
rect 489826 80336 489882 80345
rect 489826 80271 489882 80280
rect 485778 79656 485834 79665
rect 485778 79591 485834 79600
rect 491668 72276 491720 72282
rect 491668 72218 491720 72224
rect 491680 70666 491708 72218
rect 511460 70666 511488 91190
rect 512736 91180 512788 91186
rect 512736 91122 512788 91128
rect 512644 91112 512696 91118
rect 512644 91054 512696 91060
rect 491680 70638 492062 70666
rect 511382 70638 511488 70666
rect 501708 69018 501736 70108
rect 512656 69018 512684 91054
rect 512748 72146 512776 91122
rect 513378 79656 513434 79665
rect 513378 79591 513434 79600
rect 512736 72140 512788 72146
rect 512736 72082 512788 72088
rect 513392 71738 513420 79591
rect 513380 71732 513432 71738
rect 513380 71674 513432 71680
rect 474004 69012 474056 69018
rect 474004 68954 474056 68960
rect 485044 69012 485096 69018
rect 485044 68954 485096 68960
rect 501696 69012 501748 69018
rect 501696 68954 501748 68960
rect 512644 69012 512696 69018
rect 512644 68954 512696 68960
rect 463700 68876 463752 68882
rect 463700 68818 463752 68824
rect 463792 65068 463844 65074
rect 463792 65010 463844 65016
rect 485044 65068 485096 65074
rect 485044 65010 485096 65016
rect 492588 65068 492640 65074
rect 492588 65010 492640 65016
rect 462964 64932 463016 64938
rect 462964 64874 463016 64880
rect 462976 41342 463004 64874
rect 463804 55214 463832 65010
rect 464620 65000 464672 65006
rect 464620 64942 464672 64948
rect 464632 62900 464660 64942
rect 474280 64932 474332 64938
rect 474280 64874 474332 64880
rect 474292 62900 474320 64874
rect 483966 62206 484072 62234
rect 463804 55186 464200 55214
rect 464172 43738 464200 55186
rect 464172 43710 464646 43738
rect 474292 41342 474320 43044
rect 483952 41410 483980 43044
rect 484044 41410 484072 62206
rect 483940 41404 483992 41410
rect 483940 41346 483992 41352
rect 484032 41404 484084 41410
rect 484032 41346 484084 41352
rect 485056 41342 485084 65010
rect 491392 64932 491444 64938
rect 491392 64874 491444 64880
rect 485780 62144 485832 62150
rect 485780 62086 485832 62092
rect 489828 62144 489880 62150
rect 489828 62086 489880 62092
rect 485792 52737 485820 62086
rect 489840 53417 489868 62086
rect 491404 55214 491432 64874
rect 492600 62900 492628 65010
rect 502248 65000 502300 65006
rect 502248 64942 502300 64948
rect 514024 65000 514076 65006
rect 514024 64942 514076 64948
rect 502260 62900 502288 64942
rect 511934 62206 512132 62234
rect 491404 55186 492168 55214
rect 489826 53408 489882 53417
rect 489826 53343 489882 53352
rect 485778 52728 485834 52737
rect 485778 52663 485834 52672
rect 492140 43738 492168 55186
rect 492140 43710 492614 43738
rect 502260 41342 502288 43044
rect 511920 41410 511948 43044
rect 512104 41410 512132 62206
rect 513378 52728 513434 52737
rect 513378 52663 513434 52672
rect 513392 44130 513420 52663
rect 513380 44124 513432 44130
rect 513380 44066 513432 44072
rect 511908 41404 511960 41410
rect 511908 41346 511960 41352
rect 512092 41404 512144 41410
rect 512092 41346 512144 41352
rect 514036 41342 514064 64942
rect 462964 41336 463016 41342
rect 462964 41278 463016 41284
rect 474280 41336 474332 41342
rect 474280 41278 474332 41284
rect 485044 41336 485096 41342
rect 485044 41278 485096 41284
rect 502248 41336 502300 41342
rect 502248 41278 502300 41284
rect 514024 41336 514076 41342
rect 514024 41278 514076 41284
rect 462320 38276 462372 38282
rect 462320 38218 462372 38224
rect 456064 37460 456116 37466
rect 456064 37402 456116 37408
rect 473360 37460 473412 37466
rect 473360 37402 473412 37408
rect 483480 37460 483532 37466
rect 483480 37402 483532 37408
rect 501696 37460 501748 37466
rect 501696 37402 501748 37408
rect 429844 37392 429896 37398
rect 429844 37334 429896 37340
rect 445668 37392 445720 37398
rect 445668 37334 445720 37340
rect 429292 34604 429344 34610
rect 429292 34546 429344 34552
rect 429304 25673 429332 34546
rect 429290 25664 429346 25673
rect 429290 25599 429346 25608
rect 429856 16590 429884 37334
rect 445680 35972 445708 37334
rect 455328 37324 455380 37330
rect 455328 37266 455380 37272
rect 455340 35972 455368 37266
rect 434824 35278 436034 35306
rect 434628 34672 434680 34678
rect 434628 34614 434680 34620
rect 434640 26353 434668 34614
rect 434626 26344 434682 26353
rect 434626 26279 434682 26288
rect 429844 16584 429896 16590
rect 429844 16526 429896 16532
rect 429200 15156 429252 15162
rect 429200 15098 429252 15104
rect 434824 13462 434852 35278
rect 456076 26234 456104 37402
rect 464344 37392 464396 37398
rect 464344 37334 464396 37340
rect 456156 37324 456208 37330
rect 456156 37266 456208 37272
rect 455800 26206 456104 26234
rect 435732 18624 435784 18630
rect 435732 18566 435784 18572
rect 435744 16674 435772 18566
rect 455800 16674 455828 26206
rect 435744 16646 436034 16674
rect 455354 16646 455828 16674
rect 378784 13456 378836 13462
rect 378784 13398 378836 13404
rect 379612 13456 379664 13462
rect 379612 13398 379664 13404
rect 408040 13456 408092 13462
rect 408040 13398 408092 13404
rect 417700 13456 417752 13462
rect 417700 13398 417752 13404
rect 428464 13456 428516 13462
rect 428464 13398 428516 13404
rect 434812 13456 434864 13462
rect 434812 13398 434864 13404
rect 445680 13394 445708 16116
rect 456168 13394 456196 37266
rect 464356 35986 464384 37334
rect 464048 35958 464384 35986
rect 473372 35986 473400 37402
rect 483020 37324 483072 37330
rect 483020 37266 483072 37272
rect 483032 35986 483060 37266
rect 473372 35958 473708 35986
rect 483032 35958 483368 35986
rect 462228 34604 462280 34610
rect 462228 34546 462280 34552
rect 458180 34536 458232 34542
rect 458180 34478 458232 34484
rect 458192 25673 458220 34478
rect 462240 26353 462268 34546
rect 462226 26344 462282 26353
rect 462226 26279 462282 26288
rect 458178 25664 458234 25673
rect 458178 25599 458234 25608
rect 483492 16674 483520 37402
rect 483664 37392 483716 37398
rect 483664 37334 483716 37340
rect 492036 37392 492088 37398
rect 492036 37334 492088 37340
rect 483676 18018 483704 37334
rect 485044 37324 485096 37330
rect 485044 37266 485096 37272
rect 483664 18012 483716 18018
rect 483664 17954 483716 17960
rect 483368 16646 483520 16674
rect 463712 16102 464048 16130
rect 473708 16102 474044 16130
rect 463712 13462 463740 16102
rect 474016 13802 474044 16102
rect 485056 13802 485084 37266
rect 492048 35972 492076 37334
rect 501708 35972 501736 37402
rect 512736 37392 512788 37398
rect 512736 37334 512788 37340
rect 511356 37324 511408 37330
rect 511356 37266 511408 37272
rect 512644 37324 512696 37330
rect 512644 37266 512696 37272
rect 511368 35972 511396 37266
rect 485780 34672 485832 34678
rect 485780 34614 485832 34620
rect 485792 25673 485820 34614
rect 489828 34536 489880 34542
rect 489828 34478 489880 34484
rect 489840 26353 489868 34478
rect 489826 26344 489882 26353
rect 489826 26279 489882 26288
rect 485778 25664 485834 25673
rect 485778 25599 485834 25608
rect 491668 18012 491720 18018
rect 491668 17954 491720 17960
rect 491680 16674 491708 17954
rect 491680 16646 492062 16674
rect 501708 13802 501736 16116
rect 474004 13796 474056 13802
rect 474004 13738 474056 13744
rect 485044 13796 485096 13802
rect 485044 13738 485096 13744
rect 501696 13796 501748 13802
rect 501696 13738 501748 13744
rect 511368 13462 511396 16116
rect 512656 13802 512684 37266
rect 512748 18018 512776 37334
rect 513380 34604 513432 34610
rect 513380 34546 513432 34552
rect 513392 25673 513420 34546
rect 513378 25664 513434 25673
rect 513378 25599 513434 25608
rect 512736 18012 512788 18018
rect 512736 17954 512788 17960
rect 512644 13796 512696 13802
rect 512644 13738 512696 13744
rect 463700 13456 463752 13462
rect 463700 13398 463752 13404
rect 511356 13456 511408 13462
rect 511356 13398 511408 13404
rect 352012 13388 352064 13394
rect 352012 13330 352064 13336
rect 445668 13388 445720 13394
rect 445668 13330 445720 13336
rect 456156 13388 456208 13394
rect 456156 13330 456208 13336
rect 333704 13320 333756 13326
rect 333704 13262 333756 13268
rect 344284 13320 344336 13326
rect 518176 13297 518204 700334
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 529664 685976 529716 685982
rect 529664 685918 529716 685924
rect 541624 685976 541676 685982
rect 541624 685918 541676 685924
rect 557540 685976 557592 685982
rect 557540 685918 557592 685924
rect 529676 683876 529704 685918
rect 539324 685908 539376 685914
rect 539324 685850 539376 685856
rect 540244 685908 540296 685914
rect 540244 685850 540296 685856
rect 539336 683876 539364 685850
rect 519004 683318 520030 683346
rect 518806 674248 518862 674257
rect 518806 674183 518862 674192
rect 518820 665174 518848 674183
rect 518808 665168 518860 665174
rect 518808 665110 518860 665116
rect 519004 662250 519032 683318
rect 519636 665304 519688 665310
rect 519636 665246 519688 665252
rect 519648 664714 519676 665246
rect 519648 664686 520030 664714
rect 529676 662318 529704 664020
rect 539336 663746 539364 664020
rect 539324 663740 539376 663746
rect 539324 663682 539376 663688
rect 540256 662318 540284 685850
rect 541636 663746 541664 685918
rect 557552 683754 557580 685918
rect 567200 685908 567252 685914
rect 567200 685850 567252 685856
rect 567212 683754 567240 685850
rect 557552 683726 557704 683754
rect 567212 683726 567364 683754
rect 542360 683188 542412 683194
rect 542360 683130 542412 683136
rect 542372 673577 542400 683130
rect 545118 674248 545174 674257
rect 545118 674183 545174 674192
rect 545132 673810 545160 674183
rect 543004 673804 543056 673810
rect 543004 673746 543056 673752
rect 545120 673804 545172 673810
rect 545120 673746 545172 673752
rect 542358 673568 542414 673577
rect 542358 673503 542414 673512
rect 541624 663740 541676 663746
rect 541624 663682 541676 663688
rect 529664 662312 529716 662318
rect 529664 662254 529716 662260
rect 540244 662312 540296 662318
rect 540244 662254 540296 662260
rect 518992 662244 519044 662250
rect 518992 662186 519044 662192
rect 529940 658436 529992 658442
rect 529940 658378 529992 658384
rect 520280 658368 520332 658374
rect 520280 658310 520332 658316
rect 520292 656962 520320 658310
rect 529952 656962 529980 658378
rect 541624 658368 541676 658374
rect 541624 658310 541676 658316
rect 520292 656934 520628 656962
rect 529952 656934 530288 656962
rect 539948 656254 540100 656282
rect 518808 655648 518860 655654
rect 518808 655590 518860 655596
rect 518820 647465 518848 655590
rect 518806 647456 518862 647465
rect 518806 647391 518862 647400
rect 520628 637078 520964 637106
rect 530288 637078 530624 637106
rect 520936 634710 520964 637078
rect 520924 634704 520976 634710
rect 520924 634646 520976 634652
rect 530596 634642 530624 637078
rect 539612 637078 539948 637106
rect 539612 634778 539640 637078
rect 540072 634778 540100 656254
rect 539600 634772 539652 634778
rect 539600 634714 539652 634720
rect 540060 634772 540112 634778
rect 540060 634714 540112 634720
rect 541636 634710 541664 658310
rect 542360 655580 542412 655586
rect 542360 655522 542412 655528
rect 542372 646785 542400 655522
rect 542358 646776 542414 646785
rect 542358 646711 542414 646720
rect 541624 634704 541676 634710
rect 541624 634646 541676 634652
rect 530584 634636 530636 634642
rect 530584 634578 530636 634584
rect 529664 632188 529716 632194
rect 529664 632130 529716 632136
rect 541624 632188 541676 632194
rect 541624 632130 541676 632136
rect 529676 629884 529704 632130
rect 539324 632120 539376 632126
rect 539324 632062 539376 632068
rect 540244 632120 540296 632126
rect 540244 632062 540296 632068
rect 539336 629884 539364 632062
rect 519004 629326 520030 629354
rect 518806 620256 518862 620265
rect 518806 620191 518862 620200
rect 518820 611250 518848 620191
rect 518808 611244 518860 611250
rect 518808 611186 518860 611192
rect 519004 608462 519032 629326
rect 519636 611788 519688 611794
rect 519636 611730 519688 611736
rect 519648 610722 519676 611730
rect 539508 611312 539560 611318
rect 539508 611254 539560 611260
rect 539520 610722 539548 611254
rect 519648 610694 520030 610722
rect 539350 610694 539548 610722
rect 529676 608530 529704 610028
rect 540256 608530 540284 632062
rect 541636 611318 541664 632130
rect 542358 619576 542414 619585
rect 542358 619511 542414 619520
rect 541624 611312 541676 611318
rect 541624 611254 541676 611260
rect 542372 611182 542400 619511
rect 542360 611176 542412 611182
rect 542360 611118 542412 611124
rect 529664 608524 529716 608530
rect 529664 608466 529716 608472
rect 540244 608524 540296 608530
rect 540244 608466 540296 608472
rect 518992 608456 519044 608462
rect 518992 608398 519044 608404
rect 529940 604648 529992 604654
rect 529940 604590 529992 604596
rect 520280 604580 520332 604586
rect 520280 604522 520332 604528
rect 520292 602970 520320 604522
rect 529952 602970 529980 604590
rect 541624 604580 541676 604586
rect 541624 604522 541676 604528
rect 520292 602942 520628 602970
rect 529952 602942 530288 602970
rect 539948 602262 540100 602290
rect 518808 601792 518860 601798
rect 518808 601734 518860 601740
rect 518820 593473 518848 601734
rect 518806 593464 518862 593473
rect 518806 593399 518862 593408
rect 520628 583086 520964 583114
rect 530288 583086 530624 583114
rect 520936 580922 520964 583086
rect 520924 580916 520976 580922
rect 520924 580858 520976 580864
rect 530596 580854 530624 583086
rect 539612 583086 539948 583114
rect 539612 580990 539640 583086
rect 540072 580990 540100 602262
rect 539600 580984 539652 580990
rect 539600 580926 539652 580932
rect 540060 580984 540112 580990
rect 540060 580926 540112 580932
rect 541636 580922 541664 604522
rect 542360 601724 542412 601730
rect 542360 601666 542412 601672
rect 542372 592793 542400 601666
rect 542358 592784 542414 592793
rect 542358 592719 542414 592728
rect 541624 580916 541676 580922
rect 541624 580858 541676 580864
rect 530584 580848 530636 580854
rect 530584 580790 530636 580796
rect 529664 578332 529716 578338
rect 529664 578274 529716 578280
rect 541624 578332 541676 578338
rect 541624 578274 541676 578280
rect 529676 575892 529704 578274
rect 539324 578264 539376 578270
rect 539324 578206 539376 578212
rect 540244 578264 540296 578270
rect 540244 578206 540296 578212
rect 539336 575892 539364 578206
rect 519004 575334 520030 575362
rect 518806 566264 518862 566273
rect 518806 566199 518862 566208
rect 518820 557462 518848 566199
rect 518808 557456 518860 557462
rect 518808 557398 518860 557404
rect 519004 554606 519032 575334
rect 519636 558204 519688 558210
rect 519636 558146 519688 558152
rect 519648 556730 519676 558146
rect 539508 556776 539560 556782
rect 519648 556702 520030 556730
rect 539350 556724 539508 556730
rect 539350 556718 539560 556724
rect 539350 556702 539548 556718
rect 529676 554674 529704 556036
rect 540256 554674 540284 578206
rect 541636 556782 541664 578274
rect 542358 565584 542414 565593
rect 542358 565519 542414 565528
rect 542372 557530 542400 565519
rect 542360 557524 542412 557530
rect 542360 557466 542412 557472
rect 541624 556776 541676 556782
rect 541624 556718 541676 556724
rect 529664 554668 529716 554674
rect 529664 554610 529716 554616
rect 540244 554668 540296 554674
rect 540244 554610 540296 554616
rect 518992 554600 519044 554606
rect 518992 554542 519044 554548
rect 529940 550792 529992 550798
rect 529940 550734 529992 550740
rect 520280 550656 520332 550662
rect 520280 550598 520332 550604
rect 520292 548978 520320 550598
rect 529952 548978 529980 550734
rect 541624 550724 541676 550730
rect 541624 550666 541676 550672
rect 520292 548950 520628 548978
rect 529952 548950 530288 548978
rect 539948 548270 540100 548298
rect 518806 539472 518862 539481
rect 518806 539407 518862 539416
rect 518820 529854 518848 539407
rect 518808 529848 518860 529854
rect 518808 529790 518860 529796
rect 520628 529094 520964 529122
rect 530288 529094 530624 529122
rect 520936 527066 520964 529094
rect 520924 527060 520976 527066
rect 520924 527002 520976 527008
rect 530596 526998 530624 529094
rect 539612 529094 539948 529122
rect 539612 527134 539640 529094
rect 540072 527134 540100 548270
rect 539600 527128 539652 527134
rect 539600 527070 539652 527076
rect 540060 527128 540112 527134
rect 540060 527070 540112 527076
rect 541636 527066 541664 550666
rect 542358 538792 542414 538801
rect 542358 538727 542414 538736
rect 542372 529922 542400 538727
rect 542360 529916 542412 529922
rect 542360 529858 542412 529864
rect 541624 527060 541676 527066
rect 541624 527002 541676 527008
rect 530584 526992 530636 526998
rect 530584 526934 530636 526940
rect 529664 523116 529716 523122
rect 529664 523058 529716 523064
rect 541624 523116 541676 523122
rect 541624 523058 541676 523064
rect 529676 521900 529704 523058
rect 539324 523048 539376 523054
rect 539324 522990 539376 522996
rect 540244 523048 540296 523054
rect 540244 522990 540296 522996
rect 539336 521900 539364 522990
rect 519004 521206 520030 521234
rect 518806 512272 518862 512281
rect 518806 512207 518862 512216
rect 518820 503674 518848 512207
rect 518808 503668 518860 503674
rect 518808 503610 518860 503616
rect 519004 500818 519032 521206
rect 519636 504348 519688 504354
rect 519636 504290 519688 504296
rect 519648 502738 519676 504290
rect 539508 503600 539560 503606
rect 539508 503542 539560 503548
rect 539520 502738 539548 503542
rect 519648 502710 520030 502738
rect 539350 502710 539548 502738
rect 529676 500886 529704 502044
rect 540256 500886 540284 522990
rect 541636 503606 541664 523058
rect 542360 520328 542412 520334
rect 542360 520270 542412 520276
rect 542372 511601 542400 520270
rect 542358 511592 542414 511601
rect 542358 511527 542414 511536
rect 541624 503600 541676 503606
rect 541624 503542 541676 503548
rect 529664 500880 529716 500886
rect 529664 500822 529716 500828
rect 540244 500880 540296 500886
rect 540244 500822 540296 500828
rect 518992 500812 519044 500818
rect 518992 500754 519044 500760
rect 520280 496936 520332 496942
rect 520280 496878 520332 496884
rect 520292 494986 520320 496878
rect 529940 496868 529992 496874
rect 529940 496810 529992 496816
rect 541624 496868 541676 496874
rect 541624 496810 541676 496816
rect 529952 494986 529980 496810
rect 520292 494958 520628 494986
rect 529952 494958 530288 494986
rect 539948 494278 540100 494306
rect 518806 485480 518862 485489
rect 518806 485415 518862 485424
rect 518820 475998 518848 485415
rect 518808 475992 518860 475998
rect 518808 475934 518860 475940
rect 520628 475102 520964 475130
rect 530288 475102 530624 475130
rect 520936 473278 520964 475102
rect 520924 473272 520976 473278
rect 520924 473214 520976 473220
rect 530596 473210 530624 475102
rect 539612 475102 539948 475130
rect 539612 473346 539640 475102
rect 540072 473346 540100 494278
rect 539600 473340 539652 473346
rect 539600 473282 539652 473288
rect 540060 473340 540112 473346
rect 540060 473282 540112 473288
rect 541636 473278 541664 496810
rect 542358 484800 542414 484809
rect 542358 484735 542414 484744
rect 542372 476066 542400 484735
rect 542360 476060 542412 476066
rect 542360 476002 542412 476008
rect 541624 473272 541676 473278
rect 541624 473214 541676 473220
rect 530584 473204 530636 473210
rect 530584 473146 530636 473152
rect 529664 469396 529716 469402
rect 529664 469338 529716 469344
rect 529676 467908 529704 469338
rect 541624 469328 541676 469334
rect 541624 469270 541676 469276
rect 539324 469260 539376 469266
rect 539324 469202 539376 469208
rect 540244 469260 540296 469266
rect 540244 469202 540296 469208
rect 539336 467908 539364 469202
rect 519004 467214 520030 467242
rect 518808 466540 518860 466546
rect 518808 466482 518860 466488
rect 518820 458289 518848 466482
rect 518806 458280 518862 458289
rect 518806 458215 518862 458224
rect 519004 445602 519032 467214
rect 519636 450492 519688 450498
rect 519636 450434 519688 450440
rect 519648 448746 519676 450434
rect 519648 448718 520030 448746
rect 539508 448520 539560 448526
rect 539350 448468 539508 448474
rect 539350 448462 539560 448468
rect 539350 448446 539548 448462
rect 529676 445670 529704 448052
rect 540256 445670 540284 469202
rect 541636 448526 541664 469270
rect 542360 466472 542412 466478
rect 542360 466414 542412 466420
rect 542372 457609 542400 466414
rect 542358 457600 542414 457609
rect 542358 457535 542414 457544
rect 541624 448520 541676 448526
rect 541624 448462 541676 448468
rect 529664 445664 529716 445670
rect 529664 445606 529716 445612
rect 540244 445664 540296 445670
rect 540244 445606 540296 445612
rect 518992 445596 519044 445602
rect 518992 445538 519044 445544
rect 520280 443080 520332 443086
rect 520280 443022 520332 443028
rect 520292 440994 520320 443022
rect 529940 443012 529992 443018
rect 529940 442954 529992 442960
rect 541624 443012 541676 443018
rect 541624 442954 541676 442960
rect 529952 440994 529980 442954
rect 520292 440966 520628 440994
rect 529952 440966 530288 440994
rect 539948 440286 540100 440314
rect 518806 431488 518862 431497
rect 518806 431423 518862 431432
rect 518820 422278 518848 431423
rect 518808 422272 518860 422278
rect 518808 422214 518860 422220
rect 520628 421110 520964 421138
rect 530288 421110 530624 421138
rect 520936 419422 520964 421110
rect 520924 419416 520976 419422
rect 520924 419358 520976 419364
rect 530596 419354 530624 421110
rect 539612 421110 539948 421138
rect 539612 419490 539640 421110
rect 540072 419490 540100 440286
rect 539600 419484 539652 419490
rect 539600 419426 539652 419432
rect 540060 419484 540112 419490
rect 540060 419426 540112 419432
rect 541636 419422 541664 442954
rect 542360 440292 542412 440298
rect 542360 440234 542412 440240
rect 542372 430817 542400 440234
rect 542358 430808 542414 430817
rect 542358 430743 542414 430752
rect 541624 419416 541676 419422
rect 541624 419358 541676 419364
rect 530584 419348 530636 419354
rect 530584 419290 530636 419296
rect 529664 415608 529716 415614
rect 529664 415550 529716 415556
rect 529676 413916 529704 415550
rect 541624 415540 541676 415546
rect 541624 415482 541676 415488
rect 539324 415472 539376 415478
rect 539324 415414 539376 415420
rect 540244 415472 540296 415478
rect 540244 415414 540296 415420
rect 539336 413916 539364 415414
rect 519004 413222 520030 413250
rect 518806 404288 518862 404297
rect 518806 404223 518862 404232
rect 518820 394602 518848 404223
rect 518808 394596 518860 394602
rect 518808 394538 518860 394544
rect 519004 391814 519032 413222
rect 519636 395072 519688 395078
rect 519636 395014 519688 395020
rect 519648 394754 519676 395014
rect 519648 394726 520030 394754
rect 529676 391882 529704 394060
rect 539336 393310 539364 394060
rect 539324 393304 539376 393310
rect 539324 393246 539376 393252
rect 540256 391882 540284 415414
rect 541636 393310 541664 415482
rect 542358 403608 542414 403617
rect 542358 403543 542414 403552
rect 542372 394670 542400 403543
rect 542360 394664 542412 394670
rect 542360 394606 542412 394612
rect 541624 393304 541676 393310
rect 541624 393246 541676 393252
rect 529664 391876 529716 391882
rect 529664 391818 529716 391824
rect 540244 391876 540296 391882
rect 540244 391818 540296 391824
rect 518992 391808 519044 391814
rect 518992 391750 519044 391756
rect 520280 389292 520332 389298
rect 520280 389234 520332 389240
rect 520292 386866 520320 389234
rect 529940 389224 529992 389230
rect 529940 389166 529992 389172
rect 541624 389224 541676 389230
rect 541624 389166 541676 389172
rect 529952 386866 529980 389166
rect 520292 386838 520628 386866
rect 529952 386838 530288 386866
rect 518808 386504 518860 386510
rect 518808 386446 518860 386452
rect 518820 377505 518848 386446
rect 539948 386294 540100 386322
rect 518806 377496 518862 377505
rect 518806 377431 518862 377440
rect 520628 367118 520964 367146
rect 530288 367118 530624 367146
rect 520936 365634 520964 367118
rect 520924 365628 520976 365634
rect 520924 365570 520976 365576
rect 530596 365566 530624 367118
rect 539612 367118 539948 367146
rect 539612 365702 539640 367118
rect 540072 365702 540100 386294
rect 539600 365696 539652 365702
rect 539600 365638 539652 365644
rect 540060 365696 540112 365702
rect 540060 365638 540112 365644
rect 541636 365634 541664 389166
rect 542360 386436 542412 386442
rect 542360 386378 542412 386384
rect 542372 376825 542400 386378
rect 542358 376816 542414 376825
rect 542358 376751 542414 376760
rect 541624 365628 541676 365634
rect 541624 365570 541676 365576
rect 530584 365560 530636 365566
rect 530584 365502 530636 365508
rect 529664 361752 529716 361758
rect 529664 361694 529716 361700
rect 529676 359924 529704 361694
rect 541624 361684 541676 361690
rect 541624 361626 541676 361632
rect 539324 361616 539376 361622
rect 539324 361558 539376 361564
rect 540244 361616 540296 361622
rect 540244 361558 540296 361564
rect 539336 359924 539364 361558
rect 519004 359230 520030 359258
rect 518806 350296 518862 350305
rect 518806 350231 518862 350240
rect 518820 340814 518848 350231
rect 518808 340808 518860 340814
rect 518808 340750 518860 340756
rect 519004 337958 519032 359230
rect 519636 341964 519688 341970
rect 519636 341906 519688 341912
rect 519648 340762 519676 341906
rect 539508 340876 539560 340882
rect 539508 340818 539560 340824
rect 539520 340762 539548 340818
rect 519648 340734 520030 340762
rect 539350 340734 539548 340762
rect 529676 338026 529704 340068
rect 540256 338026 540284 361558
rect 541636 340882 541664 361626
rect 542358 349616 542414 349625
rect 542358 349551 542414 349560
rect 541624 340876 541676 340882
rect 541624 340818 541676 340824
rect 542372 340746 542400 349551
rect 542360 340740 542412 340746
rect 542360 340682 542412 340688
rect 529664 338020 529716 338026
rect 529664 337962 529716 337968
rect 540244 338020 540296 338026
rect 540244 337962 540296 337968
rect 518992 337952 519044 337958
rect 518992 337894 519044 337900
rect 529940 335504 529992 335510
rect 529940 335446 529992 335452
rect 520280 335436 520332 335442
rect 520280 335378 520332 335384
rect 520292 332874 520320 335378
rect 529952 332874 529980 335446
rect 541624 335368 541676 335374
rect 541624 335310 541676 335316
rect 520292 332846 520628 332874
rect 529952 332846 530288 332874
rect 539948 332302 540100 332330
rect 518806 322960 518862 322969
rect 518806 322895 518862 322904
rect 518820 314634 518848 322895
rect 518808 314628 518860 314634
rect 518808 314570 518860 314576
rect 520628 313126 520964 313154
rect 530288 313126 530624 313154
rect 520936 311778 520964 313126
rect 520924 311772 520976 311778
rect 520924 311714 520976 311720
rect 530596 311710 530624 313126
rect 539612 313126 539948 313154
rect 539612 311846 539640 313126
rect 540072 311846 540100 332302
rect 539600 311840 539652 311846
rect 539600 311782 539652 311788
rect 540060 311840 540112 311846
rect 540060 311782 540112 311788
rect 541636 311778 541664 335310
rect 542360 331288 542412 331294
rect 542360 331230 542412 331236
rect 542372 322833 542400 331230
rect 542358 322824 542414 322833
rect 542358 322759 542414 322768
rect 541624 311772 541676 311778
rect 541624 311714 541676 311720
rect 530584 311704 530636 311710
rect 530584 311646 530636 311652
rect 529664 307964 529716 307970
rect 529664 307906 529716 307912
rect 529676 305932 529704 307906
rect 541624 307896 541676 307902
rect 541624 307838 541676 307844
rect 539324 307828 539376 307834
rect 539324 307770 539376 307776
rect 540244 307828 540296 307834
rect 540244 307770 540296 307776
rect 539336 305932 539364 307770
rect 519004 305238 520030 305266
rect 518806 296304 518862 296313
rect 518806 296239 518862 296248
rect 518820 286958 518848 296239
rect 518808 286952 518860 286958
rect 518808 286894 518860 286900
rect 519004 284170 519032 305238
rect 519636 287564 519688 287570
rect 519636 287506 519688 287512
rect 519648 286770 519676 287506
rect 539508 286816 539560 286822
rect 519648 286742 520030 286770
rect 539350 286764 539508 286770
rect 539350 286758 539560 286764
rect 539350 286742 539548 286758
rect 529676 284238 529704 286076
rect 540256 284238 540284 307770
rect 541636 286822 541664 307838
rect 542358 295624 542414 295633
rect 542358 295559 542414 295568
rect 542372 287026 542400 295559
rect 542360 287020 542412 287026
rect 542360 286962 542412 286968
rect 541624 286816 541676 286822
rect 541624 286758 541676 286764
rect 529664 284232 529716 284238
rect 529664 284174 529716 284180
rect 540244 284232 540296 284238
rect 540244 284174 540296 284180
rect 518992 284164 519044 284170
rect 518992 284106 519044 284112
rect 529940 280356 529992 280362
rect 529940 280298 529992 280304
rect 520280 280220 520332 280226
rect 520280 280162 520332 280168
rect 520292 278882 520320 280162
rect 529952 278882 529980 280298
rect 541624 280288 541676 280294
rect 541624 280230 541676 280236
rect 520292 278854 520628 278882
rect 529952 278854 530288 278882
rect 539948 278310 540100 278338
rect 518808 277500 518860 277506
rect 518808 277442 518860 277448
rect 518820 269929 518848 277442
rect 518806 269920 518862 269929
rect 518806 269855 518862 269864
rect 520628 259134 520964 259162
rect 530288 259134 530624 259162
rect 520936 256630 520964 259134
rect 520924 256624 520976 256630
rect 520924 256566 520976 256572
rect 530596 256562 530624 259134
rect 539612 259134 539948 259162
rect 539612 256698 539640 259134
rect 540072 256698 540100 278310
rect 539600 256692 539652 256698
rect 539600 256634 539652 256640
rect 540060 256692 540112 256698
rect 540060 256634 540112 256640
rect 541636 256630 541664 280230
rect 542360 277432 542412 277438
rect 542360 277374 542412 277380
rect 542372 269113 542400 277374
rect 542358 269104 542414 269113
rect 542358 269039 542414 269048
rect 541624 256624 541676 256630
rect 541624 256566 541676 256572
rect 530584 256556 530636 256562
rect 530584 256498 530636 256504
rect 529664 254040 529716 254046
rect 529664 253982 529716 253988
rect 541624 254040 541676 254046
rect 541624 253982 541676 253988
rect 529676 251940 529704 253982
rect 539324 253972 539376 253978
rect 539324 253914 539376 253920
rect 540244 253972 540296 253978
rect 540244 253914 540296 253920
rect 539336 251940 539364 253914
rect 518808 251320 518860 251326
rect 518808 251262 518860 251268
rect 518820 242321 518848 251262
rect 519004 251246 520030 251274
rect 518806 242312 518862 242321
rect 518806 242247 518862 242256
rect 519004 230314 519032 251246
rect 519636 234252 519688 234258
rect 519636 234194 519688 234200
rect 519648 232778 519676 234194
rect 539508 233232 539560 233238
rect 539508 233174 539560 233180
rect 539520 232778 539548 233174
rect 519648 232750 520030 232778
rect 539350 232750 539548 232778
rect 529676 230382 529704 232084
rect 540256 230382 540284 253914
rect 541636 233238 541664 253982
rect 542360 251252 542412 251258
rect 542360 251194 542412 251200
rect 542372 241641 542400 251194
rect 542358 241632 542414 241641
rect 542358 241567 542414 241576
rect 541624 233232 541676 233238
rect 541624 233174 541676 233180
rect 529664 230376 529716 230382
rect 529664 230318 529716 230324
rect 540244 230376 540296 230382
rect 540244 230318 540296 230324
rect 518992 230308 519044 230314
rect 518992 230250 519044 230256
rect 529940 226500 529992 226506
rect 529940 226442 529992 226448
rect 520280 226432 520332 226438
rect 520280 226374 520332 226380
rect 520292 224890 520320 226374
rect 529952 224890 529980 226442
rect 541624 226432 541676 226438
rect 541624 226374 541676 226380
rect 520292 224862 520628 224890
rect 529952 224862 530288 224890
rect 539948 224318 540100 224346
rect 518808 223712 518860 223718
rect 518808 223654 518860 223660
rect 518820 215393 518848 223654
rect 518806 215384 518862 215393
rect 518806 215319 518862 215328
rect 520628 205006 520964 205034
rect 530288 205006 530624 205034
rect 520936 202774 520964 205006
rect 520924 202768 520976 202774
rect 520924 202710 520976 202716
rect 530596 202706 530624 205006
rect 539612 205006 539948 205034
rect 539612 202842 539640 205006
rect 540072 202842 540100 224318
rect 539600 202836 539652 202842
rect 539600 202778 539652 202784
rect 540060 202836 540112 202842
rect 540060 202778 540112 202784
rect 541636 202774 541664 226374
rect 542360 223644 542412 223650
rect 542360 223586 542412 223592
rect 542372 214713 542400 223586
rect 542358 214704 542414 214713
rect 542358 214639 542414 214648
rect 541624 202768 541676 202774
rect 541624 202710 541676 202716
rect 530584 202700 530636 202706
rect 530584 202642 530636 202648
rect 529664 200252 529716 200258
rect 529664 200194 529716 200200
rect 541624 200252 541676 200258
rect 541624 200194 541676 200200
rect 529676 197948 529704 200194
rect 539324 200184 539376 200190
rect 539324 200126 539376 200132
rect 540244 200184 540296 200190
rect 540244 200126 540296 200132
rect 539336 197948 539364 200126
rect 519004 197254 520030 197282
rect 518806 188320 518862 188329
rect 518806 188255 518862 188264
rect 518820 179314 518848 188255
rect 518808 179308 518860 179314
rect 518808 179250 518860 179256
rect 519004 176526 519032 197254
rect 519636 180260 519688 180266
rect 519636 180202 519688 180208
rect 519648 178786 519676 180202
rect 539508 179376 539560 179382
rect 539508 179318 539560 179324
rect 539520 178786 539548 179318
rect 519648 178758 520030 178786
rect 539350 178758 539548 178786
rect 529676 176594 529704 178092
rect 540256 176594 540284 200126
rect 541636 179382 541664 200194
rect 542358 187640 542414 187649
rect 542358 187575 542414 187584
rect 541624 179376 541676 179382
rect 541624 179318 541676 179324
rect 542372 179246 542400 187575
rect 542360 179240 542412 179246
rect 542360 179182 542412 179188
rect 529664 176588 529716 176594
rect 529664 176530 529716 176536
rect 540244 176588 540296 176594
rect 540244 176530 540296 176536
rect 518992 176520 519044 176526
rect 518992 176462 519044 176468
rect 520280 172644 520332 172650
rect 520280 172586 520332 172592
rect 541624 172644 541676 172650
rect 541624 172586 541676 172592
rect 520292 170898 520320 172586
rect 529940 172576 529992 172582
rect 529940 172518 529992 172524
rect 529952 170898 529980 172518
rect 520292 170870 520628 170898
rect 529952 170870 530288 170898
rect 539948 170326 540100 170354
rect 518806 161392 518862 161401
rect 518806 161327 518862 161336
rect 518820 151706 518848 161327
rect 518808 151700 518860 151706
rect 518808 151642 518860 151648
rect 520628 151014 520964 151042
rect 530288 151014 530624 151042
rect 520936 148986 520964 151014
rect 520924 148980 520976 148986
rect 520924 148922 520976 148928
rect 530596 148918 530624 151014
rect 539612 151014 539948 151042
rect 539612 149054 539640 151014
rect 540072 149054 540100 170326
rect 539600 149048 539652 149054
rect 539600 148990 539652 148996
rect 540060 149048 540112 149054
rect 540060 148990 540112 148996
rect 541636 148986 541664 172586
rect 542358 160712 542414 160721
rect 542358 160647 542414 160656
rect 542372 151774 542400 160647
rect 542360 151768 542412 151774
rect 542360 151710 542412 151716
rect 541624 148980 541676 148986
rect 541624 148922 541676 148928
rect 530584 148912 530636 148918
rect 530584 148854 530636 148860
rect 529664 146396 529716 146402
rect 529664 146338 529716 146344
rect 541624 146396 541676 146402
rect 541624 146338 541676 146344
rect 529676 143956 529704 146338
rect 539324 146328 539376 146334
rect 539324 146270 539376 146276
rect 540244 146328 540296 146334
rect 540244 146270 540296 146276
rect 539336 143956 539364 146270
rect 519004 143262 520030 143290
rect 518806 134328 518862 134337
rect 518806 134263 518862 134272
rect 518820 125526 518848 134263
rect 518808 125520 518860 125526
rect 518808 125462 518860 125468
rect 519004 122670 519032 143262
rect 519636 126948 519688 126954
rect 519636 126890 519688 126896
rect 519648 124794 519676 126890
rect 519648 124766 520030 124794
rect 529676 122738 529704 124100
rect 539336 122806 539364 124100
rect 539324 122800 539376 122806
rect 539324 122742 539376 122748
rect 540256 122738 540284 146270
rect 541636 122806 541664 146338
rect 542358 133648 542414 133657
rect 542358 133583 542414 133592
rect 542372 125594 542400 133583
rect 542360 125588 542412 125594
rect 542360 125530 542412 125536
rect 541624 122800 541676 122806
rect 541624 122742 541676 122748
rect 529664 122732 529716 122738
rect 529664 122674 529716 122680
rect 540244 122732 540296 122738
rect 540244 122674 540296 122680
rect 518992 122664 519044 122670
rect 518992 122606 519044 122612
rect 541624 118856 541676 118862
rect 541624 118798 541676 118804
rect 520280 118788 520332 118794
rect 520280 118730 520332 118736
rect 520292 116906 520320 118730
rect 529940 118720 529992 118726
rect 529940 118662 529992 118668
rect 529952 116906 529980 118662
rect 520292 116878 520628 116906
rect 529952 116878 530288 116906
rect 539948 116334 540100 116362
rect 518806 107400 518862 107409
rect 518806 107335 518862 107344
rect 518820 97918 518848 107335
rect 518808 97912 518860 97918
rect 518808 97854 518860 97860
rect 520628 97022 520964 97050
rect 530288 97022 530624 97050
rect 520936 95130 520964 97022
rect 520924 95124 520976 95130
rect 520924 95066 520976 95072
rect 530596 95062 530624 97022
rect 539612 97022 539948 97050
rect 539612 95198 539640 97022
rect 540072 95198 540100 116334
rect 539600 95192 539652 95198
rect 539600 95134 539652 95140
rect 540060 95192 540112 95198
rect 540060 95134 540112 95140
rect 541636 95130 541664 118798
rect 542358 106720 542414 106729
rect 542358 106655 542414 106664
rect 542372 97986 542400 106655
rect 542360 97980 542412 97986
rect 542360 97922 542412 97928
rect 541624 95124 541676 95130
rect 541624 95066 541676 95072
rect 530584 95056 530636 95062
rect 530584 94998 530636 95004
rect 529664 91248 529716 91254
rect 529664 91190 529716 91196
rect 529676 89964 529704 91190
rect 541624 91180 541676 91186
rect 541624 91122 541676 91128
rect 539324 91112 539376 91118
rect 539324 91054 539376 91060
rect 540244 91112 540296 91118
rect 540244 91054 540296 91060
rect 539336 89964 539364 91054
rect 519004 89270 520030 89298
rect 518806 80336 518862 80345
rect 518806 80271 518862 80280
rect 518820 71738 518848 80271
rect 518808 71732 518860 71738
rect 518808 71674 518860 71680
rect 519004 68882 519032 89270
rect 519636 72140 519688 72146
rect 519636 72082 519688 72088
rect 519648 70666 519676 72082
rect 539508 71664 539560 71670
rect 539508 71606 539560 71612
rect 539520 70666 539548 71606
rect 519648 70638 520030 70666
rect 539350 70638 539548 70666
rect 529676 68950 529704 70108
rect 540256 68950 540284 91054
rect 541636 71670 541664 91122
rect 542360 88392 542412 88398
rect 542360 88334 542412 88340
rect 542372 79665 542400 88334
rect 542358 79656 542414 79665
rect 542358 79591 542414 79600
rect 541624 71664 541676 71670
rect 541624 71606 541676 71612
rect 529664 68944 529716 68950
rect 529664 68886 529716 68892
rect 540244 68944 540296 68950
rect 540244 68886 540296 68892
rect 518992 68876 519044 68882
rect 518992 68818 519044 68824
rect 520280 65000 520332 65006
rect 520280 64942 520332 64948
rect 541624 65000 541676 65006
rect 541624 64942 541676 64948
rect 520292 62914 520320 64942
rect 529940 64932 529992 64938
rect 529940 64874 529992 64880
rect 529952 62914 529980 64874
rect 520292 62886 520628 62914
rect 529952 62886 530288 62914
rect 539948 62206 540100 62234
rect 518806 53408 518862 53417
rect 518806 53343 518862 53352
rect 518820 44130 518848 53343
rect 518808 44124 518860 44130
rect 518808 44066 518860 44072
rect 520628 43030 520964 43058
rect 530288 43030 530624 43058
rect 520936 41342 520964 43030
rect 520924 41336 520976 41342
rect 520924 41278 520976 41284
rect 530596 41274 530624 43030
rect 539612 43030 539948 43058
rect 539612 41410 539640 43030
rect 540072 41410 540100 62206
rect 539600 41404 539652 41410
rect 539600 41346 539652 41352
rect 540060 41404 540112 41410
rect 540060 41346 540112 41352
rect 541636 41342 541664 64942
rect 542360 62144 542412 62150
rect 542360 62086 542412 62092
rect 542372 52737 542400 62086
rect 542358 52728 542414 52737
rect 542358 52663 542414 52672
rect 541624 41336 541676 41342
rect 541624 41278 541676 41284
rect 530584 41268 530636 41274
rect 530584 41210 530636 41216
rect 543016 38146 543044 673746
rect 569958 673568 570014 673577
rect 569958 673503 570014 673512
rect 569972 665174 570000 673503
rect 569960 665168 570012 665174
rect 569960 665110 570012 665116
rect 547892 664006 548044 664034
rect 557552 664006 557704 664034
rect 547892 662250 547920 664006
rect 547880 662244 547932 662250
rect 547880 662186 547932 662192
rect 557552 661706 557580 664006
rect 557540 661700 557592 661706
rect 557540 661642 557592 661648
rect 544384 658300 544436 658306
rect 544384 658242 544436 658248
rect 548616 658300 548668 658306
rect 548616 658242 548668 658248
rect 558276 658300 558328 658306
rect 558276 658242 558328 658248
rect 544396 634642 544424 658242
rect 548628 656948 548656 658242
rect 558288 656948 558316 658242
rect 567962 656254 568068 656282
rect 546406 647456 546462 647465
rect 546406 647391 546462 647400
rect 544384 634636 544436 634642
rect 544384 634578 544436 634584
rect 546420 620265 546448 647391
rect 547892 637078 548642 637106
rect 546406 620256 546462 620265
rect 546406 620191 546462 620200
rect 547892 610706 547920 637078
rect 558288 634098 558316 637092
rect 567948 634778 567976 637092
rect 567936 634772 567988 634778
rect 567936 634714 567988 634720
rect 558276 634092 558328 634098
rect 558276 634034 558328 634040
rect 567476 634092 567528 634098
rect 567476 634034 567528 634040
rect 548340 632732 548392 632738
rect 548340 632674 548392 632680
rect 548352 629898 548380 632674
rect 557540 632188 557592 632194
rect 557540 632130 557592 632136
rect 548044 629870 548380 629898
rect 557552 629762 557580 632130
rect 567200 632120 567252 632126
rect 567200 632062 567252 632068
rect 567212 629762 567240 632062
rect 557552 629734 557704 629762
rect 567212 629734 567364 629762
rect 567488 610722 567516 634034
rect 568040 632738 568068 656254
rect 569960 655648 570012 655654
rect 569960 655590 570012 655596
rect 569972 646785 570000 655590
rect 569958 646776 570014 646785
rect 569958 646711 570014 646720
rect 568028 632732 568080 632738
rect 568028 632674 568080 632680
rect 569958 619576 570014 619585
rect 569958 619511 570014 619520
rect 569972 611250 570000 619511
rect 569960 611244 570012 611250
rect 569960 611186 570012 611192
rect 547880 610700 547932 610706
rect 547880 610642 547932 610648
rect 548156 610700 548208 610706
rect 567364 610694 567516 610722
rect 548156 610642 548208 610648
rect 547892 610014 548044 610042
rect 547892 608462 547920 610014
rect 548168 608598 548196 610642
rect 557552 610014 557704 610042
rect 557552 608598 557580 610014
rect 548156 608592 548208 608598
rect 548156 608534 548208 608540
rect 557540 608592 557592 608598
rect 557540 608534 557592 608540
rect 547880 608456 547932 608462
rect 547880 608398 547932 608404
rect 544384 604512 544436 604518
rect 544384 604454 544436 604460
rect 548616 604512 548668 604518
rect 548616 604454 548668 604460
rect 558276 604512 558328 604518
rect 558276 604454 558328 604460
rect 544396 580854 544424 604454
rect 548628 602956 548656 604454
rect 558288 602956 558316 604454
rect 567962 602262 568068 602290
rect 546406 593464 546462 593473
rect 546406 593399 546462 593408
rect 544384 580848 544436 580854
rect 544384 580790 544436 580796
rect 546420 566273 546448 593399
rect 547892 583086 548642 583114
rect 546406 566264 546462 566273
rect 546406 566199 546462 566208
rect 547892 556170 547920 583086
rect 558288 580310 558316 583100
rect 567948 580990 567976 583100
rect 567936 580984 567988 580990
rect 567936 580926 567988 580932
rect 558276 580304 558328 580310
rect 558276 580246 558328 580252
rect 567476 580304 567528 580310
rect 567476 580246 567528 580252
rect 548340 578944 548392 578950
rect 548340 578886 548392 578892
rect 548352 575906 548380 578886
rect 557540 578332 557592 578338
rect 557540 578274 557592 578280
rect 548044 575878 548380 575906
rect 557552 575906 557580 578274
rect 567200 578264 567252 578270
rect 567200 578206 567252 578212
rect 567212 575906 567240 578206
rect 557552 575878 557704 575906
rect 567212 575878 567364 575906
rect 567488 556730 567516 580246
rect 568040 578950 568068 602262
rect 569960 601792 570012 601798
rect 569960 601734 570012 601740
rect 569972 592793 570000 601734
rect 569958 592784 570014 592793
rect 569958 592719 570014 592728
rect 580262 591016 580318 591025
rect 580262 590951 580318 590960
rect 568028 578944 568080 578950
rect 568028 578886 568080 578892
rect 569958 565584 570014 565593
rect 569958 565519 570014 565528
rect 569972 557462 570000 565519
rect 569960 557456 570012 557462
rect 569960 557398 570012 557404
rect 567364 556702 567516 556730
rect 547880 556164 547932 556170
rect 547880 556106 547932 556112
rect 548156 556164 548208 556170
rect 548156 556106 548208 556112
rect 547892 556022 548044 556050
rect 547892 554606 547920 556022
rect 548168 554742 548196 556106
rect 557552 556022 557704 556050
rect 557552 554742 557580 556022
rect 548156 554736 548208 554742
rect 548156 554678 548208 554684
rect 557540 554736 557592 554742
rect 557540 554678 557592 554684
rect 547880 554600 547932 554606
rect 547880 554542 547932 554548
rect 544384 550656 544436 550662
rect 544384 550598 544436 550604
rect 548616 550656 548668 550662
rect 548616 550598 548668 550604
rect 558276 550656 558328 550662
rect 558276 550598 558328 550604
rect 544396 526998 544424 550598
rect 548628 548964 548656 550598
rect 558288 548964 558316 550598
rect 567962 548270 568068 548298
rect 546406 539472 546462 539481
rect 546406 539407 546462 539416
rect 544384 526992 544436 526998
rect 544384 526934 544436 526940
rect 546420 512281 546448 539407
rect 547892 529094 548642 529122
rect 546406 512272 546462 512281
rect 546406 512207 546462 512216
rect 547892 502722 547920 529094
rect 558288 526454 558316 529108
rect 567948 527134 567976 529108
rect 567936 527128 567988 527134
rect 567936 527070 567988 527076
rect 558276 526448 558328 526454
rect 558276 526390 558328 526396
rect 567476 526448 567528 526454
rect 567476 526390 567528 526396
rect 548340 523728 548392 523734
rect 548340 523670 548392 523676
rect 548352 521914 548380 523670
rect 557540 523116 557592 523122
rect 557540 523058 557592 523064
rect 548044 521886 548380 521914
rect 557552 521778 557580 523058
rect 567200 523048 567252 523054
rect 567200 522990 567252 522996
rect 567212 521778 567240 522990
rect 557552 521750 557704 521778
rect 567212 521750 567364 521778
rect 567488 502738 567516 526390
rect 568040 523734 568068 548270
rect 569958 538792 570014 538801
rect 569958 538727 570014 538736
rect 569972 529854 570000 538727
rect 569960 529848 570012 529854
rect 569960 529790 570012 529796
rect 568028 523728 568080 523734
rect 568028 523670 568080 523676
rect 569958 511592 570014 511601
rect 569958 511527 570014 511536
rect 569972 503674 570000 511527
rect 569960 503668 570012 503674
rect 569960 503610 570012 503616
rect 547880 502716 547932 502722
rect 547880 502658 547932 502664
rect 548156 502716 548208 502722
rect 567364 502710 567516 502738
rect 548156 502658 548208 502664
rect 547892 502030 548044 502058
rect 547892 500818 547920 502030
rect 548168 500954 548196 502658
rect 557552 502030 557704 502058
rect 557552 500954 557580 502030
rect 548156 500948 548208 500954
rect 548156 500890 548208 500896
rect 557540 500948 557592 500954
rect 557540 500890 557592 500896
rect 547880 500812 547932 500818
rect 547880 500754 547932 500760
rect 558276 496868 558328 496874
rect 558276 496810 558328 496816
rect 558288 494972 558316 496810
rect 548352 494278 548642 494306
rect 567962 494278 568068 494306
rect 548352 494086 548380 494278
rect 544384 494080 544436 494086
rect 544384 494022 544436 494028
rect 548340 494080 548392 494086
rect 548340 494022 548392 494028
rect 544396 473210 544424 494022
rect 546406 485480 546462 485489
rect 546406 485415 546462 485424
rect 544384 473204 544436 473210
rect 544384 473146 544436 473152
rect 546420 458289 546448 485415
rect 547892 475102 548642 475130
rect 546406 458280 546462 458289
rect 546406 458215 546462 458224
rect 547892 448526 547920 475102
rect 558288 472666 558316 475116
rect 567948 473346 567976 475116
rect 567936 473340 567988 473346
rect 567936 473282 567988 473288
rect 558276 472660 558328 472666
rect 558276 472602 558328 472608
rect 567476 472660 567528 472666
rect 567476 472602 567528 472608
rect 548340 469872 548392 469878
rect 548340 469814 548392 469820
rect 548352 467922 548380 469814
rect 557540 469328 557592 469334
rect 557540 469270 557592 469276
rect 548044 467894 548380 467922
rect 557552 467786 557580 469270
rect 567200 469260 567252 469266
rect 567200 469202 567252 469208
rect 567212 467786 567240 469202
rect 557552 467758 557704 467786
rect 567212 467758 567364 467786
rect 567488 448746 567516 472602
rect 568040 469878 568068 494278
rect 569958 484800 570014 484809
rect 569958 484735 570014 484744
rect 569972 475998 570000 484735
rect 569960 475992 570012 475998
rect 569960 475934 570012 475940
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 568028 469872 568080 469878
rect 568028 469814 568080 469820
rect 569960 466540 570012 466546
rect 569960 466482 570012 466488
rect 569972 457609 570000 466482
rect 569958 457600 570014 457609
rect 569958 457535 570014 457544
rect 567364 448718 567516 448746
rect 547880 448520 547932 448526
rect 547880 448462 547932 448468
rect 548156 448520 548208 448526
rect 548156 448462 548208 448468
rect 547892 448038 548044 448066
rect 547892 445602 547920 448038
rect 548168 445738 548196 448462
rect 557552 448038 557704 448066
rect 557552 445738 557580 448038
rect 548156 445732 548208 445738
rect 548156 445674 548208 445680
rect 557540 445732 557592 445738
rect 557540 445674 557592 445680
rect 547880 445596 547932 445602
rect 547880 445538 547932 445544
rect 558276 443012 558328 443018
rect 558276 442954 558328 442960
rect 558288 440980 558316 442954
rect 548352 440298 548642 440314
rect 544384 440292 544436 440298
rect 544384 440234 544436 440240
rect 548340 440292 548642 440298
rect 548392 440286 548642 440292
rect 567962 440286 568068 440314
rect 548340 440234 548392 440240
rect 544396 419354 544424 440234
rect 546406 431488 546462 431497
rect 546406 431423 546462 431432
rect 544384 419348 544436 419354
rect 544384 419290 544436 419296
rect 546420 404297 546448 431423
rect 547892 421110 548642 421138
rect 546406 404288 546462 404297
rect 546406 404223 546462 404232
rect 547892 394738 547920 421110
rect 558288 418810 558316 421124
rect 567948 419490 567976 421124
rect 567936 419484 567988 419490
rect 567936 419426 567988 419432
rect 558276 418804 558328 418810
rect 558276 418746 558328 418752
rect 567476 418804 567528 418810
rect 567476 418746 567528 418752
rect 548340 416084 548392 416090
rect 548340 416026 548392 416032
rect 548352 413930 548380 416026
rect 557540 415540 557592 415546
rect 557540 415482 557592 415488
rect 548044 413902 548380 413930
rect 557552 413794 557580 415482
rect 567200 415472 567252 415478
rect 567200 415414 567252 415420
rect 567212 413794 567240 415414
rect 557552 413766 557704 413794
rect 567212 413766 567364 413794
rect 567488 394754 567516 418746
rect 568040 416090 568068 440286
rect 569958 430808 570014 430817
rect 569958 430743 570014 430752
rect 569972 422278 570000 430743
rect 569960 422272 570012 422278
rect 569960 422214 570012 422220
rect 568028 416084 568080 416090
rect 568028 416026 568080 416032
rect 569958 403608 570014 403617
rect 569958 403543 570014 403552
rect 547880 394732 547932 394738
rect 547880 394674 547932 394680
rect 548156 394732 548208 394738
rect 567364 394726 567516 394754
rect 548156 394674 548208 394680
rect 547892 394046 548044 394074
rect 547892 391814 547920 394046
rect 548168 391950 548196 394674
rect 569972 394602 570000 403543
rect 569960 394596 570012 394602
rect 569960 394538 570012 394544
rect 557552 394046 557704 394074
rect 557552 391950 557580 394046
rect 548156 391944 548208 391950
rect 548156 391886 548208 391892
rect 557540 391944 557592 391950
rect 557540 391886 557592 391892
rect 547880 391808 547932 391814
rect 547880 391750 547932 391756
rect 558276 389224 558328 389230
rect 558276 389166 558328 389172
rect 558288 386852 558316 389166
rect 569960 386504 570012 386510
rect 548352 386442 548642 386458
rect 569960 386446 570012 386452
rect 544384 386436 544436 386442
rect 544384 386378 544436 386384
rect 548340 386436 548642 386442
rect 548392 386430 548642 386436
rect 548340 386378 548392 386384
rect 544396 365566 544424 386378
rect 567962 386294 568160 386322
rect 568132 383654 568160 386294
rect 568132 383626 568344 383654
rect 568120 378208 568172 378214
rect 568120 378150 568172 378156
rect 546406 377088 546462 377097
rect 546406 377023 546462 377032
rect 544384 365560 544436 365566
rect 544384 365502 544436 365508
rect 546420 350305 546448 377023
rect 568132 376258 568160 378150
rect 568040 376230 568160 376258
rect 547892 367118 548642 367146
rect 546406 350296 546462 350305
rect 546406 350231 546462 350240
rect 547892 340610 547920 367118
rect 558288 365022 558316 367132
rect 567948 365702 567976 367132
rect 567936 365696 567988 365702
rect 567936 365638 567988 365644
rect 558276 365016 558328 365022
rect 558276 364958 558328 364964
rect 567476 365016 567528 365022
rect 567476 364958 567528 364964
rect 548340 362228 548392 362234
rect 548340 362170 548392 362176
rect 548352 359938 548380 362170
rect 557540 361684 557592 361690
rect 557540 361626 557592 361632
rect 548044 359910 548380 359938
rect 557552 359802 557580 361626
rect 567200 361616 567252 361622
rect 567200 361558 567252 361564
rect 567212 359802 567240 361558
rect 557552 359774 557704 359802
rect 567212 359774 567364 359802
rect 567488 340762 567516 364958
rect 567364 340734 567516 340762
rect 547880 340604 547932 340610
rect 547880 340546 547932 340552
rect 548156 340604 548208 340610
rect 548156 340546 548208 340552
rect 547892 340054 548044 340082
rect 547892 337958 547920 340054
rect 548168 338094 548196 340546
rect 557552 340054 557704 340082
rect 557552 338094 557580 340054
rect 548156 338088 548208 338094
rect 548156 338030 548208 338036
rect 557540 338088 557592 338094
rect 557540 338030 557592 338036
rect 547880 337952 547932 337958
rect 547880 337894 547932 337900
rect 558276 335368 558328 335374
rect 558276 335310 558328 335316
rect 558288 332860 558316 335310
rect 548352 332586 548642 332602
rect 544384 332580 544436 332586
rect 544384 332522 544436 332528
rect 548340 332580 548642 332586
rect 548392 332574 548642 332580
rect 548340 332522 548392 332528
rect 544396 311710 544424 332522
rect 568040 332450 568068 376230
rect 568316 375986 568344 383626
rect 569972 376825 570000 386446
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 569958 376816 570014 376825
rect 569958 376751 570014 376760
rect 568132 375958 568344 375986
rect 568132 362234 568160 375958
rect 568120 362228 568172 362234
rect 568120 362170 568172 362176
rect 569958 349616 570014 349625
rect 569958 349551 570014 349560
rect 569972 340814 570000 349551
rect 569960 340808 570012 340814
rect 569960 340750 570012 340756
rect 568028 332444 568080 332450
rect 568028 332386 568080 332392
rect 567962 332302 568160 332330
rect 568028 332240 568080 332246
rect 568028 332182 568080 332188
rect 546406 322960 546462 322969
rect 546406 322895 546462 322904
rect 544384 311704 544436 311710
rect 544384 311646 544436 311652
rect 546420 296313 546448 322895
rect 547892 313126 548642 313154
rect 546406 296304 546462 296313
rect 546406 296239 546462 296248
rect 547892 286210 547920 313126
rect 558288 311166 558316 313140
rect 567948 311846 567976 313140
rect 567936 311840 567988 311846
rect 567936 311782 567988 311788
rect 558276 311160 558328 311166
rect 558276 311102 558328 311108
rect 567476 311160 567528 311166
rect 567476 311102 567528 311108
rect 548340 308440 548392 308446
rect 548340 308382 548392 308388
rect 548352 305946 548380 308382
rect 557540 307896 557592 307902
rect 557540 307838 557592 307844
rect 548044 305918 548380 305946
rect 557552 305946 557580 307838
rect 567200 307828 567252 307834
rect 567200 307770 567252 307776
rect 567212 305946 567240 307770
rect 557552 305918 557704 305946
rect 567212 305918 567364 305946
rect 567488 286770 567516 311102
rect 567364 286742 567516 286770
rect 547880 286204 547932 286210
rect 547880 286146 547932 286152
rect 548156 286204 548208 286210
rect 548156 286146 548208 286152
rect 547892 286062 548044 286090
rect 547892 284170 547920 286062
rect 548168 284306 548196 286146
rect 557552 286062 557704 286090
rect 557552 284306 557580 286062
rect 548156 284300 548208 284306
rect 548156 284242 548208 284248
rect 557540 284300 557592 284306
rect 557540 284242 557592 284248
rect 547880 284164 547932 284170
rect 547880 284106 547932 284112
rect 544384 280220 544436 280226
rect 544384 280162 544436 280168
rect 548616 280220 548668 280226
rect 548616 280162 548668 280168
rect 558276 280220 558328 280226
rect 558276 280162 558328 280168
rect 544396 256562 544424 280162
rect 548628 278868 548656 280162
rect 558288 278868 558316 280162
rect 568040 278458 568068 332182
rect 568132 308446 568160 332302
rect 579986 325272 580042 325281
rect 579986 325207 580042 325216
rect 580000 324358 580028 325207
rect 570604 324352 570656 324358
rect 570604 324294 570656 324300
rect 579988 324352 580040 324358
rect 579988 324294 580040 324300
rect 569958 322144 570014 322153
rect 569958 322079 570014 322088
rect 569972 314634 570000 322079
rect 569960 314628 570012 314634
rect 569960 314570 570012 314576
rect 568120 308440 568172 308446
rect 568120 308382 568172 308388
rect 569958 295624 570014 295633
rect 569958 295559 570014 295568
rect 569972 286958 570000 295559
rect 569960 286952 570012 286958
rect 569960 286894 570012 286900
rect 568028 278452 568080 278458
rect 568028 278394 568080 278400
rect 567962 278310 568160 278338
rect 568028 278248 568080 278254
rect 568028 278190 568080 278196
rect 546406 269240 546462 269249
rect 546406 269175 546462 269184
rect 544384 256556 544436 256562
rect 544384 256498 544436 256504
rect 546420 242321 546448 269175
rect 547892 259134 548642 259162
rect 546406 242312 546462 242321
rect 546406 242247 546462 242256
rect 547892 232762 547920 259134
rect 558288 256018 558316 259148
rect 567948 256698 567976 259148
rect 567936 256692 567988 256698
rect 567936 256634 567988 256640
rect 558276 256012 558328 256018
rect 558276 255954 558328 255960
rect 567476 256012 567528 256018
rect 567476 255954 567528 255960
rect 548340 254584 548392 254590
rect 548340 254526 548392 254532
rect 548352 251954 548380 254526
rect 557540 254040 557592 254046
rect 557540 253982 557592 253988
rect 548044 251926 548380 251954
rect 557552 251818 557580 253982
rect 567200 253972 567252 253978
rect 567200 253914 567252 253920
rect 567212 251818 567240 253914
rect 557552 251790 557704 251818
rect 567212 251790 567364 251818
rect 567488 232778 567516 255954
rect 547880 232756 547932 232762
rect 547880 232698 547932 232704
rect 548156 232756 548208 232762
rect 567364 232750 567516 232778
rect 548156 232698 548208 232704
rect 547892 232070 548044 232098
rect 547892 230314 547920 232070
rect 548168 230450 548196 232698
rect 557552 232070 557704 232098
rect 557552 230450 557580 232070
rect 548156 230444 548208 230450
rect 548156 230386 548208 230392
rect 557540 230444 557592 230450
rect 557540 230386 557592 230392
rect 547880 230308 547932 230314
rect 547880 230250 547932 230256
rect 544384 226364 544436 226370
rect 544384 226306 544436 226312
rect 548616 226364 548668 226370
rect 548616 226306 548668 226312
rect 558276 226364 558328 226370
rect 558276 226306 558328 226312
rect 544396 202706 544424 226306
rect 548628 224876 548656 226306
rect 558288 224876 558316 226306
rect 568040 224466 568068 278190
rect 568132 254590 568160 278310
rect 569960 277500 570012 277506
rect 569960 277442 570012 277448
rect 569972 269113 570000 277442
rect 569958 269104 570014 269113
rect 569958 269039 570014 269048
rect 568120 254584 568172 254590
rect 568120 254526 568172 254532
rect 569960 251320 570012 251326
rect 569960 251262 570012 251268
rect 569972 241641 570000 251262
rect 569958 241632 570014 241641
rect 569958 241567 570014 241576
rect 568028 224460 568080 224466
rect 568028 224402 568080 224408
rect 567962 224318 568160 224346
rect 568028 224256 568080 224262
rect 568028 224198 568080 224204
rect 546406 215520 546462 215529
rect 546406 215455 546462 215464
rect 544384 202700 544436 202706
rect 544384 202642 544436 202648
rect 546420 188329 546448 215455
rect 547892 205006 548642 205034
rect 546406 188320 546462 188329
rect 546406 188255 546462 188264
rect 547892 178770 547920 205006
rect 558288 202162 558316 205020
rect 567948 202842 567976 205020
rect 567936 202836 567988 202842
rect 567936 202778 567988 202784
rect 558276 202156 558328 202162
rect 558276 202098 558328 202104
rect 567476 202156 567528 202162
rect 567476 202098 567528 202104
rect 548340 200796 548392 200802
rect 548340 200738 548392 200744
rect 548352 197962 548380 200738
rect 557540 200252 557592 200258
rect 557540 200194 557592 200200
rect 548044 197934 548380 197962
rect 557552 197962 557580 200194
rect 567200 200184 567252 200190
rect 567200 200126 567252 200132
rect 567212 197962 567240 200126
rect 557552 197934 557704 197962
rect 567212 197934 567364 197962
rect 567488 178786 567516 202098
rect 547880 178764 547932 178770
rect 547880 178706 547932 178712
rect 548156 178764 548208 178770
rect 567364 178758 567516 178786
rect 548156 178706 548208 178712
rect 547892 178078 548044 178106
rect 547892 176526 547920 178078
rect 548168 176662 548196 178706
rect 557552 178078 557704 178106
rect 557552 176662 557580 178078
rect 548156 176656 548208 176662
rect 548156 176598 548208 176604
rect 557540 176656 557592 176662
rect 557540 176598 557592 176604
rect 547880 176520 547932 176526
rect 547880 176462 547932 176468
rect 544384 172576 544436 172582
rect 544384 172518 544436 172524
rect 548616 172576 548668 172582
rect 548616 172518 548668 172524
rect 558276 172576 558328 172582
rect 558276 172518 558328 172524
rect 544396 148918 544424 172518
rect 548628 170884 548656 172518
rect 558288 170884 558316 172518
rect 568040 170474 568068 224198
rect 568132 200802 568160 224318
rect 569960 223712 570012 223718
rect 569960 223654 570012 223660
rect 569972 214713 570000 223654
rect 569958 214704 570014 214713
rect 569958 214639 570014 214648
rect 568120 200796 568172 200802
rect 568120 200738 568172 200744
rect 569958 187640 570014 187649
rect 569958 187575 570014 187584
rect 569972 179314 570000 187575
rect 569960 179308 570012 179314
rect 569960 179250 570012 179256
rect 568028 170468 568080 170474
rect 568028 170410 568080 170416
rect 567962 170326 568160 170354
rect 568028 170264 568080 170270
rect 568028 170206 568080 170212
rect 546406 161392 546462 161401
rect 546406 161327 546462 161336
rect 544384 148912 544436 148918
rect 544384 148854 544436 148860
rect 546420 134337 546448 161327
rect 547892 151014 548642 151042
rect 546406 134328 546462 134337
rect 546406 134263 546462 134272
rect 547892 124710 547920 151014
rect 558288 148374 558316 151028
rect 567948 149054 567976 151028
rect 567936 149048 567988 149054
rect 567936 148990 567988 148996
rect 558276 148368 558328 148374
rect 558276 148310 558328 148316
rect 567476 148368 567528 148374
rect 567476 148310 567528 148316
rect 548340 146940 548392 146946
rect 548340 146882 548392 146888
rect 548352 143970 548380 146882
rect 557540 146396 557592 146402
rect 557540 146338 557592 146344
rect 548044 143942 548380 143970
rect 557552 143834 557580 146338
rect 567200 146328 567252 146334
rect 567200 146270 567252 146276
rect 567212 143834 567240 146270
rect 557552 143806 557704 143834
rect 567212 143806 567364 143834
rect 567488 124794 567516 148310
rect 567364 124766 567516 124794
rect 547880 124704 547932 124710
rect 547880 124646 547932 124652
rect 548156 124704 548208 124710
rect 548156 124646 548208 124652
rect 547892 124086 548044 124114
rect 547892 122670 547920 124086
rect 548168 122806 548196 124646
rect 557552 124086 557704 124114
rect 557552 122806 557580 124086
rect 548156 122800 548208 122806
rect 548156 122742 548208 122748
rect 557540 122800 557592 122806
rect 557540 122742 557592 122748
rect 547880 122664 547932 122670
rect 547880 122606 547932 122612
rect 558276 118788 558328 118794
rect 558276 118730 558328 118736
rect 544384 118720 544436 118726
rect 544384 118662 544436 118668
rect 548616 118720 548668 118726
rect 548616 118662 548668 118668
rect 544396 95062 544424 118662
rect 547972 118652 548024 118658
rect 547972 118594 548024 118600
rect 546406 107400 546462 107409
rect 546406 107335 546462 107344
rect 544384 95056 544436 95062
rect 544384 94998 544436 95004
rect 546420 80345 546448 107335
rect 547880 95464 547932 95470
rect 547880 95406 547932 95412
rect 546406 80336 546462 80345
rect 546406 80271 546462 80280
rect 547892 70718 547920 95406
rect 547984 90250 548012 118594
rect 548628 116892 548656 118662
rect 558288 116892 558316 118730
rect 567936 118720 567988 118726
rect 567936 118662 567988 118668
rect 567948 116892 567976 118662
rect 548352 97022 548642 97050
rect 548352 95470 548380 97022
rect 548340 95464 548392 95470
rect 548340 95406 548392 95412
rect 558288 94518 558316 97036
rect 567948 95198 567976 97036
rect 567936 95192 567988 95198
rect 567936 95134 567988 95140
rect 558276 94512 558328 94518
rect 558276 94454 558328 94460
rect 567476 94512 567528 94518
rect 567476 94454 567528 94460
rect 557540 91180 557592 91186
rect 557540 91122 557592 91128
rect 547984 90222 548058 90250
rect 548030 89964 548058 90222
rect 557552 89842 557580 91122
rect 567200 91112 567252 91118
rect 567200 91054 567252 91060
rect 567212 89842 567240 91054
rect 557552 89814 557704 89842
rect 567212 89814 567364 89842
rect 547880 70712 547932 70718
rect 547880 70654 547932 70660
rect 548156 70712 548208 70718
rect 567488 70666 567516 94454
rect 548156 70654 548208 70660
rect 547892 70094 548044 70122
rect 547892 68882 547920 70094
rect 548168 69018 548196 70654
rect 567364 70638 567516 70666
rect 557552 70094 557704 70122
rect 557552 69018 557580 70094
rect 548156 69012 548208 69018
rect 548156 68954 548208 68960
rect 557540 69012 557592 69018
rect 557540 68954 557592 68960
rect 547880 68876 547932 68882
rect 547880 68818 547932 68824
rect 558276 65000 558328 65006
rect 558276 64942 558328 64948
rect 547972 64932 548024 64938
rect 547972 64874 548024 64880
rect 544384 62144 544436 62150
rect 544384 62086 544436 62092
rect 544396 41274 544424 62086
rect 546406 53408 546462 53417
rect 546406 53343 546462 53352
rect 544384 41268 544436 41274
rect 544384 41210 544436 41216
rect 543004 38140 543056 38146
rect 543004 38082 543056 38088
rect 518256 37392 518308 37398
rect 518256 37334 518308 37340
rect 529664 37392 529716 37398
rect 529664 37334 529716 37340
rect 541624 37392 541676 37398
rect 541624 37334 541676 37340
rect 518268 13462 518296 37334
rect 529676 35972 529704 37334
rect 539324 37324 539376 37330
rect 539324 37266 539376 37272
rect 540244 37324 540296 37330
rect 540244 37266 540296 37272
rect 539336 35972 539364 37266
rect 519004 35278 520030 35306
rect 518808 34604 518860 34610
rect 518808 34546 518860 34552
rect 518820 26353 518848 34546
rect 518806 26344 518862 26353
rect 518806 26279 518862 26288
rect 519004 13462 519032 35278
rect 519636 18012 519688 18018
rect 519636 17954 519688 17960
rect 519648 16674 519676 17954
rect 519648 16646 520030 16674
rect 539508 16584 539560 16590
rect 539350 16532 539508 16538
rect 539350 16526 539560 16532
rect 539350 16510 539548 16526
rect 529676 13802 529704 16116
rect 540256 13802 540284 37266
rect 541636 16590 541664 37334
rect 542360 34536 542412 34542
rect 542360 34478 542412 34484
rect 542372 25673 542400 34478
rect 546420 26353 546448 53343
rect 547880 38548 547932 38554
rect 547880 38490 547932 38496
rect 546406 26344 546462 26353
rect 546406 26279 546462 26288
rect 542358 25664 542414 25673
rect 542358 25599 542414 25608
rect 541624 16584 541676 16590
rect 541624 16526 541676 16532
rect 547892 13802 547920 38490
rect 547984 36258 548012 64874
rect 558288 62900 558316 64942
rect 567936 64932 567988 64938
rect 567936 64874 567988 64880
rect 567948 62900 567976 64874
rect 548352 62206 548642 62234
rect 548352 62150 548380 62206
rect 548340 62144 548392 62150
rect 548340 62086 548392 62092
rect 548352 43030 548642 43058
rect 548352 38554 548380 43030
rect 558288 40730 558316 43044
rect 567948 41410 567976 43044
rect 567936 41404 567988 41410
rect 567936 41346 567988 41352
rect 558276 40724 558328 40730
rect 558276 40666 558328 40672
rect 567476 40724 567528 40730
rect 567476 40666 567528 40672
rect 548340 38548 548392 38554
rect 548340 38490 548392 38496
rect 557540 37392 557592 37398
rect 557540 37334 557592 37340
rect 547984 36230 548058 36258
rect 548030 35972 548058 36230
rect 557552 35986 557580 37334
rect 567200 37324 567252 37330
rect 567200 37266 567252 37272
rect 557552 35958 557704 35986
rect 567212 35894 567240 37266
rect 567350 35894 567378 35972
rect 567212 35866 567378 35894
rect 567488 16674 567516 40666
rect 568040 36786 568068 170206
rect 568132 146946 568160 170326
rect 569958 160712 570014 160721
rect 569958 160647 570014 160656
rect 569972 151706 570000 160647
rect 569960 151700 570012 151706
rect 569960 151642 570012 151648
rect 568120 146940 568172 146946
rect 568120 146882 568172 146888
rect 569958 133648 570014 133657
rect 569958 133583 570014 133592
rect 569972 125526 570000 133583
rect 569960 125520 570012 125526
rect 569960 125462 570012 125468
rect 569958 106720 570014 106729
rect 569958 106655 570014 106664
rect 569972 97918 570000 106655
rect 569960 97912 570012 97918
rect 569960 97854 570012 97860
rect 569958 79656 570014 79665
rect 569958 79591 570014 79600
rect 569972 71738 570000 79591
rect 569960 71732 570012 71738
rect 569960 71674 570012 71680
rect 569958 52728 570014 52737
rect 569958 52663 570014 52672
rect 569972 44130 570000 52663
rect 569960 44124 570012 44130
rect 569960 44066 570012 44072
rect 568028 36780 568080 36786
rect 568028 36722 568080 36728
rect 569960 34604 570012 34610
rect 569960 34546 570012 34552
rect 569972 25673 570000 34546
rect 569958 25664 570014 25673
rect 569958 25599 570014 25608
rect 567364 16646 567516 16674
rect 548030 15858 548058 16116
rect 547984 15830 548058 15858
rect 557552 16102 557704 16130
rect 529664 13796 529716 13802
rect 529664 13738 529716 13744
rect 540244 13796 540296 13802
rect 540244 13738 540296 13744
rect 547880 13796 547932 13802
rect 547880 13738 547932 13744
rect 547984 13462 548012 15830
rect 557552 13802 557580 16102
rect 557540 13796 557592 13802
rect 557540 13738 557592 13744
rect 570616 13734 570644 324294
rect 578882 272232 578938 272241
rect 578882 272167 578938 272176
rect 570696 191888 570748 191894
rect 570696 191830 570748 191836
rect 570708 38214 570736 191830
rect 570696 38208 570748 38214
rect 570696 38150 570748 38156
rect 570604 13728 570656 13734
rect 570604 13670 570656 13676
rect 518256 13456 518308 13462
rect 518256 13398 518308 13404
rect 518992 13456 519044 13462
rect 518992 13398 519044 13404
rect 547972 13456 548024 13462
rect 547972 13398 548024 13404
rect 344284 13262 344336 13268
rect 518162 13288 518218 13297
rect 238852 13252 238904 13258
rect 238852 13194 238904 13200
rect 268016 13252 268068 13258
rect 518162 13223 518218 13232
rect 268016 13194 268068 13200
rect 72056 13116 72108 13122
rect 72056 13058 72108 13064
rect 578896 13054 578924 272167
rect 579802 232384 579858 232393
rect 579802 232319 579858 232328
rect 579816 231878 579844 232319
rect 579804 231872 579856 231878
rect 579804 231814 579856 231820
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580184 191894 580212 192471
rect 580172 191888 580224 191894
rect 580172 191830 580224 191836
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580078 72992 580134 73001
rect 580078 72927 580134 72936
rect 579988 35964 580040 35970
rect 579988 35906 580040 35912
rect 580000 33153 580028 35906
rect 579986 33144 580042 33153
rect 579986 33079 580042 33088
rect 580092 13666 580120 72927
rect 580184 36718 580212 112775
rect 580172 36712 580224 36718
rect 580172 36654 580224 36660
rect 580276 36650 580304 590951
rect 580354 537840 580410 537849
rect 580354 537775 580410 537784
rect 580264 36644 580316 36650
rect 580264 36586 580316 36592
rect 580368 35222 580396 537775
rect 580446 511320 580502 511329
rect 580446 511255 580502 511264
rect 580460 38010 580488 511255
rect 580538 484664 580594 484673
rect 580538 484599 580594 484608
rect 580448 38004 580500 38010
rect 580448 37946 580500 37952
rect 580356 35216 580408 35222
rect 580356 35158 580408 35164
rect 580080 13660 580132 13666
rect 580080 13602 580132 13608
rect 580552 13598 580580 484599
rect 580630 431624 580686 431633
rect 580630 431559 580686 431568
rect 580644 36582 580672 431559
rect 580722 404968 580778 404977
rect 580722 404903 580778 404912
rect 580736 37942 580764 404903
rect 580814 351928 580870 351937
rect 580814 351863 580870 351872
rect 580724 37936 580776 37942
rect 580724 37878 580776 37884
rect 580632 36576 580684 36582
rect 580632 36518 580684 36524
rect 580540 13592 580592 13598
rect 580540 13534 580592 13540
rect 580828 13530 580856 351863
rect 580906 152688 580962 152697
rect 580906 152623 580962 152632
rect 580920 38078 580948 152623
rect 580908 38072 580960 38078
rect 580908 38014 580960 38020
rect 580816 13524 580868 13530
rect 580816 13466 580868 13472
rect 578884 13048 578936 13054
rect 578884 12990 578936 12996
rect 64420 3732 64472 3738
rect 64420 3674 64472 3680
rect 125876 3732 125928 3738
rect 125876 3674 125928 3680
rect 64236 3664 64288 3670
rect 64236 3606 64288 3612
rect 48320 3460 48372 3466
rect 48320 3402 48372 3408
rect 61476 3460 61528 3466
rect 61476 3402 61528 3408
rect 125888 480 125916 3674
rect 126980 3664 127032 3670
rect 126980 3606 127032 3612
rect 126992 480 127020 3606
rect 132960 3596 133012 3602
rect 132960 3538 133012 3544
rect 129372 3528 129424 3534
rect 129372 3470 129424 3476
rect 129384 480 129412 3470
rect 132972 480 133000 3538
rect 136456 3460 136508 3466
rect 136456 3402 136508 3408
rect 136468 480 136496 3402
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 2778 658144 2834 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3238 606056 3294 606112
rect 3422 579944 3478 580000
rect 3330 553832 3386 553888
rect 2778 527856 2834 527912
rect 2778 449520 2834 449576
rect 3146 410488 3202 410544
rect 2778 345344 2834 345400
rect 3330 293140 3386 293176
rect 3330 293120 3332 293140
rect 3332 293120 3384 293140
rect 3384 293120 3386 293140
rect 2778 254108 2834 254144
rect 2778 254088 2780 254108
rect 2780 254088 2832 254108
rect 2832 254088 2834 254108
rect 2778 241032 2834 241088
rect 3054 201864 3110 201920
rect 2962 188808 3018 188864
rect 3330 136740 3386 136776
rect 3330 136720 3332 136740
rect 3332 136720 3384 136740
rect 3384 136720 3386 136740
rect 3146 84632 3202 84688
rect 3330 58520 3386 58576
rect 2962 45464 3018 45520
rect 3514 501744 3570 501800
rect 3606 475632 3662 475688
rect 3698 397432 3754 397488
rect 3790 358400 3846 358456
rect 3882 306176 3938 306232
rect 3790 19352 3846 19408
rect 3974 149776 4030 149832
rect 4066 97552 4122 97608
rect 11886 34448 11942 34504
rect 13634 674192 13690 674248
rect 13542 620200 13598 620256
rect 13542 593408 13598 593464
rect 13542 566208 13598 566264
rect 13542 539416 13598 539472
rect 13542 512216 13598 512272
rect 13542 485424 13598 485480
rect 13542 458224 13598 458280
rect 13542 431432 13598 431488
rect 13542 404232 13598 404288
rect 13542 377440 13598 377496
rect 13542 350240 13598 350296
rect 13542 322904 13598 322960
rect 13542 296248 13598 296304
rect 13542 270000 13598 270056
rect 13542 242256 13598 242312
rect 13542 215328 13598 215384
rect 13542 188264 13598 188320
rect 13542 161336 13598 161392
rect 13542 134272 13598 134328
rect 13542 107344 13598 107400
rect 13542 80280 13598 80336
rect 13542 53352 13598 53408
rect 13450 33088 13506 33144
rect 12438 31048 12494 31104
rect 13726 647400 13782 647456
rect 17314 37848 17370 37904
rect 37278 673512 37334 673568
rect 37278 646720 37334 646776
rect 37278 619520 37334 619576
rect 37278 592728 37334 592784
rect 37278 565528 37334 565584
rect 37278 538736 37334 538792
rect 37278 511536 37334 511592
rect 37278 484744 37334 484800
rect 37278 457544 37334 457600
rect 37278 430752 37334 430808
rect 37278 403552 37334 403608
rect 37278 376760 37334 376816
rect 37278 349560 37334 349616
rect 37278 322768 37334 322824
rect 37278 295568 37334 295624
rect 37278 269048 37334 269104
rect 37278 241576 37334 241632
rect 37278 214648 37334 214704
rect 37278 187584 37334 187640
rect 37278 160656 37334 160712
rect 37278 133592 37334 133648
rect 37278 106664 37334 106720
rect 37278 79600 37334 79656
rect 37278 52672 37334 52728
rect 42706 674192 42762 674248
rect 42706 647400 42762 647456
rect 42706 620200 42762 620256
rect 42706 593408 42762 593464
rect 42706 566208 42762 566264
rect 42706 539416 42762 539472
rect 42706 512216 42762 512272
rect 42706 485424 42762 485480
rect 42706 458224 42762 458280
rect 42706 431432 42762 431488
rect 42706 404232 42762 404288
rect 42706 377440 42762 377496
rect 42706 350240 42762 350296
rect 42706 322904 42762 322960
rect 42706 296248 42762 296304
rect 42706 270000 42762 270056
rect 42706 242256 42762 242312
rect 42706 215328 42762 215384
rect 42706 188264 42762 188320
rect 42706 161336 42762 161392
rect 42706 134272 42762 134328
rect 42706 107344 42762 107400
rect 42706 80280 42762 80336
rect 42706 53352 42762 53408
rect 13726 29688 13782 29744
rect 13634 27648 13690 27704
rect 13542 26288 13598 26344
rect 13726 24112 13782 24168
rect 12438 22888 12494 22944
rect 12438 20848 12494 20904
rect 12622 19488 12678 19544
rect 12438 17448 12494 17504
rect 43442 35264 43498 35320
rect 61290 34312 61346 34368
rect 48042 16496 48098 16552
rect 19246 13232 19302 13288
rect 45006 13096 45062 13152
rect 59818 13504 59874 13560
rect 61106 13368 61162 13424
rect 63498 28328 63554 28384
rect 63498 26968 63554 27024
rect 63498 21392 63554 21448
rect 64234 35128 64290 35184
rect 64234 30232 64290 30288
rect 64142 23568 64198 23624
rect 64050 20168 64106 20224
rect 64510 31592 64566 31648
rect 64418 24928 64474 24984
rect 64326 18128 64382 18184
rect 64510 16768 64566 16824
rect 66258 673512 66314 673568
rect 70306 673784 70362 673840
rect 66258 646720 66314 646776
rect 70306 647400 70362 647456
rect 66258 619520 66314 619576
rect 70306 620200 70362 620256
rect 66258 592728 66314 592784
rect 70306 593408 70362 593464
rect 66258 565528 66314 565584
rect 70306 566208 70362 566264
rect 66258 538736 66314 538792
rect 70306 539416 70362 539472
rect 66258 511536 66314 511592
rect 70306 512216 70362 512272
rect 66258 484744 66314 484800
rect 70306 485424 70362 485480
rect 66258 457544 66314 457600
rect 70306 458224 70362 458280
rect 66258 430752 66314 430808
rect 70306 430888 70362 430944
rect 66258 403552 66314 403608
rect 70306 404232 70362 404288
rect 66258 376760 66314 376816
rect 70306 377984 70362 378040
rect 66258 349560 66314 349616
rect 70306 350240 70362 350296
rect 66258 322088 66314 322144
rect 70306 322904 70362 322960
rect 66258 295568 66314 295624
rect 70306 296248 70362 296304
rect 66258 269048 66314 269104
rect 70306 270000 70362 270056
rect 66258 241576 66314 241632
rect 70306 242256 70362 242312
rect 66258 214648 66314 214704
rect 70306 215872 70362 215928
rect 66258 187584 66314 187640
rect 70306 188264 70362 188320
rect 66258 160656 66314 160712
rect 70306 160792 70362 160848
rect 66258 133592 66314 133648
rect 70306 134272 70362 134328
rect 66258 106664 66314 106720
rect 70306 107344 70362 107400
rect 66258 79600 66314 79656
rect 70306 80280 70362 80336
rect 66258 52672 66314 52728
rect 70306 53352 70362 53408
rect 97906 674192 97962 674248
rect 93858 673512 93914 673568
rect 121458 673512 121514 673568
rect 126886 674192 126942 674248
rect 149058 673512 149114 673568
rect 97906 647400 97962 647456
rect 93858 646720 93914 646776
rect 121458 646720 121514 646776
rect 126886 647400 126942 647456
rect 149058 646720 149114 646776
rect 97906 620200 97962 620256
rect 93858 619520 93914 619576
rect 121458 619520 121514 619576
rect 126886 620200 126942 620256
rect 149058 619520 149114 619576
rect 97906 593408 97962 593464
rect 93858 592728 93914 592784
rect 121458 592728 121514 592784
rect 126886 593408 126942 593464
rect 149058 592728 149114 592784
rect 97906 566208 97962 566264
rect 93858 565528 93914 565584
rect 121458 565528 121514 565584
rect 126886 566208 126942 566264
rect 149058 565528 149114 565584
rect 97906 539416 97962 539472
rect 93858 538736 93914 538792
rect 121458 538736 121514 538792
rect 126886 539416 126942 539472
rect 149058 538736 149114 538792
rect 97906 512216 97962 512272
rect 93858 511536 93914 511592
rect 121458 511536 121514 511592
rect 126886 512216 126942 512272
rect 149058 511536 149114 511592
rect 97906 485424 97962 485480
rect 93858 484744 93914 484800
rect 121458 484744 121514 484800
rect 126886 485424 126942 485480
rect 149058 484744 149114 484800
rect 97906 458224 97962 458280
rect 93858 457544 93914 457600
rect 121458 457544 121514 457600
rect 126886 458224 126942 458280
rect 149058 457544 149114 457600
rect 97906 431432 97962 431488
rect 93858 430752 93914 430808
rect 121458 430752 121514 430808
rect 126886 431432 126942 431488
rect 149058 430752 149114 430808
rect 97906 404232 97962 404288
rect 93858 403552 93914 403608
rect 121458 403552 121514 403608
rect 126886 404232 126942 404288
rect 149058 403552 149114 403608
rect 97906 377440 97962 377496
rect 93858 376760 93914 376816
rect 121458 376760 121514 376816
rect 126886 377440 126942 377496
rect 149058 376760 149114 376816
rect 97906 350240 97962 350296
rect 93858 349560 93914 349616
rect 121458 349560 121514 349616
rect 126886 350240 126942 350296
rect 149058 349560 149114 349616
rect 97906 322904 97962 322960
rect 93858 322088 93914 322144
rect 121458 322088 121514 322144
rect 126886 322904 126942 322960
rect 149058 322088 149114 322144
rect 97906 296248 97962 296304
rect 93858 295568 93914 295624
rect 121458 295568 121514 295624
rect 126886 296248 126942 296304
rect 149058 295568 149114 295624
rect 97906 270000 97962 270056
rect 93858 269048 93914 269104
rect 121458 269048 121514 269104
rect 126886 270000 126942 270056
rect 149058 269048 149114 269104
rect 97906 242256 97962 242312
rect 93858 241576 93914 241632
rect 121458 241576 121514 241632
rect 126886 242256 126942 242312
rect 149058 241576 149114 241632
rect 97906 215328 97962 215384
rect 93858 214648 93914 214704
rect 121458 214648 121514 214704
rect 126886 215328 126942 215384
rect 149058 214648 149114 214704
rect 97906 188264 97962 188320
rect 93858 187584 93914 187640
rect 121458 187584 121514 187640
rect 126886 188264 126942 188320
rect 149058 187584 149114 187640
rect 97906 161336 97962 161392
rect 93858 160656 93914 160712
rect 121458 160656 121514 160712
rect 126886 161336 126942 161392
rect 149058 160656 149114 160712
rect 97906 134272 97962 134328
rect 93858 133592 93914 133648
rect 121458 133592 121514 133648
rect 126886 134272 126942 134328
rect 149058 133592 149114 133648
rect 97906 107344 97962 107400
rect 93858 106664 93914 106720
rect 121458 106664 121514 106720
rect 126886 107344 126942 107400
rect 149058 106664 149114 106720
rect 97906 80280 97962 80336
rect 93858 79600 93914 79656
rect 121458 79600 121514 79656
rect 126886 80280 126942 80336
rect 149058 79600 149114 79656
rect 97906 53352 97962 53408
rect 93858 52672 93914 52728
rect 121458 52672 121514 52728
rect 126886 53352 126942 53408
rect 149058 52672 149114 52728
rect 154486 674192 154542 674248
rect 178038 673512 178094 673568
rect 182086 674192 182142 674248
rect 156418 647944 156474 648000
rect 178038 646720 178094 646776
rect 184386 647944 184442 648000
rect 154486 620200 154542 620256
rect 178038 619520 178094 619576
rect 182086 620200 182142 620256
rect 154486 593408 154542 593464
rect 182086 593408 182142 593464
rect 178038 592728 178094 592784
rect 154486 566208 154542 566264
rect 178038 565528 178094 565584
rect 182086 566208 182142 566264
rect 154486 539416 154542 539472
rect 182086 539416 182142 539472
rect 178038 538736 178094 538792
rect 154486 512216 154542 512272
rect 178038 511536 178094 511592
rect 182086 512216 182142 512272
rect 154486 485424 154542 485480
rect 182086 485424 182142 485480
rect 178038 484744 178094 484800
rect 154486 458224 154542 458280
rect 178038 457544 178094 457600
rect 182086 458224 182142 458280
rect 154486 431432 154542 431488
rect 182086 431432 182142 431488
rect 178038 430752 178094 430808
rect 154486 404232 154542 404288
rect 178038 403552 178094 403608
rect 182086 404232 182142 404288
rect 154486 377440 154542 377496
rect 182086 377440 182142 377496
rect 178038 376760 178094 376816
rect 154486 350240 154542 350296
rect 178038 349560 178094 349616
rect 182086 350240 182142 350296
rect 154486 322904 154542 322960
rect 182086 322904 182142 322960
rect 178038 322088 178094 322144
rect 154486 296248 154542 296304
rect 178038 295568 178094 295624
rect 182086 296248 182142 296304
rect 154486 270000 154542 270056
rect 182086 270000 182142 270056
rect 178038 269048 178094 269104
rect 154486 242256 154542 242312
rect 178038 241576 178094 241632
rect 182086 242256 182142 242312
rect 154486 215328 154542 215384
rect 182086 215328 182142 215384
rect 178038 214648 178094 214704
rect 154486 188264 154542 188320
rect 178038 187584 178094 187640
rect 182086 188264 182142 188320
rect 154486 161336 154542 161392
rect 182086 161336 182142 161392
rect 178038 160656 178094 160712
rect 154486 134272 154542 134328
rect 178038 133592 178094 133648
rect 182086 134272 182142 134328
rect 154486 107344 154542 107400
rect 182086 107344 182142 107400
rect 178038 106664 178094 106720
rect 154486 80280 154542 80336
rect 178038 79600 178094 79656
rect 182086 80280 182142 80336
rect 154486 53352 154542 53408
rect 153842 42064 153898 42120
rect 182086 53352 182142 53408
rect 178038 52672 178094 52728
rect 209686 674192 209742 674248
rect 205638 674056 205694 674112
rect 233238 673512 233294 673568
rect 209686 647400 209742 647456
rect 205638 646720 205694 646776
rect 233238 646720 233294 646776
rect 209686 620200 209742 620256
rect 205638 619520 205694 619576
rect 233238 619520 233294 619576
rect 209686 593408 209742 593464
rect 205638 592728 205694 592784
rect 233238 592728 233294 592784
rect 209686 566208 209742 566264
rect 205638 565528 205694 565584
rect 233238 565528 233294 565584
rect 209686 539416 209742 539472
rect 205638 538736 205694 538792
rect 233238 538736 233294 538792
rect 209686 512216 209742 512272
rect 205638 511536 205694 511592
rect 233238 511536 233294 511592
rect 209686 485424 209742 485480
rect 205638 484744 205694 484800
rect 233238 484744 233294 484800
rect 209686 458224 209742 458280
rect 205638 457544 205694 457600
rect 233238 457544 233294 457600
rect 209686 431432 209742 431488
rect 205638 431296 205694 431352
rect 233238 430752 233294 430808
rect 209686 404232 209742 404288
rect 205638 403552 205694 403608
rect 233238 403552 233294 403608
rect 209686 377440 209742 377496
rect 205638 377304 205694 377360
rect 233238 376760 233294 376816
rect 209686 350240 209742 350296
rect 205638 349560 205694 349616
rect 233238 349560 233294 349616
rect 209686 323992 209742 324048
rect 205638 322088 205694 322144
rect 233238 322088 233294 322144
rect 209686 296248 209742 296304
rect 205638 295568 205694 295624
rect 233238 295568 233294 295624
rect 209686 269864 209742 269920
rect 205638 269048 205694 269104
rect 233238 269048 233294 269104
rect 209686 242256 209742 242312
rect 205638 241576 205694 241632
rect 233238 241576 233294 241632
rect 209686 215328 209742 215384
rect 205638 215192 205694 215248
rect 233238 214648 233294 214704
rect 209686 188264 209742 188320
rect 205638 187584 205694 187640
rect 233238 187584 233294 187640
rect 209686 161336 209742 161392
rect 205638 160112 205694 160168
rect 233238 160656 233294 160712
rect 209686 134272 209742 134328
rect 205638 133592 205694 133648
rect 233238 133592 233294 133648
rect 209686 107344 209742 107400
rect 205638 106664 205694 106720
rect 233238 106664 233294 106720
rect 209686 80280 209742 80336
rect 205638 79600 205694 79656
rect 233238 79600 233294 79656
rect 209686 53352 209742 53408
rect 205638 52672 205694 52728
rect 233238 52672 233294 52728
rect 70306 26832 70362 26888
rect 97906 26288 97962 26344
rect 93858 25608 93914 25664
rect 121458 25608 121514 25664
rect 126886 26288 126942 26344
rect 149058 25608 149114 25664
rect 154486 26288 154542 26344
rect 178038 25608 178094 25664
rect 182086 26288 182142 26344
rect 209686 26288 209742 26344
rect 205638 25880 205694 25936
rect 233238 25608 233294 25664
rect 238666 674192 238722 674248
rect 266266 674192 266322 674248
rect 262218 673512 262274 673568
rect 293866 674192 293922 674248
rect 289818 673512 289874 673568
rect 317418 673512 317474 673568
rect 238666 647400 238722 647456
rect 266266 647400 266322 647456
rect 262218 646720 262274 646776
rect 293866 647400 293922 647456
rect 289818 646720 289874 646776
rect 317418 646720 317474 646776
rect 238666 620200 238722 620256
rect 266266 620200 266322 620256
rect 262218 619520 262274 619576
rect 293866 620200 293922 620256
rect 289818 619520 289874 619576
rect 317418 619520 317474 619576
rect 238666 593408 238722 593464
rect 266266 593408 266322 593464
rect 262218 592728 262274 592784
rect 293866 593408 293922 593464
rect 289818 592728 289874 592784
rect 317418 592728 317474 592784
rect 238666 566208 238722 566264
rect 266266 566208 266322 566264
rect 262218 565528 262274 565584
rect 293866 566208 293922 566264
rect 289818 565528 289874 565584
rect 317418 565528 317474 565584
rect 238666 539416 238722 539472
rect 266266 539416 266322 539472
rect 262218 538736 262274 538792
rect 293866 539416 293922 539472
rect 289818 538736 289874 538792
rect 317418 538736 317474 538792
rect 238666 512216 238722 512272
rect 266266 512216 266322 512272
rect 262218 511536 262274 511592
rect 293866 512216 293922 512272
rect 289818 511536 289874 511592
rect 317418 511536 317474 511592
rect 238666 485424 238722 485480
rect 266266 485424 266322 485480
rect 262218 484744 262274 484800
rect 293866 485424 293922 485480
rect 289818 484744 289874 484800
rect 317418 484744 317474 484800
rect 238666 458224 238722 458280
rect 266266 458224 266322 458280
rect 262218 457544 262274 457600
rect 293866 458224 293922 458280
rect 289818 457544 289874 457600
rect 317418 457544 317474 457600
rect 238666 431432 238722 431488
rect 266266 431432 266322 431488
rect 262218 430752 262274 430808
rect 293866 431432 293922 431488
rect 289818 430752 289874 430808
rect 317418 430752 317474 430808
rect 238666 404232 238722 404288
rect 266266 404232 266322 404288
rect 262218 403552 262274 403608
rect 293866 404232 293922 404288
rect 289818 403552 289874 403608
rect 317418 403552 317474 403608
rect 238666 377440 238722 377496
rect 266266 377440 266322 377496
rect 262218 376760 262274 376816
rect 293866 377440 293922 377496
rect 289818 376760 289874 376816
rect 317418 376760 317474 376816
rect 238666 350240 238722 350296
rect 266266 350240 266322 350296
rect 262218 349560 262274 349616
rect 293866 350240 293922 350296
rect 289818 349560 289874 349616
rect 317418 349560 317474 349616
rect 238666 322904 238722 322960
rect 266266 322904 266322 322960
rect 262218 322768 262274 322824
rect 293866 323992 293922 324048
rect 289818 322088 289874 322144
rect 317418 322088 317474 322144
rect 238666 296248 238722 296304
rect 266266 296248 266322 296304
rect 262218 295568 262274 295624
rect 293866 296248 293922 296304
rect 289818 295568 289874 295624
rect 317418 295568 317474 295624
rect 238666 269864 238722 269920
rect 266266 269864 266322 269920
rect 262218 269048 262274 269104
rect 293866 270000 293922 270056
rect 289818 269048 289874 269104
rect 317418 269048 317474 269104
rect 238666 242256 238722 242312
rect 266266 242256 266322 242312
rect 262218 241576 262274 241632
rect 293866 242256 293922 242312
rect 289818 241576 289874 241632
rect 317418 241576 317474 241632
rect 238666 215328 238722 215384
rect 266266 215328 266322 215384
rect 262218 214648 262274 214704
rect 293866 215328 293922 215384
rect 289818 214648 289874 214704
rect 317418 214648 317474 214704
rect 238666 188264 238722 188320
rect 266266 188264 266322 188320
rect 262218 187584 262274 187640
rect 293866 188264 293922 188320
rect 289818 187584 289874 187640
rect 317418 187584 317474 187640
rect 238666 161336 238722 161392
rect 266266 161336 266322 161392
rect 262218 160656 262274 160712
rect 293866 161336 293922 161392
rect 289818 160656 289874 160712
rect 317418 160656 317474 160712
rect 238666 134272 238722 134328
rect 266266 134272 266322 134328
rect 262218 133592 262274 133648
rect 293866 134272 293922 134328
rect 289818 133592 289874 133648
rect 317418 133592 317474 133648
rect 238666 107344 238722 107400
rect 266266 107344 266322 107400
rect 262218 106664 262274 106720
rect 293866 107344 293922 107400
rect 289818 106664 289874 106720
rect 317418 106664 317474 106720
rect 238666 80280 238722 80336
rect 266266 80280 266322 80336
rect 262218 79600 262274 79656
rect 293866 80280 293922 80336
rect 289818 79600 289874 79656
rect 317418 79600 317474 79656
rect 238666 53352 238722 53408
rect 266266 53352 266322 53408
rect 262218 52672 262274 52728
rect 293866 53352 293922 53408
rect 289818 52672 289874 52728
rect 317418 52672 317474 52728
rect 322846 674192 322902 674248
rect 345018 673512 345074 673568
rect 350446 674192 350502 674248
rect 373998 673512 374054 673568
rect 378046 674192 378102 674248
rect 322846 647400 322902 647456
rect 345018 646720 345074 646776
rect 350446 647400 350502 647456
rect 378046 647400 378102 647456
rect 373998 646720 374054 646776
rect 322846 620200 322902 620256
rect 345018 619520 345074 619576
rect 350446 620200 350502 620256
rect 373998 619520 374054 619576
rect 378046 620200 378102 620256
rect 322846 593408 322902 593464
rect 345018 592728 345074 592784
rect 350446 593408 350502 593464
rect 378046 593408 378102 593464
rect 373998 592728 374054 592784
rect 322846 566208 322902 566264
rect 345018 565528 345074 565584
rect 350446 566208 350502 566264
rect 373998 565528 374054 565584
rect 378046 566208 378102 566264
rect 322846 539416 322902 539472
rect 345018 538736 345074 538792
rect 350446 539416 350502 539472
rect 378046 539416 378102 539472
rect 373998 538736 374054 538792
rect 322846 512216 322902 512272
rect 345018 511536 345074 511592
rect 350446 512216 350502 512272
rect 373998 511536 374054 511592
rect 378046 512216 378102 512272
rect 322846 485424 322902 485480
rect 345018 484744 345074 484800
rect 350446 485424 350502 485480
rect 378046 485424 378102 485480
rect 373998 484744 374054 484800
rect 322846 458224 322902 458280
rect 345018 457544 345074 457600
rect 350446 458224 350502 458280
rect 373998 457544 374054 457600
rect 378046 458224 378102 458280
rect 322846 431432 322902 431488
rect 345018 430752 345074 430808
rect 350446 431432 350502 431488
rect 378046 431432 378102 431488
rect 373998 430752 374054 430808
rect 322846 404232 322902 404288
rect 345018 403552 345074 403608
rect 350446 404232 350502 404288
rect 373998 403552 374054 403608
rect 378046 404232 378102 404288
rect 322846 377440 322902 377496
rect 345018 376760 345074 376816
rect 350446 377440 350502 377496
rect 378046 377440 378102 377496
rect 373998 377304 374054 377360
rect 322846 350240 322902 350296
rect 345018 349560 345074 349616
rect 350446 350240 350502 350296
rect 373998 349560 374054 349616
rect 378046 350240 378102 350296
rect 322846 322904 322902 322960
rect 345018 322768 345074 322824
rect 350446 322904 350502 322960
rect 378046 322904 378102 322960
rect 373998 322088 374054 322144
rect 322846 296248 322902 296304
rect 345018 295568 345074 295624
rect 350446 296248 350502 296304
rect 373998 295568 374054 295624
rect 378046 296248 378102 296304
rect 322846 270000 322902 270056
rect 345018 269048 345074 269104
rect 350446 270000 350502 270056
rect 378046 270000 378102 270056
rect 373998 269048 374054 269104
rect 322846 242256 322902 242312
rect 345018 241576 345074 241632
rect 350446 242256 350502 242312
rect 373998 241576 374054 241632
rect 378046 242256 378102 242312
rect 322846 215328 322902 215384
rect 345018 214648 345074 214704
rect 350446 215328 350502 215384
rect 378046 215328 378102 215384
rect 373998 215192 374054 215248
rect 322846 188264 322902 188320
rect 345018 187584 345074 187640
rect 350446 188264 350502 188320
rect 373998 187584 374054 187640
rect 378046 188264 378102 188320
rect 322846 161336 322902 161392
rect 345018 160656 345074 160712
rect 350446 161336 350502 161392
rect 378046 161336 378102 161392
rect 373998 160656 374054 160712
rect 322846 134272 322902 134328
rect 345018 133592 345074 133648
rect 350446 134272 350502 134328
rect 373998 133592 374054 133648
rect 378046 134272 378102 134328
rect 322846 107344 322902 107400
rect 345018 106664 345074 106720
rect 350446 107344 350502 107400
rect 378046 107344 378102 107400
rect 373998 106664 374054 106720
rect 322846 80280 322902 80336
rect 345018 79600 345074 79656
rect 350446 80280 350502 80336
rect 373998 79600 374054 79656
rect 378046 80280 378102 80336
rect 322846 53352 322902 53408
rect 345018 52672 345074 52728
rect 350446 53352 350502 53408
rect 378046 53352 378102 53408
rect 373998 52672 374054 52728
rect 238666 26288 238722 26344
rect 266266 26288 266322 26344
rect 262218 25608 262274 25664
rect 293866 26288 293922 26344
rect 289818 25608 289874 25664
rect 317418 25608 317474 25664
rect 322846 26288 322902 26344
rect 345018 25608 345074 25664
rect 350446 26288 350502 26344
rect 373998 25608 374054 25664
rect 378046 26288 378102 26344
rect 405646 674192 405702 674248
rect 401598 673512 401654 673568
rect 408406 647944 408462 648000
rect 401598 646720 401654 646776
rect 405646 620200 405702 620256
rect 401598 619520 401654 619576
rect 405646 593408 405702 593464
rect 401598 592728 401654 592784
rect 405646 566208 405702 566264
rect 401598 565528 401654 565584
rect 405646 539416 405702 539472
rect 401598 538736 401654 538792
rect 405646 512216 405702 512272
rect 401598 511536 401654 511592
rect 405646 485424 405702 485480
rect 401598 484744 401654 484800
rect 405646 458224 405702 458280
rect 401598 457544 401654 457600
rect 405646 431432 405702 431488
rect 401598 430752 401654 430808
rect 405646 404232 405702 404288
rect 401598 403552 401654 403608
rect 405646 377440 405702 377496
rect 401598 376760 401654 376816
rect 405646 350240 405702 350296
rect 401598 349560 401654 349616
rect 405646 323992 405702 324048
rect 401598 322088 401654 322144
rect 405646 296248 405702 296304
rect 401598 295568 401654 295624
rect 405646 270000 405702 270056
rect 401598 269048 401654 269104
rect 405646 242256 405702 242312
rect 401598 241576 401654 241632
rect 405646 215328 405702 215384
rect 401598 214648 401654 214704
rect 405646 188264 405702 188320
rect 401598 187584 401654 187640
rect 405646 161336 405702 161392
rect 401598 160656 401654 160712
rect 405646 134272 405702 134328
rect 401598 133592 401654 133648
rect 405646 107344 405702 107400
rect 401598 106664 401654 106720
rect 405646 80280 405702 80336
rect 401598 79600 401654 79656
rect 405646 53352 405702 53408
rect 401598 52672 401654 52728
rect 405646 26288 405702 26344
rect 401598 25608 401654 25664
rect 434626 674192 434682 674248
rect 429290 673512 429346 673568
rect 462226 674192 462282 674248
rect 458178 673512 458234 673568
rect 429290 646720 429346 646776
rect 434626 647400 434682 647456
rect 458178 646720 458234 646776
rect 434626 620200 434682 620256
rect 429290 619520 429346 619576
rect 462226 620200 462282 620256
rect 458178 619520 458234 619576
rect 429290 592728 429346 592784
rect 434626 593408 434682 593464
rect 462226 593408 462282 593464
rect 458178 592728 458234 592784
rect 434626 566208 434682 566264
rect 429290 565528 429346 565584
rect 462226 566208 462282 566264
rect 458178 565528 458234 565584
rect 429290 538736 429346 538792
rect 434626 539416 434682 539472
rect 462226 539416 462282 539472
rect 458178 538736 458234 538792
rect 434626 512216 434682 512272
rect 429290 511536 429346 511592
rect 462226 512216 462282 512272
rect 458178 511536 458234 511592
rect 429290 484744 429346 484800
rect 434626 485424 434682 485480
rect 462226 485424 462282 485480
rect 458178 484744 458234 484800
rect 434626 458224 434682 458280
rect 429290 457544 429346 457600
rect 462226 458224 462282 458280
rect 458178 457544 458234 457600
rect 429290 430752 429346 430808
rect 434626 431432 434682 431488
rect 462226 431432 462282 431488
rect 458178 430752 458234 430808
rect 434626 404232 434682 404288
rect 429290 403552 429346 403608
rect 462226 404232 462282 404288
rect 458178 403552 458234 403608
rect 429290 376760 429346 376816
rect 434626 377440 434682 377496
rect 462226 377440 462282 377496
rect 458178 376760 458234 376816
rect 434626 350240 434682 350296
rect 429290 349560 429346 349616
rect 462226 350240 462282 350296
rect 458178 349560 458234 349616
rect 429290 322088 429346 322144
rect 434626 322904 434682 322960
rect 462226 322904 462282 322960
rect 458178 322768 458234 322824
rect 434626 296248 434682 296304
rect 429290 295568 429346 295624
rect 462226 296248 462282 296304
rect 458178 295568 458234 295624
rect 429290 269048 429346 269104
rect 434626 270000 434682 270056
rect 462226 270000 462282 270056
rect 458178 269048 458234 269104
rect 434626 242256 434682 242312
rect 429290 241576 429346 241632
rect 462226 242256 462282 242312
rect 458178 241576 458234 241632
rect 429290 214648 429346 214704
rect 434626 215328 434682 215384
rect 462226 215328 462282 215384
rect 458178 214648 458234 214704
rect 434626 188264 434682 188320
rect 429290 187584 429346 187640
rect 462226 188264 462282 188320
rect 458178 187584 458234 187640
rect 429290 160656 429346 160712
rect 434626 161336 434682 161392
rect 462226 161336 462282 161392
rect 458178 160656 458234 160712
rect 434626 134272 434682 134328
rect 429290 133592 429346 133648
rect 462226 134272 462282 134328
rect 458178 133592 458234 133648
rect 429290 106664 429346 106720
rect 434626 107344 434682 107400
rect 462226 107344 462282 107400
rect 458178 106664 458234 106720
rect 434626 80280 434682 80336
rect 429290 79600 429346 79656
rect 462226 80280 462282 80336
rect 458178 79600 458234 79656
rect 429290 52672 429346 52728
rect 434626 53352 434682 53408
rect 462226 53352 462282 53408
rect 458178 52672 458234 52728
rect 489826 674192 489882 674248
rect 485778 673512 485834 673568
rect 513378 673512 513434 673568
rect 464434 647944 464490 648000
rect 489826 647400 489882 647456
rect 485778 646720 485834 646776
rect 513378 646720 513434 646776
rect 489826 620200 489882 620256
rect 485778 619520 485834 619576
rect 513378 619520 513434 619576
rect 489826 593408 489882 593464
rect 485778 592728 485834 592784
rect 513378 592728 513434 592784
rect 489826 566208 489882 566264
rect 485778 565528 485834 565584
rect 513378 565528 513434 565584
rect 489826 539416 489882 539472
rect 485778 538736 485834 538792
rect 513378 538736 513434 538792
rect 489826 512216 489882 512272
rect 485778 511536 485834 511592
rect 513378 511536 513434 511592
rect 489826 485424 489882 485480
rect 485778 484744 485834 484800
rect 513378 484744 513434 484800
rect 489826 458224 489882 458280
rect 485778 457544 485834 457600
rect 513378 457544 513434 457600
rect 489826 431432 489882 431488
rect 485778 430752 485834 430808
rect 513378 430752 513434 430808
rect 489826 404232 489882 404288
rect 485778 403552 485834 403608
rect 513378 403552 513434 403608
rect 489826 377440 489882 377496
rect 485778 376760 485834 376816
rect 513378 376760 513434 376816
rect 489826 350240 489882 350296
rect 485778 349560 485834 349616
rect 513378 349560 513434 349616
rect 489826 323992 489882 324048
rect 485778 322088 485834 322144
rect 513378 322088 513434 322144
rect 489826 296248 489882 296304
rect 485778 295568 485834 295624
rect 513378 295568 513434 295624
rect 489826 269864 489882 269920
rect 485778 269048 485834 269104
rect 513378 269048 513434 269104
rect 489826 242256 489882 242312
rect 485778 241576 485834 241632
rect 513378 241576 513434 241632
rect 489826 215328 489882 215384
rect 485778 214648 485834 214704
rect 513378 214648 513434 214704
rect 489826 188264 489882 188320
rect 485778 187584 485834 187640
rect 513378 187584 513434 187640
rect 489826 161336 489882 161392
rect 485778 160656 485834 160712
rect 513378 160656 513434 160712
rect 489826 134272 489882 134328
rect 485778 133592 485834 133648
rect 513378 133592 513434 133648
rect 489826 107344 489882 107400
rect 485778 106664 485834 106720
rect 513378 106664 513434 106720
rect 489826 80280 489882 80336
rect 485778 79600 485834 79656
rect 513378 79600 513434 79656
rect 489826 53352 489882 53408
rect 485778 52672 485834 52728
rect 513378 52672 513434 52728
rect 429290 25608 429346 25664
rect 434626 26288 434682 26344
rect 462226 26288 462282 26344
rect 458178 25608 458234 25664
rect 489826 26288 489882 26344
rect 485778 25608 485834 25664
rect 513378 25608 513434 25664
rect 580170 697176 580226 697232
rect 518806 674192 518862 674248
rect 545118 674192 545174 674248
rect 542358 673512 542414 673568
rect 518806 647400 518862 647456
rect 542358 646720 542414 646776
rect 518806 620200 518862 620256
rect 542358 619520 542414 619576
rect 518806 593408 518862 593464
rect 542358 592728 542414 592784
rect 518806 566208 518862 566264
rect 542358 565528 542414 565584
rect 518806 539416 518862 539472
rect 542358 538736 542414 538792
rect 518806 512216 518862 512272
rect 542358 511536 542414 511592
rect 518806 485424 518862 485480
rect 542358 484744 542414 484800
rect 518806 458224 518862 458280
rect 542358 457544 542414 457600
rect 518806 431432 518862 431488
rect 542358 430752 542414 430808
rect 518806 404232 518862 404288
rect 542358 403552 542414 403608
rect 518806 377440 518862 377496
rect 542358 376760 542414 376816
rect 518806 350240 518862 350296
rect 542358 349560 542414 349616
rect 518806 322904 518862 322960
rect 542358 322768 542414 322824
rect 518806 296248 518862 296304
rect 542358 295568 542414 295624
rect 518806 269864 518862 269920
rect 542358 269048 542414 269104
rect 518806 242256 518862 242312
rect 542358 241576 542414 241632
rect 518806 215328 518862 215384
rect 542358 214648 542414 214704
rect 518806 188264 518862 188320
rect 542358 187584 542414 187640
rect 518806 161336 518862 161392
rect 542358 160656 542414 160712
rect 518806 134272 518862 134328
rect 542358 133592 542414 133648
rect 518806 107344 518862 107400
rect 542358 106664 542414 106720
rect 518806 80280 518862 80336
rect 542358 79600 542414 79656
rect 518806 53352 518862 53408
rect 542358 52672 542414 52728
rect 569958 673512 570014 673568
rect 546406 647400 546462 647456
rect 546406 620200 546462 620256
rect 569958 646720 570014 646776
rect 569958 619520 570014 619576
rect 546406 593408 546462 593464
rect 546406 566208 546462 566264
rect 569958 592728 570014 592784
rect 580262 590960 580318 591016
rect 569958 565528 570014 565584
rect 546406 539416 546462 539472
rect 546406 512216 546462 512272
rect 569958 538736 570014 538792
rect 569958 511536 570014 511592
rect 546406 485424 546462 485480
rect 546406 458224 546462 458280
rect 569958 484744 570014 484800
rect 579986 471416 580042 471472
rect 569958 457544 570014 457600
rect 546406 431432 546462 431488
rect 546406 404232 546462 404288
rect 569958 430752 570014 430808
rect 569958 403552 570014 403608
rect 546406 377032 546462 377088
rect 546406 350240 546462 350296
rect 580170 378392 580226 378448
rect 569958 376760 570014 376816
rect 569958 349560 570014 349616
rect 546406 322904 546462 322960
rect 546406 296248 546462 296304
rect 579986 325216 580042 325272
rect 569958 322088 570014 322144
rect 569958 295568 570014 295624
rect 546406 269184 546462 269240
rect 546406 242256 546462 242312
rect 569958 269048 570014 269104
rect 569958 241576 570014 241632
rect 546406 215464 546462 215520
rect 546406 188264 546462 188320
rect 569958 214648 570014 214704
rect 569958 187584 570014 187640
rect 546406 161336 546462 161392
rect 546406 134272 546462 134328
rect 546406 107344 546462 107400
rect 546406 80280 546462 80336
rect 546406 53352 546462 53408
rect 518806 26288 518862 26344
rect 546406 26288 546462 26344
rect 542358 25608 542414 25664
rect 569958 160656 570014 160712
rect 569958 133592 570014 133648
rect 569958 106664 570014 106720
rect 569958 79600 570014 79656
rect 569958 52672 570014 52728
rect 569958 25608 570014 25664
rect 578882 272176 578938 272232
rect 518162 13232 518218 13288
rect 579802 232328 579858 232384
rect 580170 192480 580226 192536
rect 580170 112784 580226 112840
rect 580078 72936 580134 72992
rect 579986 33088 580042 33144
rect 580354 537784 580410 537840
rect 580446 511264 580502 511320
rect 580538 484608 580594 484664
rect 580630 431568 580686 431624
rect 580722 404912 580778 404968
rect 580814 351872 580870 351928
rect 580906 152632 580962 152688
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 583520 683756 584960 683996
rect 13629 674250 13695 674253
rect 42701 674250 42767 674253
rect 97901 674250 97967 674253
rect 126881 674250 126947 674253
rect 154481 674250 154547 674253
rect 182081 674250 182147 674253
rect 209681 674250 209747 674253
rect 238661 674250 238727 674253
rect 266261 674250 266327 674253
rect 293861 674250 293927 674253
rect 322841 674250 322907 674253
rect 350441 674250 350507 674253
rect 378041 674250 378107 674253
rect 405641 674250 405707 674253
rect 434621 674250 434687 674253
rect 462221 674250 462287 674253
rect 489821 674250 489887 674253
rect 518801 674250 518867 674253
rect 545113 674250 545179 674253
rect 13629 674248 16100 674250
rect 13629 674192 13634 674248
rect 13690 674192 16100 674248
rect 13629 674190 16100 674192
rect 42701 674248 44068 674250
rect 42701 674192 42706 674248
rect 42762 674192 44068 674248
rect 97901 674248 100188 674250
rect 42701 674190 44068 674192
rect 13629 674187 13695 674190
rect 42701 674187 42767 674190
rect 70301 673842 70367 673845
rect 72006 673842 72066 674220
rect 97901 674192 97906 674248
rect 97962 674192 100188 674248
rect 97901 674190 100188 674192
rect 126881 674248 128156 674250
rect 126881 674192 126886 674248
rect 126942 674192 128156 674248
rect 126881 674190 128156 674192
rect 154481 674248 156124 674250
rect 154481 674192 154486 674248
rect 154542 674192 156124 674248
rect 154481 674190 156124 674192
rect 182081 674248 184092 674250
rect 182081 674192 182086 674248
rect 182142 674192 184092 674248
rect 182081 674190 184092 674192
rect 209681 674248 212060 674250
rect 209681 674192 209686 674248
rect 209742 674192 212060 674248
rect 209681 674190 212060 674192
rect 238661 674248 240212 674250
rect 238661 674192 238666 674248
rect 238722 674192 240212 674248
rect 238661 674190 240212 674192
rect 266261 674248 268180 674250
rect 266261 674192 266266 674248
rect 266322 674192 268180 674248
rect 266261 674190 268180 674192
rect 293861 674248 296148 674250
rect 293861 674192 293866 674248
rect 293922 674192 296148 674248
rect 293861 674190 296148 674192
rect 322841 674248 324116 674250
rect 322841 674192 322846 674248
rect 322902 674192 324116 674248
rect 322841 674190 324116 674192
rect 350441 674248 352084 674250
rect 350441 674192 350446 674248
rect 350502 674192 352084 674248
rect 350441 674190 352084 674192
rect 378041 674248 380052 674250
rect 378041 674192 378046 674248
rect 378102 674192 380052 674248
rect 378041 674190 380052 674192
rect 405641 674248 408204 674250
rect 405641 674192 405646 674248
rect 405702 674192 408204 674248
rect 405641 674190 408204 674192
rect 434621 674248 436172 674250
rect 434621 674192 434626 674248
rect 434682 674192 436172 674248
rect 434621 674190 436172 674192
rect 462221 674248 464140 674250
rect 462221 674192 462226 674248
rect 462282 674192 464140 674248
rect 462221 674190 464140 674192
rect 489821 674248 492108 674250
rect 489821 674192 489826 674248
rect 489882 674192 492108 674248
rect 489821 674190 492108 674192
rect 518801 674248 520076 674250
rect 518801 674192 518806 674248
rect 518862 674192 520076 674248
rect 518801 674190 520076 674192
rect 545113 674248 548044 674250
rect 545113 674192 545118 674248
rect 545174 674192 548044 674248
rect 545113 674190 548044 674192
rect 97901 674187 97967 674190
rect 126881 674187 126947 674190
rect 154481 674187 154547 674190
rect 182081 674187 182147 674190
rect 209681 674187 209747 674190
rect 238661 674187 238727 674190
rect 266261 674187 266327 674190
rect 293861 674187 293927 674190
rect 322841 674187 322907 674190
rect 350441 674187 350507 674190
rect 378041 674187 378107 674190
rect 405641 674187 405707 674190
rect 434621 674187 434687 674190
rect 462221 674187 462287 674190
rect 489821 674187 489887 674190
rect 518801 674187 518867 674190
rect 545113 674187 545179 674190
rect 205633 674114 205699 674117
rect 70301 673840 72066 673842
rect 70301 673784 70306 673840
rect 70362 673784 72066 673840
rect 70301 673782 72066 673784
rect 203934 674112 205699 674114
rect 203934 674056 205638 674112
rect 205694 674056 205699 674112
rect 203934 674054 205699 674056
rect 70301 673779 70367 673782
rect 37273 673570 37339 673573
rect 66253 673570 66319 673573
rect 93853 673570 93919 673573
rect 121453 673570 121519 673573
rect 149053 673570 149119 673573
rect 178033 673570 178099 673573
rect 35788 673568 37339 673570
rect 35788 673512 37278 673568
rect 37334 673512 37339 673568
rect 35788 673510 37339 673512
rect 63940 673568 66319 673570
rect 63940 673512 66258 673568
rect 66314 673512 66319 673568
rect 63940 673510 66319 673512
rect 91908 673568 93919 673570
rect 91908 673512 93858 673568
rect 93914 673512 93919 673568
rect 91908 673510 93919 673512
rect 119876 673568 121519 673570
rect 119876 673512 121458 673568
rect 121514 673512 121519 673568
rect 119876 673510 121519 673512
rect 147844 673568 149119 673570
rect 147844 673512 149058 673568
rect 149114 673512 149119 673568
rect 147844 673510 149119 673512
rect 175812 673568 178099 673570
rect 175812 673512 178038 673568
rect 178094 673512 178099 673568
rect 203934 673540 203994 674054
rect 205633 674051 205699 674054
rect 233233 673570 233299 673573
rect 262213 673570 262279 673573
rect 289813 673570 289879 673573
rect 317413 673570 317479 673573
rect 345013 673570 345079 673573
rect 373993 673570 374059 673573
rect 401593 673570 401659 673573
rect 429285 673570 429351 673573
rect 458173 673570 458239 673573
rect 485773 673570 485839 673573
rect 513373 673570 513439 673573
rect 542353 673570 542419 673573
rect 569953 673570 570019 673573
rect 231932 673568 233299 673570
rect 175812 673510 178099 673512
rect 231932 673512 233238 673568
rect 233294 673512 233299 673568
rect 231932 673510 233299 673512
rect 259900 673568 262279 673570
rect 259900 673512 262218 673568
rect 262274 673512 262279 673568
rect 259900 673510 262279 673512
rect 287868 673568 289879 673570
rect 287868 673512 289818 673568
rect 289874 673512 289879 673568
rect 287868 673510 289879 673512
rect 315836 673568 317479 673570
rect 315836 673512 317418 673568
rect 317474 673512 317479 673568
rect 315836 673510 317479 673512
rect 343804 673568 345079 673570
rect 343804 673512 345018 673568
rect 345074 673512 345079 673568
rect 343804 673510 345079 673512
rect 371956 673568 374059 673570
rect 371956 673512 373998 673568
rect 374054 673512 374059 673568
rect 371956 673510 374059 673512
rect 399924 673568 401659 673570
rect 399924 673512 401598 673568
rect 401654 673512 401659 673568
rect 399924 673510 401659 673512
rect 427892 673568 429351 673570
rect 427892 673512 429290 673568
rect 429346 673512 429351 673568
rect 427892 673510 429351 673512
rect 455860 673568 458239 673570
rect 455860 673512 458178 673568
rect 458234 673512 458239 673568
rect 455860 673510 458239 673512
rect 483828 673568 485839 673570
rect 483828 673512 485778 673568
rect 485834 673512 485839 673568
rect 483828 673510 485839 673512
rect 511796 673568 513439 673570
rect 511796 673512 513378 673568
rect 513434 673512 513439 673568
rect 511796 673510 513439 673512
rect 539948 673568 542419 673570
rect 539948 673512 542358 673568
rect 542414 673512 542419 673568
rect 539948 673510 542419 673512
rect 567916 673568 570019 673570
rect 567916 673512 569958 673568
rect 570014 673512 570019 673568
rect 567916 673510 570019 673512
rect 37273 673507 37339 673510
rect 66253 673507 66319 673510
rect 93853 673507 93919 673510
rect 121453 673507 121519 673510
rect 149053 673507 149119 673510
rect 178033 673507 178099 673510
rect 233233 673507 233299 673510
rect 262213 673507 262279 673510
rect 289813 673507 289879 673510
rect 317413 673507 317479 673510
rect 345013 673507 345079 673510
rect 373993 673507 374059 673510
rect 401593 673507 401659 673510
rect 429285 673507 429351 673510
rect 458173 673507 458239 673510
rect 485773 673507 485839 673510
rect 513373 673507 513439 673510
rect 542353 673507 542419 673510
rect 569953 673507 570019 673510
rect -960 671108 480 671348
rect 580206 670652 580212 670716
rect 580276 670714 580282 670716
rect 583520 670714 584960 670804
rect 580276 670654 584960 670714
rect 580276 670652 580282 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 2773 658202 2839 658205
rect -960 658200 2839 658202
rect -960 658144 2778 658200
rect 2834 658144 2839 658200
rect -960 658142 2839 658144
rect -960 658052 480 658142
rect 2773 658139 2839 658142
rect 583520 657236 584960 657476
rect 156413 648002 156479 648005
rect 184381 648002 184447 648005
rect 408401 648002 408467 648005
rect 156413 648000 156522 648002
rect 156413 647944 156418 648000
rect 156474 647944 156522 648000
rect 156413 647939 156522 647944
rect 184381 648000 184490 648002
rect 184381 647944 184386 648000
rect 184442 647944 184490 648000
rect 184381 647939 184490 647944
rect 13721 647458 13787 647461
rect 42701 647458 42767 647461
rect 70301 647458 70367 647461
rect 97901 647458 97967 647461
rect 126881 647458 126947 647461
rect 13721 647456 16100 647458
rect 13721 647400 13726 647456
rect 13782 647400 16100 647456
rect 13721 647398 16100 647400
rect 42701 647456 44068 647458
rect 42701 647400 42706 647456
rect 42762 647400 44068 647456
rect 42701 647398 44068 647400
rect 70301 647456 72036 647458
rect 70301 647400 70306 647456
rect 70362 647400 72036 647456
rect 70301 647398 72036 647400
rect 97901 647456 100188 647458
rect 97901 647400 97906 647456
rect 97962 647400 100188 647456
rect 97901 647398 100188 647400
rect 126881 647456 128156 647458
rect 126881 647400 126886 647456
rect 126942 647400 128156 647456
rect 156462 647428 156522 647939
rect 184430 647428 184490 647939
rect 408358 648000 408467 648002
rect 408358 647944 408406 648000
rect 408462 647944 408467 648000
rect 408358 647939 408467 647944
rect 464429 648002 464495 648005
rect 464429 648000 464538 648002
rect 464429 647944 464434 648000
rect 464490 647944 464538 648000
rect 464429 647939 464538 647944
rect 209681 647458 209747 647461
rect 238661 647458 238727 647461
rect 266261 647458 266327 647461
rect 293861 647458 293927 647461
rect 322841 647458 322907 647461
rect 350441 647458 350507 647461
rect 378041 647458 378107 647461
rect 209681 647456 212060 647458
rect 126881 647398 128156 647400
rect 209681 647400 209686 647456
rect 209742 647400 212060 647456
rect 209681 647398 212060 647400
rect 238661 647456 240212 647458
rect 238661 647400 238666 647456
rect 238722 647400 240212 647456
rect 238661 647398 240212 647400
rect 266261 647456 268180 647458
rect 266261 647400 266266 647456
rect 266322 647400 268180 647456
rect 266261 647398 268180 647400
rect 293861 647456 296148 647458
rect 293861 647400 293866 647456
rect 293922 647400 296148 647456
rect 293861 647398 296148 647400
rect 322841 647456 324116 647458
rect 322841 647400 322846 647456
rect 322902 647400 324116 647456
rect 322841 647398 324116 647400
rect 350441 647456 352084 647458
rect 350441 647400 350446 647456
rect 350502 647400 352084 647456
rect 350441 647398 352084 647400
rect 378041 647456 380052 647458
rect 378041 647400 378046 647456
rect 378102 647400 380052 647456
rect 408358 647428 408418 647939
rect 434621 647458 434687 647461
rect 434621 647456 436172 647458
rect 378041 647398 380052 647400
rect 434621 647400 434626 647456
rect 434682 647400 436172 647456
rect 464478 647428 464538 647939
rect 489821 647458 489887 647461
rect 518801 647458 518867 647461
rect 546401 647458 546467 647461
rect 489821 647456 492108 647458
rect 434621 647398 436172 647400
rect 489821 647400 489826 647456
rect 489882 647400 492108 647456
rect 489821 647398 492108 647400
rect 518801 647456 520076 647458
rect 518801 647400 518806 647456
rect 518862 647400 520076 647456
rect 518801 647398 520076 647400
rect 546401 647456 548044 647458
rect 546401 647400 546406 647456
rect 546462 647400 548044 647456
rect 546401 647398 548044 647400
rect 13721 647395 13787 647398
rect 42701 647395 42767 647398
rect 70301 647395 70367 647398
rect 97901 647395 97967 647398
rect 126881 647395 126947 647398
rect 209681 647395 209747 647398
rect 238661 647395 238727 647398
rect 266261 647395 266327 647398
rect 293861 647395 293927 647398
rect 322841 647395 322907 647398
rect 350441 647395 350507 647398
rect 378041 647395 378107 647398
rect 434621 647395 434687 647398
rect 489821 647395 489887 647398
rect 518801 647395 518867 647398
rect 546401 647395 546467 647398
rect 37273 646778 37339 646781
rect 66253 646778 66319 646781
rect 93853 646778 93919 646781
rect 121453 646778 121519 646781
rect 149053 646778 149119 646781
rect 178033 646778 178099 646781
rect 205633 646778 205699 646781
rect 233233 646778 233299 646781
rect 262213 646778 262279 646781
rect 289813 646778 289879 646781
rect 317413 646778 317479 646781
rect 345013 646778 345079 646781
rect 373993 646778 374059 646781
rect 401593 646778 401659 646781
rect 429285 646778 429351 646781
rect 458173 646778 458239 646781
rect 485773 646778 485839 646781
rect 513373 646778 513439 646781
rect 542353 646778 542419 646781
rect 569953 646778 570019 646781
rect 35788 646776 37339 646778
rect 35788 646720 37278 646776
rect 37334 646720 37339 646776
rect 35788 646718 37339 646720
rect 63940 646776 66319 646778
rect 63940 646720 66258 646776
rect 66314 646720 66319 646776
rect 63940 646718 66319 646720
rect 91908 646776 93919 646778
rect 91908 646720 93858 646776
rect 93914 646720 93919 646776
rect 91908 646718 93919 646720
rect 119876 646776 121519 646778
rect 119876 646720 121458 646776
rect 121514 646720 121519 646776
rect 119876 646718 121519 646720
rect 147844 646776 149119 646778
rect 147844 646720 149058 646776
rect 149114 646720 149119 646776
rect 147844 646718 149119 646720
rect 175812 646776 178099 646778
rect 175812 646720 178038 646776
rect 178094 646720 178099 646776
rect 175812 646718 178099 646720
rect 203964 646776 205699 646778
rect 203964 646720 205638 646776
rect 205694 646720 205699 646776
rect 203964 646718 205699 646720
rect 231932 646776 233299 646778
rect 231932 646720 233238 646776
rect 233294 646720 233299 646776
rect 231932 646718 233299 646720
rect 259900 646776 262279 646778
rect 259900 646720 262218 646776
rect 262274 646720 262279 646776
rect 259900 646718 262279 646720
rect 287868 646776 289879 646778
rect 287868 646720 289818 646776
rect 289874 646720 289879 646776
rect 287868 646718 289879 646720
rect 315836 646776 317479 646778
rect 315836 646720 317418 646776
rect 317474 646720 317479 646776
rect 315836 646718 317479 646720
rect 343804 646776 345079 646778
rect 343804 646720 345018 646776
rect 345074 646720 345079 646776
rect 343804 646718 345079 646720
rect 371956 646776 374059 646778
rect 371956 646720 373998 646776
rect 374054 646720 374059 646776
rect 371956 646718 374059 646720
rect 399924 646776 401659 646778
rect 399924 646720 401598 646776
rect 401654 646720 401659 646776
rect 399924 646718 401659 646720
rect 427892 646776 429351 646778
rect 427892 646720 429290 646776
rect 429346 646720 429351 646776
rect 427892 646718 429351 646720
rect 455860 646776 458239 646778
rect 455860 646720 458178 646776
rect 458234 646720 458239 646776
rect 455860 646718 458239 646720
rect 483828 646776 485839 646778
rect 483828 646720 485778 646776
rect 485834 646720 485839 646776
rect 483828 646718 485839 646720
rect 511796 646776 513439 646778
rect 511796 646720 513378 646776
rect 513434 646720 513439 646776
rect 511796 646718 513439 646720
rect 539948 646776 542419 646778
rect 539948 646720 542358 646776
rect 542414 646720 542419 646776
rect 539948 646718 542419 646720
rect 567916 646776 570019 646778
rect 567916 646720 569958 646776
rect 570014 646720 570019 646776
rect 567916 646718 570019 646720
rect 37273 646715 37339 646718
rect 66253 646715 66319 646718
rect 93853 646715 93919 646718
rect 121453 646715 121519 646718
rect 149053 646715 149119 646718
rect 178033 646715 178099 646718
rect 205633 646715 205699 646718
rect 233233 646715 233299 646718
rect 262213 646715 262279 646718
rect 289813 646715 289879 646718
rect 317413 646715 317479 646718
rect 345013 646715 345079 646718
rect 373993 646715 374059 646718
rect 401593 646715 401659 646718
rect 429285 646715 429351 646718
rect 458173 646715 458239 646718
rect 485773 646715 485839 646718
rect 513373 646715 513439 646718
rect 542353 646715 542419 646718
rect 569953 646715 570019 646718
rect -960 644996 480 645236
rect 580390 643996 580396 644060
rect 580460 644058 580466 644060
rect 583520 644058 584960 644148
rect 580460 643998 584960 644058
rect 580460 643996 580466 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 583520 630716 584960 630956
rect 13537 620258 13603 620261
rect 42701 620258 42767 620261
rect 70301 620258 70367 620261
rect 97901 620258 97967 620261
rect 126881 620258 126947 620261
rect 154481 620258 154547 620261
rect 182081 620258 182147 620261
rect 209681 620258 209747 620261
rect 238661 620258 238727 620261
rect 266261 620258 266327 620261
rect 293861 620258 293927 620261
rect 322841 620258 322907 620261
rect 350441 620258 350507 620261
rect 378041 620258 378107 620261
rect 405641 620258 405707 620261
rect 434621 620258 434687 620261
rect 462221 620258 462287 620261
rect 489821 620258 489887 620261
rect 518801 620258 518867 620261
rect 546401 620258 546467 620261
rect 13537 620256 16100 620258
rect 13537 620200 13542 620256
rect 13598 620200 16100 620256
rect 13537 620198 16100 620200
rect 42701 620256 44068 620258
rect 42701 620200 42706 620256
rect 42762 620200 44068 620256
rect 42701 620198 44068 620200
rect 70301 620256 72036 620258
rect 70301 620200 70306 620256
rect 70362 620200 72036 620256
rect 70301 620198 72036 620200
rect 97901 620256 100188 620258
rect 97901 620200 97906 620256
rect 97962 620200 100188 620256
rect 97901 620198 100188 620200
rect 126881 620256 128156 620258
rect 126881 620200 126886 620256
rect 126942 620200 128156 620256
rect 126881 620198 128156 620200
rect 154481 620256 156124 620258
rect 154481 620200 154486 620256
rect 154542 620200 156124 620256
rect 154481 620198 156124 620200
rect 182081 620256 184092 620258
rect 182081 620200 182086 620256
rect 182142 620200 184092 620256
rect 182081 620198 184092 620200
rect 209681 620256 212060 620258
rect 209681 620200 209686 620256
rect 209742 620200 212060 620256
rect 209681 620198 212060 620200
rect 238661 620256 240212 620258
rect 238661 620200 238666 620256
rect 238722 620200 240212 620256
rect 238661 620198 240212 620200
rect 266261 620256 268180 620258
rect 266261 620200 266266 620256
rect 266322 620200 268180 620256
rect 266261 620198 268180 620200
rect 293861 620256 296148 620258
rect 293861 620200 293866 620256
rect 293922 620200 296148 620256
rect 293861 620198 296148 620200
rect 322841 620256 324116 620258
rect 322841 620200 322846 620256
rect 322902 620200 324116 620256
rect 322841 620198 324116 620200
rect 350441 620256 352084 620258
rect 350441 620200 350446 620256
rect 350502 620200 352084 620256
rect 350441 620198 352084 620200
rect 378041 620256 380052 620258
rect 378041 620200 378046 620256
rect 378102 620200 380052 620256
rect 378041 620198 380052 620200
rect 405641 620256 408204 620258
rect 405641 620200 405646 620256
rect 405702 620200 408204 620256
rect 405641 620198 408204 620200
rect 434621 620256 436172 620258
rect 434621 620200 434626 620256
rect 434682 620200 436172 620256
rect 434621 620198 436172 620200
rect 462221 620256 464140 620258
rect 462221 620200 462226 620256
rect 462282 620200 464140 620256
rect 462221 620198 464140 620200
rect 489821 620256 492108 620258
rect 489821 620200 489826 620256
rect 489882 620200 492108 620256
rect 489821 620198 492108 620200
rect 518801 620256 520076 620258
rect 518801 620200 518806 620256
rect 518862 620200 520076 620256
rect 518801 620198 520076 620200
rect 546401 620256 548044 620258
rect 546401 620200 546406 620256
rect 546462 620200 548044 620256
rect 546401 620198 548044 620200
rect 13537 620195 13603 620198
rect 42701 620195 42767 620198
rect 70301 620195 70367 620198
rect 97901 620195 97967 620198
rect 126881 620195 126947 620198
rect 154481 620195 154547 620198
rect 182081 620195 182147 620198
rect 209681 620195 209747 620198
rect 238661 620195 238727 620198
rect 266261 620195 266327 620198
rect 293861 620195 293927 620198
rect 322841 620195 322907 620198
rect 350441 620195 350507 620198
rect 378041 620195 378107 620198
rect 405641 620195 405707 620198
rect 434621 620195 434687 620198
rect 462221 620195 462287 620198
rect 489821 620195 489887 620198
rect 518801 620195 518867 620198
rect 546401 620195 546467 620198
rect 37273 619578 37339 619581
rect 66253 619578 66319 619581
rect 93853 619578 93919 619581
rect 121453 619578 121519 619581
rect 149053 619578 149119 619581
rect 178033 619578 178099 619581
rect 205633 619578 205699 619581
rect 233233 619578 233299 619581
rect 262213 619578 262279 619581
rect 289813 619578 289879 619581
rect 317413 619578 317479 619581
rect 345013 619578 345079 619581
rect 373993 619578 374059 619581
rect 401593 619578 401659 619581
rect 429285 619578 429351 619581
rect 458173 619578 458239 619581
rect 485773 619578 485839 619581
rect 513373 619578 513439 619581
rect 542353 619578 542419 619581
rect 569953 619578 570019 619581
rect 35788 619576 37339 619578
rect 35788 619520 37278 619576
rect 37334 619520 37339 619576
rect 35788 619518 37339 619520
rect 63940 619576 66319 619578
rect 63940 619520 66258 619576
rect 66314 619520 66319 619576
rect 63940 619518 66319 619520
rect 91908 619576 93919 619578
rect 91908 619520 93858 619576
rect 93914 619520 93919 619576
rect 91908 619518 93919 619520
rect 119876 619576 121519 619578
rect 119876 619520 121458 619576
rect 121514 619520 121519 619576
rect 119876 619518 121519 619520
rect 147844 619576 149119 619578
rect 147844 619520 149058 619576
rect 149114 619520 149119 619576
rect 147844 619518 149119 619520
rect 175812 619576 178099 619578
rect 175812 619520 178038 619576
rect 178094 619520 178099 619576
rect 175812 619518 178099 619520
rect 203964 619576 205699 619578
rect 203964 619520 205638 619576
rect 205694 619520 205699 619576
rect 203964 619518 205699 619520
rect 231932 619576 233299 619578
rect 231932 619520 233238 619576
rect 233294 619520 233299 619576
rect 231932 619518 233299 619520
rect 259900 619576 262279 619578
rect 259900 619520 262218 619576
rect 262274 619520 262279 619576
rect 259900 619518 262279 619520
rect 287868 619576 289879 619578
rect 287868 619520 289818 619576
rect 289874 619520 289879 619576
rect 287868 619518 289879 619520
rect 315836 619576 317479 619578
rect 315836 619520 317418 619576
rect 317474 619520 317479 619576
rect 315836 619518 317479 619520
rect 343804 619576 345079 619578
rect 343804 619520 345018 619576
rect 345074 619520 345079 619576
rect 343804 619518 345079 619520
rect 371956 619576 374059 619578
rect 371956 619520 373998 619576
rect 374054 619520 374059 619576
rect 371956 619518 374059 619520
rect 399924 619576 401659 619578
rect 399924 619520 401598 619576
rect 401654 619520 401659 619576
rect 399924 619518 401659 619520
rect 427892 619576 429351 619578
rect 427892 619520 429290 619576
rect 429346 619520 429351 619576
rect 427892 619518 429351 619520
rect 455860 619576 458239 619578
rect 455860 619520 458178 619576
rect 458234 619520 458239 619576
rect 455860 619518 458239 619520
rect 483828 619576 485839 619578
rect 483828 619520 485778 619576
rect 485834 619520 485839 619576
rect 483828 619518 485839 619520
rect 511796 619576 513439 619578
rect 511796 619520 513378 619576
rect 513434 619520 513439 619576
rect 511796 619518 513439 619520
rect 539948 619576 542419 619578
rect 539948 619520 542358 619576
rect 542414 619520 542419 619576
rect 539948 619518 542419 619520
rect 567916 619576 570019 619578
rect 567916 619520 569958 619576
rect 570014 619520 570019 619576
rect 567916 619518 570019 619520
rect 37273 619515 37339 619518
rect 66253 619515 66319 619518
rect 93853 619515 93919 619518
rect 121453 619515 121519 619518
rect 149053 619515 149119 619518
rect 178033 619515 178099 619518
rect 205633 619515 205699 619518
rect 233233 619515 233299 619518
rect 262213 619515 262279 619518
rect 289813 619515 289879 619518
rect 317413 619515 317479 619518
rect 345013 619515 345079 619518
rect 373993 619515 374059 619518
rect 401593 619515 401659 619518
rect 429285 619515 429351 619518
rect 458173 619515 458239 619518
rect 485773 619515 485839 619518
rect 513373 619515 513439 619518
rect 542353 619515 542419 619518
rect 569953 619515 570019 619518
rect -960 619020 480 619260
rect 580574 617476 580580 617540
rect 580644 617538 580650 617540
rect 583520 617538 584960 617628
rect 580644 617478 584960 617538
rect 580644 617476 580650 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect 13537 593466 13603 593469
rect 42701 593466 42767 593469
rect 70301 593466 70367 593469
rect 97901 593466 97967 593469
rect 126881 593466 126947 593469
rect 154481 593466 154547 593469
rect 182081 593466 182147 593469
rect 209681 593466 209747 593469
rect 238661 593466 238727 593469
rect 266261 593466 266327 593469
rect 293861 593466 293927 593469
rect 322841 593466 322907 593469
rect 350441 593466 350507 593469
rect 378041 593466 378107 593469
rect 405641 593466 405707 593469
rect 434621 593466 434687 593469
rect 462221 593466 462287 593469
rect 489821 593466 489887 593469
rect 518801 593466 518867 593469
rect 546401 593466 546467 593469
rect 13537 593464 16100 593466
rect 13537 593408 13542 593464
rect 13598 593408 16100 593464
rect 13537 593406 16100 593408
rect 42701 593464 44068 593466
rect 42701 593408 42706 593464
rect 42762 593408 44068 593464
rect 42701 593406 44068 593408
rect 70301 593464 72036 593466
rect 70301 593408 70306 593464
rect 70362 593408 72036 593464
rect 70301 593406 72036 593408
rect 97901 593464 100188 593466
rect 97901 593408 97906 593464
rect 97962 593408 100188 593464
rect 97901 593406 100188 593408
rect 126881 593464 128156 593466
rect 126881 593408 126886 593464
rect 126942 593408 128156 593464
rect 126881 593406 128156 593408
rect 154481 593464 156124 593466
rect 154481 593408 154486 593464
rect 154542 593408 156124 593464
rect 154481 593406 156124 593408
rect 182081 593464 184092 593466
rect 182081 593408 182086 593464
rect 182142 593408 184092 593464
rect 182081 593406 184092 593408
rect 209681 593464 212060 593466
rect 209681 593408 209686 593464
rect 209742 593408 212060 593464
rect 209681 593406 212060 593408
rect 238661 593464 240212 593466
rect 238661 593408 238666 593464
rect 238722 593408 240212 593464
rect 238661 593406 240212 593408
rect 266261 593464 268180 593466
rect 266261 593408 266266 593464
rect 266322 593408 268180 593464
rect 266261 593406 268180 593408
rect 293861 593464 296148 593466
rect 293861 593408 293866 593464
rect 293922 593408 296148 593464
rect 293861 593406 296148 593408
rect 322841 593464 324116 593466
rect 322841 593408 322846 593464
rect 322902 593408 324116 593464
rect 322841 593406 324116 593408
rect 350441 593464 352084 593466
rect 350441 593408 350446 593464
rect 350502 593408 352084 593464
rect 350441 593406 352084 593408
rect 378041 593464 380052 593466
rect 378041 593408 378046 593464
rect 378102 593408 380052 593464
rect 378041 593406 380052 593408
rect 405641 593464 408204 593466
rect 405641 593408 405646 593464
rect 405702 593408 408204 593464
rect 405641 593406 408204 593408
rect 434621 593464 436172 593466
rect 434621 593408 434626 593464
rect 434682 593408 436172 593464
rect 434621 593406 436172 593408
rect 462221 593464 464140 593466
rect 462221 593408 462226 593464
rect 462282 593408 464140 593464
rect 462221 593406 464140 593408
rect 489821 593464 492108 593466
rect 489821 593408 489826 593464
rect 489882 593408 492108 593464
rect 489821 593406 492108 593408
rect 518801 593464 520076 593466
rect 518801 593408 518806 593464
rect 518862 593408 520076 593464
rect 518801 593406 520076 593408
rect 546401 593464 548044 593466
rect 546401 593408 546406 593464
rect 546462 593408 548044 593464
rect 546401 593406 548044 593408
rect 13537 593403 13603 593406
rect 42701 593403 42767 593406
rect 70301 593403 70367 593406
rect 97901 593403 97967 593406
rect 126881 593403 126947 593406
rect 154481 593403 154547 593406
rect 182081 593403 182147 593406
rect 209681 593403 209747 593406
rect 238661 593403 238727 593406
rect 266261 593403 266327 593406
rect 293861 593403 293927 593406
rect 322841 593403 322907 593406
rect 350441 593403 350507 593406
rect 378041 593403 378107 593406
rect 405641 593403 405707 593406
rect 434621 593403 434687 593406
rect 462221 593403 462287 593406
rect 489821 593403 489887 593406
rect 518801 593403 518867 593406
rect 546401 593403 546467 593406
rect -960 592908 480 593148
rect 37273 592786 37339 592789
rect 66253 592786 66319 592789
rect 93853 592786 93919 592789
rect 121453 592786 121519 592789
rect 149053 592786 149119 592789
rect 178033 592786 178099 592789
rect 205633 592786 205699 592789
rect 233233 592786 233299 592789
rect 262213 592786 262279 592789
rect 289813 592786 289879 592789
rect 317413 592786 317479 592789
rect 345013 592786 345079 592789
rect 373993 592786 374059 592789
rect 401593 592786 401659 592789
rect 429285 592786 429351 592789
rect 458173 592786 458239 592789
rect 485773 592786 485839 592789
rect 513373 592786 513439 592789
rect 542353 592786 542419 592789
rect 569953 592786 570019 592789
rect 35788 592784 37339 592786
rect 35788 592728 37278 592784
rect 37334 592728 37339 592784
rect 35788 592726 37339 592728
rect 63940 592784 66319 592786
rect 63940 592728 66258 592784
rect 66314 592728 66319 592784
rect 63940 592726 66319 592728
rect 91908 592784 93919 592786
rect 91908 592728 93858 592784
rect 93914 592728 93919 592784
rect 91908 592726 93919 592728
rect 119876 592784 121519 592786
rect 119876 592728 121458 592784
rect 121514 592728 121519 592784
rect 119876 592726 121519 592728
rect 147844 592784 149119 592786
rect 147844 592728 149058 592784
rect 149114 592728 149119 592784
rect 147844 592726 149119 592728
rect 175812 592784 178099 592786
rect 175812 592728 178038 592784
rect 178094 592728 178099 592784
rect 175812 592726 178099 592728
rect 203964 592784 205699 592786
rect 203964 592728 205638 592784
rect 205694 592728 205699 592784
rect 203964 592726 205699 592728
rect 231932 592784 233299 592786
rect 231932 592728 233238 592784
rect 233294 592728 233299 592784
rect 231932 592726 233299 592728
rect 259900 592784 262279 592786
rect 259900 592728 262218 592784
rect 262274 592728 262279 592784
rect 259900 592726 262279 592728
rect 287868 592784 289879 592786
rect 287868 592728 289818 592784
rect 289874 592728 289879 592784
rect 287868 592726 289879 592728
rect 315836 592784 317479 592786
rect 315836 592728 317418 592784
rect 317474 592728 317479 592784
rect 315836 592726 317479 592728
rect 343804 592784 345079 592786
rect 343804 592728 345018 592784
rect 345074 592728 345079 592784
rect 343804 592726 345079 592728
rect 371956 592784 374059 592786
rect 371956 592728 373998 592784
rect 374054 592728 374059 592784
rect 371956 592726 374059 592728
rect 399924 592784 401659 592786
rect 399924 592728 401598 592784
rect 401654 592728 401659 592784
rect 399924 592726 401659 592728
rect 427892 592784 429351 592786
rect 427892 592728 429290 592784
rect 429346 592728 429351 592784
rect 427892 592726 429351 592728
rect 455860 592784 458239 592786
rect 455860 592728 458178 592784
rect 458234 592728 458239 592784
rect 455860 592726 458239 592728
rect 483828 592784 485839 592786
rect 483828 592728 485778 592784
rect 485834 592728 485839 592784
rect 483828 592726 485839 592728
rect 511796 592784 513439 592786
rect 511796 592728 513378 592784
rect 513434 592728 513439 592784
rect 511796 592726 513439 592728
rect 539948 592784 542419 592786
rect 539948 592728 542358 592784
rect 542414 592728 542419 592784
rect 539948 592726 542419 592728
rect 567916 592784 570019 592786
rect 567916 592728 569958 592784
rect 570014 592728 570019 592784
rect 567916 592726 570019 592728
rect 37273 592723 37339 592726
rect 66253 592723 66319 592726
rect 93853 592723 93919 592726
rect 121453 592723 121519 592726
rect 149053 592723 149119 592726
rect 178033 592723 178099 592726
rect 205633 592723 205699 592726
rect 233233 592723 233299 592726
rect 262213 592723 262279 592726
rect 289813 592723 289879 592726
rect 317413 592723 317479 592726
rect 345013 592723 345079 592726
rect 373993 592723 374059 592726
rect 401593 592723 401659 592726
rect 429285 592723 429351 592726
rect 458173 592723 458239 592726
rect 485773 592723 485839 592726
rect 513373 592723 513439 592726
rect 542353 592723 542419 592726
rect 569953 592723 570019 592726
rect 580257 591018 580323 591021
rect 583520 591018 584960 591108
rect 580257 591016 584960 591018
rect 580257 590960 580262 591016
rect 580318 590960 584960 591016
rect 580257 590958 584960 590960
rect 580257 590955 580323 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 13537 566266 13603 566269
rect 42701 566266 42767 566269
rect 70301 566266 70367 566269
rect 97901 566266 97967 566269
rect 126881 566266 126947 566269
rect 154481 566266 154547 566269
rect 182081 566266 182147 566269
rect 209681 566266 209747 566269
rect 238661 566266 238727 566269
rect 266261 566266 266327 566269
rect 293861 566266 293927 566269
rect 322841 566266 322907 566269
rect 350441 566266 350507 566269
rect 378041 566266 378107 566269
rect 405641 566266 405707 566269
rect 434621 566266 434687 566269
rect 462221 566266 462287 566269
rect 489821 566266 489887 566269
rect 518801 566266 518867 566269
rect 546401 566266 546467 566269
rect 13537 566264 16100 566266
rect 13537 566208 13542 566264
rect 13598 566208 16100 566264
rect 13537 566206 16100 566208
rect 42701 566264 44068 566266
rect 42701 566208 42706 566264
rect 42762 566208 44068 566264
rect 42701 566206 44068 566208
rect 70301 566264 72036 566266
rect 70301 566208 70306 566264
rect 70362 566208 72036 566264
rect 70301 566206 72036 566208
rect 97901 566264 100188 566266
rect 97901 566208 97906 566264
rect 97962 566208 100188 566264
rect 97901 566206 100188 566208
rect 126881 566264 128156 566266
rect 126881 566208 126886 566264
rect 126942 566208 128156 566264
rect 126881 566206 128156 566208
rect 154481 566264 156124 566266
rect 154481 566208 154486 566264
rect 154542 566208 156124 566264
rect 154481 566206 156124 566208
rect 182081 566264 184092 566266
rect 182081 566208 182086 566264
rect 182142 566208 184092 566264
rect 182081 566206 184092 566208
rect 209681 566264 212060 566266
rect 209681 566208 209686 566264
rect 209742 566208 212060 566264
rect 209681 566206 212060 566208
rect 238661 566264 240212 566266
rect 238661 566208 238666 566264
rect 238722 566208 240212 566264
rect 238661 566206 240212 566208
rect 266261 566264 268180 566266
rect 266261 566208 266266 566264
rect 266322 566208 268180 566264
rect 266261 566206 268180 566208
rect 293861 566264 296148 566266
rect 293861 566208 293866 566264
rect 293922 566208 296148 566264
rect 293861 566206 296148 566208
rect 322841 566264 324116 566266
rect 322841 566208 322846 566264
rect 322902 566208 324116 566264
rect 322841 566206 324116 566208
rect 350441 566264 352084 566266
rect 350441 566208 350446 566264
rect 350502 566208 352084 566264
rect 350441 566206 352084 566208
rect 378041 566264 380052 566266
rect 378041 566208 378046 566264
rect 378102 566208 380052 566264
rect 378041 566206 380052 566208
rect 405641 566264 408204 566266
rect 405641 566208 405646 566264
rect 405702 566208 408204 566264
rect 405641 566206 408204 566208
rect 434621 566264 436172 566266
rect 434621 566208 434626 566264
rect 434682 566208 436172 566264
rect 434621 566206 436172 566208
rect 462221 566264 464140 566266
rect 462221 566208 462226 566264
rect 462282 566208 464140 566264
rect 462221 566206 464140 566208
rect 489821 566264 492108 566266
rect 489821 566208 489826 566264
rect 489882 566208 492108 566264
rect 489821 566206 492108 566208
rect 518801 566264 520076 566266
rect 518801 566208 518806 566264
rect 518862 566208 520076 566264
rect 518801 566206 520076 566208
rect 546401 566264 548044 566266
rect 546401 566208 546406 566264
rect 546462 566208 548044 566264
rect 546401 566206 548044 566208
rect 13537 566203 13603 566206
rect 42701 566203 42767 566206
rect 70301 566203 70367 566206
rect 97901 566203 97967 566206
rect 126881 566203 126947 566206
rect 154481 566203 154547 566206
rect 182081 566203 182147 566206
rect 209681 566203 209747 566206
rect 238661 566203 238727 566206
rect 266261 566203 266327 566206
rect 293861 566203 293927 566206
rect 322841 566203 322907 566206
rect 350441 566203 350507 566206
rect 378041 566203 378107 566206
rect 405641 566203 405707 566206
rect 434621 566203 434687 566206
rect 462221 566203 462287 566206
rect 489821 566203 489887 566206
rect 518801 566203 518867 566206
rect 546401 566203 546467 566206
rect 37273 565586 37339 565589
rect 66253 565586 66319 565589
rect 93853 565586 93919 565589
rect 121453 565586 121519 565589
rect 149053 565586 149119 565589
rect 178033 565586 178099 565589
rect 205633 565586 205699 565589
rect 233233 565586 233299 565589
rect 262213 565586 262279 565589
rect 289813 565586 289879 565589
rect 317413 565586 317479 565589
rect 345013 565586 345079 565589
rect 373993 565586 374059 565589
rect 401593 565586 401659 565589
rect 429285 565586 429351 565589
rect 458173 565586 458239 565589
rect 485773 565586 485839 565589
rect 513373 565586 513439 565589
rect 542353 565586 542419 565589
rect 569953 565586 570019 565589
rect 35788 565584 37339 565586
rect 35788 565528 37278 565584
rect 37334 565528 37339 565584
rect 35788 565526 37339 565528
rect 63940 565584 66319 565586
rect 63940 565528 66258 565584
rect 66314 565528 66319 565584
rect 63940 565526 66319 565528
rect 91908 565584 93919 565586
rect 91908 565528 93858 565584
rect 93914 565528 93919 565584
rect 91908 565526 93919 565528
rect 119876 565584 121519 565586
rect 119876 565528 121458 565584
rect 121514 565528 121519 565584
rect 119876 565526 121519 565528
rect 147844 565584 149119 565586
rect 147844 565528 149058 565584
rect 149114 565528 149119 565584
rect 147844 565526 149119 565528
rect 175812 565584 178099 565586
rect 175812 565528 178038 565584
rect 178094 565528 178099 565584
rect 175812 565526 178099 565528
rect 203964 565584 205699 565586
rect 203964 565528 205638 565584
rect 205694 565528 205699 565584
rect 203964 565526 205699 565528
rect 231932 565584 233299 565586
rect 231932 565528 233238 565584
rect 233294 565528 233299 565584
rect 231932 565526 233299 565528
rect 259900 565584 262279 565586
rect 259900 565528 262218 565584
rect 262274 565528 262279 565584
rect 259900 565526 262279 565528
rect 287868 565584 289879 565586
rect 287868 565528 289818 565584
rect 289874 565528 289879 565584
rect 287868 565526 289879 565528
rect 315836 565584 317479 565586
rect 315836 565528 317418 565584
rect 317474 565528 317479 565584
rect 315836 565526 317479 565528
rect 343804 565584 345079 565586
rect 343804 565528 345018 565584
rect 345074 565528 345079 565584
rect 343804 565526 345079 565528
rect 371956 565584 374059 565586
rect 371956 565528 373998 565584
rect 374054 565528 374059 565584
rect 371956 565526 374059 565528
rect 399924 565584 401659 565586
rect 399924 565528 401598 565584
rect 401654 565528 401659 565584
rect 399924 565526 401659 565528
rect 427892 565584 429351 565586
rect 427892 565528 429290 565584
rect 429346 565528 429351 565584
rect 427892 565526 429351 565528
rect 455860 565584 458239 565586
rect 455860 565528 458178 565584
rect 458234 565528 458239 565584
rect 455860 565526 458239 565528
rect 483828 565584 485839 565586
rect 483828 565528 485778 565584
rect 485834 565528 485839 565584
rect 483828 565526 485839 565528
rect 511796 565584 513439 565586
rect 511796 565528 513378 565584
rect 513434 565528 513439 565584
rect 511796 565526 513439 565528
rect 539948 565584 542419 565586
rect 539948 565528 542358 565584
rect 542414 565528 542419 565584
rect 539948 565526 542419 565528
rect 567916 565584 570019 565586
rect 567916 565528 569958 565584
rect 570014 565528 570019 565584
rect 567916 565526 570019 565528
rect 37273 565523 37339 565526
rect 66253 565523 66319 565526
rect 93853 565523 93919 565526
rect 121453 565523 121519 565526
rect 149053 565523 149119 565526
rect 178033 565523 178099 565526
rect 205633 565523 205699 565526
rect 233233 565523 233299 565526
rect 262213 565523 262279 565526
rect 289813 565523 289879 565526
rect 317413 565523 317479 565526
rect 345013 565523 345079 565526
rect 373993 565523 374059 565526
rect 401593 565523 401659 565526
rect 429285 565523 429351 565526
rect 458173 565523 458239 565526
rect 485773 565523 485839 565526
rect 513373 565523 513439 565526
rect 542353 565523 542419 565526
rect 569953 565523 570019 565526
rect 580758 564300 580764 564364
rect 580828 564362 580834 564364
rect 583520 564362 584960 564452
rect 580828 564302 584960 564362
rect 580828 564300 580834 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 13537 539474 13603 539477
rect 42701 539474 42767 539477
rect 70301 539474 70367 539477
rect 97901 539474 97967 539477
rect 126881 539474 126947 539477
rect 154481 539474 154547 539477
rect 182081 539474 182147 539477
rect 209681 539474 209747 539477
rect 238661 539474 238727 539477
rect 266261 539474 266327 539477
rect 293861 539474 293927 539477
rect 322841 539474 322907 539477
rect 350441 539474 350507 539477
rect 378041 539474 378107 539477
rect 405641 539474 405707 539477
rect 434621 539474 434687 539477
rect 462221 539474 462287 539477
rect 489821 539474 489887 539477
rect 518801 539474 518867 539477
rect 546401 539474 546467 539477
rect 13537 539472 16100 539474
rect 13537 539416 13542 539472
rect 13598 539416 16100 539472
rect 13537 539414 16100 539416
rect 42701 539472 44068 539474
rect 42701 539416 42706 539472
rect 42762 539416 44068 539472
rect 42701 539414 44068 539416
rect 70301 539472 72036 539474
rect 70301 539416 70306 539472
rect 70362 539416 72036 539472
rect 70301 539414 72036 539416
rect 97901 539472 100188 539474
rect 97901 539416 97906 539472
rect 97962 539416 100188 539472
rect 97901 539414 100188 539416
rect 126881 539472 128156 539474
rect 126881 539416 126886 539472
rect 126942 539416 128156 539472
rect 126881 539414 128156 539416
rect 154481 539472 156124 539474
rect 154481 539416 154486 539472
rect 154542 539416 156124 539472
rect 154481 539414 156124 539416
rect 182081 539472 184092 539474
rect 182081 539416 182086 539472
rect 182142 539416 184092 539472
rect 182081 539414 184092 539416
rect 209681 539472 212060 539474
rect 209681 539416 209686 539472
rect 209742 539416 212060 539472
rect 209681 539414 212060 539416
rect 238661 539472 240212 539474
rect 238661 539416 238666 539472
rect 238722 539416 240212 539472
rect 238661 539414 240212 539416
rect 266261 539472 268180 539474
rect 266261 539416 266266 539472
rect 266322 539416 268180 539472
rect 266261 539414 268180 539416
rect 293861 539472 296148 539474
rect 293861 539416 293866 539472
rect 293922 539416 296148 539472
rect 293861 539414 296148 539416
rect 322841 539472 324116 539474
rect 322841 539416 322846 539472
rect 322902 539416 324116 539472
rect 322841 539414 324116 539416
rect 350441 539472 352084 539474
rect 350441 539416 350446 539472
rect 350502 539416 352084 539472
rect 350441 539414 352084 539416
rect 378041 539472 380052 539474
rect 378041 539416 378046 539472
rect 378102 539416 380052 539472
rect 378041 539414 380052 539416
rect 405641 539472 408204 539474
rect 405641 539416 405646 539472
rect 405702 539416 408204 539472
rect 405641 539414 408204 539416
rect 434621 539472 436172 539474
rect 434621 539416 434626 539472
rect 434682 539416 436172 539472
rect 434621 539414 436172 539416
rect 462221 539472 464140 539474
rect 462221 539416 462226 539472
rect 462282 539416 464140 539472
rect 462221 539414 464140 539416
rect 489821 539472 492108 539474
rect 489821 539416 489826 539472
rect 489882 539416 492108 539472
rect 489821 539414 492108 539416
rect 518801 539472 520076 539474
rect 518801 539416 518806 539472
rect 518862 539416 520076 539472
rect 518801 539414 520076 539416
rect 546401 539472 548044 539474
rect 546401 539416 546406 539472
rect 546462 539416 548044 539472
rect 546401 539414 548044 539416
rect 13537 539411 13603 539414
rect 42701 539411 42767 539414
rect 70301 539411 70367 539414
rect 97901 539411 97967 539414
rect 126881 539411 126947 539414
rect 154481 539411 154547 539414
rect 182081 539411 182147 539414
rect 209681 539411 209747 539414
rect 238661 539411 238727 539414
rect 266261 539411 266327 539414
rect 293861 539411 293927 539414
rect 322841 539411 322907 539414
rect 350441 539411 350507 539414
rect 378041 539411 378107 539414
rect 405641 539411 405707 539414
rect 434621 539411 434687 539414
rect 462221 539411 462287 539414
rect 489821 539411 489887 539414
rect 518801 539411 518867 539414
rect 546401 539411 546467 539414
rect 37273 538794 37339 538797
rect 66253 538794 66319 538797
rect 93853 538794 93919 538797
rect 121453 538794 121519 538797
rect 149053 538794 149119 538797
rect 178033 538794 178099 538797
rect 205633 538794 205699 538797
rect 233233 538794 233299 538797
rect 262213 538794 262279 538797
rect 289813 538794 289879 538797
rect 317413 538794 317479 538797
rect 345013 538794 345079 538797
rect 373993 538794 374059 538797
rect 401593 538794 401659 538797
rect 429285 538794 429351 538797
rect 458173 538794 458239 538797
rect 485773 538794 485839 538797
rect 513373 538794 513439 538797
rect 542353 538794 542419 538797
rect 569953 538794 570019 538797
rect 35788 538792 37339 538794
rect 35788 538736 37278 538792
rect 37334 538736 37339 538792
rect 35788 538734 37339 538736
rect 63940 538792 66319 538794
rect 63940 538736 66258 538792
rect 66314 538736 66319 538792
rect 63940 538734 66319 538736
rect 91908 538792 93919 538794
rect 91908 538736 93858 538792
rect 93914 538736 93919 538792
rect 91908 538734 93919 538736
rect 119876 538792 121519 538794
rect 119876 538736 121458 538792
rect 121514 538736 121519 538792
rect 119876 538734 121519 538736
rect 147844 538792 149119 538794
rect 147844 538736 149058 538792
rect 149114 538736 149119 538792
rect 147844 538734 149119 538736
rect 175812 538792 178099 538794
rect 175812 538736 178038 538792
rect 178094 538736 178099 538792
rect 175812 538734 178099 538736
rect 203964 538792 205699 538794
rect 203964 538736 205638 538792
rect 205694 538736 205699 538792
rect 203964 538734 205699 538736
rect 231932 538792 233299 538794
rect 231932 538736 233238 538792
rect 233294 538736 233299 538792
rect 231932 538734 233299 538736
rect 259900 538792 262279 538794
rect 259900 538736 262218 538792
rect 262274 538736 262279 538792
rect 259900 538734 262279 538736
rect 287868 538792 289879 538794
rect 287868 538736 289818 538792
rect 289874 538736 289879 538792
rect 287868 538734 289879 538736
rect 315836 538792 317479 538794
rect 315836 538736 317418 538792
rect 317474 538736 317479 538792
rect 315836 538734 317479 538736
rect 343804 538792 345079 538794
rect 343804 538736 345018 538792
rect 345074 538736 345079 538792
rect 343804 538734 345079 538736
rect 371956 538792 374059 538794
rect 371956 538736 373998 538792
rect 374054 538736 374059 538792
rect 371956 538734 374059 538736
rect 399924 538792 401659 538794
rect 399924 538736 401598 538792
rect 401654 538736 401659 538792
rect 399924 538734 401659 538736
rect 427892 538792 429351 538794
rect 427892 538736 429290 538792
rect 429346 538736 429351 538792
rect 427892 538734 429351 538736
rect 455860 538792 458239 538794
rect 455860 538736 458178 538792
rect 458234 538736 458239 538792
rect 455860 538734 458239 538736
rect 483828 538792 485839 538794
rect 483828 538736 485778 538792
rect 485834 538736 485839 538792
rect 483828 538734 485839 538736
rect 511796 538792 513439 538794
rect 511796 538736 513378 538792
rect 513434 538736 513439 538792
rect 511796 538734 513439 538736
rect 539948 538792 542419 538794
rect 539948 538736 542358 538792
rect 542414 538736 542419 538792
rect 539948 538734 542419 538736
rect 567916 538792 570019 538794
rect 567916 538736 569958 538792
rect 570014 538736 570019 538792
rect 567916 538734 570019 538736
rect 37273 538731 37339 538734
rect 66253 538731 66319 538734
rect 93853 538731 93919 538734
rect 121453 538731 121519 538734
rect 149053 538731 149119 538734
rect 178033 538731 178099 538734
rect 205633 538731 205699 538734
rect 233233 538731 233299 538734
rect 262213 538731 262279 538734
rect 289813 538731 289879 538734
rect 317413 538731 317479 538734
rect 345013 538731 345079 538734
rect 373993 538731 374059 538734
rect 401593 538731 401659 538734
rect 429285 538731 429351 538734
rect 458173 538731 458239 538734
rect 485773 538731 485839 538734
rect 513373 538731 513439 538734
rect 542353 538731 542419 538734
rect 569953 538731 570019 538734
rect 580349 537842 580415 537845
rect 583520 537842 584960 537932
rect 580349 537840 584960 537842
rect 580349 537784 580354 537840
rect 580410 537784 584960 537840
rect 580349 537782 584960 537784
rect 580349 537779 580415 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2773 527914 2839 527917
rect -960 527912 2839 527914
rect -960 527856 2778 527912
rect 2834 527856 2839 527912
rect -960 527854 2839 527856
rect -960 527764 480 527854
rect 2773 527851 2839 527854
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 13537 512274 13603 512277
rect 42701 512274 42767 512277
rect 70301 512274 70367 512277
rect 97901 512274 97967 512277
rect 126881 512274 126947 512277
rect 154481 512274 154547 512277
rect 182081 512274 182147 512277
rect 209681 512274 209747 512277
rect 238661 512274 238727 512277
rect 266261 512274 266327 512277
rect 293861 512274 293927 512277
rect 322841 512274 322907 512277
rect 350441 512274 350507 512277
rect 378041 512274 378107 512277
rect 405641 512274 405707 512277
rect 434621 512274 434687 512277
rect 462221 512274 462287 512277
rect 489821 512274 489887 512277
rect 518801 512274 518867 512277
rect 546401 512274 546467 512277
rect 13537 512272 16100 512274
rect 13537 512216 13542 512272
rect 13598 512216 16100 512272
rect 13537 512214 16100 512216
rect 42701 512272 44068 512274
rect 42701 512216 42706 512272
rect 42762 512216 44068 512272
rect 42701 512214 44068 512216
rect 70301 512272 72036 512274
rect 70301 512216 70306 512272
rect 70362 512216 72036 512272
rect 70301 512214 72036 512216
rect 97901 512272 100188 512274
rect 97901 512216 97906 512272
rect 97962 512216 100188 512272
rect 97901 512214 100188 512216
rect 126881 512272 128156 512274
rect 126881 512216 126886 512272
rect 126942 512216 128156 512272
rect 126881 512214 128156 512216
rect 154481 512272 156124 512274
rect 154481 512216 154486 512272
rect 154542 512216 156124 512272
rect 154481 512214 156124 512216
rect 182081 512272 184092 512274
rect 182081 512216 182086 512272
rect 182142 512216 184092 512272
rect 182081 512214 184092 512216
rect 209681 512272 212060 512274
rect 209681 512216 209686 512272
rect 209742 512216 212060 512272
rect 209681 512214 212060 512216
rect 238661 512272 240212 512274
rect 238661 512216 238666 512272
rect 238722 512216 240212 512272
rect 238661 512214 240212 512216
rect 266261 512272 268180 512274
rect 266261 512216 266266 512272
rect 266322 512216 268180 512272
rect 266261 512214 268180 512216
rect 293861 512272 296148 512274
rect 293861 512216 293866 512272
rect 293922 512216 296148 512272
rect 293861 512214 296148 512216
rect 322841 512272 324116 512274
rect 322841 512216 322846 512272
rect 322902 512216 324116 512272
rect 322841 512214 324116 512216
rect 350441 512272 352084 512274
rect 350441 512216 350446 512272
rect 350502 512216 352084 512272
rect 350441 512214 352084 512216
rect 378041 512272 380052 512274
rect 378041 512216 378046 512272
rect 378102 512216 380052 512272
rect 378041 512214 380052 512216
rect 405641 512272 408204 512274
rect 405641 512216 405646 512272
rect 405702 512216 408204 512272
rect 405641 512214 408204 512216
rect 434621 512272 436172 512274
rect 434621 512216 434626 512272
rect 434682 512216 436172 512272
rect 434621 512214 436172 512216
rect 462221 512272 464140 512274
rect 462221 512216 462226 512272
rect 462282 512216 464140 512272
rect 462221 512214 464140 512216
rect 489821 512272 492108 512274
rect 489821 512216 489826 512272
rect 489882 512216 492108 512272
rect 489821 512214 492108 512216
rect 518801 512272 520076 512274
rect 518801 512216 518806 512272
rect 518862 512216 520076 512272
rect 518801 512214 520076 512216
rect 546401 512272 548044 512274
rect 546401 512216 546406 512272
rect 546462 512216 548044 512272
rect 546401 512214 548044 512216
rect 13537 512211 13603 512214
rect 42701 512211 42767 512214
rect 70301 512211 70367 512214
rect 97901 512211 97967 512214
rect 126881 512211 126947 512214
rect 154481 512211 154547 512214
rect 182081 512211 182147 512214
rect 209681 512211 209747 512214
rect 238661 512211 238727 512214
rect 266261 512211 266327 512214
rect 293861 512211 293927 512214
rect 322841 512211 322907 512214
rect 350441 512211 350507 512214
rect 378041 512211 378107 512214
rect 405641 512211 405707 512214
rect 434621 512211 434687 512214
rect 462221 512211 462287 512214
rect 489821 512211 489887 512214
rect 518801 512211 518867 512214
rect 546401 512211 546467 512214
rect 37273 511594 37339 511597
rect 66253 511594 66319 511597
rect 93853 511594 93919 511597
rect 121453 511594 121519 511597
rect 149053 511594 149119 511597
rect 178033 511594 178099 511597
rect 205633 511594 205699 511597
rect 233233 511594 233299 511597
rect 262213 511594 262279 511597
rect 289813 511594 289879 511597
rect 317413 511594 317479 511597
rect 345013 511594 345079 511597
rect 373993 511594 374059 511597
rect 401593 511594 401659 511597
rect 429285 511594 429351 511597
rect 458173 511594 458239 511597
rect 485773 511594 485839 511597
rect 513373 511594 513439 511597
rect 542353 511594 542419 511597
rect 569953 511594 570019 511597
rect 35788 511592 37339 511594
rect 35788 511536 37278 511592
rect 37334 511536 37339 511592
rect 35788 511534 37339 511536
rect 63940 511592 66319 511594
rect 63940 511536 66258 511592
rect 66314 511536 66319 511592
rect 63940 511534 66319 511536
rect 91908 511592 93919 511594
rect 91908 511536 93858 511592
rect 93914 511536 93919 511592
rect 91908 511534 93919 511536
rect 119876 511592 121519 511594
rect 119876 511536 121458 511592
rect 121514 511536 121519 511592
rect 119876 511534 121519 511536
rect 147844 511592 149119 511594
rect 147844 511536 149058 511592
rect 149114 511536 149119 511592
rect 147844 511534 149119 511536
rect 175812 511592 178099 511594
rect 175812 511536 178038 511592
rect 178094 511536 178099 511592
rect 175812 511534 178099 511536
rect 203964 511592 205699 511594
rect 203964 511536 205638 511592
rect 205694 511536 205699 511592
rect 203964 511534 205699 511536
rect 231932 511592 233299 511594
rect 231932 511536 233238 511592
rect 233294 511536 233299 511592
rect 231932 511534 233299 511536
rect 259900 511592 262279 511594
rect 259900 511536 262218 511592
rect 262274 511536 262279 511592
rect 259900 511534 262279 511536
rect 287868 511592 289879 511594
rect 287868 511536 289818 511592
rect 289874 511536 289879 511592
rect 287868 511534 289879 511536
rect 315836 511592 317479 511594
rect 315836 511536 317418 511592
rect 317474 511536 317479 511592
rect 315836 511534 317479 511536
rect 343804 511592 345079 511594
rect 343804 511536 345018 511592
rect 345074 511536 345079 511592
rect 343804 511534 345079 511536
rect 371956 511592 374059 511594
rect 371956 511536 373998 511592
rect 374054 511536 374059 511592
rect 371956 511534 374059 511536
rect 399924 511592 401659 511594
rect 399924 511536 401598 511592
rect 401654 511536 401659 511592
rect 399924 511534 401659 511536
rect 427892 511592 429351 511594
rect 427892 511536 429290 511592
rect 429346 511536 429351 511592
rect 427892 511534 429351 511536
rect 455860 511592 458239 511594
rect 455860 511536 458178 511592
rect 458234 511536 458239 511592
rect 455860 511534 458239 511536
rect 483828 511592 485839 511594
rect 483828 511536 485778 511592
rect 485834 511536 485839 511592
rect 483828 511534 485839 511536
rect 511796 511592 513439 511594
rect 511796 511536 513378 511592
rect 513434 511536 513439 511592
rect 511796 511534 513439 511536
rect 539948 511592 542419 511594
rect 539948 511536 542358 511592
rect 542414 511536 542419 511592
rect 539948 511534 542419 511536
rect 567916 511592 570019 511594
rect 567916 511536 569958 511592
rect 570014 511536 570019 511592
rect 567916 511534 570019 511536
rect 37273 511531 37339 511534
rect 66253 511531 66319 511534
rect 93853 511531 93919 511534
rect 121453 511531 121519 511534
rect 149053 511531 149119 511534
rect 178033 511531 178099 511534
rect 205633 511531 205699 511534
rect 233233 511531 233299 511534
rect 262213 511531 262279 511534
rect 289813 511531 289879 511534
rect 317413 511531 317479 511534
rect 345013 511531 345079 511534
rect 373993 511531 374059 511534
rect 401593 511531 401659 511534
rect 429285 511531 429351 511534
rect 458173 511531 458239 511534
rect 485773 511531 485839 511534
rect 513373 511531 513439 511534
rect 542353 511531 542419 511534
rect 569953 511531 570019 511534
rect 580441 511322 580507 511325
rect 583520 511322 584960 511412
rect 580441 511320 584960 511322
rect 580441 511264 580446 511320
rect 580502 511264 584960 511320
rect 580441 511262 584960 511264
rect 580441 511259 580507 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3509 501802 3575 501805
rect -960 501800 3575 501802
rect -960 501744 3514 501800
rect 3570 501744 3575 501800
rect -960 501742 3575 501744
rect -960 501652 480 501742
rect 3509 501739 3575 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 13537 485482 13603 485485
rect 42701 485482 42767 485485
rect 70301 485482 70367 485485
rect 97901 485482 97967 485485
rect 126881 485482 126947 485485
rect 154481 485482 154547 485485
rect 182081 485482 182147 485485
rect 209681 485482 209747 485485
rect 238661 485482 238727 485485
rect 266261 485482 266327 485485
rect 293861 485482 293927 485485
rect 322841 485482 322907 485485
rect 350441 485482 350507 485485
rect 378041 485482 378107 485485
rect 405641 485482 405707 485485
rect 434621 485482 434687 485485
rect 462221 485482 462287 485485
rect 489821 485482 489887 485485
rect 518801 485482 518867 485485
rect 546401 485482 546467 485485
rect 13537 485480 16100 485482
rect 13537 485424 13542 485480
rect 13598 485424 16100 485480
rect 13537 485422 16100 485424
rect 42701 485480 44068 485482
rect 42701 485424 42706 485480
rect 42762 485424 44068 485480
rect 42701 485422 44068 485424
rect 70301 485480 72036 485482
rect 70301 485424 70306 485480
rect 70362 485424 72036 485480
rect 70301 485422 72036 485424
rect 97901 485480 100188 485482
rect 97901 485424 97906 485480
rect 97962 485424 100188 485480
rect 97901 485422 100188 485424
rect 126881 485480 128156 485482
rect 126881 485424 126886 485480
rect 126942 485424 128156 485480
rect 126881 485422 128156 485424
rect 154481 485480 156124 485482
rect 154481 485424 154486 485480
rect 154542 485424 156124 485480
rect 154481 485422 156124 485424
rect 182081 485480 184092 485482
rect 182081 485424 182086 485480
rect 182142 485424 184092 485480
rect 182081 485422 184092 485424
rect 209681 485480 212060 485482
rect 209681 485424 209686 485480
rect 209742 485424 212060 485480
rect 209681 485422 212060 485424
rect 238661 485480 240212 485482
rect 238661 485424 238666 485480
rect 238722 485424 240212 485480
rect 238661 485422 240212 485424
rect 266261 485480 268180 485482
rect 266261 485424 266266 485480
rect 266322 485424 268180 485480
rect 266261 485422 268180 485424
rect 293861 485480 296148 485482
rect 293861 485424 293866 485480
rect 293922 485424 296148 485480
rect 293861 485422 296148 485424
rect 322841 485480 324116 485482
rect 322841 485424 322846 485480
rect 322902 485424 324116 485480
rect 322841 485422 324116 485424
rect 350441 485480 352084 485482
rect 350441 485424 350446 485480
rect 350502 485424 352084 485480
rect 350441 485422 352084 485424
rect 378041 485480 380052 485482
rect 378041 485424 378046 485480
rect 378102 485424 380052 485480
rect 378041 485422 380052 485424
rect 405641 485480 408204 485482
rect 405641 485424 405646 485480
rect 405702 485424 408204 485480
rect 405641 485422 408204 485424
rect 434621 485480 436172 485482
rect 434621 485424 434626 485480
rect 434682 485424 436172 485480
rect 434621 485422 436172 485424
rect 462221 485480 464140 485482
rect 462221 485424 462226 485480
rect 462282 485424 464140 485480
rect 462221 485422 464140 485424
rect 489821 485480 492108 485482
rect 489821 485424 489826 485480
rect 489882 485424 492108 485480
rect 489821 485422 492108 485424
rect 518801 485480 520076 485482
rect 518801 485424 518806 485480
rect 518862 485424 520076 485480
rect 518801 485422 520076 485424
rect 546401 485480 548044 485482
rect 546401 485424 546406 485480
rect 546462 485424 548044 485480
rect 546401 485422 548044 485424
rect 13537 485419 13603 485422
rect 42701 485419 42767 485422
rect 70301 485419 70367 485422
rect 97901 485419 97967 485422
rect 126881 485419 126947 485422
rect 154481 485419 154547 485422
rect 182081 485419 182147 485422
rect 209681 485419 209747 485422
rect 238661 485419 238727 485422
rect 266261 485419 266327 485422
rect 293861 485419 293927 485422
rect 322841 485419 322907 485422
rect 350441 485419 350507 485422
rect 378041 485419 378107 485422
rect 405641 485419 405707 485422
rect 434621 485419 434687 485422
rect 462221 485419 462287 485422
rect 489821 485419 489887 485422
rect 518801 485419 518867 485422
rect 546401 485419 546467 485422
rect 37273 484802 37339 484805
rect 66253 484802 66319 484805
rect 93853 484802 93919 484805
rect 121453 484802 121519 484805
rect 149053 484802 149119 484805
rect 178033 484802 178099 484805
rect 205633 484802 205699 484805
rect 233233 484802 233299 484805
rect 262213 484802 262279 484805
rect 289813 484802 289879 484805
rect 317413 484802 317479 484805
rect 345013 484802 345079 484805
rect 373993 484802 374059 484805
rect 401593 484802 401659 484805
rect 429285 484802 429351 484805
rect 458173 484802 458239 484805
rect 485773 484802 485839 484805
rect 513373 484802 513439 484805
rect 542353 484802 542419 484805
rect 569953 484802 570019 484805
rect 35788 484800 37339 484802
rect 35788 484744 37278 484800
rect 37334 484744 37339 484800
rect 35788 484742 37339 484744
rect 63940 484800 66319 484802
rect 63940 484744 66258 484800
rect 66314 484744 66319 484800
rect 63940 484742 66319 484744
rect 91908 484800 93919 484802
rect 91908 484744 93858 484800
rect 93914 484744 93919 484800
rect 91908 484742 93919 484744
rect 119876 484800 121519 484802
rect 119876 484744 121458 484800
rect 121514 484744 121519 484800
rect 119876 484742 121519 484744
rect 147844 484800 149119 484802
rect 147844 484744 149058 484800
rect 149114 484744 149119 484800
rect 147844 484742 149119 484744
rect 175812 484800 178099 484802
rect 175812 484744 178038 484800
rect 178094 484744 178099 484800
rect 175812 484742 178099 484744
rect 203964 484800 205699 484802
rect 203964 484744 205638 484800
rect 205694 484744 205699 484800
rect 203964 484742 205699 484744
rect 231932 484800 233299 484802
rect 231932 484744 233238 484800
rect 233294 484744 233299 484800
rect 231932 484742 233299 484744
rect 259900 484800 262279 484802
rect 259900 484744 262218 484800
rect 262274 484744 262279 484800
rect 259900 484742 262279 484744
rect 287868 484800 289879 484802
rect 287868 484744 289818 484800
rect 289874 484744 289879 484800
rect 287868 484742 289879 484744
rect 315836 484800 317479 484802
rect 315836 484744 317418 484800
rect 317474 484744 317479 484800
rect 315836 484742 317479 484744
rect 343804 484800 345079 484802
rect 343804 484744 345018 484800
rect 345074 484744 345079 484800
rect 343804 484742 345079 484744
rect 371956 484800 374059 484802
rect 371956 484744 373998 484800
rect 374054 484744 374059 484800
rect 371956 484742 374059 484744
rect 399924 484800 401659 484802
rect 399924 484744 401598 484800
rect 401654 484744 401659 484800
rect 399924 484742 401659 484744
rect 427892 484800 429351 484802
rect 427892 484744 429290 484800
rect 429346 484744 429351 484800
rect 427892 484742 429351 484744
rect 455860 484800 458239 484802
rect 455860 484744 458178 484800
rect 458234 484744 458239 484800
rect 455860 484742 458239 484744
rect 483828 484800 485839 484802
rect 483828 484744 485778 484800
rect 485834 484744 485839 484800
rect 483828 484742 485839 484744
rect 511796 484800 513439 484802
rect 511796 484744 513378 484800
rect 513434 484744 513439 484800
rect 511796 484742 513439 484744
rect 539948 484800 542419 484802
rect 539948 484744 542358 484800
rect 542414 484744 542419 484800
rect 539948 484742 542419 484744
rect 567916 484800 570019 484802
rect 567916 484744 569958 484800
rect 570014 484744 570019 484800
rect 567916 484742 570019 484744
rect 37273 484739 37339 484742
rect 66253 484739 66319 484742
rect 93853 484739 93919 484742
rect 121453 484739 121519 484742
rect 149053 484739 149119 484742
rect 178033 484739 178099 484742
rect 205633 484739 205699 484742
rect 233233 484739 233299 484742
rect 262213 484739 262279 484742
rect 289813 484739 289879 484742
rect 317413 484739 317479 484742
rect 345013 484739 345079 484742
rect 373993 484739 374059 484742
rect 401593 484739 401659 484742
rect 429285 484739 429351 484742
rect 458173 484739 458239 484742
rect 485773 484739 485839 484742
rect 513373 484739 513439 484742
rect 542353 484739 542419 484742
rect 569953 484739 570019 484742
rect 580533 484666 580599 484669
rect 583520 484666 584960 484756
rect 580533 484664 584960 484666
rect 580533 484608 580538 484664
rect 580594 484608 584960 484664
rect 580533 484606 584960 484608
rect 580533 484603 580599 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3601 475690 3667 475693
rect -960 475688 3667 475690
rect -960 475632 3606 475688
rect 3662 475632 3667 475688
rect -960 475630 3667 475632
rect -960 475540 480 475630
rect 3601 475627 3667 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462484 480 462724
rect 13537 458282 13603 458285
rect 42701 458282 42767 458285
rect 70301 458282 70367 458285
rect 97901 458282 97967 458285
rect 126881 458282 126947 458285
rect 154481 458282 154547 458285
rect 182081 458282 182147 458285
rect 209681 458282 209747 458285
rect 238661 458282 238727 458285
rect 266261 458282 266327 458285
rect 293861 458282 293927 458285
rect 322841 458282 322907 458285
rect 350441 458282 350507 458285
rect 378041 458282 378107 458285
rect 405641 458282 405707 458285
rect 434621 458282 434687 458285
rect 462221 458282 462287 458285
rect 489821 458282 489887 458285
rect 518801 458282 518867 458285
rect 546401 458282 546467 458285
rect 13537 458280 16100 458282
rect 13537 458224 13542 458280
rect 13598 458224 16100 458280
rect 13537 458222 16100 458224
rect 42701 458280 44068 458282
rect 42701 458224 42706 458280
rect 42762 458224 44068 458280
rect 42701 458222 44068 458224
rect 70301 458280 72036 458282
rect 70301 458224 70306 458280
rect 70362 458224 72036 458280
rect 70301 458222 72036 458224
rect 97901 458280 100188 458282
rect 97901 458224 97906 458280
rect 97962 458224 100188 458280
rect 97901 458222 100188 458224
rect 126881 458280 128156 458282
rect 126881 458224 126886 458280
rect 126942 458224 128156 458280
rect 126881 458222 128156 458224
rect 154481 458280 156124 458282
rect 154481 458224 154486 458280
rect 154542 458224 156124 458280
rect 154481 458222 156124 458224
rect 182081 458280 184092 458282
rect 182081 458224 182086 458280
rect 182142 458224 184092 458280
rect 182081 458222 184092 458224
rect 209681 458280 212060 458282
rect 209681 458224 209686 458280
rect 209742 458224 212060 458280
rect 209681 458222 212060 458224
rect 238661 458280 240212 458282
rect 238661 458224 238666 458280
rect 238722 458224 240212 458280
rect 238661 458222 240212 458224
rect 266261 458280 268180 458282
rect 266261 458224 266266 458280
rect 266322 458224 268180 458280
rect 266261 458222 268180 458224
rect 293861 458280 296148 458282
rect 293861 458224 293866 458280
rect 293922 458224 296148 458280
rect 293861 458222 296148 458224
rect 322841 458280 324116 458282
rect 322841 458224 322846 458280
rect 322902 458224 324116 458280
rect 322841 458222 324116 458224
rect 350441 458280 352084 458282
rect 350441 458224 350446 458280
rect 350502 458224 352084 458280
rect 350441 458222 352084 458224
rect 378041 458280 380052 458282
rect 378041 458224 378046 458280
rect 378102 458224 380052 458280
rect 378041 458222 380052 458224
rect 405641 458280 408204 458282
rect 405641 458224 405646 458280
rect 405702 458224 408204 458280
rect 405641 458222 408204 458224
rect 434621 458280 436172 458282
rect 434621 458224 434626 458280
rect 434682 458224 436172 458280
rect 434621 458222 436172 458224
rect 462221 458280 464140 458282
rect 462221 458224 462226 458280
rect 462282 458224 464140 458280
rect 462221 458222 464140 458224
rect 489821 458280 492108 458282
rect 489821 458224 489826 458280
rect 489882 458224 492108 458280
rect 489821 458222 492108 458224
rect 518801 458280 520076 458282
rect 518801 458224 518806 458280
rect 518862 458224 520076 458280
rect 518801 458222 520076 458224
rect 546401 458280 548044 458282
rect 546401 458224 546406 458280
rect 546462 458224 548044 458280
rect 546401 458222 548044 458224
rect 13537 458219 13603 458222
rect 42701 458219 42767 458222
rect 70301 458219 70367 458222
rect 97901 458219 97967 458222
rect 126881 458219 126947 458222
rect 154481 458219 154547 458222
rect 182081 458219 182147 458222
rect 209681 458219 209747 458222
rect 238661 458219 238727 458222
rect 266261 458219 266327 458222
rect 293861 458219 293927 458222
rect 322841 458219 322907 458222
rect 350441 458219 350507 458222
rect 378041 458219 378107 458222
rect 405641 458219 405707 458222
rect 434621 458219 434687 458222
rect 462221 458219 462287 458222
rect 489821 458219 489887 458222
rect 518801 458219 518867 458222
rect 546401 458219 546467 458222
rect 583520 457996 584960 458236
rect 37273 457602 37339 457605
rect 66253 457602 66319 457605
rect 93853 457602 93919 457605
rect 121453 457602 121519 457605
rect 149053 457602 149119 457605
rect 178033 457602 178099 457605
rect 205633 457602 205699 457605
rect 233233 457602 233299 457605
rect 262213 457602 262279 457605
rect 289813 457602 289879 457605
rect 317413 457602 317479 457605
rect 345013 457602 345079 457605
rect 373993 457602 374059 457605
rect 401593 457602 401659 457605
rect 429285 457602 429351 457605
rect 458173 457602 458239 457605
rect 485773 457602 485839 457605
rect 513373 457602 513439 457605
rect 542353 457602 542419 457605
rect 569953 457602 570019 457605
rect 35788 457600 37339 457602
rect 35788 457544 37278 457600
rect 37334 457544 37339 457600
rect 35788 457542 37339 457544
rect 63940 457600 66319 457602
rect 63940 457544 66258 457600
rect 66314 457544 66319 457600
rect 63940 457542 66319 457544
rect 91908 457600 93919 457602
rect 91908 457544 93858 457600
rect 93914 457544 93919 457600
rect 91908 457542 93919 457544
rect 119876 457600 121519 457602
rect 119876 457544 121458 457600
rect 121514 457544 121519 457600
rect 119876 457542 121519 457544
rect 147844 457600 149119 457602
rect 147844 457544 149058 457600
rect 149114 457544 149119 457600
rect 147844 457542 149119 457544
rect 175812 457600 178099 457602
rect 175812 457544 178038 457600
rect 178094 457544 178099 457600
rect 175812 457542 178099 457544
rect 203964 457600 205699 457602
rect 203964 457544 205638 457600
rect 205694 457544 205699 457600
rect 203964 457542 205699 457544
rect 231932 457600 233299 457602
rect 231932 457544 233238 457600
rect 233294 457544 233299 457600
rect 231932 457542 233299 457544
rect 259900 457600 262279 457602
rect 259900 457544 262218 457600
rect 262274 457544 262279 457600
rect 259900 457542 262279 457544
rect 287868 457600 289879 457602
rect 287868 457544 289818 457600
rect 289874 457544 289879 457600
rect 287868 457542 289879 457544
rect 315836 457600 317479 457602
rect 315836 457544 317418 457600
rect 317474 457544 317479 457600
rect 315836 457542 317479 457544
rect 343804 457600 345079 457602
rect 343804 457544 345018 457600
rect 345074 457544 345079 457600
rect 343804 457542 345079 457544
rect 371956 457600 374059 457602
rect 371956 457544 373998 457600
rect 374054 457544 374059 457600
rect 371956 457542 374059 457544
rect 399924 457600 401659 457602
rect 399924 457544 401598 457600
rect 401654 457544 401659 457600
rect 399924 457542 401659 457544
rect 427892 457600 429351 457602
rect 427892 457544 429290 457600
rect 429346 457544 429351 457600
rect 427892 457542 429351 457544
rect 455860 457600 458239 457602
rect 455860 457544 458178 457600
rect 458234 457544 458239 457600
rect 455860 457542 458239 457544
rect 483828 457600 485839 457602
rect 483828 457544 485778 457600
rect 485834 457544 485839 457600
rect 483828 457542 485839 457544
rect 511796 457600 513439 457602
rect 511796 457544 513378 457600
rect 513434 457544 513439 457600
rect 511796 457542 513439 457544
rect 539948 457600 542419 457602
rect 539948 457544 542358 457600
rect 542414 457544 542419 457600
rect 539948 457542 542419 457544
rect 567916 457600 570019 457602
rect 567916 457544 569958 457600
rect 570014 457544 570019 457600
rect 567916 457542 570019 457544
rect 37273 457539 37339 457542
rect 66253 457539 66319 457542
rect 93853 457539 93919 457542
rect 121453 457539 121519 457542
rect 149053 457539 149119 457542
rect 178033 457539 178099 457542
rect 205633 457539 205699 457542
rect 233233 457539 233299 457542
rect 262213 457539 262279 457542
rect 289813 457539 289879 457542
rect 317413 457539 317479 457542
rect 345013 457539 345079 457542
rect 373993 457539 374059 457542
rect 401593 457539 401659 457542
rect 429285 457539 429351 457542
rect 458173 457539 458239 457542
rect 485773 457539 485839 457542
rect 513373 457539 513439 457542
rect 542353 457539 542419 457542
rect 569953 457539 570019 457542
rect -960 449578 480 449668
rect 2773 449578 2839 449581
rect -960 449576 2839 449578
rect -960 449520 2778 449576
rect 2834 449520 2839 449576
rect -960 449518 2839 449520
rect -960 449428 480 449518
rect 2773 449515 2839 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580625 431626 580691 431629
rect 583520 431626 584960 431716
rect 580625 431624 584960 431626
rect 580625 431568 580630 431624
rect 580686 431568 584960 431624
rect 580625 431566 584960 431568
rect 580625 431563 580691 431566
rect 13537 431490 13603 431493
rect 42701 431490 42767 431493
rect 97901 431490 97967 431493
rect 126881 431490 126947 431493
rect 154481 431490 154547 431493
rect 182081 431490 182147 431493
rect 209681 431490 209747 431493
rect 238661 431490 238727 431493
rect 266261 431490 266327 431493
rect 293861 431490 293927 431493
rect 322841 431490 322907 431493
rect 350441 431490 350507 431493
rect 378041 431490 378107 431493
rect 405641 431490 405707 431493
rect 434621 431490 434687 431493
rect 462221 431490 462287 431493
rect 489821 431490 489887 431493
rect 518801 431490 518867 431493
rect 546401 431490 546467 431493
rect 13537 431488 16100 431490
rect 13537 431432 13542 431488
rect 13598 431432 16100 431488
rect 13537 431430 16100 431432
rect 42701 431488 44068 431490
rect 42701 431432 42706 431488
rect 42762 431432 44068 431488
rect 97901 431488 100188 431490
rect 42701 431430 44068 431432
rect 13537 431427 13603 431430
rect 42701 431427 42767 431430
rect 70301 430946 70367 430949
rect 72006 430946 72066 431460
rect 97901 431432 97906 431488
rect 97962 431432 100188 431488
rect 97901 431430 100188 431432
rect 126881 431488 128156 431490
rect 126881 431432 126886 431488
rect 126942 431432 128156 431488
rect 126881 431430 128156 431432
rect 154481 431488 156124 431490
rect 154481 431432 154486 431488
rect 154542 431432 156124 431488
rect 154481 431430 156124 431432
rect 182081 431488 184092 431490
rect 182081 431432 182086 431488
rect 182142 431432 184092 431488
rect 182081 431430 184092 431432
rect 209681 431488 212060 431490
rect 209681 431432 209686 431488
rect 209742 431432 212060 431488
rect 209681 431430 212060 431432
rect 238661 431488 240212 431490
rect 238661 431432 238666 431488
rect 238722 431432 240212 431488
rect 238661 431430 240212 431432
rect 266261 431488 268180 431490
rect 266261 431432 266266 431488
rect 266322 431432 268180 431488
rect 266261 431430 268180 431432
rect 293861 431488 296148 431490
rect 293861 431432 293866 431488
rect 293922 431432 296148 431488
rect 293861 431430 296148 431432
rect 322841 431488 324116 431490
rect 322841 431432 322846 431488
rect 322902 431432 324116 431488
rect 322841 431430 324116 431432
rect 350441 431488 352084 431490
rect 350441 431432 350446 431488
rect 350502 431432 352084 431488
rect 350441 431430 352084 431432
rect 378041 431488 380052 431490
rect 378041 431432 378046 431488
rect 378102 431432 380052 431488
rect 378041 431430 380052 431432
rect 405641 431488 408204 431490
rect 405641 431432 405646 431488
rect 405702 431432 408204 431488
rect 405641 431430 408204 431432
rect 434621 431488 436172 431490
rect 434621 431432 434626 431488
rect 434682 431432 436172 431488
rect 434621 431430 436172 431432
rect 462221 431488 464140 431490
rect 462221 431432 462226 431488
rect 462282 431432 464140 431488
rect 462221 431430 464140 431432
rect 489821 431488 492108 431490
rect 489821 431432 489826 431488
rect 489882 431432 492108 431488
rect 489821 431430 492108 431432
rect 518801 431488 520076 431490
rect 518801 431432 518806 431488
rect 518862 431432 520076 431488
rect 518801 431430 520076 431432
rect 546401 431488 548044 431490
rect 546401 431432 546406 431488
rect 546462 431432 548044 431488
rect 583520 431476 584960 431566
rect 546401 431430 548044 431432
rect 97901 431427 97967 431430
rect 126881 431427 126947 431430
rect 154481 431427 154547 431430
rect 182081 431427 182147 431430
rect 209681 431427 209747 431430
rect 238661 431427 238727 431430
rect 266261 431427 266327 431430
rect 293861 431427 293927 431430
rect 322841 431427 322907 431430
rect 350441 431427 350507 431430
rect 378041 431427 378107 431430
rect 405641 431427 405707 431430
rect 434621 431427 434687 431430
rect 462221 431427 462287 431430
rect 489821 431427 489887 431430
rect 518801 431427 518867 431430
rect 546401 431427 546467 431430
rect 205633 431354 205699 431357
rect 70301 430944 72066 430946
rect 70301 430888 70306 430944
rect 70362 430888 72066 430944
rect 70301 430886 72066 430888
rect 203934 431352 205699 431354
rect 203934 431296 205638 431352
rect 205694 431296 205699 431352
rect 203934 431294 205699 431296
rect 70301 430883 70367 430886
rect 37273 430810 37339 430813
rect 66253 430810 66319 430813
rect 93853 430810 93919 430813
rect 121453 430810 121519 430813
rect 149053 430810 149119 430813
rect 178033 430810 178099 430813
rect 35788 430808 37339 430810
rect 35788 430752 37278 430808
rect 37334 430752 37339 430808
rect 35788 430750 37339 430752
rect 63940 430808 66319 430810
rect 63940 430752 66258 430808
rect 66314 430752 66319 430808
rect 63940 430750 66319 430752
rect 91908 430808 93919 430810
rect 91908 430752 93858 430808
rect 93914 430752 93919 430808
rect 91908 430750 93919 430752
rect 119876 430808 121519 430810
rect 119876 430752 121458 430808
rect 121514 430752 121519 430808
rect 119876 430750 121519 430752
rect 147844 430808 149119 430810
rect 147844 430752 149058 430808
rect 149114 430752 149119 430808
rect 147844 430750 149119 430752
rect 175812 430808 178099 430810
rect 175812 430752 178038 430808
rect 178094 430752 178099 430808
rect 203934 430780 203994 431294
rect 205633 431291 205699 431294
rect 233233 430810 233299 430813
rect 262213 430810 262279 430813
rect 289813 430810 289879 430813
rect 317413 430810 317479 430813
rect 345013 430810 345079 430813
rect 373993 430810 374059 430813
rect 401593 430810 401659 430813
rect 429285 430810 429351 430813
rect 458173 430810 458239 430813
rect 485773 430810 485839 430813
rect 513373 430810 513439 430813
rect 542353 430810 542419 430813
rect 569953 430810 570019 430813
rect 231932 430808 233299 430810
rect 175812 430750 178099 430752
rect 231932 430752 233238 430808
rect 233294 430752 233299 430808
rect 231932 430750 233299 430752
rect 259900 430808 262279 430810
rect 259900 430752 262218 430808
rect 262274 430752 262279 430808
rect 259900 430750 262279 430752
rect 287868 430808 289879 430810
rect 287868 430752 289818 430808
rect 289874 430752 289879 430808
rect 287868 430750 289879 430752
rect 315836 430808 317479 430810
rect 315836 430752 317418 430808
rect 317474 430752 317479 430808
rect 315836 430750 317479 430752
rect 343804 430808 345079 430810
rect 343804 430752 345018 430808
rect 345074 430752 345079 430808
rect 343804 430750 345079 430752
rect 371956 430808 374059 430810
rect 371956 430752 373998 430808
rect 374054 430752 374059 430808
rect 371956 430750 374059 430752
rect 399924 430808 401659 430810
rect 399924 430752 401598 430808
rect 401654 430752 401659 430808
rect 399924 430750 401659 430752
rect 427892 430808 429351 430810
rect 427892 430752 429290 430808
rect 429346 430752 429351 430808
rect 427892 430750 429351 430752
rect 455860 430808 458239 430810
rect 455860 430752 458178 430808
rect 458234 430752 458239 430808
rect 455860 430750 458239 430752
rect 483828 430808 485839 430810
rect 483828 430752 485778 430808
rect 485834 430752 485839 430808
rect 483828 430750 485839 430752
rect 511796 430808 513439 430810
rect 511796 430752 513378 430808
rect 513434 430752 513439 430808
rect 511796 430750 513439 430752
rect 539948 430808 542419 430810
rect 539948 430752 542358 430808
rect 542414 430752 542419 430808
rect 539948 430750 542419 430752
rect 567916 430808 570019 430810
rect 567916 430752 569958 430808
rect 570014 430752 570019 430808
rect 567916 430750 570019 430752
rect 37273 430747 37339 430750
rect 66253 430747 66319 430750
rect 93853 430747 93919 430750
rect 121453 430747 121519 430750
rect 149053 430747 149119 430750
rect 178033 430747 178099 430750
rect 233233 430747 233299 430750
rect 262213 430747 262279 430750
rect 289813 430747 289879 430750
rect 317413 430747 317479 430750
rect 345013 430747 345079 430750
rect 373993 430747 374059 430750
rect 401593 430747 401659 430750
rect 429285 430747 429351 430750
rect 458173 430747 458239 430750
rect 485773 430747 485839 430750
rect 513373 430747 513439 430750
rect 542353 430747 542419 430750
rect 569953 430747 570019 430750
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 580717 404970 580783 404973
rect 583520 404970 584960 405060
rect 580717 404968 584960 404970
rect 580717 404912 580722 404968
rect 580778 404912 584960 404968
rect 580717 404910 584960 404912
rect 580717 404907 580783 404910
rect 583520 404820 584960 404910
rect 13537 404290 13603 404293
rect 42701 404290 42767 404293
rect 70301 404290 70367 404293
rect 97901 404290 97967 404293
rect 126881 404290 126947 404293
rect 154481 404290 154547 404293
rect 182081 404290 182147 404293
rect 209681 404290 209747 404293
rect 238661 404290 238727 404293
rect 266261 404290 266327 404293
rect 293861 404290 293927 404293
rect 322841 404290 322907 404293
rect 350441 404290 350507 404293
rect 378041 404290 378107 404293
rect 405641 404290 405707 404293
rect 434621 404290 434687 404293
rect 462221 404290 462287 404293
rect 489821 404290 489887 404293
rect 518801 404290 518867 404293
rect 546401 404290 546467 404293
rect 13537 404288 16100 404290
rect 13537 404232 13542 404288
rect 13598 404232 16100 404288
rect 13537 404230 16100 404232
rect 42701 404288 44068 404290
rect 42701 404232 42706 404288
rect 42762 404232 44068 404288
rect 42701 404230 44068 404232
rect 70301 404288 72036 404290
rect 70301 404232 70306 404288
rect 70362 404232 72036 404288
rect 70301 404230 72036 404232
rect 97901 404288 100188 404290
rect 97901 404232 97906 404288
rect 97962 404232 100188 404288
rect 97901 404230 100188 404232
rect 126881 404288 128156 404290
rect 126881 404232 126886 404288
rect 126942 404232 128156 404288
rect 126881 404230 128156 404232
rect 154481 404288 156124 404290
rect 154481 404232 154486 404288
rect 154542 404232 156124 404288
rect 154481 404230 156124 404232
rect 182081 404288 184092 404290
rect 182081 404232 182086 404288
rect 182142 404232 184092 404288
rect 182081 404230 184092 404232
rect 209681 404288 212060 404290
rect 209681 404232 209686 404288
rect 209742 404232 212060 404288
rect 209681 404230 212060 404232
rect 238661 404288 240212 404290
rect 238661 404232 238666 404288
rect 238722 404232 240212 404288
rect 238661 404230 240212 404232
rect 266261 404288 268180 404290
rect 266261 404232 266266 404288
rect 266322 404232 268180 404288
rect 266261 404230 268180 404232
rect 293861 404288 296148 404290
rect 293861 404232 293866 404288
rect 293922 404232 296148 404288
rect 293861 404230 296148 404232
rect 322841 404288 324116 404290
rect 322841 404232 322846 404288
rect 322902 404232 324116 404288
rect 322841 404230 324116 404232
rect 350441 404288 352084 404290
rect 350441 404232 350446 404288
rect 350502 404232 352084 404288
rect 350441 404230 352084 404232
rect 378041 404288 380052 404290
rect 378041 404232 378046 404288
rect 378102 404232 380052 404288
rect 378041 404230 380052 404232
rect 405641 404288 408204 404290
rect 405641 404232 405646 404288
rect 405702 404232 408204 404288
rect 405641 404230 408204 404232
rect 434621 404288 436172 404290
rect 434621 404232 434626 404288
rect 434682 404232 436172 404288
rect 434621 404230 436172 404232
rect 462221 404288 464140 404290
rect 462221 404232 462226 404288
rect 462282 404232 464140 404288
rect 462221 404230 464140 404232
rect 489821 404288 492108 404290
rect 489821 404232 489826 404288
rect 489882 404232 492108 404288
rect 489821 404230 492108 404232
rect 518801 404288 520076 404290
rect 518801 404232 518806 404288
rect 518862 404232 520076 404288
rect 518801 404230 520076 404232
rect 546401 404288 548044 404290
rect 546401 404232 546406 404288
rect 546462 404232 548044 404288
rect 546401 404230 548044 404232
rect 13537 404227 13603 404230
rect 42701 404227 42767 404230
rect 70301 404227 70367 404230
rect 97901 404227 97967 404230
rect 126881 404227 126947 404230
rect 154481 404227 154547 404230
rect 182081 404227 182147 404230
rect 209681 404227 209747 404230
rect 238661 404227 238727 404230
rect 266261 404227 266327 404230
rect 293861 404227 293927 404230
rect 322841 404227 322907 404230
rect 350441 404227 350507 404230
rect 378041 404227 378107 404230
rect 405641 404227 405707 404230
rect 434621 404227 434687 404230
rect 462221 404227 462287 404230
rect 489821 404227 489887 404230
rect 518801 404227 518867 404230
rect 546401 404227 546467 404230
rect 37273 403610 37339 403613
rect 66253 403610 66319 403613
rect 93853 403610 93919 403613
rect 121453 403610 121519 403613
rect 149053 403610 149119 403613
rect 178033 403610 178099 403613
rect 205633 403610 205699 403613
rect 233233 403610 233299 403613
rect 262213 403610 262279 403613
rect 289813 403610 289879 403613
rect 317413 403610 317479 403613
rect 345013 403610 345079 403613
rect 373993 403610 374059 403613
rect 401593 403610 401659 403613
rect 429285 403610 429351 403613
rect 458173 403610 458239 403613
rect 485773 403610 485839 403613
rect 513373 403610 513439 403613
rect 542353 403610 542419 403613
rect 569953 403610 570019 403613
rect 35788 403608 37339 403610
rect 35788 403552 37278 403608
rect 37334 403552 37339 403608
rect 35788 403550 37339 403552
rect 63940 403608 66319 403610
rect 63940 403552 66258 403608
rect 66314 403552 66319 403608
rect 63940 403550 66319 403552
rect 91908 403608 93919 403610
rect 91908 403552 93858 403608
rect 93914 403552 93919 403608
rect 91908 403550 93919 403552
rect 119876 403608 121519 403610
rect 119876 403552 121458 403608
rect 121514 403552 121519 403608
rect 119876 403550 121519 403552
rect 147844 403608 149119 403610
rect 147844 403552 149058 403608
rect 149114 403552 149119 403608
rect 147844 403550 149119 403552
rect 175812 403608 178099 403610
rect 175812 403552 178038 403608
rect 178094 403552 178099 403608
rect 175812 403550 178099 403552
rect 203964 403608 205699 403610
rect 203964 403552 205638 403608
rect 205694 403552 205699 403608
rect 203964 403550 205699 403552
rect 231932 403608 233299 403610
rect 231932 403552 233238 403608
rect 233294 403552 233299 403608
rect 231932 403550 233299 403552
rect 259900 403608 262279 403610
rect 259900 403552 262218 403608
rect 262274 403552 262279 403608
rect 259900 403550 262279 403552
rect 287868 403608 289879 403610
rect 287868 403552 289818 403608
rect 289874 403552 289879 403608
rect 287868 403550 289879 403552
rect 315836 403608 317479 403610
rect 315836 403552 317418 403608
rect 317474 403552 317479 403608
rect 315836 403550 317479 403552
rect 343804 403608 345079 403610
rect 343804 403552 345018 403608
rect 345074 403552 345079 403608
rect 343804 403550 345079 403552
rect 371956 403608 374059 403610
rect 371956 403552 373998 403608
rect 374054 403552 374059 403608
rect 371956 403550 374059 403552
rect 399924 403608 401659 403610
rect 399924 403552 401598 403608
rect 401654 403552 401659 403608
rect 399924 403550 401659 403552
rect 427892 403608 429351 403610
rect 427892 403552 429290 403608
rect 429346 403552 429351 403608
rect 427892 403550 429351 403552
rect 455860 403608 458239 403610
rect 455860 403552 458178 403608
rect 458234 403552 458239 403608
rect 455860 403550 458239 403552
rect 483828 403608 485839 403610
rect 483828 403552 485778 403608
rect 485834 403552 485839 403608
rect 483828 403550 485839 403552
rect 511796 403608 513439 403610
rect 511796 403552 513378 403608
rect 513434 403552 513439 403608
rect 511796 403550 513439 403552
rect 539948 403608 542419 403610
rect 539948 403552 542358 403608
rect 542414 403552 542419 403608
rect 539948 403550 542419 403552
rect 567916 403608 570019 403610
rect 567916 403552 569958 403608
rect 570014 403552 570019 403608
rect 567916 403550 570019 403552
rect 37273 403547 37339 403550
rect 66253 403547 66319 403550
rect 93853 403547 93919 403550
rect 121453 403547 121519 403550
rect 149053 403547 149119 403550
rect 178033 403547 178099 403550
rect 205633 403547 205699 403550
rect 233233 403547 233299 403550
rect 262213 403547 262279 403550
rect 289813 403547 289879 403550
rect 317413 403547 317479 403550
rect 345013 403547 345079 403550
rect 373993 403547 374059 403550
rect 401593 403547 401659 403550
rect 429285 403547 429351 403550
rect 458173 403547 458239 403550
rect 485773 403547 485839 403550
rect 513373 403547 513439 403550
rect 542353 403547 542419 403550
rect 569953 403547 570019 403550
rect -960 397490 480 397580
rect 3693 397490 3759 397493
rect -960 397488 3759 397490
rect -960 397432 3698 397488
rect 3754 397432 3759 397488
rect -960 397430 3759 397432
rect -960 397340 480 397430
rect 3693 397427 3759 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 70301 378042 70367 378045
rect 70301 378040 72066 378042
rect 70301 377984 70306 378040
rect 70362 377984 72066 378040
rect 70301 377982 72066 377984
rect 70301 377979 70367 377982
rect 13537 377498 13603 377501
rect 42701 377498 42767 377501
rect 13537 377496 16100 377498
rect 13537 377440 13542 377496
rect 13598 377440 16100 377496
rect 13537 377438 16100 377440
rect 42701 377496 44068 377498
rect 42701 377440 42706 377496
rect 42762 377440 44068 377496
rect 72006 377468 72066 377982
rect 97901 377498 97967 377501
rect 126881 377498 126947 377501
rect 154481 377498 154547 377501
rect 182081 377498 182147 377501
rect 209681 377498 209747 377501
rect 238661 377498 238727 377501
rect 266261 377498 266327 377501
rect 293861 377498 293927 377501
rect 322841 377498 322907 377501
rect 350441 377498 350507 377501
rect 378041 377498 378107 377501
rect 405641 377498 405707 377501
rect 434621 377498 434687 377501
rect 462221 377498 462287 377501
rect 489821 377498 489887 377501
rect 518801 377498 518867 377501
rect 97901 377496 100188 377498
rect 42701 377438 44068 377440
rect 97901 377440 97906 377496
rect 97962 377440 100188 377496
rect 97901 377438 100188 377440
rect 126881 377496 128156 377498
rect 126881 377440 126886 377496
rect 126942 377440 128156 377496
rect 126881 377438 128156 377440
rect 154481 377496 156124 377498
rect 154481 377440 154486 377496
rect 154542 377440 156124 377496
rect 154481 377438 156124 377440
rect 182081 377496 184092 377498
rect 182081 377440 182086 377496
rect 182142 377440 184092 377496
rect 182081 377438 184092 377440
rect 209681 377496 212060 377498
rect 209681 377440 209686 377496
rect 209742 377440 212060 377496
rect 209681 377438 212060 377440
rect 238661 377496 240212 377498
rect 238661 377440 238666 377496
rect 238722 377440 240212 377496
rect 238661 377438 240212 377440
rect 266261 377496 268180 377498
rect 266261 377440 266266 377496
rect 266322 377440 268180 377496
rect 266261 377438 268180 377440
rect 293861 377496 296148 377498
rect 293861 377440 293866 377496
rect 293922 377440 296148 377496
rect 293861 377438 296148 377440
rect 322841 377496 324116 377498
rect 322841 377440 322846 377496
rect 322902 377440 324116 377496
rect 322841 377438 324116 377440
rect 350441 377496 352084 377498
rect 350441 377440 350446 377496
rect 350502 377440 352084 377496
rect 350441 377438 352084 377440
rect 378041 377496 380052 377498
rect 378041 377440 378046 377496
rect 378102 377440 380052 377496
rect 378041 377438 380052 377440
rect 405641 377496 408204 377498
rect 405641 377440 405646 377496
rect 405702 377440 408204 377496
rect 405641 377438 408204 377440
rect 434621 377496 436172 377498
rect 434621 377440 434626 377496
rect 434682 377440 436172 377496
rect 434621 377438 436172 377440
rect 462221 377496 464140 377498
rect 462221 377440 462226 377496
rect 462282 377440 464140 377496
rect 462221 377438 464140 377440
rect 489821 377496 492108 377498
rect 489821 377440 489826 377496
rect 489882 377440 492108 377496
rect 489821 377438 492108 377440
rect 518801 377496 520076 377498
rect 518801 377440 518806 377496
rect 518862 377440 520076 377496
rect 518801 377438 520076 377440
rect 13537 377435 13603 377438
rect 42701 377435 42767 377438
rect 97901 377435 97967 377438
rect 126881 377435 126947 377438
rect 154481 377435 154547 377438
rect 182081 377435 182147 377438
rect 209681 377435 209747 377438
rect 238661 377435 238727 377438
rect 266261 377435 266327 377438
rect 293861 377435 293927 377438
rect 322841 377435 322907 377438
rect 350441 377435 350507 377438
rect 378041 377435 378107 377438
rect 405641 377435 405707 377438
rect 434621 377435 434687 377438
rect 462221 377435 462287 377438
rect 489821 377435 489887 377438
rect 518801 377435 518867 377438
rect 205633 377362 205699 377365
rect 373993 377362 374059 377365
rect 203934 377360 205699 377362
rect 203934 377304 205638 377360
rect 205694 377304 205699 377360
rect 203934 377302 205699 377304
rect 37273 376818 37339 376821
rect 66253 376818 66319 376821
rect 93853 376818 93919 376821
rect 121453 376818 121519 376821
rect 149053 376818 149119 376821
rect 178033 376818 178099 376821
rect 35788 376816 37339 376818
rect 35788 376760 37278 376816
rect 37334 376760 37339 376816
rect 35788 376758 37339 376760
rect 63940 376816 66319 376818
rect 63940 376760 66258 376816
rect 66314 376760 66319 376816
rect 63940 376758 66319 376760
rect 91908 376816 93919 376818
rect 91908 376760 93858 376816
rect 93914 376760 93919 376816
rect 91908 376758 93919 376760
rect 119876 376816 121519 376818
rect 119876 376760 121458 376816
rect 121514 376760 121519 376816
rect 119876 376758 121519 376760
rect 147844 376816 149119 376818
rect 147844 376760 149058 376816
rect 149114 376760 149119 376816
rect 147844 376758 149119 376760
rect 175812 376816 178099 376818
rect 175812 376760 178038 376816
rect 178094 376760 178099 376816
rect 203934 376788 203994 377302
rect 205633 377299 205699 377302
rect 371926 377360 374059 377362
rect 371926 377304 373998 377360
rect 374054 377304 374059 377360
rect 371926 377302 374059 377304
rect 233233 376818 233299 376821
rect 262213 376818 262279 376821
rect 289813 376818 289879 376821
rect 317413 376818 317479 376821
rect 345013 376818 345079 376821
rect 231932 376816 233299 376818
rect 175812 376758 178099 376760
rect 231932 376760 233238 376816
rect 233294 376760 233299 376816
rect 231932 376758 233299 376760
rect 259900 376816 262279 376818
rect 259900 376760 262218 376816
rect 262274 376760 262279 376816
rect 259900 376758 262279 376760
rect 287868 376816 289879 376818
rect 287868 376760 289818 376816
rect 289874 376760 289879 376816
rect 287868 376758 289879 376760
rect 315836 376816 317479 376818
rect 315836 376760 317418 376816
rect 317474 376760 317479 376816
rect 315836 376758 317479 376760
rect 343804 376816 345079 376818
rect 343804 376760 345018 376816
rect 345074 376760 345079 376816
rect 371926 376788 371986 377302
rect 373993 377299 374059 377302
rect 546401 377090 546467 377093
rect 548014 377090 548074 377468
rect 546401 377088 548074 377090
rect 546401 377032 546406 377088
rect 546462 377032 548074 377088
rect 546401 377030 548074 377032
rect 546401 377027 546467 377030
rect 401593 376818 401659 376821
rect 429285 376818 429351 376821
rect 458173 376818 458239 376821
rect 485773 376818 485839 376821
rect 513373 376818 513439 376821
rect 542353 376818 542419 376821
rect 569953 376818 570019 376821
rect 399924 376816 401659 376818
rect 343804 376758 345079 376760
rect 399924 376760 401598 376816
rect 401654 376760 401659 376816
rect 399924 376758 401659 376760
rect 427892 376816 429351 376818
rect 427892 376760 429290 376816
rect 429346 376760 429351 376816
rect 427892 376758 429351 376760
rect 455860 376816 458239 376818
rect 455860 376760 458178 376816
rect 458234 376760 458239 376816
rect 455860 376758 458239 376760
rect 483828 376816 485839 376818
rect 483828 376760 485778 376816
rect 485834 376760 485839 376816
rect 483828 376758 485839 376760
rect 511796 376816 513439 376818
rect 511796 376760 513378 376816
rect 513434 376760 513439 376816
rect 511796 376758 513439 376760
rect 539948 376816 542419 376818
rect 539948 376760 542358 376816
rect 542414 376760 542419 376816
rect 539948 376758 542419 376760
rect 567916 376816 570019 376818
rect 567916 376760 569958 376816
rect 570014 376760 570019 376816
rect 567916 376758 570019 376760
rect 37273 376755 37339 376758
rect 66253 376755 66319 376758
rect 93853 376755 93919 376758
rect 121453 376755 121519 376758
rect 149053 376755 149119 376758
rect 178033 376755 178099 376758
rect 233233 376755 233299 376758
rect 262213 376755 262279 376758
rect 289813 376755 289879 376758
rect 317413 376755 317479 376758
rect 345013 376755 345079 376758
rect 401593 376755 401659 376758
rect 429285 376755 429351 376758
rect 458173 376755 458239 376758
rect 485773 376755 485839 376758
rect 513373 376755 513439 376758
rect 542353 376755 542419 376758
rect 569953 376755 570019 376758
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358458 480 358548
rect 3785 358458 3851 358461
rect -960 358456 3851 358458
rect -960 358400 3790 358456
rect 3846 358400 3851 358456
rect -960 358398 3851 358400
rect -960 358308 480 358398
rect 3785 358395 3851 358398
rect 580809 351930 580875 351933
rect 583520 351930 584960 352020
rect 580809 351928 584960 351930
rect 580809 351872 580814 351928
rect 580870 351872 584960 351928
rect 580809 351870 584960 351872
rect 580809 351867 580875 351870
rect 583520 351780 584960 351870
rect 13537 350298 13603 350301
rect 42701 350298 42767 350301
rect 70301 350298 70367 350301
rect 97901 350298 97967 350301
rect 126881 350298 126947 350301
rect 154481 350298 154547 350301
rect 182081 350298 182147 350301
rect 209681 350298 209747 350301
rect 238661 350298 238727 350301
rect 266261 350298 266327 350301
rect 293861 350298 293927 350301
rect 322841 350298 322907 350301
rect 350441 350298 350507 350301
rect 378041 350298 378107 350301
rect 405641 350298 405707 350301
rect 434621 350298 434687 350301
rect 462221 350298 462287 350301
rect 489821 350298 489887 350301
rect 518801 350298 518867 350301
rect 546401 350298 546467 350301
rect 13537 350296 16100 350298
rect 13537 350240 13542 350296
rect 13598 350240 16100 350296
rect 13537 350238 16100 350240
rect 42701 350296 44068 350298
rect 42701 350240 42706 350296
rect 42762 350240 44068 350296
rect 42701 350238 44068 350240
rect 70301 350296 72036 350298
rect 70301 350240 70306 350296
rect 70362 350240 72036 350296
rect 70301 350238 72036 350240
rect 97901 350296 100188 350298
rect 97901 350240 97906 350296
rect 97962 350240 100188 350296
rect 97901 350238 100188 350240
rect 126881 350296 128156 350298
rect 126881 350240 126886 350296
rect 126942 350240 128156 350296
rect 126881 350238 128156 350240
rect 154481 350296 156124 350298
rect 154481 350240 154486 350296
rect 154542 350240 156124 350296
rect 154481 350238 156124 350240
rect 182081 350296 184092 350298
rect 182081 350240 182086 350296
rect 182142 350240 184092 350296
rect 182081 350238 184092 350240
rect 209681 350296 212060 350298
rect 209681 350240 209686 350296
rect 209742 350240 212060 350296
rect 209681 350238 212060 350240
rect 238661 350296 240212 350298
rect 238661 350240 238666 350296
rect 238722 350240 240212 350296
rect 238661 350238 240212 350240
rect 266261 350296 268180 350298
rect 266261 350240 266266 350296
rect 266322 350240 268180 350296
rect 266261 350238 268180 350240
rect 293861 350296 296148 350298
rect 293861 350240 293866 350296
rect 293922 350240 296148 350296
rect 293861 350238 296148 350240
rect 322841 350296 324116 350298
rect 322841 350240 322846 350296
rect 322902 350240 324116 350296
rect 322841 350238 324116 350240
rect 350441 350296 352084 350298
rect 350441 350240 350446 350296
rect 350502 350240 352084 350296
rect 350441 350238 352084 350240
rect 378041 350296 380052 350298
rect 378041 350240 378046 350296
rect 378102 350240 380052 350296
rect 378041 350238 380052 350240
rect 405641 350296 408204 350298
rect 405641 350240 405646 350296
rect 405702 350240 408204 350296
rect 405641 350238 408204 350240
rect 434621 350296 436172 350298
rect 434621 350240 434626 350296
rect 434682 350240 436172 350296
rect 434621 350238 436172 350240
rect 462221 350296 464140 350298
rect 462221 350240 462226 350296
rect 462282 350240 464140 350296
rect 462221 350238 464140 350240
rect 489821 350296 492108 350298
rect 489821 350240 489826 350296
rect 489882 350240 492108 350296
rect 489821 350238 492108 350240
rect 518801 350296 520076 350298
rect 518801 350240 518806 350296
rect 518862 350240 520076 350296
rect 518801 350238 520076 350240
rect 546401 350296 548044 350298
rect 546401 350240 546406 350296
rect 546462 350240 548044 350296
rect 546401 350238 548044 350240
rect 13537 350235 13603 350238
rect 42701 350235 42767 350238
rect 70301 350235 70367 350238
rect 97901 350235 97967 350238
rect 126881 350235 126947 350238
rect 154481 350235 154547 350238
rect 182081 350235 182147 350238
rect 209681 350235 209747 350238
rect 238661 350235 238727 350238
rect 266261 350235 266327 350238
rect 293861 350235 293927 350238
rect 322841 350235 322907 350238
rect 350441 350235 350507 350238
rect 378041 350235 378107 350238
rect 405641 350235 405707 350238
rect 434621 350235 434687 350238
rect 462221 350235 462287 350238
rect 489821 350235 489887 350238
rect 518801 350235 518867 350238
rect 546401 350235 546467 350238
rect 37273 349618 37339 349621
rect 66253 349618 66319 349621
rect 93853 349618 93919 349621
rect 121453 349618 121519 349621
rect 149053 349618 149119 349621
rect 178033 349618 178099 349621
rect 205633 349618 205699 349621
rect 233233 349618 233299 349621
rect 262213 349618 262279 349621
rect 289813 349618 289879 349621
rect 317413 349618 317479 349621
rect 345013 349618 345079 349621
rect 373993 349618 374059 349621
rect 401593 349618 401659 349621
rect 429285 349618 429351 349621
rect 458173 349618 458239 349621
rect 485773 349618 485839 349621
rect 513373 349618 513439 349621
rect 542353 349618 542419 349621
rect 569953 349618 570019 349621
rect 35788 349616 37339 349618
rect 35788 349560 37278 349616
rect 37334 349560 37339 349616
rect 35788 349558 37339 349560
rect 63940 349616 66319 349618
rect 63940 349560 66258 349616
rect 66314 349560 66319 349616
rect 63940 349558 66319 349560
rect 91908 349616 93919 349618
rect 91908 349560 93858 349616
rect 93914 349560 93919 349616
rect 91908 349558 93919 349560
rect 119876 349616 121519 349618
rect 119876 349560 121458 349616
rect 121514 349560 121519 349616
rect 119876 349558 121519 349560
rect 147844 349616 149119 349618
rect 147844 349560 149058 349616
rect 149114 349560 149119 349616
rect 147844 349558 149119 349560
rect 175812 349616 178099 349618
rect 175812 349560 178038 349616
rect 178094 349560 178099 349616
rect 175812 349558 178099 349560
rect 203964 349616 205699 349618
rect 203964 349560 205638 349616
rect 205694 349560 205699 349616
rect 203964 349558 205699 349560
rect 231932 349616 233299 349618
rect 231932 349560 233238 349616
rect 233294 349560 233299 349616
rect 231932 349558 233299 349560
rect 259900 349616 262279 349618
rect 259900 349560 262218 349616
rect 262274 349560 262279 349616
rect 259900 349558 262279 349560
rect 287868 349616 289879 349618
rect 287868 349560 289818 349616
rect 289874 349560 289879 349616
rect 287868 349558 289879 349560
rect 315836 349616 317479 349618
rect 315836 349560 317418 349616
rect 317474 349560 317479 349616
rect 315836 349558 317479 349560
rect 343804 349616 345079 349618
rect 343804 349560 345018 349616
rect 345074 349560 345079 349616
rect 343804 349558 345079 349560
rect 371956 349616 374059 349618
rect 371956 349560 373998 349616
rect 374054 349560 374059 349616
rect 371956 349558 374059 349560
rect 399924 349616 401659 349618
rect 399924 349560 401598 349616
rect 401654 349560 401659 349616
rect 399924 349558 401659 349560
rect 427892 349616 429351 349618
rect 427892 349560 429290 349616
rect 429346 349560 429351 349616
rect 427892 349558 429351 349560
rect 455860 349616 458239 349618
rect 455860 349560 458178 349616
rect 458234 349560 458239 349616
rect 455860 349558 458239 349560
rect 483828 349616 485839 349618
rect 483828 349560 485778 349616
rect 485834 349560 485839 349616
rect 483828 349558 485839 349560
rect 511796 349616 513439 349618
rect 511796 349560 513378 349616
rect 513434 349560 513439 349616
rect 511796 349558 513439 349560
rect 539948 349616 542419 349618
rect 539948 349560 542358 349616
rect 542414 349560 542419 349616
rect 539948 349558 542419 349560
rect 567916 349616 570019 349618
rect 567916 349560 569958 349616
rect 570014 349560 570019 349616
rect 567916 349558 570019 349560
rect 37273 349555 37339 349558
rect 66253 349555 66319 349558
rect 93853 349555 93919 349558
rect 121453 349555 121519 349558
rect 149053 349555 149119 349558
rect 178033 349555 178099 349558
rect 205633 349555 205699 349558
rect 233233 349555 233299 349558
rect 262213 349555 262279 349558
rect 289813 349555 289879 349558
rect 317413 349555 317479 349558
rect 345013 349555 345079 349558
rect 373993 349555 374059 349558
rect 401593 349555 401659 349558
rect 429285 349555 429351 349558
rect 458173 349555 458239 349558
rect 485773 349555 485839 349558
rect 513373 349555 513439 349558
rect 542353 349555 542419 349558
rect 569953 349555 570019 349558
rect -960 345402 480 345492
rect 2773 345402 2839 345405
rect -960 345400 2839 345402
rect -960 345344 2778 345400
rect 2834 345344 2839 345400
rect -960 345342 2839 345344
rect -960 345252 480 345342
rect 2773 345339 2839 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579981 325274 580047 325277
rect 583520 325274 584960 325364
rect 579981 325272 584960 325274
rect 579981 325216 579986 325272
rect 580042 325216 584960 325272
rect 579981 325214 584960 325216
rect 579981 325211 580047 325214
rect 583520 325124 584960 325214
rect 209681 324050 209747 324053
rect 293861 324050 293927 324053
rect 405641 324050 405707 324053
rect 489821 324050 489887 324053
rect 209681 324048 212090 324050
rect 209681 323992 209686 324048
rect 209742 323992 212090 324048
rect 209681 323990 212090 323992
rect 209681 323987 209747 323990
rect 212030 323408 212090 323990
rect 293861 324048 296178 324050
rect 293861 323992 293866 324048
rect 293922 323992 296178 324048
rect 293861 323990 296178 323992
rect 293861 323987 293927 323990
rect 296118 323408 296178 323990
rect 405641 324048 408234 324050
rect 405641 323992 405646 324048
rect 405702 323992 408234 324048
rect 405641 323990 408234 323992
rect 405641 323987 405707 323990
rect 408174 323408 408234 323990
rect 489821 324048 492138 324050
rect 489821 323992 489826 324048
rect 489882 323992 492138 324048
rect 489821 323990 492138 323992
rect 489821 323987 489887 323990
rect 492078 323408 492138 323990
rect 13537 322962 13603 322965
rect 16070 322962 16130 323408
rect 13537 322960 16130 322962
rect 13537 322904 13542 322960
rect 13598 322904 16130 322960
rect 13537 322902 16130 322904
rect 42701 322962 42767 322965
rect 44038 322962 44098 323408
rect 42701 322960 44098 322962
rect 42701 322904 42706 322960
rect 42762 322904 44098 322960
rect 42701 322902 44098 322904
rect 70301 322962 70367 322965
rect 72006 322962 72066 323408
rect 70301 322960 72066 322962
rect 70301 322904 70306 322960
rect 70362 322904 72066 322960
rect 70301 322902 72066 322904
rect 97901 322962 97967 322965
rect 100158 322962 100218 323408
rect 97901 322960 100218 322962
rect 97901 322904 97906 322960
rect 97962 322904 100218 322960
rect 97901 322902 100218 322904
rect 126881 322962 126947 322965
rect 128126 322962 128186 323408
rect 126881 322960 128186 322962
rect 126881 322904 126886 322960
rect 126942 322904 128186 322960
rect 126881 322902 128186 322904
rect 154481 322962 154547 322965
rect 156094 322962 156154 323408
rect 154481 322960 156154 322962
rect 154481 322904 154486 322960
rect 154542 322904 156154 322960
rect 154481 322902 156154 322904
rect 182081 322962 182147 322965
rect 184062 322962 184122 323408
rect 182081 322960 184122 322962
rect 182081 322904 182086 322960
rect 182142 322904 184122 322960
rect 182081 322902 184122 322904
rect 238661 322962 238727 322965
rect 240182 322962 240242 323408
rect 238661 322960 240242 322962
rect 238661 322904 238666 322960
rect 238722 322904 240242 322960
rect 238661 322902 240242 322904
rect 266261 322962 266327 322965
rect 268150 322962 268210 323408
rect 266261 322960 268210 322962
rect 266261 322904 266266 322960
rect 266322 322904 268210 322960
rect 266261 322902 268210 322904
rect 322841 322962 322907 322965
rect 324086 322962 324146 323408
rect 322841 322960 324146 322962
rect 322841 322904 322846 322960
rect 322902 322904 324146 322960
rect 322841 322902 324146 322904
rect 350441 322962 350507 322965
rect 352054 322962 352114 323408
rect 350441 322960 352114 322962
rect 350441 322904 350446 322960
rect 350502 322904 352114 322960
rect 350441 322902 352114 322904
rect 378041 322962 378107 322965
rect 380022 322962 380082 323408
rect 378041 322960 380082 322962
rect 378041 322904 378046 322960
rect 378102 322904 380082 322960
rect 378041 322902 380082 322904
rect 434621 322962 434687 322965
rect 436142 322962 436202 323408
rect 434621 322960 436202 322962
rect 434621 322904 434626 322960
rect 434682 322904 436202 322960
rect 434621 322902 436202 322904
rect 462221 322962 462287 322965
rect 464110 322962 464170 323408
rect 462221 322960 464170 322962
rect 462221 322904 462226 322960
rect 462282 322904 464170 322960
rect 462221 322902 464170 322904
rect 518801 322962 518867 322965
rect 520046 322962 520106 323408
rect 518801 322960 520106 322962
rect 518801 322904 518806 322960
rect 518862 322904 520106 322960
rect 518801 322902 520106 322904
rect 546401 322962 546467 322965
rect 548014 322962 548074 323408
rect 546401 322960 548074 322962
rect 546401 322904 546406 322960
rect 546462 322904 548074 322960
rect 546401 322902 548074 322904
rect 13537 322899 13603 322902
rect 42701 322899 42767 322902
rect 70301 322899 70367 322902
rect 97901 322899 97967 322902
rect 126881 322899 126947 322902
rect 154481 322899 154547 322902
rect 182081 322899 182147 322902
rect 238661 322899 238727 322902
rect 266261 322899 266327 322902
rect 322841 322899 322907 322902
rect 350441 322899 350507 322902
rect 378041 322899 378107 322902
rect 434621 322899 434687 322902
rect 462221 322899 462287 322902
rect 518801 322899 518867 322902
rect 546401 322899 546467 322902
rect 37273 322826 37339 322829
rect 262213 322826 262279 322829
rect 345013 322826 345079 322829
rect 458173 322826 458239 322829
rect 542353 322826 542419 322829
rect 35758 322824 37339 322826
rect 35758 322768 37278 322824
rect 37334 322768 37339 322824
rect 35758 322766 37339 322768
rect 35758 322728 35818 322766
rect 37273 322763 37339 322766
rect 259870 322824 262279 322826
rect 259870 322768 262218 322824
rect 262274 322768 262279 322824
rect 259870 322766 262279 322768
rect 259870 322728 259930 322766
rect 262213 322763 262279 322766
rect 343774 322824 345079 322826
rect 343774 322768 345018 322824
rect 345074 322768 345079 322824
rect 343774 322766 345079 322768
rect 343774 322728 343834 322766
rect 345013 322763 345079 322766
rect 455830 322824 458239 322826
rect 455830 322768 458178 322824
rect 458234 322768 458239 322824
rect 455830 322766 458239 322768
rect 455830 322728 455890 322766
rect 458173 322763 458239 322766
rect 539918 322824 542419 322826
rect 539918 322768 542358 322824
rect 542414 322768 542419 322824
rect 539918 322766 542419 322768
rect 539918 322728 539978 322766
rect 542353 322763 542419 322766
rect 63910 322146 63970 322728
rect 66253 322146 66319 322149
rect 63910 322144 66319 322146
rect 63910 322088 66258 322144
rect 66314 322088 66319 322144
rect 63910 322086 66319 322088
rect 91878 322146 91938 322728
rect 93853 322146 93919 322149
rect 91878 322144 93919 322146
rect 91878 322088 93858 322144
rect 93914 322088 93919 322144
rect 91878 322086 93919 322088
rect 119846 322146 119906 322728
rect 121453 322146 121519 322149
rect 119846 322144 121519 322146
rect 119846 322088 121458 322144
rect 121514 322088 121519 322144
rect 119846 322086 121519 322088
rect 147814 322146 147874 322728
rect 149053 322146 149119 322149
rect 147814 322144 149119 322146
rect 147814 322088 149058 322144
rect 149114 322088 149119 322144
rect 147814 322086 149119 322088
rect 175782 322146 175842 322728
rect 178033 322146 178099 322149
rect 175782 322144 178099 322146
rect 175782 322088 178038 322144
rect 178094 322088 178099 322144
rect 175782 322086 178099 322088
rect 203934 322146 203994 322728
rect 205633 322146 205699 322149
rect 203934 322144 205699 322146
rect 203934 322088 205638 322144
rect 205694 322088 205699 322144
rect 203934 322086 205699 322088
rect 231902 322146 231962 322728
rect 233233 322146 233299 322149
rect 231902 322144 233299 322146
rect 231902 322088 233238 322144
rect 233294 322088 233299 322144
rect 231902 322086 233299 322088
rect 287838 322146 287898 322728
rect 289813 322146 289879 322149
rect 287838 322144 289879 322146
rect 287838 322088 289818 322144
rect 289874 322088 289879 322144
rect 287838 322086 289879 322088
rect 315806 322146 315866 322728
rect 317413 322146 317479 322149
rect 315806 322144 317479 322146
rect 315806 322088 317418 322144
rect 317474 322088 317479 322144
rect 315806 322086 317479 322088
rect 371926 322146 371986 322728
rect 373993 322146 374059 322149
rect 371926 322144 374059 322146
rect 371926 322088 373998 322144
rect 374054 322088 374059 322144
rect 371926 322086 374059 322088
rect 399894 322146 399954 322728
rect 401593 322146 401659 322149
rect 399894 322144 401659 322146
rect 399894 322088 401598 322144
rect 401654 322088 401659 322144
rect 399894 322086 401659 322088
rect 427862 322146 427922 322728
rect 429285 322146 429351 322149
rect 427862 322144 429351 322146
rect 427862 322088 429290 322144
rect 429346 322088 429351 322144
rect 427862 322086 429351 322088
rect 483798 322146 483858 322728
rect 485773 322146 485839 322149
rect 483798 322144 485839 322146
rect 483798 322088 485778 322144
rect 485834 322088 485839 322144
rect 483798 322086 485839 322088
rect 511766 322146 511826 322728
rect 513373 322146 513439 322149
rect 511766 322144 513439 322146
rect 511766 322088 513378 322144
rect 513434 322088 513439 322144
rect 511766 322086 513439 322088
rect 567886 322146 567946 322728
rect 569953 322146 570019 322149
rect 567886 322144 570019 322146
rect 567886 322088 569958 322144
rect 570014 322088 570019 322144
rect 567886 322086 570019 322088
rect 66253 322083 66319 322086
rect 93853 322083 93919 322086
rect 121453 322083 121519 322086
rect 149053 322083 149119 322086
rect 178033 322083 178099 322086
rect 205633 322083 205699 322086
rect 233233 322083 233299 322086
rect 289813 322083 289879 322086
rect 317413 322083 317479 322086
rect 373993 322083 374059 322086
rect 401593 322083 401659 322086
rect 429285 322083 429351 322086
rect 485773 322083 485839 322086
rect 513373 322083 513439 322086
rect 569953 322083 570019 322086
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306234 480 306324
rect 3877 306234 3943 306237
rect -960 306232 3943 306234
rect -960 306176 3882 306232
rect 3938 306176 3943 306232
rect -960 306174 3943 306176
rect -960 306084 480 306174
rect 3877 306171 3943 306174
rect 583520 298604 584960 298844
rect 13537 296306 13603 296309
rect 42701 296306 42767 296309
rect 70301 296306 70367 296309
rect 97901 296306 97967 296309
rect 126881 296306 126947 296309
rect 154481 296306 154547 296309
rect 182081 296306 182147 296309
rect 209681 296306 209747 296309
rect 238661 296306 238727 296309
rect 266261 296306 266327 296309
rect 293861 296306 293927 296309
rect 322841 296306 322907 296309
rect 350441 296306 350507 296309
rect 378041 296306 378107 296309
rect 405641 296306 405707 296309
rect 434621 296306 434687 296309
rect 462221 296306 462287 296309
rect 489821 296306 489887 296309
rect 518801 296306 518867 296309
rect 546401 296306 546467 296309
rect 13537 296304 16100 296306
rect 13537 296248 13542 296304
rect 13598 296248 16100 296304
rect 13537 296246 16100 296248
rect 42701 296304 44068 296306
rect 42701 296248 42706 296304
rect 42762 296248 44068 296304
rect 42701 296246 44068 296248
rect 70301 296304 72036 296306
rect 70301 296248 70306 296304
rect 70362 296248 72036 296304
rect 70301 296246 72036 296248
rect 97901 296304 100188 296306
rect 97901 296248 97906 296304
rect 97962 296248 100188 296304
rect 97901 296246 100188 296248
rect 126881 296304 128156 296306
rect 126881 296248 126886 296304
rect 126942 296248 128156 296304
rect 126881 296246 128156 296248
rect 154481 296304 156124 296306
rect 154481 296248 154486 296304
rect 154542 296248 156124 296304
rect 154481 296246 156124 296248
rect 182081 296304 184092 296306
rect 182081 296248 182086 296304
rect 182142 296248 184092 296304
rect 182081 296246 184092 296248
rect 209681 296304 212060 296306
rect 209681 296248 209686 296304
rect 209742 296248 212060 296304
rect 209681 296246 212060 296248
rect 238661 296304 240212 296306
rect 238661 296248 238666 296304
rect 238722 296248 240212 296304
rect 238661 296246 240212 296248
rect 266261 296304 268180 296306
rect 266261 296248 266266 296304
rect 266322 296248 268180 296304
rect 266261 296246 268180 296248
rect 293861 296304 296148 296306
rect 293861 296248 293866 296304
rect 293922 296248 296148 296304
rect 293861 296246 296148 296248
rect 322841 296304 324116 296306
rect 322841 296248 322846 296304
rect 322902 296248 324116 296304
rect 322841 296246 324116 296248
rect 350441 296304 352084 296306
rect 350441 296248 350446 296304
rect 350502 296248 352084 296304
rect 350441 296246 352084 296248
rect 378041 296304 380052 296306
rect 378041 296248 378046 296304
rect 378102 296248 380052 296304
rect 378041 296246 380052 296248
rect 405641 296304 408204 296306
rect 405641 296248 405646 296304
rect 405702 296248 408204 296304
rect 405641 296246 408204 296248
rect 434621 296304 436172 296306
rect 434621 296248 434626 296304
rect 434682 296248 436172 296304
rect 434621 296246 436172 296248
rect 462221 296304 464140 296306
rect 462221 296248 462226 296304
rect 462282 296248 464140 296304
rect 462221 296246 464140 296248
rect 489821 296304 492108 296306
rect 489821 296248 489826 296304
rect 489882 296248 492108 296304
rect 489821 296246 492108 296248
rect 518801 296304 520076 296306
rect 518801 296248 518806 296304
rect 518862 296248 520076 296304
rect 518801 296246 520076 296248
rect 546401 296304 548044 296306
rect 546401 296248 546406 296304
rect 546462 296248 548044 296304
rect 546401 296246 548044 296248
rect 13537 296243 13603 296246
rect 42701 296243 42767 296246
rect 70301 296243 70367 296246
rect 97901 296243 97967 296246
rect 126881 296243 126947 296246
rect 154481 296243 154547 296246
rect 182081 296243 182147 296246
rect 209681 296243 209747 296246
rect 238661 296243 238727 296246
rect 266261 296243 266327 296246
rect 293861 296243 293927 296246
rect 322841 296243 322907 296246
rect 350441 296243 350507 296246
rect 378041 296243 378107 296246
rect 405641 296243 405707 296246
rect 434621 296243 434687 296246
rect 462221 296243 462287 296246
rect 489821 296243 489887 296246
rect 518801 296243 518867 296246
rect 546401 296243 546467 296246
rect 37273 295626 37339 295629
rect 66253 295626 66319 295629
rect 93853 295626 93919 295629
rect 121453 295626 121519 295629
rect 149053 295626 149119 295629
rect 178033 295626 178099 295629
rect 205633 295626 205699 295629
rect 233233 295626 233299 295629
rect 262213 295626 262279 295629
rect 289813 295626 289879 295629
rect 317413 295626 317479 295629
rect 345013 295626 345079 295629
rect 373993 295626 374059 295629
rect 401593 295626 401659 295629
rect 429285 295626 429351 295629
rect 458173 295626 458239 295629
rect 485773 295626 485839 295629
rect 513373 295626 513439 295629
rect 542353 295626 542419 295629
rect 569953 295626 570019 295629
rect 35788 295624 37339 295626
rect 35788 295568 37278 295624
rect 37334 295568 37339 295624
rect 35788 295566 37339 295568
rect 63940 295624 66319 295626
rect 63940 295568 66258 295624
rect 66314 295568 66319 295624
rect 63940 295566 66319 295568
rect 91908 295624 93919 295626
rect 91908 295568 93858 295624
rect 93914 295568 93919 295624
rect 91908 295566 93919 295568
rect 119876 295624 121519 295626
rect 119876 295568 121458 295624
rect 121514 295568 121519 295624
rect 119876 295566 121519 295568
rect 147844 295624 149119 295626
rect 147844 295568 149058 295624
rect 149114 295568 149119 295624
rect 147844 295566 149119 295568
rect 175812 295624 178099 295626
rect 175812 295568 178038 295624
rect 178094 295568 178099 295624
rect 175812 295566 178099 295568
rect 203964 295624 205699 295626
rect 203964 295568 205638 295624
rect 205694 295568 205699 295624
rect 203964 295566 205699 295568
rect 231932 295624 233299 295626
rect 231932 295568 233238 295624
rect 233294 295568 233299 295624
rect 231932 295566 233299 295568
rect 259900 295624 262279 295626
rect 259900 295568 262218 295624
rect 262274 295568 262279 295624
rect 259900 295566 262279 295568
rect 287868 295624 289879 295626
rect 287868 295568 289818 295624
rect 289874 295568 289879 295624
rect 287868 295566 289879 295568
rect 315836 295624 317479 295626
rect 315836 295568 317418 295624
rect 317474 295568 317479 295624
rect 315836 295566 317479 295568
rect 343804 295624 345079 295626
rect 343804 295568 345018 295624
rect 345074 295568 345079 295624
rect 343804 295566 345079 295568
rect 371956 295624 374059 295626
rect 371956 295568 373998 295624
rect 374054 295568 374059 295624
rect 371956 295566 374059 295568
rect 399924 295624 401659 295626
rect 399924 295568 401598 295624
rect 401654 295568 401659 295624
rect 399924 295566 401659 295568
rect 427892 295624 429351 295626
rect 427892 295568 429290 295624
rect 429346 295568 429351 295624
rect 427892 295566 429351 295568
rect 455860 295624 458239 295626
rect 455860 295568 458178 295624
rect 458234 295568 458239 295624
rect 455860 295566 458239 295568
rect 483828 295624 485839 295626
rect 483828 295568 485778 295624
rect 485834 295568 485839 295624
rect 483828 295566 485839 295568
rect 511796 295624 513439 295626
rect 511796 295568 513378 295624
rect 513434 295568 513439 295624
rect 511796 295566 513439 295568
rect 539948 295624 542419 295626
rect 539948 295568 542358 295624
rect 542414 295568 542419 295624
rect 539948 295566 542419 295568
rect 567916 295624 570019 295626
rect 567916 295568 569958 295624
rect 570014 295568 570019 295624
rect 567916 295566 570019 295568
rect 37273 295563 37339 295566
rect 66253 295563 66319 295566
rect 93853 295563 93919 295566
rect 121453 295563 121519 295566
rect 149053 295563 149119 295566
rect 178033 295563 178099 295566
rect 205633 295563 205699 295566
rect 233233 295563 233299 295566
rect 262213 295563 262279 295566
rect 289813 295563 289879 295566
rect 317413 295563 317479 295566
rect 345013 295563 345079 295566
rect 373993 295563 374059 295566
rect 401593 295563 401659 295566
rect 429285 295563 429351 295566
rect 458173 295563 458239 295566
rect 485773 295563 485839 295566
rect 513373 295563 513439 295566
rect 542353 295563 542419 295566
rect 569953 295563 570019 295566
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 578877 272234 578943 272237
rect 583520 272234 584960 272324
rect 578877 272232 584960 272234
rect 578877 272176 578882 272232
rect 578938 272176 584960 272232
rect 578877 272174 584960 272176
rect 578877 272171 578943 272174
rect 583520 272084 584960 272174
rect 13537 270058 13603 270061
rect 42701 270058 42767 270061
rect 70301 270058 70367 270061
rect 97901 270058 97967 270061
rect 126881 270058 126947 270061
rect 154481 270058 154547 270061
rect 182081 270058 182147 270061
rect 293861 270058 293927 270061
rect 322841 270058 322907 270061
rect 350441 270058 350507 270061
rect 378041 270058 378107 270061
rect 405641 270058 405707 270061
rect 434621 270058 434687 270061
rect 462221 270058 462287 270061
rect 13537 270056 16130 270058
rect 13537 270000 13542 270056
rect 13598 270000 16130 270056
rect 13537 269998 16130 270000
rect 13537 269995 13603 269998
rect 16070 269416 16130 269998
rect 42701 270056 44098 270058
rect 42701 270000 42706 270056
rect 42762 270000 44098 270056
rect 42701 269998 44098 270000
rect 42701 269995 42767 269998
rect 44038 269416 44098 269998
rect 70301 270056 72066 270058
rect 70301 270000 70306 270056
rect 70362 270000 72066 270056
rect 70301 269998 72066 270000
rect 70301 269995 70367 269998
rect 72006 269416 72066 269998
rect 97901 270056 100218 270058
rect 97901 270000 97906 270056
rect 97962 270000 100218 270056
rect 97901 269998 100218 270000
rect 97901 269995 97967 269998
rect 100158 269416 100218 269998
rect 126881 270056 128186 270058
rect 126881 270000 126886 270056
rect 126942 270000 128186 270056
rect 126881 269998 128186 270000
rect 126881 269995 126947 269998
rect 128126 269416 128186 269998
rect 154481 270056 156154 270058
rect 154481 270000 154486 270056
rect 154542 270000 156154 270056
rect 154481 269998 156154 270000
rect 154481 269995 154547 269998
rect 156094 269416 156154 269998
rect 182081 270056 184122 270058
rect 182081 270000 182086 270056
rect 182142 270000 184122 270056
rect 182081 269998 184122 270000
rect 182081 269995 182147 269998
rect 184062 269416 184122 269998
rect 293861 270056 296178 270058
rect 293861 270000 293866 270056
rect 293922 270000 296178 270056
rect 293861 269998 296178 270000
rect 293861 269995 293927 269998
rect 209681 269922 209747 269925
rect 238661 269922 238727 269925
rect 266261 269922 266327 269925
rect 209681 269920 212090 269922
rect 209681 269864 209686 269920
rect 209742 269864 212090 269920
rect 209681 269862 212090 269864
rect 209681 269859 209747 269862
rect 212030 269416 212090 269862
rect 238661 269920 240242 269922
rect 238661 269864 238666 269920
rect 238722 269864 240242 269920
rect 238661 269862 240242 269864
rect 238661 269859 238727 269862
rect 240182 269416 240242 269862
rect 266261 269920 268210 269922
rect 266261 269864 266266 269920
rect 266322 269864 268210 269920
rect 266261 269862 268210 269864
rect 266261 269859 266327 269862
rect 268150 269416 268210 269862
rect 296118 269416 296178 269998
rect 322841 270056 324146 270058
rect 322841 270000 322846 270056
rect 322902 270000 324146 270056
rect 322841 269998 324146 270000
rect 322841 269995 322907 269998
rect 324086 269416 324146 269998
rect 350441 270056 352114 270058
rect 350441 270000 350446 270056
rect 350502 270000 352114 270056
rect 350441 269998 352114 270000
rect 350441 269995 350507 269998
rect 352054 269416 352114 269998
rect 378041 270056 380082 270058
rect 378041 270000 378046 270056
rect 378102 270000 380082 270056
rect 378041 269998 380082 270000
rect 378041 269995 378107 269998
rect 380022 269416 380082 269998
rect 405641 270056 408234 270058
rect 405641 270000 405646 270056
rect 405702 270000 408234 270056
rect 405641 269998 408234 270000
rect 405641 269995 405707 269998
rect 408174 269416 408234 269998
rect 434621 270056 436202 270058
rect 434621 270000 434626 270056
rect 434682 270000 436202 270056
rect 434621 269998 436202 270000
rect 434621 269995 434687 269998
rect 436142 269416 436202 269998
rect 462221 270056 464170 270058
rect 462221 270000 462226 270056
rect 462282 270000 464170 270056
rect 462221 269998 464170 270000
rect 462221 269995 462287 269998
rect 464110 269416 464170 269998
rect 489821 269922 489887 269925
rect 518801 269922 518867 269925
rect 489821 269920 492138 269922
rect 489821 269864 489826 269920
rect 489882 269864 492138 269920
rect 489821 269862 492138 269864
rect 489821 269859 489887 269862
rect 492078 269416 492138 269862
rect 518801 269920 520106 269922
rect 518801 269864 518806 269920
rect 518862 269864 520106 269920
rect 518801 269862 520106 269864
rect 518801 269859 518867 269862
rect 520046 269416 520106 269862
rect 546401 269242 546467 269245
rect 548014 269242 548074 269416
rect 546401 269240 548074 269242
rect 546401 269184 546406 269240
rect 546462 269184 548074 269240
rect 546401 269182 548074 269184
rect 546401 269179 546467 269182
rect 37273 269106 37339 269109
rect 66253 269106 66319 269109
rect 93853 269106 93919 269109
rect 121453 269106 121519 269109
rect 149053 269106 149119 269109
rect 178033 269106 178099 269109
rect 205633 269106 205699 269109
rect 233233 269106 233299 269109
rect 262213 269106 262279 269109
rect 289813 269106 289879 269109
rect 317413 269106 317479 269109
rect 345013 269106 345079 269109
rect 373993 269106 374059 269109
rect 401593 269106 401659 269109
rect 429285 269106 429351 269109
rect 458173 269106 458239 269109
rect 485773 269106 485839 269109
rect 513373 269106 513439 269109
rect 542353 269106 542419 269109
rect 569953 269106 570019 269109
rect 35758 269104 37339 269106
rect 35758 269048 37278 269104
rect 37334 269048 37339 269104
rect 35758 269046 37339 269048
rect 35758 268736 35818 269046
rect 37273 269043 37339 269046
rect 63910 269104 66319 269106
rect 63910 269048 66258 269104
rect 66314 269048 66319 269104
rect 63910 269046 66319 269048
rect 63910 268736 63970 269046
rect 66253 269043 66319 269046
rect 91878 269104 93919 269106
rect 91878 269048 93858 269104
rect 93914 269048 93919 269104
rect 91878 269046 93919 269048
rect 91878 268736 91938 269046
rect 93853 269043 93919 269046
rect 119846 269104 121519 269106
rect 119846 269048 121458 269104
rect 121514 269048 121519 269104
rect 119846 269046 121519 269048
rect 119846 268736 119906 269046
rect 121453 269043 121519 269046
rect 147814 269104 149119 269106
rect 147814 269048 149058 269104
rect 149114 269048 149119 269104
rect 147814 269046 149119 269048
rect 147814 268736 147874 269046
rect 149053 269043 149119 269046
rect 175782 269104 178099 269106
rect 175782 269048 178038 269104
rect 178094 269048 178099 269104
rect 175782 269046 178099 269048
rect 175782 268736 175842 269046
rect 178033 269043 178099 269046
rect 203934 269104 205699 269106
rect 203934 269048 205638 269104
rect 205694 269048 205699 269104
rect 203934 269046 205699 269048
rect 203934 268736 203994 269046
rect 205633 269043 205699 269046
rect 231902 269104 233299 269106
rect 231902 269048 233238 269104
rect 233294 269048 233299 269104
rect 231902 269046 233299 269048
rect 231902 268736 231962 269046
rect 233233 269043 233299 269046
rect 259870 269104 262279 269106
rect 259870 269048 262218 269104
rect 262274 269048 262279 269104
rect 259870 269046 262279 269048
rect 259870 268736 259930 269046
rect 262213 269043 262279 269046
rect 287838 269104 289879 269106
rect 287838 269048 289818 269104
rect 289874 269048 289879 269104
rect 287838 269046 289879 269048
rect 287838 268736 287898 269046
rect 289813 269043 289879 269046
rect 315806 269104 317479 269106
rect 315806 269048 317418 269104
rect 317474 269048 317479 269104
rect 315806 269046 317479 269048
rect 315806 268736 315866 269046
rect 317413 269043 317479 269046
rect 343774 269104 345079 269106
rect 343774 269048 345018 269104
rect 345074 269048 345079 269104
rect 343774 269046 345079 269048
rect 343774 268736 343834 269046
rect 345013 269043 345079 269046
rect 371926 269104 374059 269106
rect 371926 269048 373998 269104
rect 374054 269048 374059 269104
rect 371926 269046 374059 269048
rect 371926 268736 371986 269046
rect 373993 269043 374059 269046
rect 399894 269104 401659 269106
rect 399894 269048 401598 269104
rect 401654 269048 401659 269104
rect 399894 269046 401659 269048
rect 399894 268736 399954 269046
rect 401593 269043 401659 269046
rect 427862 269104 429351 269106
rect 427862 269048 429290 269104
rect 429346 269048 429351 269104
rect 427862 269046 429351 269048
rect 427862 268736 427922 269046
rect 429285 269043 429351 269046
rect 455830 269104 458239 269106
rect 455830 269048 458178 269104
rect 458234 269048 458239 269104
rect 455830 269046 458239 269048
rect 455830 268736 455890 269046
rect 458173 269043 458239 269046
rect 483798 269104 485839 269106
rect 483798 269048 485778 269104
rect 485834 269048 485839 269104
rect 483798 269046 485839 269048
rect 483798 268736 483858 269046
rect 485773 269043 485839 269046
rect 511766 269104 513439 269106
rect 511766 269048 513378 269104
rect 513434 269048 513439 269104
rect 511766 269046 513439 269048
rect 511766 268736 511826 269046
rect 513373 269043 513439 269046
rect 539918 269104 542419 269106
rect 539918 269048 542358 269104
rect 542414 269048 542419 269104
rect 539918 269046 542419 269048
rect 539918 268736 539978 269046
rect 542353 269043 542419 269046
rect 567886 269104 570019 269106
rect 567886 269048 569958 269104
rect 570014 269048 570019 269104
rect 567886 269046 570019 269048
rect 567886 268736 567946 269046
rect 569953 269043 570019 269046
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 254146 480 254236
rect 2773 254146 2839 254149
rect -960 254144 2839 254146
rect -960 254088 2778 254144
rect 2834 254088 2839 254144
rect -960 254086 2839 254088
rect -960 253996 480 254086
rect 2773 254083 2839 254086
rect 583520 245428 584960 245668
rect 13537 242314 13603 242317
rect 42701 242314 42767 242317
rect 70301 242314 70367 242317
rect 97901 242314 97967 242317
rect 126881 242314 126947 242317
rect 154481 242314 154547 242317
rect 182081 242314 182147 242317
rect 209681 242314 209747 242317
rect 238661 242314 238727 242317
rect 266261 242314 266327 242317
rect 293861 242314 293927 242317
rect 322841 242314 322907 242317
rect 350441 242314 350507 242317
rect 378041 242314 378107 242317
rect 405641 242314 405707 242317
rect 434621 242314 434687 242317
rect 462221 242314 462287 242317
rect 489821 242314 489887 242317
rect 518801 242314 518867 242317
rect 546401 242314 546467 242317
rect 13537 242312 16100 242314
rect 13537 242256 13542 242312
rect 13598 242256 16100 242312
rect 13537 242254 16100 242256
rect 42701 242312 44068 242314
rect 42701 242256 42706 242312
rect 42762 242256 44068 242312
rect 42701 242254 44068 242256
rect 70301 242312 72036 242314
rect 70301 242256 70306 242312
rect 70362 242256 72036 242312
rect 70301 242254 72036 242256
rect 97901 242312 100188 242314
rect 97901 242256 97906 242312
rect 97962 242256 100188 242312
rect 97901 242254 100188 242256
rect 126881 242312 128156 242314
rect 126881 242256 126886 242312
rect 126942 242256 128156 242312
rect 126881 242254 128156 242256
rect 154481 242312 156124 242314
rect 154481 242256 154486 242312
rect 154542 242256 156124 242312
rect 154481 242254 156124 242256
rect 182081 242312 184092 242314
rect 182081 242256 182086 242312
rect 182142 242256 184092 242312
rect 182081 242254 184092 242256
rect 209681 242312 212060 242314
rect 209681 242256 209686 242312
rect 209742 242256 212060 242312
rect 209681 242254 212060 242256
rect 238661 242312 240212 242314
rect 238661 242256 238666 242312
rect 238722 242256 240212 242312
rect 238661 242254 240212 242256
rect 266261 242312 268180 242314
rect 266261 242256 266266 242312
rect 266322 242256 268180 242312
rect 266261 242254 268180 242256
rect 293861 242312 296148 242314
rect 293861 242256 293866 242312
rect 293922 242256 296148 242312
rect 293861 242254 296148 242256
rect 322841 242312 324116 242314
rect 322841 242256 322846 242312
rect 322902 242256 324116 242312
rect 322841 242254 324116 242256
rect 350441 242312 352084 242314
rect 350441 242256 350446 242312
rect 350502 242256 352084 242312
rect 350441 242254 352084 242256
rect 378041 242312 380052 242314
rect 378041 242256 378046 242312
rect 378102 242256 380052 242312
rect 378041 242254 380052 242256
rect 405641 242312 408204 242314
rect 405641 242256 405646 242312
rect 405702 242256 408204 242312
rect 405641 242254 408204 242256
rect 434621 242312 436172 242314
rect 434621 242256 434626 242312
rect 434682 242256 436172 242312
rect 434621 242254 436172 242256
rect 462221 242312 464140 242314
rect 462221 242256 462226 242312
rect 462282 242256 464140 242312
rect 462221 242254 464140 242256
rect 489821 242312 492108 242314
rect 489821 242256 489826 242312
rect 489882 242256 492108 242312
rect 489821 242254 492108 242256
rect 518801 242312 520076 242314
rect 518801 242256 518806 242312
rect 518862 242256 520076 242312
rect 518801 242254 520076 242256
rect 546401 242312 548044 242314
rect 546401 242256 546406 242312
rect 546462 242256 548044 242312
rect 546401 242254 548044 242256
rect 13537 242251 13603 242254
rect 42701 242251 42767 242254
rect 70301 242251 70367 242254
rect 97901 242251 97967 242254
rect 126881 242251 126947 242254
rect 154481 242251 154547 242254
rect 182081 242251 182147 242254
rect 209681 242251 209747 242254
rect 238661 242251 238727 242254
rect 266261 242251 266327 242254
rect 293861 242251 293927 242254
rect 322841 242251 322907 242254
rect 350441 242251 350507 242254
rect 378041 242251 378107 242254
rect 405641 242251 405707 242254
rect 434621 242251 434687 242254
rect 462221 242251 462287 242254
rect 489821 242251 489887 242254
rect 518801 242251 518867 242254
rect 546401 242251 546467 242254
rect 37273 241634 37339 241637
rect 66253 241634 66319 241637
rect 93853 241634 93919 241637
rect 121453 241634 121519 241637
rect 149053 241634 149119 241637
rect 178033 241634 178099 241637
rect 205633 241634 205699 241637
rect 233233 241634 233299 241637
rect 262213 241634 262279 241637
rect 289813 241634 289879 241637
rect 317413 241634 317479 241637
rect 345013 241634 345079 241637
rect 373993 241634 374059 241637
rect 401593 241634 401659 241637
rect 429285 241634 429351 241637
rect 458173 241634 458239 241637
rect 485773 241634 485839 241637
rect 513373 241634 513439 241637
rect 542353 241634 542419 241637
rect 569953 241634 570019 241637
rect 35788 241632 37339 241634
rect 35788 241576 37278 241632
rect 37334 241576 37339 241632
rect 35788 241574 37339 241576
rect 63940 241632 66319 241634
rect 63940 241576 66258 241632
rect 66314 241576 66319 241632
rect 63940 241574 66319 241576
rect 91908 241632 93919 241634
rect 91908 241576 93858 241632
rect 93914 241576 93919 241632
rect 91908 241574 93919 241576
rect 119876 241632 121519 241634
rect 119876 241576 121458 241632
rect 121514 241576 121519 241632
rect 119876 241574 121519 241576
rect 147844 241632 149119 241634
rect 147844 241576 149058 241632
rect 149114 241576 149119 241632
rect 147844 241574 149119 241576
rect 175812 241632 178099 241634
rect 175812 241576 178038 241632
rect 178094 241576 178099 241632
rect 175812 241574 178099 241576
rect 203964 241632 205699 241634
rect 203964 241576 205638 241632
rect 205694 241576 205699 241632
rect 203964 241574 205699 241576
rect 231932 241632 233299 241634
rect 231932 241576 233238 241632
rect 233294 241576 233299 241632
rect 231932 241574 233299 241576
rect 259900 241632 262279 241634
rect 259900 241576 262218 241632
rect 262274 241576 262279 241632
rect 259900 241574 262279 241576
rect 287868 241632 289879 241634
rect 287868 241576 289818 241632
rect 289874 241576 289879 241632
rect 287868 241574 289879 241576
rect 315836 241632 317479 241634
rect 315836 241576 317418 241632
rect 317474 241576 317479 241632
rect 315836 241574 317479 241576
rect 343804 241632 345079 241634
rect 343804 241576 345018 241632
rect 345074 241576 345079 241632
rect 343804 241574 345079 241576
rect 371956 241632 374059 241634
rect 371956 241576 373998 241632
rect 374054 241576 374059 241632
rect 371956 241574 374059 241576
rect 399924 241632 401659 241634
rect 399924 241576 401598 241632
rect 401654 241576 401659 241632
rect 399924 241574 401659 241576
rect 427892 241632 429351 241634
rect 427892 241576 429290 241632
rect 429346 241576 429351 241632
rect 427892 241574 429351 241576
rect 455860 241632 458239 241634
rect 455860 241576 458178 241632
rect 458234 241576 458239 241632
rect 455860 241574 458239 241576
rect 483828 241632 485839 241634
rect 483828 241576 485778 241632
rect 485834 241576 485839 241632
rect 483828 241574 485839 241576
rect 511796 241632 513439 241634
rect 511796 241576 513378 241632
rect 513434 241576 513439 241632
rect 511796 241574 513439 241576
rect 539948 241632 542419 241634
rect 539948 241576 542358 241632
rect 542414 241576 542419 241632
rect 539948 241574 542419 241576
rect 567916 241632 570019 241634
rect 567916 241576 569958 241632
rect 570014 241576 570019 241632
rect 567916 241574 570019 241576
rect 37273 241571 37339 241574
rect 66253 241571 66319 241574
rect 93853 241571 93919 241574
rect 121453 241571 121519 241574
rect 149053 241571 149119 241574
rect 178033 241571 178099 241574
rect 205633 241571 205699 241574
rect 233233 241571 233299 241574
rect 262213 241571 262279 241574
rect 289813 241571 289879 241574
rect 317413 241571 317479 241574
rect 345013 241571 345079 241574
rect 373993 241571 374059 241574
rect 401593 241571 401659 241574
rect 429285 241571 429351 241574
rect 458173 241571 458239 241574
rect 485773 241571 485839 241574
rect 513373 241571 513439 241574
rect 542353 241571 542419 241574
rect 569953 241571 570019 241574
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 579797 232386 579863 232389
rect 583520 232386 584960 232476
rect 579797 232384 584960 232386
rect 579797 232328 579802 232384
rect 579858 232328 584960 232384
rect 579797 232326 584960 232328
rect 579797 232323 579863 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect 70301 215930 70367 215933
rect 70301 215928 72066 215930
rect 70301 215872 70306 215928
rect 70362 215872 72066 215928
rect 70301 215870 72066 215872
rect 70301 215867 70367 215870
rect 13537 215386 13603 215389
rect 42701 215386 42767 215389
rect 13537 215384 16100 215386
rect 13537 215328 13542 215384
rect 13598 215328 16100 215384
rect 13537 215326 16100 215328
rect 42701 215384 44068 215386
rect 42701 215328 42706 215384
rect 42762 215328 44068 215384
rect 72006 215356 72066 215870
rect 546401 215522 546467 215525
rect 546401 215520 548074 215522
rect 546401 215464 546406 215520
rect 546462 215464 548074 215520
rect 546401 215462 548074 215464
rect 546401 215459 546467 215462
rect 97901 215386 97967 215389
rect 126881 215386 126947 215389
rect 154481 215386 154547 215389
rect 182081 215386 182147 215389
rect 209681 215386 209747 215389
rect 238661 215386 238727 215389
rect 266261 215386 266327 215389
rect 293861 215386 293927 215389
rect 322841 215386 322907 215389
rect 350441 215386 350507 215389
rect 378041 215386 378107 215389
rect 405641 215386 405707 215389
rect 434621 215386 434687 215389
rect 462221 215386 462287 215389
rect 489821 215386 489887 215389
rect 518801 215386 518867 215389
rect 97901 215384 100188 215386
rect 42701 215326 44068 215328
rect 97901 215328 97906 215384
rect 97962 215328 100188 215384
rect 97901 215326 100188 215328
rect 126881 215384 128156 215386
rect 126881 215328 126886 215384
rect 126942 215328 128156 215384
rect 126881 215326 128156 215328
rect 154481 215384 156124 215386
rect 154481 215328 154486 215384
rect 154542 215328 156124 215384
rect 154481 215326 156124 215328
rect 182081 215384 184092 215386
rect 182081 215328 182086 215384
rect 182142 215328 184092 215384
rect 182081 215326 184092 215328
rect 209681 215384 212060 215386
rect 209681 215328 209686 215384
rect 209742 215328 212060 215384
rect 209681 215326 212060 215328
rect 238661 215384 240212 215386
rect 238661 215328 238666 215384
rect 238722 215328 240212 215384
rect 238661 215326 240212 215328
rect 266261 215384 268180 215386
rect 266261 215328 266266 215384
rect 266322 215328 268180 215384
rect 266261 215326 268180 215328
rect 293861 215384 296148 215386
rect 293861 215328 293866 215384
rect 293922 215328 296148 215384
rect 293861 215326 296148 215328
rect 322841 215384 324116 215386
rect 322841 215328 322846 215384
rect 322902 215328 324116 215384
rect 322841 215326 324116 215328
rect 350441 215384 352084 215386
rect 350441 215328 350446 215384
rect 350502 215328 352084 215384
rect 350441 215326 352084 215328
rect 378041 215384 380052 215386
rect 378041 215328 378046 215384
rect 378102 215328 380052 215384
rect 378041 215326 380052 215328
rect 405641 215384 408204 215386
rect 405641 215328 405646 215384
rect 405702 215328 408204 215384
rect 405641 215326 408204 215328
rect 434621 215384 436172 215386
rect 434621 215328 434626 215384
rect 434682 215328 436172 215384
rect 434621 215326 436172 215328
rect 462221 215384 464140 215386
rect 462221 215328 462226 215384
rect 462282 215328 464140 215384
rect 462221 215326 464140 215328
rect 489821 215384 492108 215386
rect 489821 215328 489826 215384
rect 489882 215328 492108 215384
rect 489821 215326 492108 215328
rect 518801 215384 520076 215386
rect 518801 215328 518806 215384
rect 518862 215328 520076 215384
rect 548014 215356 548074 215462
rect 518801 215326 520076 215328
rect 13537 215323 13603 215326
rect 42701 215323 42767 215326
rect 97901 215323 97967 215326
rect 126881 215323 126947 215326
rect 154481 215323 154547 215326
rect 182081 215323 182147 215326
rect 209681 215323 209747 215326
rect 238661 215323 238727 215326
rect 266261 215323 266327 215326
rect 293861 215323 293927 215326
rect 322841 215323 322907 215326
rect 350441 215323 350507 215326
rect 378041 215323 378107 215326
rect 405641 215323 405707 215326
rect 434621 215323 434687 215326
rect 462221 215323 462287 215326
rect 489821 215323 489887 215326
rect 518801 215323 518867 215326
rect 205633 215250 205699 215253
rect 373993 215250 374059 215253
rect 203934 215248 205699 215250
rect 203934 215192 205638 215248
rect 205694 215192 205699 215248
rect 203934 215190 205699 215192
rect -960 214828 480 215068
rect 37273 214706 37339 214709
rect 66253 214706 66319 214709
rect 93853 214706 93919 214709
rect 121453 214706 121519 214709
rect 149053 214706 149119 214709
rect 178033 214706 178099 214709
rect 35788 214704 37339 214706
rect 35788 214648 37278 214704
rect 37334 214648 37339 214704
rect 35788 214646 37339 214648
rect 63940 214704 66319 214706
rect 63940 214648 66258 214704
rect 66314 214648 66319 214704
rect 63940 214646 66319 214648
rect 91908 214704 93919 214706
rect 91908 214648 93858 214704
rect 93914 214648 93919 214704
rect 91908 214646 93919 214648
rect 119876 214704 121519 214706
rect 119876 214648 121458 214704
rect 121514 214648 121519 214704
rect 119876 214646 121519 214648
rect 147844 214704 149119 214706
rect 147844 214648 149058 214704
rect 149114 214648 149119 214704
rect 147844 214646 149119 214648
rect 175812 214704 178099 214706
rect 175812 214648 178038 214704
rect 178094 214648 178099 214704
rect 203934 214676 203994 215190
rect 205633 215187 205699 215190
rect 371926 215248 374059 215250
rect 371926 215192 373998 215248
rect 374054 215192 374059 215248
rect 371926 215190 374059 215192
rect 233233 214706 233299 214709
rect 262213 214706 262279 214709
rect 289813 214706 289879 214709
rect 317413 214706 317479 214709
rect 345013 214706 345079 214709
rect 231932 214704 233299 214706
rect 175812 214646 178099 214648
rect 231932 214648 233238 214704
rect 233294 214648 233299 214704
rect 231932 214646 233299 214648
rect 259900 214704 262279 214706
rect 259900 214648 262218 214704
rect 262274 214648 262279 214704
rect 259900 214646 262279 214648
rect 287868 214704 289879 214706
rect 287868 214648 289818 214704
rect 289874 214648 289879 214704
rect 287868 214646 289879 214648
rect 315836 214704 317479 214706
rect 315836 214648 317418 214704
rect 317474 214648 317479 214704
rect 315836 214646 317479 214648
rect 343804 214704 345079 214706
rect 343804 214648 345018 214704
rect 345074 214648 345079 214704
rect 371926 214676 371986 215190
rect 373993 215187 374059 215190
rect 401593 214706 401659 214709
rect 429285 214706 429351 214709
rect 458173 214706 458239 214709
rect 485773 214706 485839 214709
rect 513373 214706 513439 214709
rect 542353 214706 542419 214709
rect 569953 214706 570019 214709
rect 399924 214704 401659 214706
rect 343804 214646 345079 214648
rect 399924 214648 401598 214704
rect 401654 214648 401659 214704
rect 399924 214646 401659 214648
rect 427892 214704 429351 214706
rect 427892 214648 429290 214704
rect 429346 214648 429351 214704
rect 427892 214646 429351 214648
rect 455860 214704 458239 214706
rect 455860 214648 458178 214704
rect 458234 214648 458239 214704
rect 455860 214646 458239 214648
rect 483828 214704 485839 214706
rect 483828 214648 485778 214704
rect 485834 214648 485839 214704
rect 483828 214646 485839 214648
rect 511796 214704 513439 214706
rect 511796 214648 513378 214704
rect 513434 214648 513439 214704
rect 511796 214646 513439 214648
rect 539948 214704 542419 214706
rect 539948 214648 542358 214704
rect 542414 214648 542419 214704
rect 539948 214646 542419 214648
rect 567916 214704 570019 214706
rect 567916 214648 569958 214704
rect 570014 214648 570019 214704
rect 567916 214646 570019 214648
rect 37273 214643 37339 214646
rect 66253 214643 66319 214646
rect 93853 214643 93919 214646
rect 121453 214643 121519 214646
rect 149053 214643 149119 214646
rect 178033 214643 178099 214646
rect 233233 214643 233299 214646
rect 262213 214643 262279 214646
rect 289813 214643 289879 214646
rect 317413 214643 317479 214646
rect 345013 214643 345079 214646
rect 401593 214643 401659 214646
rect 429285 214643 429351 214646
rect 458173 214643 458239 214646
rect 485773 214643 485839 214646
rect 513373 214643 513439 214646
rect 542353 214643 542419 214646
rect 569953 214643 570019 214646
rect 583520 205580 584960 205820
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 2957 188866 3023 188869
rect -960 188864 3023 188866
rect -960 188808 2962 188864
rect 3018 188808 3023 188864
rect -960 188806 3023 188808
rect -960 188716 480 188806
rect 2957 188803 3023 188806
rect 13537 188322 13603 188325
rect 42701 188322 42767 188325
rect 70301 188322 70367 188325
rect 97901 188322 97967 188325
rect 126881 188322 126947 188325
rect 154481 188322 154547 188325
rect 182081 188322 182147 188325
rect 209681 188322 209747 188325
rect 238661 188322 238727 188325
rect 266261 188322 266327 188325
rect 293861 188322 293927 188325
rect 322841 188322 322907 188325
rect 350441 188322 350507 188325
rect 378041 188322 378107 188325
rect 405641 188322 405707 188325
rect 434621 188322 434687 188325
rect 462221 188322 462287 188325
rect 489821 188322 489887 188325
rect 518801 188322 518867 188325
rect 546401 188322 546467 188325
rect 13537 188320 16100 188322
rect 13537 188264 13542 188320
rect 13598 188264 16100 188320
rect 13537 188262 16100 188264
rect 42701 188320 44068 188322
rect 42701 188264 42706 188320
rect 42762 188264 44068 188320
rect 42701 188262 44068 188264
rect 70301 188320 72036 188322
rect 70301 188264 70306 188320
rect 70362 188264 72036 188320
rect 70301 188262 72036 188264
rect 97901 188320 100188 188322
rect 97901 188264 97906 188320
rect 97962 188264 100188 188320
rect 97901 188262 100188 188264
rect 126881 188320 128156 188322
rect 126881 188264 126886 188320
rect 126942 188264 128156 188320
rect 126881 188262 128156 188264
rect 154481 188320 156124 188322
rect 154481 188264 154486 188320
rect 154542 188264 156124 188320
rect 154481 188262 156124 188264
rect 182081 188320 184092 188322
rect 182081 188264 182086 188320
rect 182142 188264 184092 188320
rect 182081 188262 184092 188264
rect 209681 188320 212060 188322
rect 209681 188264 209686 188320
rect 209742 188264 212060 188320
rect 209681 188262 212060 188264
rect 238661 188320 240212 188322
rect 238661 188264 238666 188320
rect 238722 188264 240212 188320
rect 238661 188262 240212 188264
rect 266261 188320 268180 188322
rect 266261 188264 266266 188320
rect 266322 188264 268180 188320
rect 266261 188262 268180 188264
rect 293861 188320 296148 188322
rect 293861 188264 293866 188320
rect 293922 188264 296148 188320
rect 293861 188262 296148 188264
rect 322841 188320 324116 188322
rect 322841 188264 322846 188320
rect 322902 188264 324116 188320
rect 322841 188262 324116 188264
rect 350441 188320 352084 188322
rect 350441 188264 350446 188320
rect 350502 188264 352084 188320
rect 350441 188262 352084 188264
rect 378041 188320 380052 188322
rect 378041 188264 378046 188320
rect 378102 188264 380052 188320
rect 378041 188262 380052 188264
rect 405641 188320 408204 188322
rect 405641 188264 405646 188320
rect 405702 188264 408204 188320
rect 405641 188262 408204 188264
rect 434621 188320 436172 188322
rect 434621 188264 434626 188320
rect 434682 188264 436172 188320
rect 434621 188262 436172 188264
rect 462221 188320 464140 188322
rect 462221 188264 462226 188320
rect 462282 188264 464140 188320
rect 462221 188262 464140 188264
rect 489821 188320 492108 188322
rect 489821 188264 489826 188320
rect 489882 188264 492108 188320
rect 489821 188262 492108 188264
rect 518801 188320 520076 188322
rect 518801 188264 518806 188320
rect 518862 188264 520076 188320
rect 518801 188262 520076 188264
rect 546401 188320 548044 188322
rect 546401 188264 546406 188320
rect 546462 188264 548044 188320
rect 546401 188262 548044 188264
rect 13537 188259 13603 188262
rect 42701 188259 42767 188262
rect 70301 188259 70367 188262
rect 97901 188259 97967 188262
rect 126881 188259 126947 188262
rect 154481 188259 154547 188262
rect 182081 188259 182147 188262
rect 209681 188259 209747 188262
rect 238661 188259 238727 188262
rect 266261 188259 266327 188262
rect 293861 188259 293927 188262
rect 322841 188259 322907 188262
rect 350441 188259 350507 188262
rect 378041 188259 378107 188262
rect 405641 188259 405707 188262
rect 434621 188259 434687 188262
rect 462221 188259 462287 188262
rect 489821 188259 489887 188262
rect 518801 188259 518867 188262
rect 546401 188259 546467 188262
rect 37273 187642 37339 187645
rect 66253 187642 66319 187645
rect 93853 187642 93919 187645
rect 121453 187642 121519 187645
rect 149053 187642 149119 187645
rect 178033 187642 178099 187645
rect 205633 187642 205699 187645
rect 233233 187642 233299 187645
rect 262213 187642 262279 187645
rect 289813 187642 289879 187645
rect 317413 187642 317479 187645
rect 345013 187642 345079 187645
rect 373993 187642 374059 187645
rect 401593 187642 401659 187645
rect 429285 187642 429351 187645
rect 458173 187642 458239 187645
rect 485773 187642 485839 187645
rect 513373 187642 513439 187645
rect 542353 187642 542419 187645
rect 569953 187642 570019 187645
rect 35788 187640 37339 187642
rect 35788 187584 37278 187640
rect 37334 187584 37339 187640
rect 35788 187582 37339 187584
rect 63940 187640 66319 187642
rect 63940 187584 66258 187640
rect 66314 187584 66319 187640
rect 63940 187582 66319 187584
rect 91908 187640 93919 187642
rect 91908 187584 93858 187640
rect 93914 187584 93919 187640
rect 91908 187582 93919 187584
rect 119876 187640 121519 187642
rect 119876 187584 121458 187640
rect 121514 187584 121519 187640
rect 119876 187582 121519 187584
rect 147844 187640 149119 187642
rect 147844 187584 149058 187640
rect 149114 187584 149119 187640
rect 147844 187582 149119 187584
rect 175812 187640 178099 187642
rect 175812 187584 178038 187640
rect 178094 187584 178099 187640
rect 175812 187582 178099 187584
rect 203964 187640 205699 187642
rect 203964 187584 205638 187640
rect 205694 187584 205699 187640
rect 203964 187582 205699 187584
rect 231932 187640 233299 187642
rect 231932 187584 233238 187640
rect 233294 187584 233299 187640
rect 231932 187582 233299 187584
rect 259900 187640 262279 187642
rect 259900 187584 262218 187640
rect 262274 187584 262279 187640
rect 259900 187582 262279 187584
rect 287868 187640 289879 187642
rect 287868 187584 289818 187640
rect 289874 187584 289879 187640
rect 287868 187582 289879 187584
rect 315836 187640 317479 187642
rect 315836 187584 317418 187640
rect 317474 187584 317479 187640
rect 315836 187582 317479 187584
rect 343804 187640 345079 187642
rect 343804 187584 345018 187640
rect 345074 187584 345079 187640
rect 343804 187582 345079 187584
rect 371956 187640 374059 187642
rect 371956 187584 373998 187640
rect 374054 187584 374059 187640
rect 371956 187582 374059 187584
rect 399924 187640 401659 187642
rect 399924 187584 401598 187640
rect 401654 187584 401659 187640
rect 399924 187582 401659 187584
rect 427892 187640 429351 187642
rect 427892 187584 429290 187640
rect 429346 187584 429351 187640
rect 427892 187582 429351 187584
rect 455860 187640 458239 187642
rect 455860 187584 458178 187640
rect 458234 187584 458239 187640
rect 455860 187582 458239 187584
rect 483828 187640 485839 187642
rect 483828 187584 485778 187640
rect 485834 187584 485839 187640
rect 483828 187582 485839 187584
rect 511796 187640 513439 187642
rect 511796 187584 513378 187640
rect 513434 187584 513439 187640
rect 511796 187582 513439 187584
rect 539948 187640 542419 187642
rect 539948 187584 542358 187640
rect 542414 187584 542419 187640
rect 539948 187582 542419 187584
rect 567916 187640 570019 187642
rect 567916 187584 569958 187640
rect 570014 187584 570019 187640
rect 567916 187582 570019 187584
rect 37273 187579 37339 187582
rect 66253 187579 66319 187582
rect 93853 187579 93919 187582
rect 121453 187579 121519 187582
rect 149053 187579 149119 187582
rect 178033 187579 178099 187582
rect 205633 187579 205699 187582
rect 233233 187579 233299 187582
rect 262213 187579 262279 187582
rect 289813 187579 289879 187582
rect 317413 187579 317479 187582
rect 345013 187579 345079 187582
rect 373993 187579 374059 187582
rect 401593 187579 401659 187582
rect 429285 187579 429351 187582
rect 458173 187579 458239 187582
rect 485773 187579 485839 187582
rect 513373 187579 513439 187582
rect 542353 187579 542419 187582
rect 569953 187579 570019 187582
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 13537 161394 13603 161397
rect 42701 161394 42767 161397
rect 97901 161394 97967 161397
rect 126881 161394 126947 161397
rect 154481 161394 154547 161397
rect 182081 161394 182147 161397
rect 209681 161394 209747 161397
rect 238661 161394 238727 161397
rect 266261 161394 266327 161397
rect 293861 161394 293927 161397
rect 322841 161394 322907 161397
rect 350441 161394 350507 161397
rect 378041 161394 378107 161397
rect 405641 161394 405707 161397
rect 434621 161394 434687 161397
rect 462221 161394 462287 161397
rect 489821 161394 489887 161397
rect 518801 161394 518867 161397
rect 546401 161394 546467 161397
rect 13537 161392 16100 161394
rect 13537 161336 13542 161392
rect 13598 161336 16100 161392
rect 13537 161334 16100 161336
rect 42701 161392 44068 161394
rect 42701 161336 42706 161392
rect 42762 161336 44068 161392
rect 97901 161392 100188 161394
rect 42701 161334 44068 161336
rect 13537 161331 13603 161334
rect 42701 161331 42767 161334
rect 70301 160850 70367 160853
rect 72006 160850 72066 161364
rect 97901 161336 97906 161392
rect 97962 161336 100188 161392
rect 97901 161334 100188 161336
rect 126881 161392 128156 161394
rect 126881 161336 126886 161392
rect 126942 161336 128156 161392
rect 126881 161334 128156 161336
rect 154481 161392 156124 161394
rect 154481 161336 154486 161392
rect 154542 161336 156124 161392
rect 154481 161334 156124 161336
rect 182081 161392 184092 161394
rect 182081 161336 182086 161392
rect 182142 161336 184092 161392
rect 182081 161334 184092 161336
rect 209681 161392 212060 161394
rect 209681 161336 209686 161392
rect 209742 161336 212060 161392
rect 209681 161334 212060 161336
rect 238661 161392 240212 161394
rect 238661 161336 238666 161392
rect 238722 161336 240212 161392
rect 238661 161334 240212 161336
rect 266261 161392 268180 161394
rect 266261 161336 266266 161392
rect 266322 161336 268180 161392
rect 266261 161334 268180 161336
rect 293861 161392 296148 161394
rect 293861 161336 293866 161392
rect 293922 161336 296148 161392
rect 293861 161334 296148 161336
rect 322841 161392 324116 161394
rect 322841 161336 322846 161392
rect 322902 161336 324116 161392
rect 322841 161334 324116 161336
rect 350441 161392 352084 161394
rect 350441 161336 350446 161392
rect 350502 161336 352084 161392
rect 350441 161334 352084 161336
rect 378041 161392 380052 161394
rect 378041 161336 378046 161392
rect 378102 161336 380052 161392
rect 378041 161334 380052 161336
rect 405641 161392 408204 161394
rect 405641 161336 405646 161392
rect 405702 161336 408204 161392
rect 405641 161334 408204 161336
rect 434621 161392 436172 161394
rect 434621 161336 434626 161392
rect 434682 161336 436172 161392
rect 434621 161334 436172 161336
rect 462221 161392 464140 161394
rect 462221 161336 462226 161392
rect 462282 161336 464140 161392
rect 462221 161334 464140 161336
rect 489821 161392 492108 161394
rect 489821 161336 489826 161392
rect 489882 161336 492108 161392
rect 489821 161334 492108 161336
rect 518801 161392 520076 161394
rect 518801 161336 518806 161392
rect 518862 161336 520076 161392
rect 518801 161334 520076 161336
rect 546401 161392 548044 161394
rect 546401 161336 546406 161392
rect 546462 161336 548044 161392
rect 546401 161334 548044 161336
rect 97901 161331 97967 161334
rect 126881 161331 126947 161334
rect 154481 161331 154547 161334
rect 182081 161331 182147 161334
rect 209681 161331 209747 161334
rect 238661 161331 238727 161334
rect 266261 161331 266327 161334
rect 293861 161331 293927 161334
rect 322841 161331 322907 161334
rect 350441 161331 350507 161334
rect 378041 161331 378107 161334
rect 405641 161331 405707 161334
rect 434621 161331 434687 161334
rect 462221 161331 462287 161334
rect 489821 161331 489887 161334
rect 518801 161331 518867 161334
rect 546401 161331 546467 161334
rect 70301 160848 72066 160850
rect 70301 160792 70306 160848
rect 70362 160792 72066 160848
rect 70301 160790 72066 160792
rect 70301 160787 70367 160790
rect 37273 160714 37339 160717
rect 66253 160714 66319 160717
rect 93853 160714 93919 160717
rect 121453 160714 121519 160717
rect 149053 160714 149119 160717
rect 178033 160714 178099 160717
rect 233233 160714 233299 160717
rect 262213 160714 262279 160717
rect 289813 160714 289879 160717
rect 317413 160714 317479 160717
rect 345013 160714 345079 160717
rect 373993 160714 374059 160717
rect 401593 160714 401659 160717
rect 429285 160714 429351 160717
rect 458173 160714 458239 160717
rect 485773 160714 485839 160717
rect 513373 160714 513439 160717
rect 542353 160714 542419 160717
rect 569953 160714 570019 160717
rect 35788 160712 37339 160714
rect 35788 160656 37278 160712
rect 37334 160656 37339 160712
rect 35788 160654 37339 160656
rect 63940 160712 66319 160714
rect 63940 160656 66258 160712
rect 66314 160656 66319 160712
rect 63940 160654 66319 160656
rect 91908 160712 93919 160714
rect 91908 160656 93858 160712
rect 93914 160656 93919 160712
rect 91908 160654 93919 160656
rect 119876 160712 121519 160714
rect 119876 160656 121458 160712
rect 121514 160656 121519 160712
rect 119876 160654 121519 160656
rect 147844 160712 149119 160714
rect 147844 160656 149058 160712
rect 149114 160656 149119 160712
rect 147844 160654 149119 160656
rect 175812 160712 178099 160714
rect 175812 160656 178038 160712
rect 178094 160656 178099 160712
rect 231932 160712 233299 160714
rect 175812 160654 178099 160656
rect 37273 160651 37339 160654
rect 66253 160651 66319 160654
rect 93853 160651 93919 160654
rect 121453 160651 121519 160654
rect 149053 160651 149119 160654
rect 178033 160651 178099 160654
rect 203934 160170 203994 160684
rect 231932 160656 233238 160712
rect 233294 160656 233299 160712
rect 231932 160654 233299 160656
rect 259900 160712 262279 160714
rect 259900 160656 262218 160712
rect 262274 160656 262279 160712
rect 259900 160654 262279 160656
rect 287868 160712 289879 160714
rect 287868 160656 289818 160712
rect 289874 160656 289879 160712
rect 287868 160654 289879 160656
rect 315836 160712 317479 160714
rect 315836 160656 317418 160712
rect 317474 160656 317479 160712
rect 315836 160654 317479 160656
rect 343804 160712 345079 160714
rect 343804 160656 345018 160712
rect 345074 160656 345079 160712
rect 343804 160654 345079 160656
rect 371956 160712 374059 160714
rect 371956 160656 373998 160712
rect 374054 160656 374059 160712
rect 371956 160654 374059 160656
rect 399924 160712 401659 160714
rect 399924 160656 401598 160712
rect 401654 160656 401659 160712
rect 399924 160654 401659 160656
rect 427892 160712 429351 160714
rect 427892 160656 429290 160712
rect 429346 160656 429351 160712
rect 427892 160654 429351 160656
rect 455860 160712 458239 160714
rect 455860 160656 458178 160712
rect 458234 160656 458239 160712
rect 455860 160654 458239 160656
rect 483828 160712 485839 160714
rect 483828 160656 485778 160712
rect 485834 160656 485839 160712
rect 483828 160654 485839 160656
rect 511796 160712 513439 160714
rect 511796 160656 513378 160712
rect 513434 160656 513439 160712
rect 511796 160654 513439 160656
rect 539948 160712 542419 160714
rect 539948 160656 542358 160712
rect 542414 160656 542419 160712
rect 539948 160654 542419 160656
rect 567916 160712 570019 160714
rect 567916 160656 569958 160712
rect 570014 160656 570019 160712
rect 567916 160654 570019 160656
rect 233233 160651 233299 160654
rect 262213 160651 262279 160654
rect 289813 160651 289879 160654
rect 317413 160651 317479 160654
rect 345013 160651 345079 160654
rect 373993 160651 374059 160654
rect 401593 160651 401659 160654
rect 429285 160651 429351 160654
rect 458173 160651 458239 160654
rect 485773 160651 485839 160654
rect 513373 160651 513439 160654
rect 542353 160651 542419 160654
rect 569953 160651 570019 160654
rect 205633 160170 205699 160173
rect 203934 160168 205699 160170
rect 203934 160112 205638 160168
rect 205694 160112 205699 160168
rect 203934 160110 205699 160112
rect 205633 160107 205699 160110
rect 580901 152690 580967 152693
rect 583520 152690 584960 152780
rect 580901 152688 584960 152690
rect 580901 152632 580906 152688
rect 580962 152632 584960 152688
rect 580901 152630 584960 152632
rect 580901 152627 580967 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3969 149834 4035 149837
rect -960 149832 4035 149834
rect -960 149776 3974 149832
rect 4030 149776 4035 149832
rect -960 149774 4035 149776
rect -960 149684 480 149774
rect 3969 149771 4035 149774
rect 583520 139212 584960 139452
rect -960 136778 480 136868
rect 3325 136778 3391 136781
rect -960 136776 3391 136778
rect -960 136720 3330 136776
rect 3386 136720 3391 136776
rect -960 136718 3391 136720
rect -960 136628 480 136718
rect 3325 136715 3391 136718
rect 13537 134330 13603 134333
rect 42701 134330 42767 134333
rect 70301 134330 70367 134333
rect 97901 134330 97967 134333
rect 126881 134330 126947 134333
rect 154481 134330 154547 134333
rect 182081 134330 182147 134333
rect 209681 134330 209747 134333
rect 238661 134330 238727 134333
rect 266261 134330 266327 134333
rect 293861 134330 293927 134333
rect 322841 134330 322907 134333
rect 350441 134330 350507 134333
rect 378041 134330 378107 134333
rect 405641 134330 405707 134333
rect 434621 134330 434687 134333
rect 462221 134330 462287 134333
rect 489821 134330 489887 134333
rect 518801 134330 518867 134333
rect 546401 134330 546467 134333
rect 13537 134328 16100 134330
rect 13537 134272 13542 134328
rect 13598 134272 16100 134328
rect 13537 134270 16100 134272
rect 42701 134328 44068 134330
rect 42701 134272 42706 134328
rect 42762 134272 44068 134328
rect 42701 134270 44068 134272
rect 70301 134328 72036 134330
rect 70301 134272 70306 134328
rect 70362 134272 72036 134328
rect 70301 134270 72036 134272
rect 97901 134328 100188 134330
rect 97901 134272 97906 134328
rect 97962 134272 100188 134328
rect 97901 134270 100188 134272
rect 126881 134328 128156 134330
rect 126881 134272 126886 134328
rect 126942 134272 128156 134328
rect 126881 134270 128156 134272
rect 154481 134328 156124 134330
rect 154481 134272 154486 134328
rect 154542 134272 156124 134328
rect 154481 134270 156124 134272
rect 182081 134328 184092 134330
rect 182081 134272 182086 134328
rect 182142 134272 184092 134328
rect 182081 134270 184092 134272
rect 209681 134328 212060 134330
rect 209681 134272 209686 134328
rect 209742 134272 212060 134328
rect 209681 134270 212060 134272
rect 238661 134328 240212 134330
rect 238661 134272 238666 134328
rect 238722 134272 240212 134328
rect 238661 134270 240212 134272
rect 266261 134328 268180 134330
rect 266261 134272 266266 134328
rect 266322 134272 268180 134328
rect 266261 134270 268180 134272
rect 293861 134328 296148 134330
rect 293861 134272 293866 134328
rect 293922 134272 296148 134328
rect 293861 134270 296148 134272
rect 322841 134328 324116 134330
rect 322841 134272 322846 134328
rect 322902 134272 324116 134328
rect 322841 134270 324116 134272
rect 350441 134328 352084 134330
rect 350441 134272 350446 134328
rect 350502 134272 352084 134328
rect 350441 134270 352084 134272
rect 378041 134328 380052 134330
rect 378041 134272 378046 134328
rect 378102 134272 380052 134328
rect 378041 134270 380052 134272
rect 405641 134328 408204 134330
rect 405641 134272 405646 134328
rect 405702 134272 408204 134328
rect 405641 134270 408204 134272
rect 434621 134328 436172 134330
rect 434621 134272 434626 134328
rect 434682 134272 436172 134328
rect 434621 134270 436172 134272
rect 462221 134328 464140 134330
rect 462221 134272 462226 134328
rect 462282 134272 464140 134328
rect 462221 134270 464140 134272
rect 489821 134328 492108 134330
rect 489821 134272 489826 134328
rect 489882 134272 492108 134328
rect 489821 134270 492108 134272
rect 518801 134328 520076 134330
rect 518801 134272 518806 134328
rect 518862 134272 520076 134328
rect 518801 134270 520076 134272
rect 546401 134328 548044 134330
rect 546401 134272 546406 134328
rect 546462 134272 548044 134328
rect 546401 134270 548044 134272
rect 13537 134267 13603 134270
rect 42701 134267 42767 134270
rect 70301 134267 70367 134270
rect 97901 134267 97967 134270
rect 126881 134267 126947 134270
rect 154481 134267 154547 134270
rect 182081 134267 182147 134270
rect 209681 134267 209747 134270
rect 238661 134267 238727 134270
rect 266261 134267 266327 134270
rect 293861 134267 293927 134270
rect 322841 134267 322907 134270
rect 350441 134267 350507 134270
rect 378041 134267 378107 134270
rect 405641 134267 405707 134270
rect 434621 134267 434687 134270
rect 462221 134267 462287 134270
rect 489821 134267 489887 134270
rect 518801 134267 518867 134270
rect 546401 134267 546467 134270
rect 37273 133650 37339 133653
rect 66253 133650 66319 133653
rect 93853 133650 93919 133653
rect 121453 133650 121519 133653
rect 149053 133650 149119 133653
rect 178033 133650 178099 133653
rect 205633 133650 205699 133653
rect 233233 133650 233299 133653
rect 262213 133650 262279 133653
rect 289813 133650 289879 133653
rect 317413 133650 317479 133653
rect 345013 133650 345079 133653
rect 373993 133650 374059 133653
rect 401593 133650 401659 133653
rect 429285 133650 429351 133653
rect 458173 133650 458239 133653
rect 485773 133650 485839 133653
rect 513373 133650 513439 133653
rect 542353 133650 542419 133653
rect 569953 133650 570019 133653
rect 35788 133648 37339 133650
rect 35788 133592 37278 133648
rect 37334 133592 37339 133648
rect 35788 133590 37339 133592
rect 63940 133648 66319 133650
rect 63940 133592 66258 133648
rect 66314 133592 66319 133648
rect 63940 133590 66319 133592
rect 91908 133648 93919 133650
rect 91908 133592 93858 133648
rect 93914 133592 93919 133648
rect 91908 133590 93919 133592
rect 119876 133648 121519 133650
rect 119876 133592 121458 133648
rect 121514 133592 121519 133648
rect 119876 133590 121519 133592
rect 147844 133648 149119 133650
rect 147844 133592 149058 133648
rect 149114 133592 149119 133648
rect 147844 133590 149119 133592
rect 175812 133648 178099 133650
rect 175812 133592 178038 133648
rect 178094 133592 178099 133648
rect 175812 133590 178099 133592
rect 203964 133648 205699 133650
rect 203964 133592 205638 133648
rect 205694 133592 205699 133648
rect 203964 133590 205699 133592
rect 231932 133648 233299 133650
rect 231932 133592 233238 133648
rect 233294 133592 233299 133648
rect 231932 133590 233299 133592
rect 259900 133648 262279 133650
rect 259900 133592 262218 133648
rect 262274 133592 262279 133648
rect 259900 133590 262279 133592
rect 287868 133648 289879 133650
rect 287868 133592 289818 133648
rect 289874 133592 289879 133648
rect 287868 133590 289879 133592
rect 315836 133648 317479 133650
rect 315836 133592 317418 133648
rect 317474 133592 317479 133648
rect 315836 133590 317479 133592
rect 343804 133648 345079 133650
rect 343804 133592 345018 133648
rect 345074 133592 345079 133648
rect 343804 133590 345079 133592
rect 371956 133648 374059 133650
rect 371956 133592 373998 133648
rect 374054 133592 374059 133648
rect 371956 133590 374059 133592
rect 399924 133648 401659 133650
rect 399924 133592 401598 133648
rect 401654 133592 401659 133648
rect 399924 133590 401659 133592
rect 427892 133648 429351 133650
rect 427892 133592 429290 133648
rect 429346 133592 429351 133648
rect 427892 133590 429351 133592
rect 455860 133648 458239 133650
rect 455860 133592 458178 133648
rect 458234 133592 458239 133648
rect 455860 133590 458239 133592
rect 483828 133648 485839 133650
rect 483828 133592 485778 133648
rect 485834 133592 485839 133648
rect 483828 133590 485839 133592
rect 511796 133648 513439 133650
rect 511796 133592 513378 133648
rect 513434 133592 513439 133648
rect 511796 133590 513439 133592
rect 539948 133648 542419 133650
rect 539948 133592 542358 133648
rect 542414 133592 542419 133648
rect 539948 133590 542419 133592
rect 567916 133648 570019 133650
rect 567916 133592 569958 133648
rect 570014 133592 570019 133648
rect 567916 133590 570019 133592
rect 37273 133587 37339 133590
rect 66253 133587 66319 133590
rect 93853 133587 93919 133590
rect 121453 133587 121519 133590
rect 149053 133587 149119 133590
rect 178033 133587 178099 133590
rect 205633 133587 205699 133590
rect 233233 133587 233299 133590
rect 262213 133587 262279 133590
rect 289813 133587 289879 133590
rect 317413 133587 317479 133590
rect 345013 133587 345079 133590
rect 373993 133587 374059 133590
rect 401593 133587 401659 133590
rect 429285 133587 429351 133590
rect 458173 133587 458239 133590
rect 485773 133587 485839 133590
rect 513373 133587 513439 133590
rect 542353 133587 542419 133590
rect 569953 133587 570019 133590
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect -960 110516 480 110756
rect 13537 107402 13603 107405
rect 42701 107402 42767 107405
rect 70301 107402 70367 107405
rect 97901 107402 97967 107405
rect 126881 107402 126947 107405
rect 154481 107402 154547 107405
rect 182081 107402 182147 107405
rect 209681 107402 209747 107405
rect 238661 107402 238727 107405
rect 266261 107402 266327 107405
rect 293861 107402 293927 107405
rect 322841 107402 322907 107405
rect 350441 107402 350507 107405
rect 378041 107402 378107 107405
rect 405641 107402 405707 107405
rect 434621 107402 434687 107405
rect 462221 107402 462287 107405
rect 489821 107402 489887 107405
rect 518801 107402 518867 107405
rect 546401 107402 546467 107405
rect 13537 107400 16100 107402
rect 13537 107344 13542 107400
rect 13598 107344 16100 107400
rect 13537 107342 16100 107344
rect 42701 107400 44068 107402
rect 42701 107344 42706 107400
rect 42762 107344 44068 107400
rect 42701 107342 44068 107344
rect 70301 107400 72036 107402
rect 70301 107344 70306 107400
rect 70362 107344 72036 107400
rect 70301 107342 72036 107344
rect 97901 107400 100188 107402
rect 97901 107344 97906 107400
rect 97962 107344 100188 107400
rect 97901 107342 100188 107344
rect 126881 107400 128156 107402
rect 126881 107344 126886 107400
rect 126942 107344 128156 107400
rect 126881 107342 128156 107344
rect 154481 107400 156124 107402
rect 154481 107344 154486 107400
rect 154542 107344 156124 107400
rect 154481 107342 156124 107344
rect 182081 107400 184092 107402
rect 182081 107344 182086 107400
rect 182142 107344 184092 107400
rect 182081 107342 184092 107344
rect 209681 107400 212060 107402
rect 209681 107344 209686 107400
rect 209742 107344 212060 107400
rect 209681 107342 212060 107344
rect 238661 107400 240212 107402
rect 238661 107344 238666 107400
rect 238722 107344 240212 107400
rect 238661 107342 240212 107344
rect 266261 107400 268180 107402
rect 266261 107344 266266 107400
rect 266322 107344 268180 107400
rect 266261 107342 268180 107344
rect 293861 107400 296148 107402
rect 293861 107344 293866 107400
rect 293922 107344 296148 107400
rect 293861 107342 296148 107344
rect 322841 107400 324116 107402
rect 322841 107344 322846 107400
rect 322902 107344 324116 107400
rect 322841 107342 324116 107344
rect 350441 107400 352084 107402
rect 350441 107344 350446 107400
rect 350502 107344 352084 107400
rect 350441 107342 352084 107344
rect 378041 107400 380052 107402
rect 378041 107344 378046 107400
rect 378102 107344 380052 107400
rect 378041 107342 380052 107344
rect 405641 107400 408204 107402
rect 405641 107344 405646 107400
rect 405702 107344 408204 107400
rect 405641 107342 408204 107344
rect 434621 107400 436172 107402
rect 434621 107344 434626 107400
rect 434682 107344 436172 107400
rect 434621 107342 436172 107344
rect 462221 107400 464140 107402
rect 462221 107344 462226 107400
rect 462282 107344 464140 107400
rect 462221 107342 464140 107344
rect 489821 107400 492108 107402
rect 489821 107344 489826 107400
rect 489882 107344 492108 107400
rect 489821 107342 492108 107344
rect 518801 107400 520076 107402
rect 518801 107344 518806 107400
rect 518862 107344 520076 107400
rect 518801 107342 520076 107344
rect 546401 107400 548044 107402
rect 546401 107344 546406 107400
rect 546462 107344 548044 107400
rect 546401 107342 548044 107344
rect 13537 107339 13603 107342
rect 42701 107339 42767 107342
rect 70301 107339 70367 107342
rect 97901 107339 97967 107342
rect 126881 107339 126947 107342
rect 154481 107339 154547 107342
rect 182081 107339 182147 107342
rect 209681 107339 209747 107342
rect 238661 107339 238727 107342
rect 266261 107339 266327 107342
rect 293861 107339 293927 107342
rect 322841 107339 322907 107342
rect 350441 107339 350507 107342
rect 378041 107339 378107 107342
rect 405641 107339 405707 107342
rect 434621 107339 434687 107342
rect 462221 107339 462287 107342
rect 489821 107339 489887 107342
rect 518801 107339 518867 107342
rect 546401 107339 546467 107342
rect 147844 106730 148242 106790
rect 37273 106722 37339 106725
rect 66253 106722 66319 106725
rect 93853 106722 93919 106725
rect 121453 106722 121519 106725
rect 35788 106720 37339 106722
rect 35788 106664 37278 106720
rect 37334 106664 37339 106720
rect 35788 106662 37339 106664
rect 63940 106720 66319 106722
rect 63940 106664 66258 106720
rect 66314 106664 66319 106720
rect 63940 106662 66319 106664
rect 91908 106720 93919 106722
rect 91908 106664 93858 106720
rect 93914 106664 93919 106720
rect 91908 106662 93919 106664
rect 119876 106720 121519 106722
rect 119876 106664 121458 106720
rect 121514 106664 121519 106720
rect 119876 106662 121519 106664
rect 148182 106722 148242 106730
rect 149053 106722 149119 106725
rect 178033 106722 178099 106725
rect 205633 106722 205699 106725
rect 233233 106722 233299 106725
rect 262213 106722 262279 106725
rect 289813 106722 289879 106725
rect 317413 106722 317479 106725
rect 345013 106722 345079 106725
rect 373993 106722 374059 106725
rect 401593 106722 401659 106725
rect 429285 106722 429351 106725
rect 458173 106722 458239 106725
rect 485773 106722 485839 106725
rect 513373 106722 513439 106725
rect 542353 106722 542419 106725
rect 569953 106722 570019 106725
rect 148182 106720 149119 106722
rect 148182 106664 149058 106720
rect 149114 106664 149119 106720
rect 148182 106662 149119 106664
rect 175812 106720 178099 106722
rect 175812 106664 178038 106720
rect 178094 106664 178099 106720
rect 175812 106662 178099 106664
rect 203964 106720 205699 106722
rect 203964 106664 205638 106720
rect 205694 106664 205699 106720
rect 203964 106662 205699 106664
rect 231932 106720 233299 106722
rect 231932 106664 233238 106720
rect 233294 106664 233299 106720
rect 231932 106662 233299 106664
rect 259900 106720 262279 106722
rect 259900 106664 262218 106720
rect 262274 106664 262279 106720
rect 259900 106662 262279 106664
rect 287868 106720 289879 106722
rect 287868 106664 289818 106720
rect 289874 106664 289879 106720
rect 287868 106662 289879 106664
rect 315836 106720 317479 106722
rect 315836 106664 317418 106720
rect 317474 106664 317479 106720
rect 315836 106662 317479 106664
rect 343804 106720 345079 106722
rect 343804 106664 345018 106720
rect 345074 106664 345079 106720
rect 343804 106662 345079 106664
rect 371956 106720 374059 106722
rect 371956 106664 373998 106720
rect 374054 106664 374059 106720
rect 371956 106662 374059 106664
rect 399924 106720 401659 106722
rect 399924 106664 401598 106720
rect 401654 106664 401659 106720
rect 399924 106662 401659 106664
rect 427892 106720 429351 106722
rect 427892 106664 429290 106720
rect 429346 106664 429351 106720
rect 427892 106662 429351 106664
rect 455860 106720 458239 106722
rect 455860 106664 458178 106720
rect 458234 106664 458239 106720
rect 455860 106662 458239 106664
rect 483828 106720 485839 106722
rect 483828 106664 485778 106720
rect 485834 106664 485839 106720
rect 483828 106662 485839 106664
rect 511796 106720 513439 106722
rect 511796 106664 513378 106720
rect 513434 106664 513439 106720
rect 511796 106662 513439 106664
rect 539948 106720 542419 106722
rect 539948 106664 542358 106720
rect 542414 106664 542419 106720
rect 539948 106662 542419 106664
rect 567916 106720 570019 106722
rect 567916 106664 569958 106720
rect 570014 106664 570019 106720
rect 567916 106662 570019 106664
rect 37273 106659 37339 106662
rect 66253 106659 66319 106662
rect 93853 106659 93919 106662
rect 121453 106659 121519 106662
rect 149053 106659 149119 106662
rect 178033 106659 178099 106662
rect 205633 106659 205699 106662
rect 233233 106659 233299 106662
rect 262213 106659 262279 106662
rect 289813 106659 289879 106662
rect 317413 106659 317479 106662
rect 345013 106659 345079 106662
rect 373993 106659 374059 106662
rect 401593 106659 401659 106662
rect 429285 106659 429351 106662
rect 458173 106659 458239 106662
rect 485773 106659 485839 106662
rect 513373 106659 513439 106662
rect 542353 106659 542419 106662
rect 569953 106659 570019 106662
rect 583520 99364 584960 99604
rect -960 97610 480 97700
rect 4061 97610 4127 97613
rect -960 97608 4127 97610
rect -960 97552 4066 97608
rect 4122 97552 4127 97608
rect -960 97550 4127 97552
rect -960 97460 480 97550
rect 4061 97547 4127 97550
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 13537 80338 13603 80341
rect 42701 80338 42767 80341
rect 70301 80338 70367 80341
rect 97901 80338 97967 80341
rect 126881 80338 126947 80341
rect 154481 80338 154547 80341
rect 182081 80338 182147 80341
rect 209681 80338 209747 80341
rect 238661 80338 238727 80341
rect 266261 80338 266327 80341
rect 293861 80338 293927 80341
rect 322841 80338 322907 80341
rect 350441 80338 350507 80341
rect 378041 80338 378107 80341
rect 405641 80338 405707 80341
rect 434621 80338 434687 80341
rect 462221 80338 462287 80341
rect 489821 80338 489887 80341
rect 518801 80338 518867 80341
rect 546401 80338 546467 80341
rect 13537 80336 16100 80338
rect 13537 80280 13542 80336
rect 13598 80280 16100 80336
rect 13537 80278 16100 80280
rect 42701 80336 44068 80338
rect 42701 80280 42706 80336
rect 42762 80280 44068 80336
rect 42701 80278 44068 80280
rect 70301 80336 72036 80338
rect 70301 80280 70306 80336
rect 70362 80280 72036 80336
rect 70301 80278 72036 80280
rect 97901 80336 100188 80338
rect 97901 80280 97906 80336
rect 97962 80280 100188 80336
rect 97901 80278 100188 80280
rect 126881 80336 128156 80338
rect 126881 80280 126886 80336
rect 126942 80280 128156 80336
rect 126881 80278 128156 80280
rect 154481 80336 156124 80338
rect 154481 80280 154486 80336
rect 154542 80280 156124 80336
rect 154481 80278 156124 80280
rect 182081 80336 184092 80338
rect 182081 80280 182086 80336
rect 182142 80280 184092 80336
rect 182081 80278 184092 80280
rect 209681 80336 212060 80338
rect 209681 80280 209686 80336
rect 209742 80280 212060 80336
rect 209681 80278 212060 80280
rect 238661 80336 240212 80338
rect 238661 80280 238666 80336
rect 238722 80280 240212 80336
rect 238661 80278 240212 80280
rect 266261 80336 268180 80338
rect 266261 80280 266266 80336
rect 266322 80280 268180 80336
rect 266261 80278 268180 80280
rect 293861 80336 296148 80338
rect 293861 80280 293866 80336
rect 293922 80280 296148 80336
rect 293861 80278 296148 80280
rect 322841 80336 324116 80338
rect 322841 80280 322846 80336
rect 322902 80280 324116 80336
rect 322841 80278 324116 80280
rect 350441 80336 352084 80338
rect 350441 80280 350446 80336
rect 350502 80280 352084 80336
rect 350441 80278 352084 80280
rect 378041 80336 380052 80338
rect 378041 80280 378046 80336
rect 378102 80280 380052 80336
rect 378041 80278 380052 80280
rect 405641 80336 408204 80338
rect 405641 80280 405646 80336
rect 405702 80280 408204 80336
rect 405641 80278 408204 80280
rect 434621 80336 436172 80338
rect 434621 80280 434626 80336
rect 434682 80280 436172 80336
rect 434621 80278 436172 80280
rect 462221 80336 464140 80338
rect 462221 80280 462226 80336
rect 462282 80280 464140 80336
rect 462221 80278 464140 80280
rect 489821 80336 492108 80338
rect 489821 80280 489826 80336
rect 489882 80280 492108 80336
rect 489821 80278 492108 80280
rect 518801 80336 520076 80338
rect 518801 80280 518806 80336
rect 518862 80280 520076 80336
rect 518801 80278 520076 80280
rect 546401 80336 548044 80338
rect 546401 80280 546406 80336
rect 546462 80280 548044 80336
rect 546401 80278 548044 80280
rect 13537 80275 13603 80278
rect 42701 80275 42767 80278
rect 70301 80275 70367 80278
rect 97901 80275 97967 80278
rect 126881 80275 126947 80278
rect 154481 80275 154547 80278
rect 182081 80275 182147 80278
rect 209681 80275 209747 80278
rect 238661 80275 238727 80278
rect 266261 80275 266327 80278
rect 293861 80275 293927 80278
rect 322841 80275 322907 80278
rect 350441 80275 350507 80278
rect 378041 80275 378107 80278
rect 405641 80275 405707 80278
rect 434621 80275 434687 80278
rect 462221 80275 462287 80278
rect 489821 80275 489887 80278
rect 518801 80275 518867 80278
rect 546401 80275 546467 80278
rect 37273 79658 37339 79661
rect 66253 79658 66319 79661
rect 93853 79658 93919 79661
rect 121453 79658 121519 79661
rect 149053 79658 149119 79661
rect 178033 79658 178099 79661
rect 205633 79658 205699 79661
rect 233233 79658 233299 79661
rect 262213 79658 262279 79661
rect 289813 79658 289879 79661
rect 317413 79658 317479 79661
rect 345013 79658 345079 79661
rect 373993 79658 374059 79661
rect 401593 79658 401659 79661
rect 429285 79658 429351 79661
rect 458173 79658 458239 79661
rect 485773 79658 485839 79661
rect 513373 79658 513439 79661
rect 542353 79658 542419 79661
rect 569953 79658 570019 79661
rect 35788 79656 37339 79658
rect 35788 79600 37278 79656
rect 37334 79600 37339 79656
rect 35788 79598 37339 79600
rect 63940 79656 66319 79658
rect 63940 79600 66258 79656
rect 66314 79600 66319 79656
rect 63940 79598 66319 79600
rect 91908 79656 93919 79658
rect 91908 79600 93858 79656
rect 93914 79600 93919 79656
rect 91908 79598 93919 79600
rect 119876 79656 121519 79658
rect 119876 79600 121458 79656
rect 121514 79600 121519 79656
rect 119876 79598 121519 79600
rect 147844 79656 149119 79658
rect 147844 79600 149058 79656
rect 149114 79600 149119 79656
rect 147844 79598 149119 79600
rect 175812 79656 178099 79658
rect 175812 79600 178038 79656
rect 178094 79600 178099 79656
rect 175812 79598 178099 79600
rect 203964 79656 205699 79658
rect 203964 79600 205638 79656
rect 205694 79600 205699 79656
rect 203964 79598 205699 79600
rect 231932 79656 233299 79658
rect 231932 79600 233238 79656
rect 233294 79600 233299 79656
rect 231932 79598 233299 79600
rect 259900 79656 262279 79658
rect 259900 79600 262218 79656
rect 262274 79600 262279 79656
rect 259900 79598 262279 79600
rect 287868 79656 289879 79658
rect 287868 79600 289818 79656
rect 289874 79600 289879 79656
rect 287868 79598 289879 79600
rect 315836 79656 317479 79658
rect 315836 79600 317418 79656
rect 317474 79600 317479 79656
rect 315836 79598 317479 79600
rect 343804 79656 345079 79658
rect 343804 79600 345018 79656
rect 345074 79600 345079 79656
rect 343804 79598 345079 79600
rect 371956 79656 374059 79658
rect 371956 79600 373998 79656
rect 374054 79600 374059 79656
rect 371956 79598 374059 79600
rect 399924 79656 401659 79658
rect 399924 79600 401598 79656
rect 401654 79600 401659 79656
rect 399924 79598 401659 79600
rect 427892 79656 429351 79658
rect 427892 79600 429290 79656
rect 429346 79600 429351 79656
rect 427892 79598 429351 79600
rect 455860 79656 458239 79658
rect 455860 79600 458178 79656
rect 458234 79600 458239 79656
rect 455860 79598 458239 79600
rect 483828 79656 485839 79658
rect 483828 79600 485778 79656
rect 485834 79600 485839 79656
rect 483828 79598 485839 79600
rect 511796 79656 513439 79658
rect 511796 79600 513378 79656
rect 513434 79600 513439 79656
rect 511796 79598 513439 79600
rect 539948 79656 542419 79658
rect 539948 79600 542358 79656
rect 542414 79600 542419 79656
rect 539948 79598 542419 79600
rect 567916 79656 570019 79658
rect 567916 79600 569958 79656
rect 570014 79600 570019 79656
rect 567916 79598 570019 79600
rect 37273 79595 37339 79598
rect 66253 79595 66319 79598
rect 93853 79595 93919 79598
rect 121453 79595 121519 79598
rect 149053 79595 149119 79598
rect 178033 79595 178099 79598
rect 205633 79595 205699 79598
rect 233233 79595 233299 79598
rect 262213 79595 262279 79598
rect 289813 79595 289879 79598
rect 317413 79595 317479 79598
rect 345013 79595 345079 79598
rect 373993 79595 374059 79598
rect 401593 79595 401659 79598
rect 429285 79595 429351 79598
rect 458173 79595 458239 79598
rect 485773 79595 485839 79598
rect 513373 79595 513439 79598
rect 542353 79595 542419 79598
rect 569953 79595 570019 79598
rect 580073 72994 580139 72997
rect 583520 72994 584960 73084
rect 580073 72992 584960 72994
rect 580073 72936 580078 72992
rect 580134 72936 584960 72992
rect 580073 72934 584960 72936
rect 580073 72931 580139 72934
rect 583520 72844 584960 72934
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58578 480 58668
rect 3325 58578 3391 58581
rect -960 58576 3391 58578
rect -960 58520 3330 58576
rect 3386 58520 3391 58576
rect -960 58518 3391 58520
rect -960 58428 480 58518
rect 3325 58515 3391 58518
rect 13537 53410 13603 53413
rect 42701 53410 42767 53413
rect 70301 53410 70367 53413
rect 97901 53410 97967 53413
rect 126881 53410 126947 53413
rect 154481 53410 154547 53413
rect 182081 53410 182147 53413
rect 209681 53410 209747 53413
rect 238661 53410 238727 53413
rect 266261 53410 266327 53413
rect 293861 53410 293927 53413
rect 322841 53410 322907 53413
rect 350441 53410 350507 53413
rect 378041 53410 378107 53413
rect 405641 53410 405707 53413
rect 434621 53410 434687 53413
rect 462221 53410 462287 53413
rect 489821 53410 489887 53413
rect 518801 53410 518867 53413
rect 546401 53410 546467 53413
rect 13537 53408 16100 53410
rect 13537 53352 13542 53408
rect 13598 53352 16100 53408
rect 13537 53350 16100 53352
rect 42701 53408 44068 53410
rect 42701 53352 42706 53408
rect 42762 53352 44068 53408
rect 42701 53350 44068 53352
rect 70301 53408 72036 53410
rect 70301 53352 70306 53408
rect 70362 53352 72036 53408
rect 70301 53350 72036 53352
rect 97901 53408 100188 53410
rect 97901 53352 97906 53408
rect 97962 53352 100188 53408
rect 97901 53350 100188 53352
rect 126881 53408 128156 53410
rect 126881 53352 126886 53408
rect 126942 53352 128156 53408
rect 126881 53350 128156 53352
rect 154481 53408 156124 53410
rect 154481 53352 154486 53408
rect 154542 53352 156124 53408
rect 154481 53350 156124 53352
rect 182081 53408 184092 53410
rect 182081 53352 182086 53408
rect 182142 53352 184092 53408
rect 182081 53350 184092 53352
rect 209681 53408 212060 53410
rect 209681 53352 209686 53408
rect 209742 53352 212060 53408
rect 209681 53350 212060 53352
rect 238661 53408 240212 53410
rect 238661 53352 238666 53408
rect 238722 53352 240212 53408
rect 238661 53350 240212 53352
rect 266261 53408 268180 53410
rect 266261 53352 266266 53408
rect 266322 53352 268180 53408
rect 266261 53350 268180 53352
rect 293861 53408 296148 53410
rect 293861 53352 293866 53408
rect 293922 53352 296148 53408
rect 293861 53350 296148 53352
rect 322841 53408 324116 53410
rect 322841 53352 322846 53408
rect 322902 53352 324116 53408
rect 322841 53350 324116 53352
rect 350441 53408 352084 53410
rect 350441 53352 350446 53408
rect 350502 53352 352084 53408
rect 350441 53350 352084 53352
rect 378041 53408 380052 53410
rect 378041 53352 378046 53408
rect 378102 53352 380052 53408
rect 378041 53350 380052 53352
rect 405641 53408 408204 53410
rect 405641 53352 405646 53408
rect 405702 53352 408204 53408
rect 405641 53350 408204 53352
rect 434621 53408 436172 53410
rect 434621 53352 434626 53408
rect 434682 53352 436172 53408
rect 434621 53350 436172 53352
rect 462221 53408 464140 53410
rect 462221 53352 462226 53408
rect 462282 53352 464140 53408
rect 462221 53350 464140 53352
rect 489821 53408 492108 53410
rect 489821 53352 489826 53408
rect 489882 53352 492108 53408
rect 489821 53350 492108 53352
rect 518801 53408 520076 53410
rect 518801 53352 518806 53408
rect 518862 53352 520076 53408
rect 518801 53350 520076 53352
rect 546401 53408 548044 53410
rect 546401 53352 546406 53408
rect 546462 53352 548044 53408
rect 546401 53350 548044 53352
rect 13537 53347 13603 53350
rect 42701 53347 42767 53350
rect 70301 53347 70367 53350
rect 97901 53347 97967 53350
rect 126881 53347 126947 53350
rect 154481 53347 154547 53350
rect 182081 53347 182147 53350
rect 209681 53347 209747 53350
rect 238661 53347 238727 53350
rect 266261 53347 266327 53350
rect 293861 53347 293927 53350
rect 322841 53347 322907 53350
rect 350441 53347 350507 53350
rect 378041 53347 378107 53350
rect 405641 53347 405707 53350
rect 434621 53347 434687 53350
rect 462221 53347 462287 53350
rect 489821 53347 489887 53350
rect 518801 53347 518867 53350
rect 546401 53347 546467 53350
rect 37273 52730 37339 52733
rect 66253 52730 66319 52733
rect 93853 52730 93919 52733
rect 121453 52730 121519 52733
rect 149053 52730 149119 52733
rect 178033 52730 178099 52733
rect 205633 52730 205699 52733
rect 233233 52730 233299 52733
rect 262213 52730 262279 52733
rect 289813 52730 289879 52733
rect 317413 52730 317479 52733
rect 345013 52730 345079 52733
rect 373993 52730 374059 52733
rect 401593 52730 401659 52733
rect 429285 52730 429351 52733
rect 458173 52730 458239 52733
rect 485773 52730 485839 52733
rect 513373 52730 513439 52733
rect 542353 52730 542419 52733
rect 569953 52730 570019 52733
rect 35788 52728 37339 52730
rect 35788 52672 37278 52728
rect 37334 52672 37339 52728
rect 35788 52670 37339 52672
rect 63940 52728 66319 52730
rect 63940 52672 66258 52728
rect 66314 52672 66319 52728
rect 63940 52670 66319 52672
rect 91908 52728 93919 52730
rect 91908 52672 93858 52728
rect 93914 52672 93919 52728
rect 91908 52670 93919 52672
rect 119876 52728 121519 52730
rect 119876 52672 121458 52728
rect 121514 52672 121519 52728
rect 119876 52670 121519 52672
rect 147844 52728 149119 52730
rect 147844 52672 149058 52728
rect 149114 52672 149119 52728
rect 147844 52670 149119 52672
rect 175812 52728 178099 52730
rect 175812 52672 178038 52728
rect 178094 52672 178099 52728
rect 175812 52670 178099 52672
rect 203964 52728 205699 52730
rect 203964 52672 205638 52728
rect 205694 52672 205699 52728
rect 203964 52670 205699 52672
rect 231932 52728 233299 52730
rect 231932 52672 233238 52728
rect 233294 52672 233299 52728
rect 231932 52670 233299 52672
rect 259900 52728 262279 52730
rect 259900 52672 262218 52728
rect 262274 52672 262279 52728
rect 259900 52670 262279 52672
rect 287868 52728 289879 52730
rect 287868 52672 289818 52728
rect 289874 52672 289879 52728
rect 287868 52670 289879 52672
rect 315836 52728 317479 52730
rect 315836 52672 317418 52728
rect 317474 52672 317479 52728
rect 315836 52670 317479 52672
rect 343804 52728 345079 52730
rect 343804 52672 345018 52728
rect 345074 52672 345079 52728
rect 343804 52670 345079 52672
rect 371956 52728 374059 52730
rect 371956 52672 373998 52728
rect 374054 52672 374059 52728
rect 371956 52670 374059 52672
rect 399924 52728 401659 52730
rect 399924 52672 401598 52728
rect 401654 52672 401659 52728
rect 399924 52670 401659 52672
rect 427892 52728 429351 52730
rect 427892 52672 429290 52728
rect 429346 52672 429351 52728
rect 427892 52670 429351 52672
rect 455860 52728 458239 52730
rect 455860 52672 458178 52728
rect 458234 52672 458239 52728
rect 455860 52670 458239 52672
rect 483828 52728 485839 52730
rect 483828 52672 485778 52728
rect 485834 52672 485839 52728
rect 483828 52670 485839 52672
rect 511796 52728 513439 52730
rect 511796 52672 513378 52728
rect 513434 52672 513439 52728
rect 511796 52670 513439 52672
rect 539948 52728 542419 52730
rect 539948 52672 542358 52728
rect 542414 52672 542419 52728
rect 539948 52670 542419 52672
rect 567916 52728 570019 52730
rect 567916 52672 569958 52728
rect 570014 52672 570019 52728
rect 567916 52670 570019 52672
rect 37273 52667 37339 52670
rect 66253 52667 66319 52670
rect 93853 52667 93919 52670
rect 121453 52667 121519 52670
rect 149053 52667 149119 52670
rect 178033 52667 178099 52670
rect 205633 52667 205699 52670
rect 233233 52667 233299 52670
rect 262213 52667 262279 52670
rect 289813 52667 289879 52670
rect 317413 52667 317479 52670
rect 345013 52667 345079 52670
rect 373993 52667 374059 52670
rect 401593 52667 401659 52670
rect 429285 52667 429351 52670
rect 458173 52667 458239 52670
rect 485773 52667 485839 52670
rect 513373 52667 513439 52670
rect 542353 52667 542419 52670
rect 569953 52667 570019 52670
rect 583520 46188 584960 46428
rect -960 45522 480 45612
rect 2957 45522 3023 45525
rect -960 45520 3023 45522
rect -960 45464 2962 45520
rect 3018 45464 3023 45520
rect -960 45462 3023 45464
rect -960 45372 480 45462
rect 2957 45459 3023 45462
rect 48078 42060 48084 42124
rect 48148 42122 48154 42124
rect 153837 42122 153903 42125
rect 48148 42120 153903 42122
rect 48148 42064 153842 42120
rect 153898 42064 153903 42120
rect 48148 42062 153903 42064
rect 48148 42060 48154 42062
rect 153837 42059 153903 42062
rect 17309 37906 17375 37909
rect 580758 37906 580764 37908
rect 17309 37904 580764 37906
rect 17309 37848 17314 37904
rect 17370 37848 580764 37904
rect 17309 37846 580764 37848
rect 17309 37843 17375 37846
rect 580758 37844 580764 37846
rect 580828 37844 580834 37908
rect 42742 35260 42748 35324
rect 42812 35322 42818 35324
rect 43437 35322 43503 35325
rect 42812 35320 43503 35322
rect 42812 35264 43442 35320
rect 43498 35264 43503 35320
rect 42812 35262 43503 35264
rect 42812 35260 42818 35262
rect 43437 35259 43503 35262
rect 64229 35186 64295 35189
rect 61916 35184 64295 35186
rect 61916 35128 64234 35184
rect 64290 35128 64295 35184
rect 61916 35126 64295 35128
rect 64229 35123 64295 35126
rect 11881 34506 11947 34509
rect 11881 34504 16100 34506
rect 11881 34448 11886 34504
rect 11942 34448 16100 34504
rect 11881 34446 16100 34448
rect 11881 34443 11947 34446
rect 61285 34370 61351 34373
rect 61285 34368 61394 34370
rect 61285 34312 61290 34368
rect 61346 34312 61394 34368
rect 61285 34307 61394 34312
rect 61334 33796 61394 34307
rect 13445 33146 13511 33149
rect 579981 33146 580047 33149
rect 583520 33146 584960 33236
rect 13445 33144 16100 33146
rect 13445 33088 13450 33144
rect 13506 33088 16100 33144
rect 13445 33086 16100 33088
rect 579981 33144 584960 33146
rect 579981 33088 579986 33144
rect 580042 33088 584960 33144
rect 579981 33086 584960 33088
rect 13445 33083 13511 33086
rect 579981 33083 580047 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 64505 31650 64571 31653
rect 61916 31648 64571 31650
rect 61916 31592 64510 31648
rect 64566 31592 64571 31648
rect 61916 31590 64571 31592
rect 64505 31587 64571 31590
rect 12433 31106 12499 31109
rect 12433 31104 16100 31106
rect 12433 31048 12438 31104
rect 12494 31048 16100 31104
rect 12433 31046 16100 31048
rect 12433 31043 12499 31046
rect 64229 30290 64295 30293
rect 61916 30288 64295 30290
rect 61916 30232 64234 30288
rect 64290 30232 64295 30288
rect 61916 30230 64295 30232
rect 64229 30227 64295 30230
rect 13721 29746 13787 29749
rect 13721 29744 16100 29746
rect 13721 29688 13726 29744
rect 13782 29688 16100 29744
rect 13721 29686 16100 29688
rect 13721 29683 13787 29686
rect 63493 28386 63559 28389
rect 61916 28384 63559 28386
rect 61916 28328 63498 28384
rect 63554 28328 63559 28384
rect 61916 28326 63559 28328
rect 63493 28323 63559 28326
rect 13629 27706 13695 27709
rect 13629 27704 16100 27706
rect 13629 27648 13634 27704
rect 13690 27648 16100 27704
rect 13629 27646 16100 27648
rect 13629 27643 13695 27646
rect 63493 27026 63559 27029
rect 61916 27024 63559 27026
rect 61916 26968 63498 27024
rect 63554 26968 63559 27024
rect 61916 26966 63559 26968
rect 63493 26963 63559 26966
rect 70301 26890 70367 26893
rect 70301 26888 72066 26890
rect 70301 26832 70306 26888
rect 70362 26832 72066 26888
rect 70301 26830 72066 26832
rect 70301 26827 70367 26830
rect 13537 26346 13603 26349
rect 13537 26344 16100 26346
rect 13537 26288 13542 26344
rect 13598 26288 16100 26344
rect 72006 26316 72066 26830
rect 97901 26346 97967 26349
rect 126881 26346 126947 26349
rect 154481 26346 154547 26349
rect 182081 26346 182147 26349
rect 209681 26346 209747 26349
rect 238661 26346 238727 26349
rect 266261 26346 266327 26349
rect 293861 26346 293927 26349
rect 322841 26346 322907 26349
rect 350441 26346 350507 26349
rect 378041 26346 378107 26349
rect 405641 26346 405707 26349
rect 434621 26346 434687 26349
rect 462221 26346 462287 26349
rect 489821 26346 489887 26349
rect 518801 26346 518867 26349
rect 546401 26346 546467 26349
rect 97901 26344 100188 26346
rect 13537 26286 16100 26288
rect 97901 26288 97906 26344
rect 97962 26288 100188 26344
rect 97901 26286 100188 26288
rect 126881 26344 128156 26346
rect 126881 26288 126886 26344
rect 126942 26288 128156 26344
rect 126881 26286 128156 26288
rect 154481 26344 156124 26346
rect 154481 26288 154486 26344
rect 154542 26288 156124 26344
rect 154481 26286 156124 26288
rect 182081 26344 184092 26346
rect 182081 26288 182086 26344
rect 182142 26288 184092 26344
rect 182081 26286 184092 26288
rect 209681 26344 212060 26346
rect 209681 26288 209686 26344
rect 209742 26288 212060 26344
rect 209681 26286 212060 26288
rect 238661 26344 240212 26346
rect 238661 26288 238666 26344
rect 238722 26288 240212 26344
rect 238661 26286 240212 26288
rect 266261 26344 268180 26346
rect 266261 26288 266266 26344
rect 266322 26288 268180 26344
rect 266261 26286 268180 26288
rect 293861 26344 296148 26346
rect 293861 26288 293866 26344
rect 293922 26288 296148 26344
rect 293861 26286 296148 26288
rect 322841 26344 324116 26346
rect 322841 26288 322846 26344
rect 322902 26288 324116 26344
rect 322841 26286 324116 26288
rect 350441 26344 352084 26346
rect 350441 26288 350446 26344
rect 350502 26288 352084 26344
rect 350441 26286 352084 26288
rect 378041 26344 380052 26346
rect 378041 26288 378046 26344
rect 378102 26288 380052 26344
rect 378041 26286 380052 26288
rect 405641 26344 408204 26346
rect 405641 26288 405646 26344
rect 405702 26288 408204 26344
rect 405641 26286 408204 26288
rect 434621 26344 436172 26346
rect 434621 26288 434626 26344
rect 434682 26288 436172 26344
rect 434621 26286 436172 26288
rect 462221 26344 464140 26346
rect 462221 26288 462226 26344
rect 462282 26288 464140 26344
rect 462221 26286 464140 26288
rect 489821 26344 492108 26346
rect 489821 26288 489826 26344
rect 489882 26288 492108 26344
rect 489821 26286 492108 26288
rect 518801 26344 520076 26346
rect 518801 26288 518806 26344
rect 518862 26288 520076 26344
rect 518801 26286 520076 26288
rect 546401 26344 548044 26346
rect 546401 26288 546406 26344
rect 546462 26288 548044 26344
rect 546401 26286 548044 26288
rect 13537 26283 13603 26286
rect 97901 26283 97967 26286
rect 126881 26283 126947 26286
rect 154481 26283 154547 26286
rect 182081 26283 182147 26286
rect 209681 26283 209747 26286
rect 238661 26283 238727 26286
rect 266261 26283 266327 26286
rect 293861 26283 293927 26286
rect 322841 26283 322907 26286
rect 350441 26283 350507 26286
rect 378041 26283 378107 26286
rect 405641 26283 405707 26286
rect 434621 26283 434687 26286
rect 462221 26283 462287 26286
rect 489821 26283 489887 26286
rect 518801 26283 518867 26286
rect 546401 26283 546467 26286
rect 205633 25938 205699 25941
rect 203934 25936 205699 25938
rect 203934 25880 205638 25936
rect 205694 25880 205699 25936
rect 203934 25878 205699 25880
rect 93853 25666 93919 25669
rect 121453 25666 121519 25669
rect 149053 25666 149119 25669
rect 178033 25666 178099 25669
rect 91908 25664 93919 25666
rect 91908 25608 93858 25664
rect 93914 25608 93919 25664
rect 91908 25606 93919 25608
rect 119876 25664 121519 25666
rect 119876 25608 121458 25664
rect 121514 25608 121519 25664
rect 119876 25606 121519 25608
rect 147844 25664 149119 25666
rect 147844 25608 149058 25664
rect 149114 25608 149119 25664
rect 147844 25606 149119 25608
rect 175812 25664 178099 25666
rect 175812 25608 178038 25664
rect 178094 25608 178099 25664
rect 203934 25636 203994 25878
rect 205633 25875 205699 25878
rect 233233 25666 233299 25669
rect 262213 25666 262279 25669
rect 289813 25666 289879 25669
rect 317413 25666 317479 25669
rect 345013 25666 345079 25669
rect 373993 25666 374059 25669
rect 401593 25666 401659 25669
rect 429285 25666 429351 25669
rect 458173 25666 458239 25669
rect 485773 25666 485839 25669
rect 513373 25666 513439 25669
rect 542353 25666 542419 25669
rect 569953 25666 570019 25669
rect 231932 25664 233299 25666
rect 175812 25606 178099 25608
rect 231932 25608 233238 25664
rect 233294 25608 233299 25664
rect 231932 25606 233299 25608
rect 259900 25664 262279 25666
rect 259900 25608 262218 25664
rect 262274 25608 262279 25664
rect 259900 25606 262279 25608
rect 287868 25664 289879 25666
rect 287868 25608 289818 25664
rect 289874 25608 289879 25664
rect 287868 25606 289879 25608
rect 315836 25664 317479 25666
rect 315836 25608 317418 25664
rect 317474 25608 317479 25664
rect 315836 25606 317479 25608
rect 343804 25664 345079 25666
rect 343804 25608 345018 25664
rect 345074 25608 345079 25664
rect 343804 25606 345079 25608
rect 371956 25664 374059 25666
rect 371956 25608 373998 25664
rect 374054 25608 374059 25664
rect 371956 25606 374059 25608
rect 399924 25664 401659 25666
rect 399924 25608 401598 25664
rect 401654 25608 401659 25664
rect 399924 25606 401659 25608
rect 427892 25664 429351 25666
rect 427892 25608 429290 25664
rect 429346 25608 429351 25664
rect 427892 25606 429351 25608
rect 455860 25664 458239 25666
rect 455860 25608 458178 25664
rect 458234 25608 458239 25664
rect 455860 25606 458239 25608
rect 483828 25664 485839 25666
rect 483828 25608 485778 25664
rect 485834 25608 485839 25664
rect 483828 25606 485839 25608
rect 511796 25664 513439 25666
rect 511796 25608 513378 25664
rect 513434 25608 513439 25664
rect 511796 25606 513439 25608
rect 539948 25664 542419 25666
rect 539948 25608 542358 25664
rect 542414 25608 542419 25664
rect 539948 25606 542419 25608
rect 567916 25664 570019 25666
rect 567916 25608 569958 25664
rect 570014 25608 570019 25664
rect 567916 25606 570019 25608
rect 93853 25603 93919 25606
rect 121453 25603 121519 25606
rect 149053 25603 149119 25606
rect 178033 25603 178099 25606
rect 233233 25603 233299 25606
rect 262213 25603 262279 25606
rect 289813 25603 289879 25606
rect 317413 25603 317479 25606
rect 345013 25603 345079 25606
rect 373993 25603 374059 25606
rect 401593 25603 401659 25606
rect 429285 25603 429351 25606
rect 458173 25603 458239 25606
rect 485773 25603 485839 25606
rect 513373 25603 513439 25606
rect 542353 25603 542419 25606
rect 569953 25603 570019 25606
rect 64413 24986 64479 24989
rect 61916 24984 64479 24986
rect 61916 24928 64418 24984
rect 64474 24928 64479 24984
rect 61916 24926 64479 24928
rect 64413 24923 64479 24926
rect 13721 24170 13787 24173
rect 13721 24168 16100 24170
rect 13721 24112 13726 24168
rect 13782 24112 16100 24168
rect 13721 24110 16100 24112
rect 13721 24107 13787 24110
rect 64137 23626 64203 23629
rect 61916 23624 64203 23626
rect 61916 23568 64142 23624
rect 64198 23568 64203 23624
rect 61916 23566 64203 23568
rect 64137 23563 64203 23566
rect 12433 22946 12499 22949
rect 12433 22944 16100 22946
rect 12433 22888 12438 22944
rect 12494 22888 16100 22944
rect 12433 22886 16100 22888
rect 12433 22883 12499 22886
rect 63493 21450 63559 21453
rect 61916 21448 63559 21450
rect 61916 21392 63498 21448
rect 63554 21392 63559 21448
rect 61916 21390 63559 21392
rect 63493 21387 63559 21390
rect 12433 20906 12499 20909
rect 12433 20904 16100 20906
rect 12433 20848 12438 20904
rect 12494 20848 16100 20904
rect 12433 20846 16100 20848
rect 12433 20843 12499 20846
rect 64045 20226 64111 20229
rect 61916 20224 64111 20226
rect 61916 20168 64050 20224
rect 64106 20168 64111 20224
rect 61916 20166 64111 20168
rect 64045 20163 64111 20166
rect 583520 19668 584960 19908
rect 12617 19546 12683 19549
rect 12617 19544 16100 19546
rect -960 19410 480 19500
rect 12617 19488 12622 19544
rect 12678 19488 16100 19544
rect 12617 19486 16100 19488
rect 12617 19483 12683 19486
rect 3785 19410 3851 19413
rect -960 19408 3851 19410
rect -960 19352 3790 19408
rect 3846 19352 3851 19408
rect -960 19350 3851 19352
rect -960 19260 480 19350
rect 3785 19347 3851 19350
rect 64321 18186 64387 18189
rect 61916 18184 64387 18186
rect 61916 18128 64326 18184
rect 64382 18128 64387 18184
rect 61916 18126 64387 18128
rect 64321 18123 64387 18126
rect 12433 17506 12499 17509
rect 12433 17504 16100 17506
rect 12433 17448 12438 17504
rect 12494 17448 16100 17504
rect 12433 17446 16100 17448
rect 12433 17443 12499 17446
rect 64505 16826 64571 16829
rect 61916 16824 64571 16826
rect 61916 16768 64510 16824
rect 64566 16768 64571 16824
rect 61916 16766 64571 16768
rect 64505 16763 64571 16766
rect 48037 16556 48103 16557
rect 48037 16554 48084 16556
rect 47992 16552 48084 16554
rect 47992 16496 48042 16552
rect 47992 16494 48084 16496
rect 48037 16492 48084 16494
rect 48148 16492 48154 16556
rect 48037 16491 48103 16492
rect 59813 13562 59879 13565
rect 580574 13562 580580 13564
rect 59813 13560 580580 13562
rect 59813 13504 59818 13560
rect 59874 13504 580580 13560
rect 59813 13502 580580 13504
rect 59813 13499 59879 13502
rect 580574 13500 580580 13502
rect 580644 13500 580650 13564
rect 61101 13426 61167 13429
rect 580206 13426 580212 13428
rect 61101 13424 580212 13426
rect 61101 13368 61106 13424
rect 61162 13368 580212 13424
rect 61101 13366 580212 13368
rect 61101 13363 61167 13366
rect 580206 13364 580212 13366
rect 580276 13364 580282 13428
rect 19241 13290 19307 13293
rect 518157 13290 518223 13293
rect 19241 13288 518223 13290
rect 19241 13232 19246 13288
rect 19302 13232 518162 13288
rect 518218 13232 518223 13288
rect 19241 13230 518223 13232
rect 19241 13227 19307 13230
rect 518157 13227 518223 13230
rect 45001 13154 45067 13157
rect 580390 13154 580396 13156
rect 45001 13152 580396 13154
rect 45001 13096 45006 13152
rect 45062 13096 580396 13152
rect 45001 13094 580396 13096
rect 45001 13091 45067 13094
rect 580390 13092 580396 13094
rect 580460 13092 580466 13156
rect -960 6490 480 6580
rect -960 6430 674 6490
rect 583520 6476 584960 6716
rect -960 6354 480 6430
rect 614 6354 674 6430
rect -960 6340 674 6354
rect 246 6294 674 6340
rect 246 5810 306 6294
rect 246 5750 6930 5810
rect 6870 5674 6930 5750
rect 42742 5674 42748 5676
rect 6870 5614 42748 5674
rect 42742 5612 42748 5614
rect 42812 5612 42818 5676
<< via3 >>
rect 580212 670652 580276 670716
rect 580396 643996 580460 644060
rect 580580 617476 580644 617540
rect 580764 564300 580828 564364
rect 48084 42060 48148 42124
rect 580764 37844 580828 37908
rect 42748 35260 42812 35324
rect 48084 16552 48148 16556
rect 48084 16496 48098 16552
rect 48098 16496 48148 16552
rect 48084 16492 48148 16496
rect 580580 13500 580644 13564
rect 580212 13364 580276 13428
rect 580396 13092 580460 13156
rect 42748 5612 42812 5676
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 -7066 -8106 711002
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 -6106 -7146 710042
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 -5146 -6186 709082
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 -4186 -5226 708122
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 -3226 -4266 707162
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 -2266 -3306 706202
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 698454 -2346 705242
rect 37994 705798 38614 711590
rect 37994 705562 38026 705798
rect 38262 705562 38346 705798
rect 38582 705562 38614 705798
rect 37994 705478 38614 705562
rect 37994 705242 38026 705478
rect 38262 705242 38346 705478
rect 38582 705242 38614 705478
rect -2966 698218 -2934 698454
rect -2698 698218 -2614 698454
rect -2378 698218 -2346 698454
rect -2966 698134 -2346 698218
rect -2966 697898 -2934 698134
rect -2698 697898 -2614 698134
rect -2378 697898 -2346 698134
rect -2966 671454 -2346 697898
rect -2966 671218 -2934 671454
rect -2698 671218 -2614 671454
rect -2378 671218 -2346 671454
rect -2966 671134 -2346 671218
rect -2966 670898 -2934 671134
rect -2698 670898 -2614 671134
rect -2378 670898 -2346 671134
rect -2966 644454 -2346 670898
rect -2966 644218 -2934 644454
rect -2698 644218 -2614 644454
rect -2378 644218 -2346 644454
rect -2966 644134 -2346 644218
rect -2966 643898 -2934 644134
rect -2698 643898 -2614 644134
rect -2378 643898 -2346 644134
rect -2966 617454 -2346 643898
rect -2966 617218 -2934 617454
rect -2698 617218 -2614 617454
rect -2378 617218 -2346 617454
rect -2966 617134 -2346 617218
rect -2966 616898 -2934 617134
rect -2698 616898 -2614 617134
rect -2378 616898 -2346 617134
rect -2966 590454 -2346 616898
rect -2966 590218 -2934 590454
rect -2698 590218 -2614 590454
rect -2378 590218 -2346 590454
rect -2966 590134 -2346 590218
rect -2966 589898 -2934 590134
rect -2698 589898 -2614 590134
rect -2378 589898 -2346 590134
rect -2966 563454 -2346 589898
rect -2966 563218 -2934 563454
rect -2698 563218 -2614 563454
rect -2378 563218 -2346 563454
rect -2966 563134 -2346 563218
rect -2966 562898 -2934 563134
rect -2698 562898 -2614 563134
rect -2378 562898 -2346 563134
rect -2966 536454 -2346 562898
rect -2966 536218 -2934 536454
rect -2698 536218 -2614 536454
rect -2378 536218 -2346 536454
rect -2966 536134 -2346 536218
rect -2966 535898 -2934 536134
rect -2698 535898 -2614 536134
rect -2378 535898 -2346 536134
rect -2966 509454 -2346 535898
rect -2966 509218 -2934 509454
rect -2698 509218 -2614 509454
rect -2378 509218 -2346 509454
rect -2966 509134 -2346 509218
rect -2966 508898 -2934 509134
rect -2698 508898 -2614 509134
rect -2378 508898 -2346 509134
rect -2966 482454 -2346 508898
rect -2966 482218 -2934 482454
rect -2698 482218 -2614 482454
rect -2378 482218 -2346 482454
rect -2966 482134 -2346 482218
rect -2966 481898 -2934 482134
rect -2698 481898 -2614 482134
rect -2378 481898 -2346 482134
rect -2966 455454 -2346 481898
rect -2966 455218 -2934 455454
rect -2698 455218 -2614 455454
rect -2378 455218 -2346 455454
rect -2966 455134 -2346 455218
rect -2966 454898 -2934 455134
rect -2698 454898 -2614 455134
rect -2378 454898 -2346 455134
rect -2966 428454 -2346 454898
rect -2966 428218 -2934 428454
rect -2698 428218 -2614 428454
rect -2378 428218 -2346 428454
rect -2966 428134 -2346 428218
rect -2966 427898 -2934 428134
rect -2698 427898 -2614 428134
rect -2378 427898 -2346 428134
rect -2966 401454 -2346 427898
rect -2966 401218 -2934 401454
rect -2698 401218 -2614 401454
rect -2378 401218 -2346 401454
rect -2966 401134 -2346 401218
rect -2966 400898 -2934 401134
rect -2698 400898 -2614 401134
rect -2378 400898 -2346 401134
rect -2966 374454 -2346 400898
rect -2966 374218 -2934 374454
rect -2698 374218 -2614 374454
rect -2378 374218 -2346 374454
rect -2966 374134 -2346 374218
rect -2966 373898 -2934 374134
rect -2698 373898 -2614 374134
rect -2378 373898 -2346 374134
rect -2966 347454 -2346 373898
rect -2966 347218 -2934 347454
rect -2698 347218 -2614 347454
rect -2378 347218 -2346 347454
rect -2966 347134 -2346 347218
rect -2966 346898 -2934 347134
rect -2698 346898 -2614 347134
rect -2378 346898 -2346 347134
rect -2966 320454 -2346 346898
rect -2966 320218 -2934 320454
rect -2698 320218 -2614 320454
rect -2378 320218 -2346 320454
rect -2966 320134 -2346 320218
rect -2966 319898 -2934 320134
rect -2698 319898 -2614 320134
rect -2378 319898 -2346 320134
rect -2966 293454 -2346 319898
rect -2966 293218 -2934 293454
rect -2698 293218 -2614 293454
rect -2378 293218 -2346 293454
rect -2966 293134 -2346 293218
rect -2966 292898 -2934 293134
rect -2698 292898 -2614 293134
rect -2378 292898 -2346 293134
rect -2966 266454 -2346 292898
rect -2966 266218 -2934 266454
rect -2698 266218 -2614 266454
rect -2378 266218 -2346 266454
rect -2966 266134 -2346 266218
rect -2966 265898 -2934 266134
rect -2698 265898 -2614 266134
rect -2378 265898 -2346 266134
rect -2966 239454 -2346 265898
rect -2966 239218 -2934 239454
rect -2698 239218 -2614 239454
rect -2378 239218 -2346 239454
rect -2966 239134 -2346 239218
rect -2966 238898 -2934 239134
rect -2698 238898 -2614 239134
rect -2378 238898 -2346 239134
rect -2966 212454 -2346 238898
rect -2966 212218 -2934 212454
rect -2698 212218 -2614 212454
rect -2378 212218 -2346 212454
rect -2966 212134 -2346 212218
rect -2966 211898 -2934 212134
rect -2698 211898 -2614 212134
rect -2378 211898 -2346 212134
rect -2966 185454 -2346 211898
rect -2966 185218 -2934 185454
rect -2698 185218 -2614 185454
rect -2378 185218 -2346 185454
rect -2966 185134 -2346 185218
rect -2966 184898 -2934 185134
rect -2698 184898 -2614 185134
rect -2378 184898 -2346 185134
rect -2966 158454 -2346 184898
rect -2966 158218 -2934 158454
rect -2698 158218 -2614 158454
rect -2378 158218 -2346 158454
rect -2966 158134 -2346 158218
rect -2966 157898 -2934 158134
rect -2698 157898 -2614 158134
rect -2378 157898 -2346 158134
rect -2966 131454 -2346 157898
rect -2966 131218 -2934 131454
rect -2698 131218 -2614 131454
rect -2378 131218 -2346 131454
rect -2966 131134 -2346 131218
rect -2966 130898 -2934 131134
rect -2698 130898 -2614 131134
rect -2378 130898 -2346 131134
rect -2966 104454 -2346 130898
rect -2966 104218 -2934 104454
rect -2698 104218 -2614 104454
rect -2378 104218 -2346 104454
rect -2966 104134 -2346 104218
rect -2966 103898 -2934 104134
rect -2698 103898 -2614 104134
rect -2378 103898 -2346 104134
rect -2966 77454 -2346 103898
rect -2966 77218 -2934 77454
rect -2698 77218 -2614 77454
rect -2378 77218 -2346 77454
rect -2966 77134 -2346 77218
rect -2966 76898 -2934 77134
rect -2698 76898 -2614 77134
rect -2378 76898 -2346 77134
rect -2966 50454 -2346 76898
rect -2966 50218 -2934 50454
rect -2698 50218 -2614 50454
rect -2378 50218 -2346 50454
rect -2966 50134 -2346 50218
rect -2966 49898 -2934 50134
rect -2698 49898 -2614 50134
rect -2378 49898 -2346 50134
rect -2966 23454 -2346 49898
rect -2966 23218 -2934 23454
rect -2698 23218 -2614 23454
rect -2378 23218 -2346 23454
rect -2966 23134 -2346 23218
rect -2966 22898 -2934 23134
rect -2698 22898 -2614 23134
rect -2378 22898 -2346 23134
rect -2966 -1306 -2346 22898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 701829 -1386 704282
rect -2006 701593 -1974 701829
rect -1738 701593 -1654 701829
rect -1418 701593 -1386 701829
rect -2006 701509 -1386 701593
rect -2006 701273 -1974 701509
rect -1738 701273 -1654 701509
rect -1418 701273 -1386 701509
rect -2006 674829 -1386 701273
rect 37994 698454 38614 705242
rect 37994 698218 38026 698454
rect 38262 698218 38346 698454
rect 38582 698218 38614 698454
rect 37994 698134 38614 698218
rect 37994 697898 38026 698134
rect 38262 697898 38346 698134
rect 38582 697898 38614 698134
rect 37994 686000 38614 697898
rect 41494 704838 42114 711590
rect 41494 704602 41526 704838
rect 41762 704602 41846 704838
rect 42082 704602 42114 704838
rect 41494 704518 42114 704602
rect 41494 704282 41526 704518
rect 41762 704282 41846 704518
rect 42082 704282 42114 704518
rect 41494 701829 42114 704282
rect 41494 701593 41526 701829
rect 41762 701593 41846 701829
rect 42082 701593 42114 701829
rect 41494 701509 42114 701593
rect 41494 701273 41526 701509
rect 41762 701273 41846 701509
rect 42082 701273 42114 701509
rect 41494 686000 42114 701273
rect 65994 705798 66614 711590
rect 65994 705562 66026 705798
rect 66262 705562 66346 705798
rect 66582 705562 66614 705798
rect 65994 705478 66614 705562
rect 65994 705242 66026 705478
rect 66262 705242 66346 705478
rect 66582 705242 66614 705478
rect 65994 698454 66614 705242
rect 65994 698218 66026 698454
rect 66262 698218 66346 698454
rect 66582 698218 66614 698454
rect 65994 698134 66614 698218
rect 65994 697898 66026 698134
rect 66262 697898 66346 698134
rect 66582 697898 66614 698134
rect 65994 686000 66614 697898
rect 69494 704838 70114 711590
rect 69494 704602 69526 704838
rect 69762 704602 69846 704838
rect 70082 704602 70114 704838
rect 69494 704518 70114 704602
rect 69494 704282 69526 704518
rect 69762 704282 69846 704518
rect 70082 704282 70114 704518
rect 69494 701829 70114 704282
rect 69494 701593 69526 701829
rect 69762 701593 69846 701829
rect 70082 701593 70114 701829
rect 69494 701509 70114 701593
rect 69494 701273 69526 701509
rect 69762 701273 69846 701509
rect 70082 701273 70114 701509
rect 69494 686000 70114 701273
rect 93994 705798 94614 711590
rect 93994 705562 94026 705798
rect 94262 705562 94346 705798
rect 94582 705562 94614 705798
rect 93994 705478 94614 705562
rect 93994 705242 94026 705478
rect 94262 705242 94346 705478
rect 94582 705242 94614 705478
rect 93994 698454 94614 705242
rect 93994 698218 94026 698454
rect 94262 698218 94346 698454
rect 94582 698218 94614 698454
rect 93994 698134 94614 698218
rect 93994 697898 94026 698134
rect 94262 697898 94346 698134
rect 94582 697898 94614 698134
rect 93994 686000 94614 697898
rect 97494 704838 98114 711590
rect 97494 704602 97526 704838
rect 97762 704602 97846 704838
rect 98082 704602 98114 704838
rect 97494 704518 98114 704602
rect 97494 704282 97526 704518
rect 97762 704282 97846 704518
rect 98082 704282 98114 704518
rect 97494 701829 98114 704282
rect 97494 701593 97526 701829
rect 97762 701593 97846 701829
rect 98082 701593 98114 701829
rect 97494 701509 98114 701593
rect 97494 701273 97526 701509
rect 97762 701273 97846 701509
rect 98082 701273 98114 701509
rect 97494 686000 98114 701273
rect 121994 705798 122614 711590
rect 121994 705562 122026 705798
rect 122262 705562 122346 705798
rect 122582 705562 122614 705798
rect 121994 705478 122614 705562
rect 121994 705242 122026 705478
rect 122262 705242 122346 705478
rect 122582 705242 122614 705478
rect 121994 698454 122614 705242
rect 121994 698218 122026 698454
rect 122262 698218 122346 698454
rect 122582 698218 122614 698454
rect 121994 698134 122614 698218
rect 121994 697898 122026 698134
rect 122262 697898 122346 698134
rect 122582 697898 122614 698134
rect 121994 686000 122614 697898
rect 125494 704838 126114 711590
rect 125494 704602 125526 704838
rect 125762 704602 125846 704838
rect 126082 704602 126114 704838
rect 125494 704518 126114 704602
rect 125494 704282 125526 704518
rect 125762 704282 125846 704518
rect 126082 704282 126114 704518
rect 125494 701829 126114 704282
rect 125494 701593 125526 701829
rect 125762 701593 125846 701829
rect 126082 701593 126114 701829
rect 125494 701509 126114 701593
rect 125494 701273 125526 701509
rect 125762 701273 125846 701509
rect 126082 701273 126114 701509
rect 125494 686000 126114 701273
rect 149994 705798 150614 711590
rect 149994 705562 150026 705798
rect 150262 705562 150346 705798
rect 150582 705562 150614 705798
rect 149994 705478 150614 705562
rect 149994 705242 150026 705478
rect 150262 705242 150346 705478
rect 150582 705242 150614 705478
rect 149994 698454 150614 705242
rect 149994 698218 150026 698454
rect 150262 698218 150346 698454
rect 150582 698218 150614 698454
rect 149994 698134 150614 698218
rect 149994 697898 150026 698134
rect 150262 697898 150346 698134
rect 150582 697898 150614 698134
rect 149994 686000 150614 697898
rect 153494 704838 154114 711590
rect 153494 704602 153526 704838
rect 153762 704602 153846 704838
rect 154082 704602 154114 704838
rect 153494 704518 154114 704602
rect 153494 704282 153526 704518
rect 153762 704282 153846 704518
rect 154082 704282 154114 704518
rect 153494 701829 154114 704282
rect 153494 701593 153526 701829
rect 153762 701593 153846 701829
rect 154082 701593 154114 701829
rect 153494 701509 154114 701593
rect 153494 701273 153526 701509
rect 153762 701273 153846 701509
rect 154082 701273 154114 701509
rect 153494 686000 154114 701273
rect 177994 705798 178614 711590
rect 177994 705562 178026 705798
rect 178262 705562 178346 705798
rect 178582 705562 178614 705798
rect 177994 705478 178614 705562
rect 177994 705242 178026 705478
rect 178262 705242 178346 705478
rect 178582 705242 178614 705478
rect 177994 698454 178614 705242
rect 177994 698218 178026 698454
rect 178262 698218 178346 698454
rect 178582 698218 178614 698454
rect 177994 698134 178614 698218
rect 177994 697898 178026 698134
rect 178262 697898 178346 698134
rect 178582 697898 178614 698134
rect 177994 686000 178614 697898
rect 181494 704838 182114 711590
rect 181494 704602 181526 704838
rect 181762 704602 181846 704838
rect 182082 704602 182114 704838
rect 181494 704518 182114 704602
rect 181494 704282 181526 704518
rect 181762 704282 181846 704518
rect 182082 704282 182114 704518
rect 181494 701829 182114 704282
rect 181494 701593 181526 701829
rect 181762 701593 181846 701829
rect 182082 701593 182114 701829
rect 181494 701509 182114 701593
rect 181494 701273 181526 701509
rect 181762 701273 181846 701509
rect 182082 701273 182114 701509
rect 181494 686000 182114 701273
rect 205994 705798 206614 711590
rect 205994 705562 206026 705798
rect 206262 705562 206346 705798
rect 206582 705562 206614 705798
rect 205994 705478 206614 705562
rect 205994 705242 206026 705478
rect 206262 705242 206346 705478
rect 206582 705242 206614 705478
rect 205994 698454 206614 705242
rect 205994 698218 206026 698454
rect 206262 698218 206346 698454
rect 206582 698218 206614 698454
rect 205994 698134 206614 698218
rect 205994 697898 206026 698134
rect 206262 697898 206346 698134
rect 206582 697898 206614 698134
rect 205994 686000 206614 697898
rect 209494 704838 210114 711590
rect 209494 704602 209526 704838
rect 209762 704602 209846 704838
rect 210082 704602 210114 704838
rect 209494 704518 210114 704602
rect 209494 704282 209526 704518
rect 209762 704282 209846 704518
rect 210082 704282 210114 704518
rect 209494 701829 210114 704282
rect 209494 701593 209526 701829
rect 209762 701593 209846 701829
rect 210082 701593 210114 701829
rect 209494 701509 210114 701593
rect 209494 701273 209526 701509
rect 209762 701273 209846 701509
rect 210082 701273 210114 701509
rect 209494 686000 210114 701273
rect 233994 705798 234614 711590
rect 233994 705562 234026 705798
rect 234262 705562 234346 705798
rect 234582 705562 234614 705798
rect 233994 705478 234614 705562
rect 233994 705242 234026 705478
rect 234262 705242 234346 705478
rect 234582 705242 234614 705478
rect 233994 698454 234614 705242
rect 233994 698218 234026 698454
rect 234262 698218 234346 698454
rect 234582 698218 234614 698454
rect 233994 698134 234614 698218
rect 233994 697898 234026 698134
rect 234262 697898 234346 698134
rect 234582 697898 234614 698134
rect 233994 686000 234614 697898
rect 237494 704838 238114 711590
rect 237494 704602 237526 704838
rect 237762 704602 237846 704838
rect 238082 704602 238114 704838
rect 237494 704518 238114 704602
rect 237494 704282 237526 704518
rect 237762 704282 237846 704518
rect 238082 704282 238114 704518
rect 237494 701829 238114 704282
rect 237494 701593 237526 701829
rect 237762 701593 237846 701829
rect 238082 701593 238114 701829
rect 237494 701509 238114 701593
rect 237494 701273 237526 701509
rect 237762 701273 237846 701509
rect 238082 701273 238114 701509
rect 237494 686000 238114 701273
rect 261994 705798 262614 711590
rect 261994 705562 262026 705798
rect 262262 705562 262346 705798
rect 262582 705562 262614 705798
rect 261994 705478 262614 705562
rect 261994 705242 262026 705478
rect 262262 705242 262346 705478
rect 262582 705242 262614 705478
rect 261994 698454 262614 705242
rect 261994 698218 262026 698454
rect 262262 698218 262346 698454
rect 262582 698218 262614 698454
rect 261994 698134 262614 698218
rect 261994 697898 262026 698134
rect 262262 697898 262346 698134
rect 262582 697898 262614 698134
rect 261994 686000 262614 697898
rect 265494 704838 266114 711590
rect 265494 704602 265526 704838
rect 265762 704602 265846 704838
rect 266082 704602 266114 704838
rect 265494 704518 266114 704602
rect 265494 704282 265526 704518
rect 265762 704282 265846 704518
rect 266082 704282 266114 704518
rect 265494 701829 266114 704282
rect 265494 701593 265526 701829
rect 265762 701593 265846 701829
rect 266082 701593 266114 701829
rect 265494 701509 266114 701593
rect 265494 701273 265526 701509
rect 265762 701273 265846 701509
rect 266082 701273 266114 701509
rect 265494 686000 266114 701273
rect 289994 705798 290614 711590
rect 289994 705562 290026 705798
rect 290262 705562 290346 705798
rect 290582 705562 290614 705798
rect 289994 705478 290614 705562
rect 289994 705242 290026 705478
rect 290262 705242 290346 705478
rect 290582 705242 290614 705478
rect 289994 698454 290614 705242
rect 289994 698218 290026 698454
rect 290262 698218 290346 698454
rect 290582 698218 290614 698454
rect 289994 698134 290614 698218
rect 289994 697898 290026 698134
rect 290262 697898 290346 698134
rect 290582 697898 290614 698134
rect 289994 686000 290614 697898
rect 293494 704838 294114 711590
rect 293494 704602 293526 704838
rect 293762 704602 293846 704838
rect 294082 704602 294114 704838
rect 293494 704518 294114 704602
rect 293494 704282 293526 704518
rect 293762 704282 293846 704518
rect 294082 704282 294114 704518
rect 293494 701829 294114 704282
rect 293494 701593 293526 701829
rect 293762 701593 293846 701829
rect 294082 701593 294114 701829
rect 293494 701509 294114 701593
rect 293494 701273 293526 701509
rect 293762 701273 293846 701509
rect 294082 701273 294114 701509
rect 293494 686000 294114 701273
rect 317994 705798 318614 711590
rect 317994 705562 318026 705798
rect 318262 705562 318346 705798
rect 318582 705562 318614 705798
rect 317994 705478 318614 705562
rect 317994 705242 318026 705478
rect 318262 705242 318346 705478
rect 318582 705242 318614 705478
rect 317994 698454 318614 705242
rect 317994 698218 318026 698454
rect 318262 698218 318346 698454
rect 318582 698218 318614 698454
rect 317994 698134 318614 698218
rect 317994 697898 318026 698134
rect 318262 697898 318346 698134
rect 318582 697898 318614 698134
rect 317994 686000 318614 697898
rect 321494 704838 322114 711590
rect 321494 704602 321526 704838
rect 321762 704602 321846 704838
rect 322082 704602 322114 704838
rect 321494 704518 322114 704602
rect 321494 704282 321526 704518
rect 321762 704282 321846 704518
rect 322082 704282 322114 704518
rect 321494 701829 322114 704282
rect 321494 701593 321526 701829
rect 321762 701593 321846 701829
rect 322082 701593 322114 701829
rect 321494 701509 322114 701593
rect 321494 701273 321526 701509
rect 321762 701273 321846 701509
rect 322082 701273 322114 701509
rect 321494 686000 322114 701273
rect 345994 705798 346614 711590
rect 345994 705562 346026 705798
rect 346262 705562 346346 705798
rect 346582 705562 346614 705798
rect 345994 705478 346614 705562
rect 345994 705242 346026 705478
rect 346262 705242 346346 705478
rect 346582 705242 346614 705478
rect 345994 698454 346614 705242
rect 345994 698218 346026 698454
rect 346262 698218 346346 698454
rect 346582 698218 346614 698454
rect 345994 698134 346614 698218
rect 345994 697898 346026 698134
rect 346262 697898 346346 698134
rect 346582 697898 346614 698134
rect 345994 686000 346614 697898
rect 349494 704838 350114 711590
rect 349494 704602 349526 704838
rect 349762 704602 349846 704838
rect 350082 704602 350114 704838
rect 349494 704518 350114 704602
rect 349494 704282 349526 704518
rect 349762 704282 349846 704518
rect 350082 704282 350114 704518
rect 349494 701829 350114 704282
rect 349494 701593 349526 701829
rect 349762 701593 349846 701829
rect 350082 701593 350114 701829
rect 349494 701509 350114 701593
rect 349494 701273 349526 701509
rect 349762 701273 349846 701509
rect 350082 701273 350114 701509
rect 349494 686000 350114 701273
rect 373994 705798 374614 711590
rect 373994 705562 374026 705798
rect 374262 705562 374346 705798
rect 374582 705562 374614 705798
rect 373994 705478 374614 705562
rect 373994 705242 374026 705478
rect 374262 705242 374346 705478
rect 374582 705242 374614 705478
rect 373994 698454 374614 705242
rect 373994 698218 374026 698454
rect 374262 698218 374346 698454
rect 374582 698218 374614 698454
rect 373994 698134 374614 698218
rect 373994 697898 374026 698134
rect 374262 697898 374346 698134
rect 374582 697898 374614 698134
rect 373994 686000 374614 697898
rect 377494 704838 378114 711590
rect 377494 704602 377526 704838
rect 377762 704602 377846 704838
rect 378082 704602 378114 704838
rect 377494 704518 378114 704602
rect 377494 704282 377526 704518
rect 377762 704282 377846 704518
rect 378082 704282 378114 704518
rect 377494 701829 378114 704282
rect 377494 701593 377526 701829
rect 377762 701593 377846 701829
rect 378082 701593 378114 701829
rect 377494 701509 378114 701593
rect 377494 701273 377526 701509
rect 377762 701273 377846 701509
rect 378082 701273 378114 701509
rect 377494 686000 378114 701273
rect 401994 705798 402614 711590
rect 401994 705562 402026 705798
rect 402262 705562 402346 705798
rect 402582 705562 402614 705798
rect 401994 705478 402614 705562
rect 401994 705242 402026 705478
rect 402262 705242 402346 705478
rect 402582 705242 402614 705478
rect 401994 698454 402614 705242
rect 401994 698218 402026 698454
rect 402262 698218 402346 698454
rect 402582 698218 402614 698454
rect 401994 698134 402614 698218
rect 401994 697898 402026 698134
rect 402262 697898 402346 698134
rect 402582 697898 402614 698134
rect 401994 686000 402614 697898
rect 405494 704838 406114 711590
rect 405494 704602 405526 704838
rect 405762 704602 405846 704838
rect 406082 704602 406114 704838
rect 405494 704518 406114 704602
rect 405494 704282 405526 704518
rect 405762 704282 405846 704518
rect 406082 704282 406114 704518
rect 405494 701829 406114 704282
rect 405494 701593 405526 701829
rect 405762 701593 405846 701829
rect 406082 701593 406114 701829
rect 405494 701509 406114 701593
rect 405494 701273 405526 701509
rect 405762 701273 405846 701509
rect 406082 701273 406114 701509
rect 405494 686000 406114 701273
rect 429994 705798 430614 711590
rect 429994 705562 430026 705798
rect 430262 705562 430346 705798
rect 430582 705562 430614 705798
rect 429994 705478 430614 705562
rect 429994 705242 430026 705478
rect 430262 705242 430346 705478
rect 430582 705242 430614 705478
rect 429994 698454 430614 705242
rect 429994 698218 430026 698454
rect 430262 698218 430346 698454
rect 430582 698218 430614 698454
rect 429994 698134 430614 698218
rect 429994 697898 430026 698134
rect 430262 697898 430346 698134
rect 430582 697898 430614 698134
rect 429994 686000 430614 697898
rect 433494 704838 434114 711590
rect 433494 704602 433526 704838
rect 433762 704602 433846 704838
rect 434082 704602 434114 704838
rect 433494 704518 434114 704602
rect 433494 704282 433526 704518
rect 433762 704282 433846 704518
rect 434082 704282 434114 704518
rect 433494 701829 434114 704282
rect 433494 701593 433526 701829
rect 433762 701593 433846 701829
rect 434082 701593 434114 701829
rect 433494 701509 434114 701593
rect 433494 701273 433526 701509
rect 433762 701273 433846 701509
rect 434082 701273 434114 701509
rect 433494 686000 434114 701273
rect 457994 705798 458614 711590
rect 457994 705562 458026 705798
rect 458262 705562 458346 705798
rect 458582 705562 458614 705798
rect 457994 705478 458614 705562
rect 457994 705242 458026 705478
rect 458262 705242 458346 705478
rect 458582 705242 458614 705478
rect 457994 698454 458614 705242
rect 457994 698218 458026 698454
rect 458262 698218 458346 698454
rect 458582 698218 458614 698454
rect 457994 698134 458614 698218
rect 457994 697898 458026 698134
rect 458262 697898 458346 698134
rect 458582 697898 458614 698134
rect 457994 686000 458614 697898
rect 461494 704838 462114 711590
rect 461494 704602 461526 704838
rect 461762 704602 461846 704838
rect 462082 704602 462114 704838
rect 461494 704518 462114 704602
rect 461494 704282 461526 704518
rect 461762 704282 461846 704518
rect 462082 704282 462114 704518
rect 461494 701829 462114 704282
rect 461494 701593 461526 701829
rect 461762 701593 461846 701829
rect 462082 701593 462114 701829
rect 461494 701509 462114 701593
rect 461494 701273 461526 701509
rect 461762 701273 461846 701509
rect 462082 701273 462114 701509
rect 461494 686000 462114 701273
rect 485994 705798 486614 711590
rect 485994 705562 486026 705798
rect 486262 705562 486346 705798
rect 486582 705562 486614 705798
rect 485994 705478 486614 705562
rect 485994 705242 486026 705478
rect 486262 705242 486346 705478
rect 486582 705242 486614 705478
rect 485994 698454 486614 705242
rect 485994 698218 486026 698454
rect 486262 698218 486346 698454
rect 486582 698218 486614 698454
rect 485994 698134 486614 698218
rect 485994 697898 486026 698134
rect 486262 697898 486346 698134
rect 486582 697898 486614 698134
rect 485994 686000 486614 697898
rect 489494 704838 490114 711590
rect 489494 704602 489526 704838
rect 489762 704602 489846 704838
rect 490082 704602 490114 704838
rect 489494 704518 490114 704602
rect 489494 704282 489526 704518
rect 489762 704282 489846 704518
rect 490082 704282 490114 704518
rect 489494 701829 490114 704282
rect 489494 701593 489526 701829
rect 489762 701593 489846 701829
rect 490082 701593 490114 701829
rect 489494 701509 490114 701593
rect 489494 701273 489526 701509
rect 489762 701273 489846 701509
rect 490082 701273 490114 701509
rect 489494 686000 490114 701273
rect 513994 705798 514614 711590
rect 513994 705562 514026 705798
rect 514262 705562 514346 705798
rect 514582 705562 514614 705798
rect 513994 705478 514614 705562
rect 513994 705242 514026 705478
rect 514262 705242 514346 705478
rect 514582 705242 514614 705478
rect 513994 698454 514614 705242
rect 513994 698218 514026 698454
rect 514262 698218 514346 698454
rect 514582 698218 514614 698454
rect 513994 698134 514614 698218
rect 513994 697898 514026 698134
rect 514262 697898 514346 698134
rect 514582 697898 514614 698134
rect 513994 686000 514614 697898
rect 517494 704838 518114 711590
rect 517494 704602 517526 704838
rect 517762 704602 517846 704838
rect 518082 704602 518114 704838
rect 517494 704518 518114 704602
rect 517494 704282 517526 704518
rect 517762 704282 517846 704518
rect 518082 704282 518114 704518
rect 517494 701829 518114 704282
rect 517494 701593 517526 701829
rect 517762 701593 517846 701829
rect 518082 701593 518114 701829
rect 517494 701509 518114 701593
rect 517494 701273 517526 701509
rect 517762 701273 517846 701509
rect 518082 701273 518114 701509
rect 517494 686000 518114 701273
rect 541994 705798 542614 711590
rect 541994 705562 542026 705798
rect 542262 705562 542346 705798
rect 542582 705562 542614 705798
rect 541994 705478 542614 705562
rect 541994 705242 542026 705478
rect 542262 705242 542346 705478
rect 542582 705242 542614 705478
rect 541994 698454 542614 705242
rect 541994 698218 542026 698454
rect 542262 698218 542346 698454
rect 542582 698218 542614 698454
rect 541994 698134 542614 698218
rect 541994 697898 542026 698134
rect 542262 697898 542346 698134
rect 542582 697898 542614 698134
rect 541994 686000 542614 697898
rect 545494 704838 546114 711590
rect 545494 704602 545526 704838
rect 545762 704602 545846 704838
rect 546082 704602 546114 704838
rect 545494 704518 546114 704602
rect 545494 704282 545526 704518
rect 545762 704282 545846 704518
rect 546082 704282 546114 704518
rect 545494 701829 546114 704282
rect 545494 701593 545526 701829
rect 545762 701593 545846 701829
rect 546082 701593 546114 701829
rect 545494 701509 546114 701593
rect 545494 701273 545526 701509
rect 545762 701273 545846 701509
rect 546082 701273 546114 701509
rect 545494 686000 546114 701273
rect 569994 705798 570614 711590
rect 569994 705562 570026 705798
rect 570262 705562 570346 705798
rect 570582 705562 570614 705798
rect 569994 705478 570614 705562
rect 569994 705242 570026 705478
rect 570262 705242 570346 705478
rect 570582 705242 570614 705478
rect 569994 698454 570614 705242
rect 569994 698218 570026 698454
rect 570262 698218 570346 698454
rect 570582 698218 570614 698454
rect 569994 698134 570614 698218
rect 569994 697898 570026 698134
rect 570262 697898 570346 698134
rect 570582 697898 570614 698134
rect 569994 686000 570614 697898
rect 573494 704838 574114 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 573494 704602 573526 704838
rect 573762 704602 573846 704838
rect 574082 704602 574114 704838
rect 573494 704518 574114 704602
rect 573494 704282 573526 704518
rect 573762 704282 573846 704518
rect 574082 704282 574114 704518
rect 573494 701829 574114 704282
rect 573494 701593 573526 701829
rect 573762 701593 573846 701829
rect 574082 701593 574114 701829
rect 573494 701509 574114 701593
rect 573494 701273 573526 701509
rect 573762 701273 573846 701509
rect 574082 701273 574114 701509
rect -2006 674593 -1974 674829
rect -1738 674593 -1654 674829
rect -1418 674593 -1386 674829
rect -2006 674509 -1386 674593
rect -2006 674273 -1974 674509
rect -1738 674273 -1654 674509
rect -1418 674273 -1386 674509
rect -2006 647829 -1386 674273
rect 19910 674829 20230 674861
rect 19910 674593 19952 674829
rect 20188 674593 20230 674829
rect 19910 674509 20230 674593
rect 19910 674273 19952 674509
rect 20188 674273 20230 674509
rect 19910 674241 20230 674273
rect 25840 674829 26160 674861
rect 25840 674593 25882 674829
rect 26118 674593 26160 674829
rect 25840 674509 26160 674593
rect 25840 674273 25882 674509
rect 26118 674273 26160 674509
rect 25840 674241 26160 674273
rect 31771 674829 32091 674861
rect 31771 674593 31813 674829
rect 32049 674593 32091 674829
rect 31771 674509 32091 674593
rect 31771 674273 31813 674509
rect 32049 674273 32091 674509
rect 31771 674241 32091 674273
rect 47910 674829 48230 674861
rect 47910 674593 47952 674829
rect 48188 674593 48230 674829
rect 47910 674509 48230 674593
rect 47910 674273 47952 674509
rect 48188 674273 48230 674509
rect 47910 674241 48230 674273
rect 53840 674829 54160 674861
rect 53840 674593 53882 674829
rect 54118 674593 54160 674829
rect 53840 674509 54160 674593
rect 53840 674273 53882 674509
rect 54118 674273 54160 674509
rect 53840 674241 54160 674273
rect 59771 674829 60091 674861
rect 59771 674593 59813 674829
rect 60049 674593 60091 674829
rect 59771 674509 60091 674593
rect 59771 674273 59813 674509
rect 60049 674273 60091 674509
rect 59771 674241 60091 674273
rect 75910 674829 76230 674861
rect 75910 674593 75952 674829
rect 76188 674593 76230 674829
rect 75910 674509 76230 674593
rect 75910 674273 75952 674509
rect 76188 674273 76230 674509
rect 75910 674241 76230 674273
rect 81840 674829 82160 674861
rect 81840 674593 81882 674829
rect 82118 674593 82160 674829
rect 81840 674509 82160 674593
rect 81840 674273 81882 674509
rect 82118 674273 82160 674509
rect 81840 674241 82160 674273
rect 87771 674829 88091 674861
rect 87771 674593 87813 674829
rect 88049 674593 88091 674829
rect 87771 674509 88091 674593
rect 87771 674273 87813 674509
rect 88049 674273 88091 674509
rect 87771 674241 88091 674273
rect 103910 674829 104230 674861
rect 103910 674593 103952 674829
rect 104188 674593 104230 674829
rect 103910 674509 104230 674593
rect 103910 674273 103952 674509
rect 104188 674273 104230 674509
rect 103910 674241 104230 674273
rect 109840 674829 110160 674861
rect 109840 674593 109882 674829
rect 110118 674593 110160 674829
rect 109840 674509 110160 674593
rect 109840 674273 109882 674509
rect 110118 674273 110160 674509
rect 109840 674241 110160 674273
rect 115771 674829 116091 674861
rect 115771 674593 115813 674829
rect 116049 674593 116091 674829
rect 115771 674509 116091 674593
rect 115771 674273 115813 674509
rect 116049 674273 116091 674509
rect 115771 674241 116091 674273
rect 131910 674829 132230 674861
rect 131910 674593 131952 674829
rect 132188 674593 132230 674829
rect 131910 674509 132230 674593
rect 131910 674273 131952 674509
rect 132188 674273 132230 674509
rect 131910 674241 132230 674273
rect 137840 674829 138160 674861
rect 137840 674593 137882 674829
rect 138118 674593 138160 674829
rect 137840 674509 138160 674593
rect 137840 674273 137882 674509
rect 138118 674273 138160 674509
rect 137840 674241 138160 674273
rect 143771 674829 144091 674861
rect 143771 674593 143813 674829
rect 144049 674593 144091 674829
rect 143771 674509 144091 674593
rect 143771 674273 143813 674509
rect 144049 674273 144091 674509
rect 143771 674241 144091 674273
rect 159910 674829 160230 674861
rect 159910 674593 159952 674829
rect 160188 674593 160230 674829
rect 159910 674509 160230 674593
rect 159910 674273 159952 674509
rect 160188 674273 160230 674509
rect 159910 674241 160230 674273
rect 165840 674829 166160 674861
rect 165840 674593 165882 674829
rect 166118 674593 166160 674829
rect 165840 674509 166160 674593
rect 165840 674273 165882 674509
rect 166118 674273 166160 674509
rect 165840 674241 166160 674273
rect 171771 674829 172091 674861
rect 171771 674593 171813 674829
rect 172049 674593 172091 674829
rect 171771 674509 172091 674593
rect 171771 674273 171813 674509
rect 172049 674273 172091 674509
rect 171771 674241 172091 674273
rect 187910 674829 188230 674861
rect 187910 674593 187952 674829
rect 188188 674593 188230 674829
rect 187910 674509 188230 674593
rect 187910 674273 187952 674509
rect 188188 674273 188230 674509
rect 187910 674241 188230 674273
rect 193840 674829 194160 674861
rect 193840 674593 193882 674829
rect 194118 674593 194160 674829
rect 193840 674509 194160 674593
rect 193840 674273 193882 674509
rect 194118 674273 194160 674509
rect 193840 674241 194160 674273
rect 199771 674829 200091 674861
rect 199771 674593 199813 674829
rect 200049 674593 200091 674829
rect 199771 674509 200091 674593
rect 199771 674273 199813 674509
rect 200049 674273 200091 674509
rect 199771 674241 200091 674273
rect 215910 674829 216230 674861
rect 215910 674593 215952 674829
rect 216188 674593 216230 674829
rect 215910 674509 216230 674593
rect 215910 674273 215952 674509
rect 216188 674273 216230 674509
rect 215910 674241 216230 674273
rect 221840 674829 222160 674861
rect 221840 674593 221882 674829
rect 222118 674593 222160 674829
rect 221840 674509 222160 674593
rect 221840 674273 221882 674509
rect 222118 674273 222160 674509
rect 221840 674241 222160 674273
rect 227771 674829 228091 674861
rect 227771 674593 227813 674829
rect 228049 674593 228091 674829
rect 227771 674509 228091 674593
rect 227771 674273 227813 674509
rect 228049 674273 228091 674509
rect 227771 674241 228091 674273
rect 243910 674829 244230 674861
rect 243910 674593 243952 674829
rect 244188 674593 244230 674829
rect 243910 674509 244230 674593
rect 243910 674273 243952 674509
rect 244188 674273 244230 674509
rect 243910 674241 244230 674273
rect 249840 674829 250160 674861
rect 249840 674593 249882 674829
rect 250118 674593 250160 674829
rect 249840 674509 250160 674593
rect 249840 674273 249882 674509
rect 250118 674273 250160 674509
rect 249840 674241 250160 674273
rect 255771 674829 256091 674861
rect 255771 674593 255813 674829
rect 256049 674593 256091 674829
rect 255771 674509 256091 674593
rect 255771 674273 255813 674509
rect 256049 674273 256091 674509
rect 255771 674241 256091 674273
rect 271910 674829 272230 674861
rect 271910 674593 271952 674829
rect 272188 674593 272230 674829
rect 271910 674509 272230 674593
rect 271910 674273 271952 674509
rect 272188 674273 272230 674509
rect 271910 674241 272230 674273
rect 277840 674829 278160 674861
rect 277840 674593 277882 674829
rect 278118 674593 278160 674829
rect 277840 674509 278160 674593
rect 277840 674273 277882 674509
rect 278118 674273 278160 674509
rect 277840 674241 278160 674273
rect 283771 674829 284091 674861
rect 283771 674593 283813 674829
rect 284049 674593 284091 674829
rect 283771 674509 284091 674593
rect 283771 674273 283813 674509
rect 284049 674273 284091 674509
rect 283771 674241 284091 674273
rect 299910 674829 300230 674861
rect 299910 674593 299952 674829
rect 300188 674593 300230 674829
rect 299910 674509 300230 674593
rect 299910 674273 299952 674509
rect 300188 674273 300230 674509
rect 299910 674241 300230 674273
rect 305840 674829 306160 674861
rect 305840 674593 305882 674829
rect 306118 674593 306160 674829
rect 305840 674509 306160 674593
rect 305840 674273 305882 674509
rect 306118 674273 306160 674509
rect 305840 674241 306160 674273
rect 311771 674829 312091 674861
rect 311771 674593 311813 674829
rect 312049 674593 312091 674829
rect 311771 674509 312091 674593
rect 311771 674273 311813 674509
rect 312049 674273 312091 674509
rect 311771 674241 312091 674273
rect 327910 674829 328230 674861
rect 327910 674593 327952 674829
rect 328188 674593 328230 674829
rect 327910 674509 328230 674593
rect 327910 674273 327952 674509
rect 328188 674273 328230 674509
rect 327910 674241 328230 674273
rect 333840 674829 334160 674861
rect 333840 674593 333882 674829
rect 334118 674593 334160 674829
rect 333840 674509 334160 674593
rect 333840 674273 333882 674509
rect 334118 674273 334160 674509
rect 333840 674241 334160 674273
rect 339771 674829 340091 674861
rect 339771 674593 339813 674829
rect 340049 674593 340091 674829
rect 339771 674509 340091 674593
rect 339771 674273 339813 674509
rect 340049 674273 340091 674509
rect 339771 674241 340091 674273
rect 355910 674829 356230 674861
rect 355910 674593 355952 674829
rect 356188 674593 356230 674829
rect 355910 674509 356230 674593
rect 355910 674273 355952 674509
rect 356188 674273 356230 674509
rect 355910 674241 356230 674273
rect 361840 674829 362160 674861
rect 361840 674593 361882 674829
rect 362118 674593 362160 674829
rect 361840 674509 362160 674593
rect 361840 674273 361882 674509
rect 362118 674273 362160 674509
rect 361840 674241 362160 674273
rect 367771 674829 368091 674861
rect 367771 674593 367813 674829
rect 368049 674593 368091 674829
rect 367771 674509 368091 674593
rect 367771 674273 367813 674509
rect 368049 674273 368091 674509
rect 367771 674241 368091 674273
rect 383910 674829 384230 674861
rect 383910 674593 383952 674829
rect 384188 674593 384230 674829
rect 383910 674509 384230 674593
rect 383910 674273 383952 674509
rect 384188 674273 384230 674509
rect 383910 674241 384230 674273
rect 389840 674829 390160 674861
rect 389840 674593 389882 674829
rect 390118 674593 390160 674829
rect 389840 674509 390160 674593
rect 389840 674273 389882 674509
rect 390118 674273 390160 674509
rect 389840 674241 390160 674273
rect 395771 674829 396091 674861
rect 395771 674593 395813 674829
rect 396049 674593 396091 674829
rect 395771 674509 396091 674593
rect 395771 674273 395813 674509
rect 396049 674273 396091 674509
rect 395771 674241 396091 674273
rect 411910 674829 412230 674861
rect 411910 674593 411952 674829
rect 412188 674593 412230 674829
rect 411910 674509 412230 674593
rect 411910 674273 411952 674509
rect 412188 674273 412230 674509
rect 411910 674241 412230 674273
rect 417840 674829 418160 674861
rect 417840 674593 417882 674829
rect 418118 674593 418160 674829
rect 417840 674509 418160 674593
rect 417840 674273 417882 674509
rect 418118 674273 418160 674509
rect 417840 674241 418160 674273
rect 423771 674829 424091 674861
rect 423771 674593 423813 674829
rect 424049 674593 424091 674829
rect 423771 674509 424091 674593
rect 423771 674273 423813 674509
rect 424049 674273 424091 674509
rect 423771 674241 424091 674273
rect 439910 674829 440230 674861
rect 439910 674593 439952 674829
rect 440188 674593 440230 674829
rect 439910 674509 440230 674593
rect 439910 674273 439952 674509
rect 440188 674273 440230 674509
rect 439910 674241 440230 674273
rect 445840 674829 446160 674861
rect 445840 674593 445882 674829
rect 446118 674593 446160 674829
rect 445840 674509 446160 674593
rect 445840 674273 445882 674509
rect 446118 674273 446160 674509
rect 445840 674241 446160 674273
rect 451771 674829 452091 674861
rect 451771 674593 451813 674829
rect 452049 674593 452091 674829
rect 451771 674509 452091 674593
rect 451771 674273 451813 674509
rect 452049 674273 452091 674509
rect 451771 674241 452091 674273
rect 467910 674829 468230 674861
rect 467910 674593 467952 674829
rect 468188 674593 468230 674829
rect 467910 674509 468230 674593
rect 467910 674273 467952 674509
rect 468188 674273 468230 674509
rect 467910 674241 468230 674273
rect 473840 674829 474160 674861
rect 473840 674593 473882 674829
rect 474118 674593 474160 674829
rect 473840 674509 474160 674593
rect 473840 674273 473882 674509
rect 474118 674273 474160 674509
rect 473840 674241 474160 674273
rect 479771 674829 480091 674861
rect 479771 674593 479813 674829
rect 480049 674593 480091 674829
rect 479771 674509 480091 674593
rect 479771 674273 479813 674509
rect 480049 674273 480091 674509
rect 479771 674241 480091 674273
rect 495910 674829 496230 674861
rect 495910 674593 495952 674829
rect 496188 674593 496230 674829
rect 495910 674509 496230 674593
rect 495910 674273 495952 674509
rect 496188 674273 496230 674509
rect 495910 674241 496230 674273
rect 501840 674829 502160 674861
rect 501840 674593 501882 674829
rect 502118 674593 502160 674829
rect 501840 674509 502160 674593
rect 501840 674273 501882 674509
rect 502118 674273 502160 674509
rect 501840 674241 502160 674273
rect 507771 674829 508091 674861
rect 507771 674593 507813 674829
rect 508049 674593 508091 674829
rect 507771 674509 508091 674593
rect 507771 674273 507813 674509
rect 508049 674273 508091 674509
rect 507771 674241 508091 674273
rect 523910 674829 524230 674861
rect 523910 674593 523952 674829
rect 524188 674593 524230 674829
rect 523910 674509 524230 674593
rect 523910 674273 523952 674509
rect 524188 674273 524230 674509
rect 523910 674241 524230 674273
rect 529840 674829 530160 674861
rect 529840 674593 529882 674829
rect 530118 674593 530160 674829
rect 529840 674509 530160 674593
rect 529840 674273 529882 674509
rect 530118 674273 530160 674509
rect 529840 674241 530160 674273
rect 535771 674829 536091 674861
rect 535771 674593 535813 674829
rect 536049 674593 536091 674829
rect 535771 674509 536091 674593
rect 535771 674273 535813 674509
rect 536049 674273 536091 674509
rect 535771 674241 536091 674273
rect 551910 674829 552230 674861
rect 551910 674593 551952 674829
rect 552188 674593 552230 674829
rect 551910 674509 552230 674593
rect 551910 674273 551952 674509
rect 552188 674273 552230 674509
rect 551910 674241 552230 674273
rect 557840 674829 558160 674861
rect 557840 674593 557882 674829
rect 558118 674593 558160 674829
rect 557840 674509 558160 674593
rect 557840 674273 557882 674509
rect 558118 674273 558160 674509
rect 557840 674241 558160 674273
rect 563771 674829 564091 674861
rect 563771 674593 563813 674829
rect 564049 674593 564091 674829
rect 563771 674509 564091 674593
rect 563771 674273 563813 674509
rect 564049 674273 564091 674509
rect 563771 674241 564091 674273
rect 573494 674829 574114 701273
rect 573494 674593 573526 674829
rect 573762 674593 573846 674829
rect 574082 674593 574114 674829
rect 573494 674509 574114 674593
rect 573494 674273 573526 674509
rect 573762 674273 573846 674509
rect 574082 674273 574114 674509
rect 22874 671454 23194 671486
rect 22874 671218 22916 671454
rect 23152 671218 23194 671454
rect 22874 671134 23194 671218
rect 22874 670898 22916 671134
rect 23152 670898 23194 671134
rect 22874 670866 23194 670898
rect 28805 671454 29125 671486
rect 28805 671218 28847 671454
rect 29083 671218 29125 671454
rect 28805 671134 29125 671218
rect 28805 670898 28847 671134
rect 29083 670898 29125 671134
rect 28805 670866 29125 670898
rect 50874 671454 51194 671486
rect 50874 671218 50916 671454
rect 51152 671218 51194 671454
rect 50874 671134 51194 671218
rect 50874 670898 50916 671134
rect 51152 670898 51194 671134
rect 50874 670866 51194 670898
rect 56805 671454 57125 671486
rect 56805 671218 56847 671454
rect 57083 671218 57125 671454
rect 56805 671134 57125 671218
rect 56805 670898 56847 671134
rect 57083 670898 57125 671134
rect 56805 670866 57125 670898
rect 78874 671454 79194 671486
rect 78874 671218 78916 671454
rect 79152 671218 79194 671454
rect 78874 671134 79194 671218
rect 78874 670898 78916 671134
rect 79152 670898 79194 671134
rect 78874 670866 79194 670898
rect 84805 671454 85125 671486
rect 84805 671218 84847 671454
rect 85083 671218 85125 671454
rect 84805 671134 85125 671218
rect 84805 670898 84847 671134
rect 85083 670898 85125 671134
rect 84805 670866 85125 670898
rect 106874 671454 107194 671486
rect 106874 671218 106916 671454
rect 107152 671218 107194 671454
rect 106874 671134 107194 671218
rect 106874 670898 106916 671134
rect 107152 670898 107194 671134
rect 106874 670866 107194 670898
rect 112805 671454 113125 671486
rect 112805 671218 112847 671454
rect 113083 671218 113125 671454
rect 112805 671134 113125 671218
rect 112805 670898 112847 671134
rect 113083 670898 113125 671134
rect 112805 670866 113125 670898
rect 134874 671454 135194 671486
rect 134874 671218 134916 671454
rect 135152 671218 135194 671454
rect 134874 671134 135194 671218
rect 134874 670898 134916 671134
rect 135152 670898 135194 671134
rect 134874 670866 135194 670898
rect 140805 671454 141125 671486
rect 140805 671218 140847 671454
rect 141083 671218 141125 671454
rect 140805 671134 141125 671218
rect 140805 670898 140847 671134
rect 141083 670898 141125 671134
rect 140805 670866 141125 670898
rect 162874 671454 163194 671486
rect 162874 671218 162916 671454
rect 163152 671218 163194 671454
rect 162874 671134 163194 671218
rect 162874 670898 162916 671134
rect 163152 670898 163194 671134
rect 162874 670866 163194 670898
rect 168805 671454 169125 671486
rect 168805 671218 168847 671454
rect 169083 671218 169125 671454
rect 168805 671134 169125 671218
rect 168805 670898 168847 671134
rect 169083 670898 169125 671134
rect 168805 670866 169125 670898
rect 190874 671454 191194 671486
rect 190874 671218 190916 671454
rect 191152 671218 191194 671454
rect 190874 671134 191194 671218
rect 190874 670898 190916 671134
rect 191152 670898 191194 671134
rect 190874 670866 191194 670898
rect 196805 671454 197125 671486
rect 196805 671218 196847 671454
rect 197083 671218 197125 671454
rect 196805 671134 197125 671218
rect 196805 670898 196847 671134
rect 197083 670898 197125 671134
rect 196805 670866 197125 670898
rect 218874 671454 219194 671486
rect 218874 671218 218916 671454
rect 219152 671218 219194 671454
rect 218874 671134 219194 671218
rect 218874 670898 218916 671134
rect 219152 670898 219194 671134
rect 218874 670866 219194 670898
rect 224805 671454 225125 671486
rect 224805 671218 224847 671454
rect 225083 671218 225125 671454
rect 224805 671134 225125 671218
rect 224805 670898 224847 671134
rect 225083 670898 225125 671134
rect 224805 670866 225125 670898
rect 246874 671454 247194 671486
rect 246874 671218 246916 671454
rect 247152 671218 247194 671454
rect 246874 671134 247194 671218
rect 246874 670898 246916 671134
rect 247152 670898 247194 671134
rect 246874 670866 247194 670898
rect 252805 671454 253125 671486
rect 252805 671218 252847 671454
rect 253083 671218 253125 671454
rect 252805 671134 253125 671218
rect 252805 670898 252847 671134
rect 253083 670898 253125 671134
rect 252805 670866 253125 670898
rect 274874 671454 275194 671486
rect 274874 671218 274916 671454
rect 275152 671218 275194 671454
rect 274874 671134 275194 671218
rect 274874 670898 274916 671134
rect 275152 670898 275194 671134
rect 274874 670866 275194 670898
rect 280805 671454 281125 671486
rect 280805 671218 280847 671454
rect 281083 671218 281125 671454
rect 280805 671134 281125 671218
rect 280805 670898 280847 671134
rect 281083 670898 281125 671134
rect 280805 670866 281125 670898
rect 302874 671454 303194 671486
rect 302874 671218 302916 671454
rect 303152 671218 303194 671454
rect 302874 671134 303194 671218
rect 302874 670898 302916 671134
rect 303152 670898 303194 671134
rect 302874 670866 303194 670898
rect 308805 671454 309125 671486
rect 308805 671218 308847 671454
rect 309083 671218 309125 671454
rect 308805 671134 309125 671218
rect 308805 670898 308847 671134
rect 309083 670898 309125 671134
rect 308805 670866 309125 670898
rect 330874 671454 331194 671486
rect 330874 671218 330916 671454
rect 331152 671218 331194 671454
rect 330874 671134 331194 671218
rect 330874 670898 330916 671134
rect 331152 670898 331194 671134
rect 330874 670866 331194 670898
rect 336805 671454 337125 671486
rect 336805 671218 336847 671454
rect 337083 671218 337125 671454
rect 336805 671134 337125 671218
rect 336805 670898 336847 671134
rect 337083 670898 337125 671134
rect 336805 670866 337125 670898
rect 358874 671454 359194 671486
rect 358874 671218 358916 671454
rect 359152 671218 359194 671454
rect 358874 671134 359194 671218
rect 358874 670898 358916 671134
rect 359152 670898 359194 671134
rect 358874 670866 359194 670898
rect 364805 671454 365125 671486
rect 364805 671218 364847 671454
rect 365083 671218 365125 671454
rect 364805 671134 365125 671218
rect 364805 670898 364847 671134
rect 365083 670898 365125 671134
rect 364805 670866 365125 670898
rect 386874 671454 387194 671486
rect 386874 671218 386916 671454
rect 387152 671218 387194 671454
rect 386874 671134 387194 671218
rect 386874 670898 386916 671134
rect 387152 670898 387194 671134
rect 386874 670866 387194 670898
rect 392805 671454 393125 671486
rect 392805 671218 392847 671454
rect 393083 671218 393125 671454
rect 392805 671134 393125 671218
rect 392805 670898 392847 671134
rect 393083 670898 393125 671134
rect 392805 670866 393125 670898
rect 414874 671454 415194 671486
rect 414874 671218 414916 671454
rect 415152 671218 415194 671454
rect 414874 671134 415194 671218
rect 414874 670898 414916 671134
rect 415152 670898 415194 671134
rect 414874 670866 415194 670898
rect 420805 671454 421125 671486
rect 420805 671218 420847 671454
rect 421083 671218 421125 671454
rect 420805 671134 421125 671218
rect 420805 670898 420847 671134
rect 421083 670898 421125 671134
rect 420805 670866 421125 670898
rect 442874 671454 443194 671486
rect 442874 671218 442916 671454
rect 443152 671218 443194 671454
rect 442874 671134 443194 671218
rect 442874 670898 442916 671134
rect 443152 670898 443194 671134
rect 442874 670866 443194 670898
rect 448805 671454 449125 671486
rect 448805 671218 448847 671454
rect 449083 671218 449125 671454
rect 448805 671134 449125 671218
rect 448805 670898 448847 671134
rect 449083 670898 449125 671134
rect 448805 670866 449125 670898
rect 470874 671454 471194 671486
rect 470874 671218 470916 671454
rect 471152 671218 471194 671454
rect 470874 671134 471194 671218
rect 470874 670898 470916 671134
rect 471152 670898 471194 671134
rect 470874 670866 471194 670898
rect 476805 671454 477125 671486
rect 476805 671218 476847 671454
rect 477083 671218 477125 671454
rect 476805 671134 477125 671218
rect 476805 670898 476847 671134
rect 477083 670898 477125 671134
rect 476805 670866 477125 670898
rect 498874 671454 499194 671486
rect 498874 671218 498916 671454
rect 499152 671218 499194 671454
rect 498874 671134 499194 671218
rect 498874 670898 498916 671134
rect 499152 670898 499194 671134
rect 498874 670866 499194 670898
rect 504805 671454 505125 671486
rect 504805 671218 504847 671454
rect 505083 671218 505125 671454
rect 504805 671134 505125 671218
rect 504805 670898 504847 671134
rect 505083 670898 505125 671134
rect 504805 670866 505125 670898
rect 526874 671454 527194 671486
rect 526874 671218 526916 671454
rect 527152 671218 527194 671454
rect 526874 671134 527194 671218
rect 526874 670898 526916 671134
rect 527152 670898 527194 671134
rect 526874 670866 527194 670898
rect 532805 671454 533125 671486
rect 532805 671218 532847 671454
rect 533083 671218 533125 671454
rect 532805 671134 533125 671218
rect 532805 670898 532847 671134
rect 533083 670898 533125 671134
rect 532805 670866 533125 670898
rect 554874 671454 555194 671486
rect 554874 671218 554916 671454
rect 555152 671218 555194 671454
rect 554874 671134 555194 671218
rect 554874 670898 554916 671134
rect 555152 670898 555194 671134
rect 554874 670866 555194 670898
rect 560805 671454 561125 671486
rect 560805 671218 560847 671454
rect 561083 671218 561125 671454
rect 560805 671134 561125 671218
rect 560805 670898 560847 671134
rect 561083 670898 561125 671134
rect 560805 670866 561125 670898
rect -2006 647593 -1974 647829
rect -1738 647593 -1654 647829
rect -1418 647593 -1386 647829
rect -2006 647509 -1386 647593
rect -2006 647273 -1974 647509
rect -1738 647273 -1654 647509
rect -1418 647273 -1386 647509
rect -2006 620829 -1386 647273
rect 19909 647829 20229 647861
rect 19909 647593 19951 647829
rect 20187 647593 20229 647829
rect 19909 647509 20229 647593
rect 19909 647273 19951 647509
rect 20187 647273 20229 647509
rect 19909 647241 20229 647273
rect 25840 647829 26160 647861
rect 25840 647593 25882 647829
rect 26118 647593 26160 647829
rect 25840 647509 26160 647593
rect 25840 647273 25882 647509
rect 26118 647273 26160 647509
rect 25840 647241 26160 647273
rect 31770 647829 32090 647861
rect 31770 647593 31812 647829
rect 32048 647593 32090 647829
rect 31770 647509 32090 647593
rect 31770 647273 31812 647509
rect 32048 647273 32090 647509
rect 31770 647241 32090 647273
rect 47909 647829 48229 647861
rect 47909 647593 47951 647829
rect 48187 647593 48229 647829
rect 47909 647509 48229 647593
rect 47909 647273 47951 647509
rect 48187 647273 48229 647509
rect 47909 647241 48229 647273
rect 53840 647829 54160 647861
rect 53840 647593 53882 647829
rect 54118 647593 54160 647829
rect 53840 647509 54160 647593
rect 53840 647273 53882 647509
rect 54118 647273 54160 647509
rect 53840 647241 54160 647273
rect 59770 647829 60090 647861
rect 59770 647593 59812 647829
rect 60048 647593 60090 647829
rect 59770 647509 60090 647593
rect 59770 647273 59812 647509
rect 60048 647273 60090 647509
rect 59770 647241 60090 647273
rect 75909 647829 76229 647861
rect 75909 647593 75951 647829
rect 76187 647593 76229 647829
rect 75909 647509 76229 647593
rect 75909 647273 75951 647509
rect 76187 647273 76229 647509
rect 75909 647241 76229 647273
rect 81840 647829 82160 647861
rect 81840 647593 81882 647829
rect 82118 647593 82160 647829
rect 81840 647509 82160 647593
rect 81840 647273 81882 647509
rect 82118 647273 82160 647509
rect 81840 647241 82160 647273
rect 87770 647829 88090 647861
rect 87770 647593 87812 647829
rect 88048 647593 88090 647829
rect 87770 647509 88090 647593
rect 87770 647273 87812 647509
rect 88048 647273 88090 647509
rect 87770 647241 88090 647273
rect 103909 647829 104229 647861
rect 103909 647593 103951 647829
rect 104187 647593 104229 647829
rect 103909 647509 104229 647593
rect 103909 647273 103951 647509
rect 104187 647273 104229 647509
rect 103909 647241 104229 647273
rect 109840 647829 110160 647861
rect 109840 647593 109882 647829
rect 110118 647593 110160 647829
rect 109840 647509 110160 647593
rect 109840 647273 109882 647509
rect 110118 647273 110160 647509
rect 109840 647241 110160 647273
rect 115770 647829 116090 647861
rect 115770 647593 115812 647829
rect 116048 647593 116090 647829
rect 115770 647509 116090 647593
rect 115770 647273 115812 647509
rect 116048 647273 116090 647509
rect 115770 647241 116090 647273
rect 131909 647829 132229 647861
rect 131909 647593 131951 647829
rect 132187 647593 132229 647829
rect 131909 647509 132229 647593
rect 131909 647273 131951 647509
rect 132187 647273 132229 647509
rect 131909 647241 132229 647273
rect 137840 647829 138160 647861
rect 137840 647593 137882 647829
rect 138118 647593 138160 647829
rect 137840 647509 138160 647593
rect 137840 647273 137882 647509
rect 138118 647273 138160 647509
rect 137840 647241 138160 647273
rect 143770 647829 144090 647861
rect 143770 647593 143812 647829
rect 144048 647593 144090 647829
rect 143770 647509 144090 647593
rect 143770 647273 143812 647509
rect 144048 647273 144090 647509
rect 143770 647241 144090 647273
rect 159909 647829 160229 647861
rect 159909 647593 159951 647829
rect 160187 647593 160229 647829
rect 159909 647509 160229 647593
rect 159909 647273 159951 647509
rect 160187 647273 160229 647509
rect 159909 647241 160229 647273
rect 165840 647829 166160 647861
rect 165840 647593 165882 647829
rect 166118 647593 166160 647829
rect 165840 647509 166160 647593
rect 165840 647273 165882 647509
rect 166118 647273 166160 647509
rect 165840 647241 166160 647273
rect 171770 647829 172090 647861
rect 171770 647593 171812 647829
rect 172048 647593 172090 647829
rect 171770 647509 172090 647593
rect 171770 647273 171812 647509
rect 172048 647273 172090 647509
rect 171770 647241 172090 647273
rect 187909 647829 188229 647861
rect 187909 647593 187951 647829
rect 188187 647593 188229 647829
rect 187909 647509 188229 647593
rect 187909 647273 187951 647509
rect 188187 647273 188229 647509
rect 187909 647241 188229 647273
rect 193840 647829 194160 647861
rect 193840 647593 193882 647829
rect 194118 647593 194160 647829
rect 193840 647509 194160 647593
rect 193840 647273 193882 647509
rect 194118 647273 194160 647509
rect 193840 647241 194160 647273
rect 199770 647829 200090 647861
rect 199770 647593 199812 647829
rect 200048 647593 200090 647829
rect 199770 647509 200090 647593
rect 199770 647273 199812 647509
rect 200048 647273 200090 647509
rect 199770 647241 200090 647273
rect 215909 647829 216229 647861
rect 215909 647593 215951 647829
rect 216187 647593 216229 647829
rect 215909 647509 216229 647593
rect 215909 647273 215951 647509
rect 216187 647273 216229 647509
rect 215909 647241 216229 647273
rect 221840 647829 222160 647861
rect 221840 647593 221882 647829
rect 222118 647593 222160 647829
rect 221840 647509 222160 647593
rect 221840 647273 221882 647509
rect 222118 647273 222160 647509
rect 221840 647241 222160 647273
rect 227770 647829 228090 647861
rect 227770 647593 227812 647829
rect 228048 647593 228090 647829
rect 227770 647509 228090 647593
rect 227770 647273 227812 647509
rect 228048 647273 228090 647509
rect 227770 647241 228090 647273
rect 243909 647829 244229 647861
rect 243909 647593 243951 647829
rect 244187 647593 244229 647829
rect 243909 647509 244229 647593
rect 243909 647273 243951 647509
rect 244187 647273 244229 647509
rect 243909 647241 244229 647273
rect 249840 647829 250160 647861
rect 249840 647593 249882 647829
rect 250118 647593 250160 647829
rect 249840 647509 250160 647593
rect 249840 647273 249882 647509
rect 250118 647273 250160 647509
rect 249840 647241 250160 647273
rect 255770 647829 256090 647861
rect 255770 647593 255812 647829
rect 256048 647593 256090 647829
rect 255770 647509 256090 647593
rect 255770 647273 255812 647509
rect 256048 647273 256090 647509
rect 255770 647241 256090 647273
rect 271909 647829 272229 647861
rect 271909 647593 271951 647829
rect 272187 647593 272229 647829
rect 271909 647509 272229 647593
rect 271909 647273 271951 647509
rect 272187 647273 272229 647509
rect 271909 647241 272229 647273
rect 277840 647829 278160 647861
rect 277840 647593 277882 647829
rect 278118 647593 278160 647829
rect 277840 647509 278160 647593
rect 277840 647273 277882 647509
rect 278118 647273 278160 647509
rect 277840 647241 278160 647273
rect 283770 647829 284090 647861
rect 283770 647593 283812 647829
rect 284048 647593 284090 647829
rect 283770 647509 284090 647593
rect 283770 647273 283812 647509
rect 284048 647273 284090 647509
rect 283770 647241 284090 647273
rect 299909 647829 300229 647861
rect 299909 647593 299951 647829
rect 300187 647593 300229 647829
rect 299909 647509 300229 647593
rect 299909 647273 299951 647509
rect 300187 647273 300229 647509
rect 299909 647241 300229 647273
rect 305840 647829 306160 647861
rect 305840 647593 305882 647829
rect 306118 647593 306160 647829
rect 305840 647509 306160 647593
rect 305840 647273 305882 647509
rect 306118 647273 306160 647509
rect 305840 647241 306160 647273
rect 311770 647829 312090 647861
rect 311770 647593 311812 647829
rect 312048 647593 312090 647829
rect 311770 647509 312090 647593
rect 311770 647273 311812 647509
rect 312048 647273 312090 647509
rect 311770 647241 312090 647273
rect 327909 647829 328229 647861
rect 327909 647593 327951 647829
rect 328187 647593 328229 647829
rect 327909 647509 328229 647593
rect 327909 647273 327951 647509
rect 328187 647273 328229 647509
rect 327909 647241 328229 647273
rect 333840 647829 334160 647861
rect 333840 647593 333882 647829
rect 334118 647593 334160 647829
rect 333840 647509 334160 647593
rect 333840 647273 333882 647509
rect 334118 647273 334160 647509
rect 333840 647241 334160 647273
rect 339770 647829 340090 647861
rect 339770 647593 339812 647829
rect 340048 647593 340090 647829
rect 339770 647509 340090 647593
rect 339770 647273 339812 647509
rect 340048 647273 340090 647509
rect 339770 647241 340090 647273
rect 355909 647829 356229 647861
rect 355909 647593 355951 647829
rect 356187 647593 356229 647829
rect 355909 647509 356229 647593
rect 355909 647273 355951 647509
rect 356187 647273 356229 647509
rect 355909 647241 356229 647273
rect 361840 647829 362160 647861
rect 361840 647593 361882 647829
rect 362118 647593 362160 647829
rect 361840 647509 362160 647593
rect 361840 647273 361882 647509
rect 362118 647273 362160 647509
rect 361840 647241 362160 647273
rect 367770 647829 368090 647861
rect 367770 647593 367812 647829
rect 368048 647593 368090 647829
rect 367770 647509 368090 647593
rect 367770 647273 367812 647509
rect 368048 647273 368090 647509
rect 367770 647241 368090 647273
rect 383909 647829 384229 647861
rect 383909 647593 383951 647829
rect 384187 647593 384229 647829
rect 383909 647509 384229 647593
rect 383909 647273 383951 647509
rect 384187 647273 384229 647509
rect 383909 647241 384229 647273
rect 389840 647829 390160 647861
rect 389840 647593 389882 647829
rect 390118 647593 390160 647829
rect 389840 647509 390160 647593
rect 389840 647273 389882 647509
rect 390118 647273 390160 647509
rect 389840 647241 390160 647273
rect 395770 647829 396090 647861
rect 395770 647593 395812 647829
rect 396048 647593 396090 647829
rect 395770 647509 396090 647593
rect 395770 647273 395812 647509
rect 396048 647273 396090 647509
rect 395770 647241 396090 647273
rect 411909 647829 412229 647861
rect 411909 647593 411951 647829
rect 412187 647593 412229 647829
rect 411909 647509 412229 647593
rect 411909 647273 411951 647509
rect 412187 647273 412229 647509
rect 411909 647241 412229 647273
rect 417840 647829 418160 647861
rect 417840 647593 417882 647829
rect 418118 647593 418160 647829
rect 417840 647509 418160 647593
rect 417840 647273 417882 647509
rect 418118 647273 418160 647509
rect 417840 647241 418160 647273
rect 423770 647829 424090 647861
rect 423770 647593 423812 647829
rect 424048 647593 424090 647829
rect 423770 647509 424090 647593
rect 423770 647273 423812 647509
rect 424048 647273 424090 647509
rect 423770 647241 424090 647273
rect 439909 647829 440229 647861
rect 439909 647593 439951 647829
rect 440187 647593 440229 647829
rect 439909 647509 440229 647593
rect 439909 647273 439951 647509
rect 440187 647273 440229 647509
rect 439909 647241 440229 647273
rect 445840 647829 446160 647861
rect 445840 647593 445882 647829
rect 446118 647593 446160 647829
rect 445840 647509 446160 647593
rect 445840 647273 445882 647509
rect 446118 647273 446160 647509
rect 445840 647241 446160 647273
rect 451770 647829 452090 647861
rect 451770 647593 451812 647829
rect 452048 647593 452090 647829
rect 451770 647509 452090 647593
rect 451770 647273 451812 647509
rect 452048 647273 452090 647509
rect 451770 647241 452090 647273
rect 467909 647829 468229 647861
rect 467909 647593 467951 647829
rect 468187 647593 468229 647829
rect 467909 647509 468229 647593
rect 467909 647273 467951 647509
rect 468187 647273 468229 647509
rect 467909 647241 468229 647273
rect 473840 647829 474160 647861
rect 473840 647593 473882 647829
rect 474118 647593 474160 647829
rect 473840 647509 474160 647593
rect 473840 647273 473882 647509
rect 474118 647273 474160 647509
rect 473840 647241 474160 647273
rect 479770 647829 480090 647861
rect 479770 647593 479812 647829
rect 480048 647593 480090 647829
rect 479770 647509 480090 647593
rect 479770 647273 479812 647509
rect 480048 647273 480090 647509
rect 479770 647241 480090 647273
rect 495909 647829 496229 647861
rect 495909 647593 495951 647829
rect 496187 647593 496229 647829
rect 495909 647509 496229 647593
rect 495909 647273 495951 647509
rect 496187 647273 496229 647509
rect 495909 647241 496229 647273
rect 501840 647829 502160 647861
rect 501840 647593 501882 647829
rect 502118 647593 502160 647829
rect 501840 647509 502160 647593
rect 501840 647273 501882 647509
rect 502118 647273 502160 647509
rect 501840 647241 502160 647273
rect 507770 647829 508090 647861
rect 507770 647593 507812 647829
rect 508048 647593 508090 647829
rect 507770 647509 508090 647593
rect 507770 647273 507812 647509
rect 508048 647273 508090 647509
rect 507770 647241 508090 647273
rect 523909 647829 524229 647861
rect 523909 647593 523951 647829
rect 524187 647593 524229 647829
rect 523909 647509 524229 647593
rect 523909 647273 523951 647509
rect 524187 647273 524229 647509
rect 523909 647241 524229 647273
rect 529840 647829 530160 647861
rect 529840 647593 529882 647829
rect 530118 647593 530160 647829
rect 529840 647509 530160 647593
rect 529840 647273 529882 647509
rect 530118 647273 530160 647509
rect 529840 647241 530160 647273
rect 535770 647829 536090 647861
rect 535770 647593 535812 647829
rect 536048 647593 536090 647829
rect 535770 647509 536090 647593
rect 535770 647273 535812 647509
rect 536048 647273 536090 647509
rect 535770 647241 536090 647273
rect 551909 647829 552229 647861
rect 551909 647593 551951 647829
rect 552187 647593 552229 647829
rect 551909 647509 552229 647593
rect 551909 647273 551951 647509
rect 552187 647273 552229 647509
rect 551909 647241 552229 647273
rect 557840 647829 558160 647861
rect 557840 647593 557882 647829
rect 558118 647593 558160 647829
rect 557840 647509 558160 647593
rect 557840 647273 557882 647509
rect 558118 647273 558160 647509
rect 557840 647241 558160 647273
rect 563770 647829 564090 647861
rect 563770 647593 563812 647829
rect 564048 647593 564090 647829
rect 563770 647509 564090 647593
rect 563770 647273 563812 647509
rect 564048 647273 564090 647509
rect 563770 647241 564090 647273
rect 573494 647829 574114 674273
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 701829 585930 704282
rect 585310 701593 585342 701829
rect 585578 701593 585662 701829
rect 585898 701593 585930 701829
rect 585310 701509 585930 701593
rect 585310 701273 585342 701509
rect 585578 701273 585662 701509
rect 585898 701273 585930 701509
rect 585310 674829 585930 701273
rect 585310 674593 585342 674829
rect 585578 674593 585662 674829
rect 585898 674593 585930 674829
rect 585310 674509 585930 674593
rect 585310 674273 585342 674509
rect 585578 674273 585662 674509
rect 585898 674273 585930 674509
rect 580211 670716 580277 670717
rect 580211 670652 580212 670716
rect 580276 670652 580277 670716
rect 580211 670651 580277 670652
rect 573494 647593 573526 647829
rect 573762 647593 573846 647829
rect 574082 647593 574114 647829
rect 573494 647509 574114 647593
rect 573494 647273 573526 647509
rect 573762 647273 573846 647509
rect 574082 647273 574114 647509
rect 22875 644454 23195 644486
rect 22875 644218 22917 644454
rect 23153 644218 23195 644454
rect 22875 644134 23195 644218
rect 22875 643898 22917 644134
rect 23153 643898 23195 644134
rect 22875 643866 23195 643898
rect 28806 644454 29126 644486
rect 28806 644218 28848 644454
rect 29084 644218 29126 644454
rect 28806 644134 29126 644218
rect 28806 643898 28848 644134
rect 29084 643898 29126 644134
rect 28806 643866 29126 643898
rect 50875 644454 51195 644486
rect 50875 644218 50917 644454
rect 51153 644218 51195 644454
rect 50875 644134 51195 644218
rect 50875 643898 50917 644134
rect 51153 643898 51195 644134
rect 50875 643866 51195 643898
rect 56806 644454 57126 644486
rect 56806 644218 56848 644454
rect 57084 644218 57126 644454
rect 56806 644134 57126 644218
rect 56806 643898 56848 644134
rect 57084 643898 57126 644134
rect 56806 643866 57126 643898
rect 78875 644454 79195 644486
rect 78875 644218 78917 644454
rect 79153 644218 79195 644454
rect 78875 644134 79195 644218
rect 78875 643898 78917 644134
rect 79153 643898 79195 644134
rect 78875 643866 79195 643898
rect 84806 644454 85126 644486
rect 84806 644218 84848 644454
rect 85084 644218 85126 644454
rect 84806 644134 85126 644218
rect 84806 643898 84848 644134
rect 85084 643898 85126 644134
rect 84806 643866 85126 643898
rect 106875 644454 107195 644486
rect 106875 644218 106917 644454
rect 107153 644218 107195 644454
rect 106875 644134 107195 644218
rect 106875 643898 106917 644134
rect 107153 643898 107195 644134
rect 106875 643866 107195 643898
rect 112806 644454 113126 644486
rect 112806 644218 112848 644454
rect 113084 644218 113126 644454
rect 112806 644134 113126 644218
rect 112806 643898 112848 644134
rect 113084 643898 113126 644134
rect 112806 643866 113126 643898
rect 134875 644454 135195 644486
rect 134875 644218 134917 644454
rect 135153 644218 135195 644454
rect 134875 644134 135195 644218
rect 134875 643898 134917 644134
rect 135153 643898 135195 644134
rect 134875 643866 135195 643898
rect 140806 644454 141126 644486
rect 140806 644218 140848 644454
rect 141084 644218 141126 644454
rect 140806 644134 141126 644218
rect 140806 643898 140848 644134
rect 141084 643898 141126 644134
rect 140806 643866 141126 643898
rect 162875 644454 163195 644486
rect 162875 644218 162917 644454
rect 163153 644218 163195 644454
rect 162875 644134 163195 644218
rect 162875 643898 162917 644134
rect 163153 643898 163195 644134
rect 162875 643866 163195 643898
rect 168806 644454 169126 644486
rect 168806 644218 168848 644454
rect 169084 644218 169126 644454
rect 168806 644134 169126 644218
rect 168806 643898 168848 644134
rect 169084 643898 169126 644134
rect 168806 643866 169126 643898
rect 190875 644454 191195 644486
rect 190875 644218 190917 644454
rect 191153 644218 191195 644454
rect 190875 644134 191195 644218
rect 190875 643898 190917 644134
rect 191153 643898 191195 644134
rect 190875 643866 191195 643898
rect 196806 644454 197126 644486
rect 196806 644218 196848 644454
rect 197084 644218 197126 644454
rect 196806 644134 197126 644218
rect 196806 643898 196848 644134
rect 197084 643898 197126 644134
rect 196806 643866 197126 643898
rect 218875 644454 219195 644486
rect 218875 644218 218917 644454
rect 219153 644218 219195 644454
rect 218875 644134 219195 644218
rect 218875 643898 218917 644134
rect 219153 643898 219195 644134
rect 218875 643866 219195 643898
rect 224806 644454 225126 644486
rect 224806 644218 224848 644454
rect 225084 644218 225126 644454
rect 224806 644134 225126 644218
rect 224806 643898 224848 644134
rect 225084 643898 225126 644134
rect 224806 643866 225126 643898
rect 246875 644454 247195 644486
rect 246875 644218 246917 644454
rect 247153 644218 247195 644454
rect 246875 644134 247195 644218
rect 246875 643898 246917 644134
rect 247153 643898 247195 644134
rect 246875 643866 247195 643898
rect 252806 644454 253126 644486
rect 252806 644218 252848 644454
rect 253084 644218 253126 644454
rect 252806 644134 253126 644218
rect 252806 643898 252848 644134
rect 253084 643898 253126 644134
rect 252806 643866 253126 643898
rect 274875 644454 275195 644486
rect 274875 644218 274917 644454
rect 275153 644218 275195 644454
rect 274875 644134 275195 644218
rect 274875 643898 274917 644134
rect 275153 643898 275195 644134
rect 274875 643866 275195 643898
rect 280806 644454 281126 644486
rect 280806 644218 280848 644454
rect 281084 644218 281126 644454
rect 280806 644134 281126 644218
rect 280806 643898 280848 644134
rect 281084 643898 281126 644134
rect 280806 643866 281126 643898
rect 302875 644454 303195 644486
rect 302875 644218 302917 644454
rect 303153 644218 303195 644454
rect 302875 644134 303195 644218
rect 302875 643898 302917 644134
rect 303153 643898 303195 644134
rect 302875 643866 303195 643898
rect 308806 644454 309126 644486
rect 308806 644218 308848 644454
rect 309084 644218 309126 644454
rect 308806 644134 309126 644218
rect 308806 643898 308848 644134
rect 309084 643898 309126 644134
rect 308806 643866 309126 643898
rect 330875 644454 331195 644486
rect 330875 644218 330917 644454
rect 331153 644218 331195 644454
rect 330875 644134 331195 644218
rect 330875 643898 330917 644134
rect 331153 643898 331195 644134
rect 330875 643866 331195 643898
rect 336806 644454 337126 644486
rect 336806 644218 336848 644454
rect 337084 644218 337126 644454
rect 336806 644134 337126 644218
rect 336806 643898 336848 644134
rect 337084 643898 337126 644134
rect 336806 643866 337126 643898
rect 358875 644454 359195 644486
rect 358875 644218 358917 644454
rect 359153 644218 359195 644454
rect 358875 644134 359195 644218
rect 358875 643898 358917 644134
rect 359153 643898 359195 644134
rect 358875 643866 359195 643898
rect 364806 644454 365126 644486
rect 364806 644218 364848 644454
rect 365084 644218 365126 644454
rect 364806 644134 365126 644218
rect 364806 643898 364848 644134
rect 365084 643898 365126 644134
rect 364806 643866 365126 643898
rect 386875 644454 387195 644486
rect 386875 644218 386917 644454
rect 387153 644218 387195 644454
rect 386875 644134 387195 644218
rect 386875 643898 386917 644134
rect 387153 643898 387195 644134
rect 386875 643866 387195 643898
rect 392806 644454 393126 644486
rect 392806 644218 392848 644454
rect 393084 644218 393126 644454
rect 392806 644134 393126 644218
rect 392806 643898 392848 644134
rect 393084 643898 393126 644134
rect 392806 643866 393126 643898
rect 414875 644454 415195 644486
rect 414875 644218 414917 644454
rect 415153 644218 415195 644454
rect 414875 644134 415195 644218
rect 414875 643898 414917 644134
rect 415153 643898 415195 644134
rect 414875 643866 415195 643898
rect 420806 644454 421126 644486
rect 420806 644218 420848 644454
rect 421084 644218 421126 644454
rect 420806 644134 421126 644218
rect 420806 643898 420848 644134
rect 421084 643898 421126 644134
rect 420806 643866 421126 643898
rect 442875 644454 443195 644486
rect 442875 644218 442917 644454
rect 443153 644218 443195 644454
rect 442875 644134 443195 644218
rect 442875 643898 442917 644134
rect 443153 643898 443195 644134
rect 442875 643866 443195 643898
rect 448806 644454 449126 644486
rect 448806 644218 448848 644454
rect 449084 644218 449126 644454
rect 448806 644134 449126 644218
rect 448806 643898 448848 644134
rect 449084 643898 449126 644134
rect 448806 643866 449126 643898
rect 470875 644454 471195 644486
rect 470875 644218 470917 644454
rect 471153 644218 471195 644454
rect 470875 644134 471195 644218
rect 470875 643898 470917 644134
rect 471153 643898 471195 644134
rect 470875 643866 471195 643898
rect 476806 644454 477126 644486
rect 476806 644218 476848 644454
rect 477084 644218 477126 644454
rect 476806 644134 477126 644218
rect 476806 643898 476848 644134
rect 477084 643898 477126 644134
rect 476806 643866 477126 643898
rect 498875 644454 499195 644486
rect 498875 644218 498917 644454
rect 499153 644218 499195 644454
rect 498875 644134 499195 644218
rect 498875 643898 498917 644134
rect 499153 643898 499195 644134
rect 498875 643866 499195 643898
rect 504806 644454 505126 644486
rect 504806 644218 504848 644454
rect 505084 644218 505126 644454
rect 504806 644134 505126 644218
rect 504806 643898 504848 644134
rect 505084 643898 505126 644134
rect 504806 643866 505126 643898
rect 526875 644454 527195 644486
rect 526875 644218 526917 644454
rect 527153 644218 527195 644454
rect 526875 644134 527195 644218
rect 526875 643898 526917 644134
rect 527153 643898 527195 644134
rect 526875 643866 527195 643898
rect 532806 644454 533126 644486
rect 532806 644218 532848 644454
rect 533084 644218 533126 644454
rect 532806 644134 533126 644218
rect 532806 643898 532848 644134
rect 533084 643898 533126 644134
rect 532806 643866 533126 643898
rect 554875 644454 555195 644486
rect 554875 644218 554917 644454
rect 555153 644218 555195 644454
rect 554875 644134 555195 644218
rect 554875 643898 554917 644134
rect 555153 643898 555195 644134
rect 554875 643866 555195 643898
rect 560806 644454 561126 644486
rect 560806 644218 560848 644454
rect 561084 644218 561126 644454
rect 560806 644134 561126 644218
rect 560806 643898 560848 644134
rect 561084 643898 561126 644134
rect 560806 643866 561126 643898
rect -2006 620593 -1974 620829
rect -1738 620593 -1654 620829
rect -1418 620593 -1386 620829
rect -2006 620509 -1386 620593
rect -2006 620273 -1974 620509
rect -1738 620273 -1654 620509
rect -1418 620273 -1386 620509
rect -2006 593829 -1386 620273
rect 19910 620829 20230 620861
rect 19910 620593 19952 620829
rect 20188 620593 20230 620829
rect 19910 620509 20230 620593
rect 19910 620273 19952 620509
rect 20188 620273 20230 620509
rect 19910 620241 20230 620273
rect 25840 620829 26160 620861
rect 25840 620593 25882 620829
rect 26118 620593 26160 620829
rect 25840 620509 26160 620593
rect 25840 620273 25882 620509
rect 26118 620273 26160 620509
rect 25840 620241 26160 620273
rect 31771 620829 32091 620861
rect 31771 620593 31813 620829
rect 32049 620593 32091 620829
rect 31771 620509 32091 620593
rect 31771 620273 31813 620509
rect 32049 620273 32091 620509
rect 31771 620241 32091 620273
rect 47910 620829 48230 620861
rect 47910 620593 47952 620829
rect 48188 620593 48230 620829
rect 47910 620509 48230 620593
rect 47910 620273 47952 620509
rect 48188 620273 48230 620509
rect 47910 620241 48230 620273
rect 53840 620829 54160 620861
rect 53840 620593 53882 620829
rect 54118 620593 54160 620829
rect 53840 620509 54160 620593
rect 53840 620273 53882 620509
rect 54118 620273 54160 620509
rect 53840 620241 54160 620273
rect 59771 620829 60091 620861
rect 59771 620593 59813 620829
rect 60049 620593 60091 620829
rect 59771 620509 60091 620593
rect 59771 620273 59813 620509
rect 60049 620273 60091 620509
rect 59771 620241 60091 620273
rect 75910 620829 76230 620861
rect 75910 620593 75952 620829
rect 76188 620593 76230 620829
rect 75910 620509 76230 620593
rect 75910 620273 75952 620509
rect 76188 620273 76230 620509
rect 75910 620241 76230 620273
rect 81840 620829 82160 620861
rect 81840 620593 81882 620829
rect 82118 620593 82160 620829
rect 81840 620509 82160 620593
rect 81840 620273 81882 620509
rect 82118 620273 82160 620509
rect 81840 620241 82160 620273
rect 87771 620829 88091 620861
rect 87771 620593 87813 620829
rect 88049 620593 88091 620829
rect 87771 620509 88091 620593
rect 87771 620273 87813 620509
rect 88049 620273 88091 620509
rect 87771 620241 88091 620273
rect 103910 620829 104230 620861
rect 103910 620593 103952 620829
rect 104188 620593 104230 620829
rect 103910 620509 104230 620593
rect 103910 620273 103952 620509
rect 104188 620273 104230 620509
rect 103910 620241 104230 620273
rect 109840 620829 110160 620861
rect 109840 620593 109882 620829
rect 110118 620593 110160 620829
rect 109840 620509 110160 620593
rect 109840 620273 109882 620509
rect 110118 620273 110160 620509
rect 109840 620241 110160 620273
rect 115771 620829 116091 620861
rect 115771 620593 115813 620829
rect 116049 620593 116091 620829
rect 115771 620509 116091 620593
rect 115771 620273 115813 620509
rect 116049 620273 116091 620509
rect 115771 620241 116091 620273
rect 131910 620829 132230 620861
rect 131910 620593 131952 620829
rect 132188 620593 132230 620829
rect 131910 620509 132230 620593
rect 131910 620273 131952 620509
rect 132188 620273 132230 620509
rect 131910 620241 132230 620273
rect 137840 620829 138160 620861
rect 137840 620593 137882 620829
rect 138118 620593 138160 620829
rect 137840 620509 138160 620593
rect 137840 620273 137882 620509
rect 138118 620273 138160 620509
rect 137840 620241 138160 620273
rect 143771 620829 144091 620861
rect 143771 620593 143813 620829
rect 144049 620593 144091 620829
rect 143771 620509 144091 620593
rect 143771 620273 143813 620509
rect 144049 620273 144091 620509
rect 143771 620241 144091 620273
rect 159910 620829 160230 620861
rect 159910 620593 159952 620829
rect 160188 620593 160230 620829
rect 159910 620509 160230 620593
rect 159910 620273 159952 620509
rect 160188 620273 160230 620509
rect 159910 620241 160230 620273
rect 165840 620829 166160 620861
rect 165840 620593 165882 620829
rect 166118 620593 166160 620829
rect 165840 620509 166160 620593
rect 165840 620273 165882 620509
rect 166118 620273 166160 620509
rect 165840 620241 166160 620273
rect 171771 620829 172091 620861
rect 171771 620593 171813 620829
rect 172049 620593 172091 620829
rect 171771 620509 172091 620593
rect 171771 620273 171813 620509
rect 172049 620273 172091 620509
rect 171771 620241 172091 620273
rect 187910 620829 188230 620861
rect 187910 620593 187952 620829
rect 188188 620593 188230 620829
rect 187910 620509 188230 620593
rect 187910 620273 187952 620509
rect 188188 620273 188230 620509
rect 187910 620241 188230 620273
rect 193840 620829 194160 620861
rect 193840 620593 193882 620829
rect 194118 620593 194160 620829
rect 193840 620509 194160 620593
rect 193840 620273 193882 620509
rect 194118 620273 194160 620509
rect 193840 620241 194160 620273
rect 199771 620829 200091 620861
rect 199771 620593 199813 620829
rect 200049 620593 200091 620829
rect 199771 620509 200091 620593
rect 199771 620273 199813 620509
rect 200049 620273 200091 620509
rect 199771 620241 200091 620273
rect 215910 620829 216230 620861
rect 215910 620593 215952 620829
rect 216188 620593 216230 620829
rect 215910 620509 216230 620593
rect 215910 620273 215952 620509
rect 216188 620273 216230 620509
rect 215910 620241 216230 620273
rect 221840 620829 222160 620861
rect 221840 620593 221882 620829
rect 222118 620593 222160 620829
rect 221840 620509 222160 620593
rect 221840 620273 221882 620509
rect 222118 620273 222160 620509
rect 221840 620241 222160 620273
rect 227771 620829 228091 620861
rect 227771 620593 227813 620829
rect 228049 620593 228091 620829
rect 227771 620509 228091 620593
rect 227771 620273 227813 620509
rect 228049 620273 228091 620509
rect 227771 620241 228091 620273
rect 243910 620829 244230 620861
rect 243910 620593 243952 620829
rect 244188 620593 244230 620829
rect 243910 620509 244230 620593
rect 243910 620273 243952 620509
rect 244188 620273 244230 620509
rect 243910 620241 244230 620273
rect 249840 620829 250160 620861
rect 249840 620593 249882 620829
rect 250118 620593 250160 620829
rect 249840 620509 250160 620593
rect 249840 620273 249882 620509
rect 250118 620273 250160 620509
rect 249840 620241 250160 620273
rect 255771 620829 256091 620861
rect 255771 620593 255813 620829
rect 256049 620593 256091 620829
rect 255771 620509 256091 620593
rect 255771 620273 255813 620509
rect 256049 620273 256091 620509
rect 255771 620241 256091 620273
rect 271910 620829 272230 620861
rect 271910 620593 271952 620829
rect 272188 620593 272230 620829
rect 271910 620509 272230 620593
rect 271910 620273 271952 620509
rect 272188 620273 272230 620509
rect 271910 620241 272230 620273
rect 277840 620829 278160 620861
rect 277840 620593 277882 620829
rect 278118 620593 278160 620829
rect 277840 620509 278160 620593
rect 277840 620273 277882 620509
rect 278118 620273 278160 620509
rect 277840 620241 278160 620273
rect 283771 620829 284091 620861
rect 283771 620593 283813 620829
rect 284049 620593 284091 620829
rect 283771 620509 284091 620593
rect 283771 620273 283813 620509
rect 284049 620273 284091 620509
rect 283771 620241 284091 620273
rect 299910 620829 300230 620861
rect 299910 620593 299952 620829
rect 300188 620593 300230 620829
rect 299910 620509 300230 620593
rect 299910 620273 299952 620509
rect 300188 620273 300230 620509
rect 299910 620241 300230 620273
rect 305840 620829 306160 620861
rect 305840 620593 305882 620829
rect 306118 620593 306160 620829
rect 305840 620509 306160 620593
rect 305840 620273 305882 620509
rect 306118 620273 306160 620509
rect 305840 620241 306160 620273
rect 311771 620829 312091 620861
rect 311771 620593 311813 620829
rect 312049 620593 312091 620829
rect 311771 620509 312091 620593
rect 311771 620273 311813 620509
rect 312049 620273 312091 620509
rect 311771 620241 312091 620273
rect 327910 620829 328230 620861
rect 327910 620593 327952 620829
rect 328188 620593 328230 620829
rect 327910 620509 328230 620593
rect 327910 620273 327952 620509
rect 328188 620273 328230 620509
rect 327910 620241 328230 620273
rect 333840 620829 334160 620861
rect 333840 620593 333882 620829
rect 334118 620593 334160 620829
rect 333840 620509 334160 620593
rect 333840 620273 333882 620509
rect 334118 620273 334160 620509
rect 333840 620241 334160 620273
rect 339771 620829 340091 620861
rect 339771 620593 339813 620829
rect 340049 620593 340091 620829
rect 339771 620509 340091 620593
rect 339771 620273 339813 620509
rect 340049 620273 340091 620509
rect 339771 620241 340091 620273
rect 355910 620829 356230 620861
rect 355910 620593 355952 620829
rect 356188 620593 356230 620829
rect 355910 620509 356230 620593
rect 355910 620273 355952 620509
rect 356188 620273 356230 620509
rect 355910 620241 356230 620273
rect 361840 620829 362160 620861
rect 361840 620593 361882 620829
rect 362118 620593 362160 620829
rect 361840 620509 362160 620593
rect 361840 620273 361882 620509
rect 362118 620273 362160 620509
rect 361840 620241 362160 620273
rect 367771 620829 368091 620861
rect 367771 620593 367813 620829
rect 368049 620593 368091 620829
rect 367771 620509 368091 620593
rect 367771 620273 367813 620509
rect 368049 620273 368091 620509
rect 367771 620241 368091 620273
rect 383910 620829 384230 620861
rect 383910 620593 383952 620829
rect 384188 620593 384230 620829
rect 383910 620509 384230 620593
rect 383910 620273 383952 620509
rect 384188 620273 384230 620509
rect 383910 620241 384230 620273
rect 389840 620829 390160 620861
rect 389840 620593 389882 620829
rect 390118 620593 390160 620829
rect 389840 620509 390160 620593
rect 389840 620273 389882 620509
rect 390118 620273 390160 620509
rect 389840 620241 390160 620273
rect 395771 620829 396091 620861
rect 395771 620593 395813 620829
rect 396049 620593 396091 620829
rect 395771 620509 396091 620593
rect 395771 620273 395813 620509
rect 396049 620273 396091 620509
rect 395771 620241 396091 620273
rect 411910 620829 412230 620861
rect 411910 620593 411952 620829
rect 412188 620593 412230 620829
rect 411910 620509 412230 620593
rect 411910 620273 411952 620509
rect 412188 620273 412230 620509
rect 411910 620241 412230 620273
rect 417840 620829 418160 620861
rect 417840 620593 417882 620829
rect 418118 620593 418160 620829
rect 417840 620509 418160 620593
rect 417840 620273 417882 620509
rect 418118 620273 418160 620509
rect 417840 620241 418160 620273
rect 423771 620829 424091 620861
rect 423771 620593 423813 620829
rect 424049 620593 424091 620829
rect 423771 620509 424091 620593
rect 423771 620273 423813 620509
rect 424049 620273 424091 620509
rect 423771 620241 424091 620273
rect 439910 620829 440230 620861
rect 439910 620593 439952 620829
rect 440188 620593 440230 620829
rect 439910 620509 440230 620593
rect 439910 620273 439952 620509
rect 440188 620273 440230 620509
rect 439910 620241 440230 620273
rect 445840 620829 446160 620861
rect 445840 620593 445882 620829
rect 446118 620593 446160 620829
rect 445840 620509 446160 620593
rect 445840 620273 445882 620509
rect 446118 620273 446160 620509
rect 445840 620241 446160 620273
rect 451771 620829 452091 620861
rect 451771 620593 451813 620829
rect 452049 620593 452091 620829
rect 451771 620509 452091 620593
rect 451771 620273 451813 620509
rect 452049 620273 452091 620509
rect 451771 620241 452091 620273
rect 467910 620829 468230 620861
rect 467910 620593 467952 620829
rect 468188 620593 468230 620829
rect 467910 620509 468230 620593
rect 467910 620273 467952 620509
rect 468188 620273 468230 620509
rect 467910 620241 468230 620273
rect 473840 620829 474160 620861
rect 473840 620593 473882 620829
rect 474118 620593 474160 620829
rect 473840 620509 474160 620593
rect 473840 620273 473882 620509
rect 474118 620273 474160 620509
rect 473840 620241 474160 620273
rect 479771 620829 480091 620861
rect 479771 620593 479813 620829
rect 480049 620593 480091 620829
rect 479771 620509 480091 620593
rect 479771 620273 479813 620509
rect 480049 620273 480091 620509
rect 479771 620241 480091 620273
rect 495910 620829 496230 620861
rect 495910 620593 495952 620829
rect 496188 620593 496230 620829
rect 495910 620509 496230 620593
rect 495910 620273 495952 620509
rect 496188 620273 496230 620509
rect 495910 620241 496230 620273
rect 501840 620829 502160 620861
rect 501840 620593 501882 620829
rect 502118 620593 502160 620829
rect 501840 620509 502160 620593
rect 501840 620273 501882 620509
rect 502118 620273 502160 620509
rect 501840 620241 502160 620273
rect 507771 620829 508091 620861
rect 507771 620593 507813 620829
rect 508049 620593 508091 620829
rect 507771 620509 508091 620593
rect 507771 620273 507813 620509
rect 508049 620273 508091 620509
rect 507771 620241 508091 620273
rect 523910 620829 524230 620861
rect 523910 620593 523952 620829
rect 524188 620593 524230 620829
rect 523910 620509 524230 620593
rect 523910 620273 523952 620509
rect 524188 620273 524230 620509
rect 523910 620241 524230 620273
rect 529840 620829 530160 620861
rect 529840 620593 529882 620829
rect 530118 620593 530160 620829
rect 529840 620509 530160 620593
rect 529840 620273 529882 620509
rect 530118 620273 530160 620509
rect 529840 620241 530160 620273
rect 535771 620829 536091 620861
rect 535771 620593 535813 620829
rect 536049 620593 536091 620829
rect 535771 620509 536091 620593
rect 535771 620273 535813 620509
rect 536049 620273 536091 620509
rect 535771 620241 536091 620273
rect 551910 620829 552230 620861
rect 551910 620593 551952 620829
rect 552188 620593 552230 620829
rect 551910 620509 552230 620593
rect 551910 620273 551952 620509
rect 552188 620273 552230 620509
rect 551910 620241 552230 620273
rect 557840 620829 558160 620861
rect 557840 620593 557882 620829
rect 558118 620593 558160 620829
rect 557840 620509 558160 620593
rect 557840 620273 557882 620509
rect 558118 620273 558160 620509
rect 557840 620241 558160 620273
rect 563771 620829 564091 620861
rect 563771 620593 563813 620829
rect 564049 620593 564091 620829
rect 563771 620509 564091 620593
rect 563771 620273 563813 620509
rect 564049 620273 564091 620509
rect 563771 620241 564091 620273
rect 573494 620829 574114 647273
rect 573494 620593 573526 620829
rect 573762 620593 573846 620829
rect 574082 620593 574114 620829
rect 573494 620509 574114 620593
rect 573494 620273 573526 620509
rect 573762 620273 573846 620509
rect 574082 620273 574114 620509
rect 22874 617454 23194 617486
rect 22874 617218 22916 617454
rect 23152 617218 23194 617454
rect 22874 617134 23194 617218
rect 22874 616898 22916 617134
rect 23152 616898 23194 617134
rect 22874 616866 23194 616898
rect 28805 617454 29125 617486
rect 28805 617218 28847 617454
rect 29083 617218 29125 617454
rect 28805 617134 29125 617218
rect 28805 616898 28847 617134
rect 29083 616898 29125 617134
rect 28805 616866 29125 616898
rect 50874 617454 51194 617486
rect 50874 617218 50916 617454
rect 51152 617218 51194 617454
rect 50874 617134 51194 617218
rect 50874 616898 50916 617134
rect 51152 616898 51194 617134
rect 50874 616866 51194 616898
rect 56805 617454 57125 617486
rect 56805 617218 56847 617454
rect 57083 617218 57125 617454
rect 56805 617134 57125 617218
rect 56805 616898 56847 617134
rect 57083 616898 57125 617134
rect 56805 616866 57125 616898
rect 78874 617454 79194 617486
rect 78874 617218 78916 617454
rect 79152 617218 79194 617454
rect 78874 617134 79194 617218
rect 78874 616898 78916 617134
rect 79152 616898 79194 617134
rect 78874 616866 79194 616898
rect 84805 617454 85125 617486
rect 84805 617218 84847 617454
rect 85083 617218 85125 617454
rect 84805 617134 85125 617218
rect 84805 616898 84847 617134
rect 85083 616898 85125 617134
rect 84805 616866 85125 616898
rect 106874 617454 107194 617486
rect 106874 617218 106916 617454
rect 107152 617218 107194 617454
rect 106874 617134 107194 617218
rect 106874 616898 106916 617134
rect 107152 616898 107194 617134
rect 106874 616866 107194 616898
rect 112805 617454 113125 617486
rect 112805 617218 112847 617454
rect 113083 617218 113125 617454
rect 112805 617134 113125 617218
rect 112805 616898 112847 617134
rect 113083 616898 113125 617134
rect 112805 616866 113125 616898
rect 134874 617454 135194 617486
rect 134874 617218 134916 617454
rect 135152 617218 135194 617454
rect 134874 617134 135194 617218
rect 134874 616898 134916 617134
rect 135152 616898 135194 617134
rect 134874 616866 135194 616898
rect 140805 617454 141125 617486
rect 140805 617218 140847 617454
rect 141083 617218 141125 617454
rect 140805 617134 141125 617218
rect 140805 616898 140847 617134
rect 141083 616898 141125 617134
rect 140805 616866 141125 616898
rect 162874 617454 163194 617486
rect 162874 617218 162916 617454
rect 163152 617218 163194 617454
rect 162874 617134 163194 617218
rect 162874 616898 162916 617134
rect 163152 616898 163194 617134
rect 162874 616866 163194 616898
rect 168805 617454 169125 617486
rect 168805 617218 168847 617454
rect 169083 617218 169125 617454
rect 168805 617134 169125 617218
rect 168805 616898 168847 617134
rect 169083 616898 169125 617134
rect 168805 616866 169125 616898
rect 190874 617454 191194 617486
rect 190874 617218 190916 617454
rect 191152 617218 191194 617454
rect 190874 617134 191194 617218
rect 190874 616898 190916 617134
rect 191152 616898 191194 617134
rect 190874 616866 191194 616898
rect 196805 617454 197125 617486
rect 196805 617218 196847 617454
rect 197083 617218 197125 617454
rect 196805 617134 197125 617218
rect 196805 616898 196847 617134
rect 197083 616898 197125 617134
rect 196805 616866 197125 616898
rect 218874 617454 219194 617486
rect 218874 617218 218916 617454
rect 219152 617218 219194 617454
rect 218874 617134 219194 617218
rect 218874 616898 218916 617134
rect 219152 616898 219194 617134
rect 218874 616866 219194 616898
rect 224805 617454 225125 617486
rect 224805 617218 224847 617454
rect 225083 617218 225125 617454
rect 224805 617134 225125 617218
rect 224805 616898 224847 617134
rect 225083 616898 225125 617134
rect 224805 616866 225125 616898
rect 246874 617454 247194 617486
rect 246874 617218 246916 617454
rect 247152 617218 247194 617454
rect 246874 617134 247194 617218
rect 246874 616898 246916 617134
rect 247152 616898 247194 617134
rect 246874 616866 247194 616898
rect 252805 617454 253125 617486
rect 252805 617218 252847 617454
rect 253083 617218 253125 617454
rect 252805 617134 253125 617218
rect 252805 616898 252847 617134
rect 253083 616898 253125 617134
rect 252805 616866 253125 616898
rect 274874 617454 275194 617486
rect 274874 617218 274916 617454
rect 275152 617218 275194 617454
rect 274874 617134 275194 617218
rect 274874 616898 274916 617134
rect 275152 616898 275194 617134
rect 274874 616866 275194 616898
rect 280805 617454 281125 617486
rect 280805 617218 280847 617454
rect 281083 617218 281125 617454
rect 280805 617134 281125 617218
rect 280805 616898 280847 617134
rect 281083 616898 281125 617134
rect 280805 616866 281125 616898
rect 302874 617454 303194 617486
rect 302874 617218 302916 617454
rect 303152 617218 303194 617454
rect 302874 617134 303194 617218
rect 302874 616898 302916 617134
rect 303152 616898 303194 617134
rect 302874 616866 303194 616898
rect 308805 617454 309125 617486
rect 308805 617218 308847 617454
rect 309083 617218 309125 617454
rect 308805 617134 309125 617218
rect 308805 616898 308847 617134
rect 309083 616898 309125 617134
rect 308805 616866 309125 616898
rect 330874 617454 331194 617486
rect 330874 617218 330916 617454
rect 331152 617218 331194 617454
rect 330874 617134 331194 617218
rect 330874 616898 330916 617134
rect 331152 616898 331194 617134
rect 330874 616866 331194 616898
rect 336805 617454 337125 617486
rect 336805 617218 336847 617454
rect 337083 617218 337125 617454
rect 336805 617134 337125 617218
rect 336805 616898 336847 617134
rect 337083 616898 337125 617134
rect 336805 616866 337125 616898
rect 358874 617454 359194 617486
rect 358874 617218 358916 617454
rect 359152 617218 359194 617454
rect 358874 617134 359194 617218
rect 358874 616898 358916 617134
rect 359152 616898 359194 617134
rect 358874 616866 359194 616898
rect 364805 617454 365125 617486
rect 364805 617218 364847 617454
rect 365083 617218 365125 617454
rect 364805 617134 365125 617218
rect 364805 616898 364847 617134
rect 365083 616898 365125 617134
rect 364805 616866 365125 616898
rect 386874 617454 387194 617486
rect 386874 617218 386916 617454
rect 387152 617218 387194 617454
rect 386874 617134 387194 617218
rect 386874 616898 386916 617134
rect 387152 616898 387194 617134
rect 386874 616866 387194 616898
rect 392805 617454 393125 617486
rect 392805 617218 392847 617454
rect 393083 617218 393125 617454
rect 392805 617134 393125 617218
rect 392805 616898 392847 617134
rect 393083 616898 393125 617134
rect 392805 616866 393125 616898
rect 414874 617454 415194 617486
rect 414874 617218 414916 617454
rect 415152 617218 415194 617454
rect 414874 617134 415194 617218
rect 414874 616898 414916 617134
rect 415152 616898 415194 617134
rect 414874 616866 415194 616898
rect 420805 617454 421125 617486
rect 420805 617218 420847 617454
rect 421083 617218 421125 617454
rect 420805 617134 421125 617218
rect 420805 616898 420847 617134
rect 421083 616898 421125 617134
rect 420805 616866 421125 616898
rect 442874 617454 443194 617486
rect 442874 617218 442916 617454
rect 443152 617218 443194 617454
rect 442874 617134 443194 617218
rect 442874 616898 442916 617134
rect 443152 616898 443194 617134
rect 442874 616866 443194 616898
rect 448805 617454 449125 617486
rect 448805 617218 448847 617454
rect 449083 617218 449125 617454
rect 448805 617134 449125 617218
rect 448805 616898 448847 617134
rect 449083 616898 449125 617134
rect 448805 616866 449125 616898
rect 470874 617454 471194 617486
rect 470874 617218 470916 617454
rect 471152 617218 471194 617454
rect 470874 617134 471194 617218
rect 470874 616898 470916 617134
rect 471152 616898 471194 617134
rect 470874 616866 471194 616898
rect 476805 617454 477125 617486
rect 476805 617218 476847 617454
rect 477083 617218 477125 617454
rect 476805 617134 477125 617218
rect 476805 616898 476847 617134
rect 477083 616898 477125 617134
rect 476805 616866 477125 616898
rect 498874 617454 499194 617486
rect 498874 617218 498916 617454
rect 499152 617218 499194 617454
rect 498874 617134 499194 617218
rect 498874 616898 498916 617134
rect 499152 616898 499194 617134
rect 498874 616866 499194 616898
rect 504805 617454 505125 617486
rect 504805 617218 504847 617454
rect 505083 617218 505125 617454
rect 504805 617134 505125 617218
rect 504805 616898 504847 617134
rect 505083 616898 505125 617134
rect 504805 616866 505125 616898
rect 526874 617454 527194 617486
rect 526874 617218 526916 617454
rect 527152 617218 527194 617454
rect 526874 617134 527194 617218
rect 526874 616898 526916 617134
rect 527152 616898 527194 617134
rect 526874 616866 527194 616898
rect 532805 617454 533125 617486
rect 532805 617218 532847 617454
rect 533083 617218 533125 617454
rect 532805 617134 533125 617218
rect 532805 616898 532847 617134
rect 533083 616898 533125 617134
rect 532805 616866 533125 616898
rect 554874 617454 555194 617486
rect 554874 617218 554916 617454
rect 555152 617218 555194 617454
rect 554874 617134 555194 617218
rect 554874 616898 554916 617134
rect 555152 616898 555194 617134
rect 554874 616866 555194 616898
rect 560805 617454 561125 617486
rect 560805 617218 560847 617454
rect 561083 617218 561125 617454
rect 560805 617134 561125 617218
rect 560805 616898 560847 617134
rect 561083 616898 561125 617134
rect 560805 616866 561125 616898
rect -2006 593593 -1974 593829
rect -1738 593593 -1654 593829
rect -1418 593593 -1386 593829
rect -2006 593509 -1386 593593
rect -2006 593273 -1974 593509
rect -1738 593273 -1654 593509
rect -1418 593273 -1386 593509
rect -2006 566829 -1386 593273
rect 19909 593829 20229 593861
rect 19909 593593 19951 593829
rect 20187 593593 20229 593829
rect 19909 593509 20229 593593
rect 19909 593273 19951 593509
rect 20187 593273 20229 593509
rect 19909 593241 20229 593273
rect 25840 593829 26160 593861
rect 25840 593593 25882 593829
rect 26118 593593 26160 593829
rect 25840 593509 26160 593593
rect 25840 593273 25882 593509
rect 26118 593273 26160 593509
rect 25840 593241 26160 593273
rect 31770 593829 32090 593861
rect 31770 593593 31812 593829
rect 32048 593593 32090 593829
rect 31770 593509 32090 593593
rect 31770 593273 31812 593509
rect 32048 593273 32090 593509
rect 31770 593241 32090 593273
rect 47909 593829 48229 593861
rect 47909 593593 47951 593829
rect 48187 593593 48229 593829
rect 47909 593509 48229 593593
rect 47909 593273 47951 593509
rect 48187 593273 48229 593509
rect 47909 593241 48229 593273
rect 53840 593829 54160 593861
rect 53840 593593 53882 593829
rect 54118 593593 54160 593829
rect 53840 593509 54160 593593
rect 53840 593273 53882 593509
rect 54118 593273 54160 593509
rect 53840 593241 54160 593273
rect 59770 593829 60090 593861
rect 59770 593593 59812 593829
rect 60048 593593 60090 593829
rect 59770 593509 60090 593593
rect 59770 593273 59812 593509
rect 60048 593273 60090 593509
rect 59770 593241 60090 593273
rect 75909 593829 76229 593861
rect 75909 593593 75951 593829
rect 76187 593593 76229 593829
rect 75909 593509 76229 593593
rect 75909 593273 75951 593509
rect 76187 593273 76229 593509
rect 75909 593241 76229 593273
rect 81840 593829 82160 593861
rect 81840 593593 81882 593829
rect 82118 593593 82160 593829
rect 81840 593509 82160 593593
rect 81840 593273 81882 593509
rect 82118 593273 82160 593509
rect 81840 593241 82160 593273
rect 87770 593829 88090 593861
rect 87770 593593 87812 593829
rect 88048 593593 88090 593829
rect 87770 593509 88090 593593
rect 87770 593273 87812 593509
rect 88048 593273 88090 593509
rect 87770 593241 88090 593273
rect 103909 593829 104229 593861
rect 103909 593593 103951 593829
rect 104187 593593 104229 593829
rect 103909 593509 104229 593593
rect 103909 593273 103951 593509
rect 104187 593273 104229 593509
rect 103909 593241 104229 593273
rect 109840 593829 110160 593861
rect 109840 593593 109882 593829
rect 110118 593593 110160 593829
rect 109840 593509 110160 593593
rect 109840 593273 109882 593509
rect 110118 593273 110160 593509
rect 109840 593241 110160 593273
rect 115770 593829 116090 593861
rect 115770 593593 115812 593829
rect 116048 593593 116090 593829
rect 115770 593509 116090 593593
rect 115770 593273 115812 593509
rect 116048 593273 116090 593509
rect 115770 593241 116090 593273
rect 131909 593829 132229 593861
rect 131909 593593 131951 593829
rect 132187 593593 132229 593829
rect 131909 593509 132229 593593
rect 131909 593273 131951 593509
rect 132187 593273 132229 593509
rect 131909 593241 132229 593273
rect 137840 593829 138160 593861
rect 137840 593593 137882 593829
rect 138118 593593 138160 593829
rect 137840 593509 138160 593593
rect 137840 593273 137882 593509
rect 138118 593273 138160 593509
rect 137840 593241 138160 593273
rect 143770 593829 144090 593861
rect 143770 593593 143812 593829
rect 144048 593593 144090 593829
rect 143770 593509 144090 593593
rect 143770 593273 143812 593509
rect 144048 593273 144090 593509
rect 143770 593241 144090 593273
rect 159909 593829 160229 593861
rect 159909 593593 159951 593829
rect 160187 593593 160229 593829
rect 159909 593509 160229 593593
rect 159909 593273 159951 593509
rect 160187 593273 160229 593509
rect 159909 593241 160229 593273
rect 165840 593829 166160 593861
rect 165840 593593 165882 593829
rect 166118 593593 166160 593829
rect 165840 593509 166160 593593
rect 165840 593273 165882 593509
rect 166118 593273 166160 593509
rect 165840 593241 166160 593273
rect 171770 593829 172090 593861
rect 171770 593593 171812 593829
rect 172048 593593 172090 593829
rect 171770 593509 172090 593593
rect 171770 593273 171812 593509
rect 172048 593273 172090 593509
rect 171770 593241 172090 593273
rect 187909 593829 188229 593861
rect 187909 593593 187951 593829
rect 188187 593593 188229 593829
rect 187909 593509 188229 593593
rect 187909 593273 187951 593509
rect 188187 593273 188229 593509
rect 187909 593241 188229 593273
rect 193840 593829 194160 593861
rect 193840 593593 193882 593829
rect 194118 593593 194160 593829
rect 193840 593509 194160 593593
rect 193840 593273 193882 593509
rect 194118 593273 194160 593509
rect 193840 593241 194160 593273
rect 199770 593829 200090 593861
rect 199770 593593 199812 593829
rect 200048 593593 200090 593829
rect 199770 593509 200090 593593
rect 199770 593273 199812 593509
rect 200048 593273 200090 593509
rect 199770 593241 200090 593273
rect 215909 593829 216229 593861
rect 215909 593593 215951 593829
rect 216187 593593 216229 593829
rect 215909 593509 216229 593593
rect 215909 593273 215951 593509
rect 216187 593273 216229 593509
rect 215909 593241 216229 593273
rect 221840 593829 222160 593861
rect 221840 593593 221882 593829
rect 222118 593593 222160 593829
rect 221840 593509 222160 593593
rect 221840 593273 221882 593509
rect 222118 593273 222160 593509
rect 221840 593241 222160 593273
rect 227770 593829 228090 593861
rect 227770 593593 227812 593829
rect 228048 593593 228090 593829
rect 227770 593509 228090 593593
rect 227770 593273 227812 593509
rect 228048 593273 228090 593509
rect 227770 593241 228090 593273
rect 243909 593829 244229 593861
rect 243909 593593 243951 593829
rect 244187 593593 244229 593829
rect 243909 593509 244229 593593
rect 243909 593273 243951 593509
rect 244187 593273 244229 593509
rect 243909 593241 244229 593273
rect 249840 593829 250160 593861
rect 249840 593593 249882 593829
rect 250118 593593 250160 593829
rect 249840 593509 250160 593593
rect 249840 593273 249882 593509
rect 250118 593273 250160 593509
rect 249840 593241 250160 593273
rect 255770 593829 256090 593861
rect 255770 593593 255812 593829
rect 256048 593593 256090 593829
rect 255770 593509 256090 593593
rect 255770 593273 255812 593509
rect 256048 593273 256090 593509
rect 255770 593241 256090 593273
rect 271909 593829 272229 593861
rect 271909 593593 271951 593829
rect 272187 593593 272229 593829
rect 271909 593509 272229 593593
rect 271909 593273 271951 593509
rect 272187 593273 272229 593509
rect 271909 593241 272229 593273
rect 277840 593829 278160 593861
rect 277840 593593 277882 593829
rect 278118 593593 278160 593829
rect 277840 593509 278160 593593
rect 277840 593273 277882 593509
rect 278118 593273 278160 593509
rect 277840 593241 278160 593273
rect 283770 593829 284090 593861
rect 283770 593593 283812 593829
rect 284048 593593 284090 593829
rect 283770 593509 284090 593593
rect 283770 593273 283812 593509
rect 284048 593273 284090 593509
rect 283770 593241 284090 593273
rect 299909 593829 300229 593861
rect 299909 593593 299951 593829
rect 300187 593593 300229 593829
rect 299909 593509 300229 593593
rect 299909 593273 299951 593509
rect 300187 593273 300229 593509
rect 299909 593241 300229 593273
rect 305840 593829 306160 593861
rect 305840 593593 305882 593829
rect 306118 593593 306160 593829
rect 305840 593509 306160 593593
rect 305840 593273 305882 593509
rect 306118 593273 306160 593509
rect 305840 593241 306160 593273
rect 311770 593829 312090 593861
rect 311770 593593 311812 593829
rect 312048 593593 312090 593829
rect 311770 593509 312090 593593
rect 311770 593273 311812 593509
rect 312048 593273 312090 593509
rect 311770 593241 312090 593273
rect 327909 593829 328229 593861
rect 327909 593593 327951 593829
rect 328187 593593 328229 593829
rect 327909 593509 328229 593593
rect 327909 593273 327951 593509
rect 328187 593273 328229 593509
rect 327909 593241 328229 593273
rect 333840 593829 334160 593861
rect 333840 593593 333882 593829
rect 334118 593593 334160 593829
rect 333840 593509 334160 593593
rect 333840 593273 333882 593509
rect 334118 593273 334160 593509
rect 333840 593241 334160 593273
rect 339770 593829 340090 593861
rect 339770 593593 339812 593829
rect 340048 593593 340090 593829
rect 339770 593509 340090 593593
rect 339770 593273 339812 593509
rect 340048 593273 340090 593509
rect 339770 593241 340090 593273
rect 355909 593829 356229 593861
rect 355909 593593 355951 593829
rect 356187 593593 356229 593829
rect 355909 593509 356229 593593
rect 355909 593273 355951 593509
rect 356187 593273 356229 593509
rect 355909 593241 356229 593273
rect 361840 593829 362160 593861
rect 361840 593593 361882 593829
rect 362118 593593 362160 593829
rect 361840 593509 362160 593593
rect 361840 593273 361882 593509
rect 362118 593273 362160 593509
rect 361840 593241 362160 593273
rect 367770 593829 368090 593861
rect 367770 593593 367812 593829
rect 368048 593593 368090 593829
rect 367770 593509 368090 593593
rect 367770 593273 367812 593509
rect 368048 593273 368090 593509
rect 367770 593241 368090 593273
rect 383909 593829 384229 593861
rect 383909 593593 383951 593829
rect 384187 593593 384229 593829
rect 383909 593509 384229 593593
rect 383909 593273 383951 593509
rect 384187 593273 384229 593509
rect 383909 593241 384229 593273
rect 389840 593829 390160 593861
rect 389840 593593 389882 593829
rect 390118 593593 390160 593829
rect 389840 593509 390160 593593
rect 389840 593273 389882 593509
rect 390118 593273 390160 593509
rect 389840 593241 390160 593273
rect 395770 593829 396090 593861
rect 395770 593593 395812 593829
rect 396048 593593 396090 593829
rect 395770 593509 396090 593593
rect 395770 593273 395812 593509
rect 396048 593273 396090 593509
rect 395770 593241 396090 593273
rect 411909 593829 412229 593861
rect 411909 593593 411951 593829
rect 412187 593593 412229 593829
rect 411909 593509 412229 593593
rect 411909 593273 411951 593509
rect 412187 593273 412229 593509
rect 411909 593241 412229 593273
rect 417840 593829 418160 593861
rect 417840 593593 417882 593829
rect 418118 593593 418160 593829
rect 417840 593509 418160 593593
rect 417840 593273 417882 593509
rect 418118 593273 418160 593509
rect 417840 593241 418160 593273
rect 423770 593829 424090 593861
rect 423770 593593 423812 593829
rect 424048 593593 424090 593829
rect 423770 593509 424090 593593
rect 423770 593273 423812 593509
rect 424048 593273 424090 593509
rect 423770 593241 424090 593273
rect 439909 593829 440229 593861
rect 439909 593593 439951 593829
rect 440187 593593 440229 593829
rect 439909 593509 440229 593593
rect 439909 593273 439951 593509
rect 440187 593273 440229 593509
rect 439909 593241 440229 593273
rect 445840 593829 446160 593861
rect 445840 593593 445882 593829
rect 446118 593593 446160 593829
rect 445840 593509 446160 593593
rect 445840 593273 445882 593509
rect 446118 593273 446160 593509
rect 445840 593241 446160 593273
rect 451770 593829 452090 593861
rect 451770 593593 451812 593829
rect 452048 593593 452090 593829
rect 451770 593509 452090 593593
rect 451770 593273 451812 593509
rect 452048 593273 452090 593509
rect 451770 593241 452090 593273
rect 467909 593829 468229 593861
rect 467909 593593 467951 593829
rect 468187 593593 468229 593829
rect 467909 593509 468229 593593
rect 467909 593273 467951 593509
rect 468187 593273 468229 593509
rect 467909 593241 468229 593273
rect 473840 593829 474160 593861
rect 473840 593593 473882 593829
rect 474118 593593 474160 593829
rect 473840 593509 474160 593593
rect 473840 593273 473882 593509
rect 474118 593273 474160 593509
rect 473840 593241 474160 593273
rect 479770 593829 480090 593861
rect 479770 593593 479812 593829
rect 480048 593593 480090 593829
rect 479770 593509 480090 593593
rect 479770 593273 479812 593509
rect 480048 593273 480090 593509
rect 479770 593241 480090 593273
rect 495909 593829 496229 593861
rect 495909 593593 495951 593829
rect 496187 593593 496229 593829
rect 495909 593509 496229 593593
rect 495909 593273 495951 593509
rect 496187 593273 496229 593509
rect 495909 593241 496229 593273
rect 501840 593829 502160 593861
rect 501840 593593 501882 593829
rect 502118 593593 502160 593829
rect 501840 593509 502160 593593
rect 501840 593273 501882 593509
rect 502118 593273 502160 593509
rect 501840 593241 502160 593273
rect 507770 593829 508090 593861
rect 507770 593593 507812 593829
rect 508048 593593 508090 593829
rect 507770 593509 508090 593593
rect 507770 593273 507812 593509
rect 508048 593273 508090 593509
rect 507770 593241 508090 593273
rect 523909 593829 524229 593861
rect 523909 593593 523951 593829
rect 524187 593593 524229 593829
rect 523909 593509 524229 593593
rect 523909 593273 523951 593509
rect 524187 593273 524229 593509
rect 523909 593241 524229 593273
rect 529840 593829 530160 593861
rect 529840 593593 529882 593829
rect 530118 593593 530160 593829
rect 529840 593509 530160 593593
rect 529840 593273 529882 593509
rect 530118 593273 530160 593509
rect 529840 593241 530160 593273
rect 535770 593829 536090 593861
rect 535770 593593 535812 593829
rect 536048 593593 536090 593829
rect 535770 593509 536090 593593
rect 535770 593273 535812 593509
rect 536048 593273 536090 593509
rect 535770 593241 536090 593273
rect 551909 593829 552229 593861
rect 551909 593593 551951 593829
rect 552187 593593 552229 593829
rect 551909 593509 552229 593593
rect 551909 593273 551951 593509
rect 552187 593273 552229 593509
rect 551909 593241 552229 593273
rect 557840 593829 558160 593861
rect 557840 593593 557882 593829
rect 558118 593593 558160 593829
rect 557840 593509 558160 593593
rect 557840 593273 557882 593509
rect 558118 593273 558160 593509
rect 557840 593241 558160 593273
rect 563770 593829 564090 593861
rect 563770 593593 563812 593829
rect 564048 593593 564090 593829
rect 563770 593509 564090 593593
rect 563770 593273 563812 593509
rect 564048 593273 564090 593509
rect 563770 593241 564090 593273
rect 573494 593829 574114 620273
rect 573494 593593 573526 593829
rect 573762 593593 573846 593829
rect 574082 593593 574114 593829
rect 573494 593509 574114 593593
rect 573494 593273 573526 593509
rect 573762 593273 573846 593509
rect 574082 593273 574114 593509
rect 22875 590454 23195 590486
rect 22875 590218 22917 590454
rect 23153 590218 23195 590454
rect 22875 590134 23195 590218
rect 22875 589898 22917 590134
rect 23153 589898 23195 590134
rect 22875 589866 23195 589898
rect 28806 590454 29126 590486
rect 28806 590218 28848 590454
rect 29084 590218 29126 590454
rect 28806 590134 29126 590218
rect 28806 589898 28848 590134
rect 29084 589898 29126 590134
rect 28806 589866 29126 589898
rect 50875 590454 51195 590486
rect 50875 590218 50917 590454
rect 51153 590218 51195 590454
rect 50875 590134 51195 590218
rect 50875 589898 50917 590134
rect 51153 589898 51195 590134
rect 50875 589866 51195 589898
rect 56806 590454 57126 590486
rect 56806 590218 56848 590454
rect 57084 590218 57126 590454
rect 56806 590134 57126 590218
rect 56806 589898 56848 590134
rect 57084 589898 57126 590134
rect 56806 589866 57126 589898
rect 78875 590454 79195 590486
rect 78875 590218 78917 590454
rect 79153 590218 79195 590454
rect 78875 590134 79195 590218
rect 78875 589898 78917 590134
rect 79153 589898 79195 590134
rect 78875 589866 79195 589898
rect 84806 590454 85126 590486
rect 84806 590218 84848 590454
rect 85084 590218 85126 590454
rect 84806 590134 85126 590218
rect 84806 589898 84848 590134
rect 85084 589898 85126 590134
rect 84806 589866 85126 589898
rect 106875 590454 107195 590486
rect 106875 590218 106917 590454
rect 107153 590218 107195 590454
rect 106875 590134 107195 590218
rect 106875 589898 106917 590134
rect 107153 589898 107195 590134
rect 106875 589866 107195 589898
rect 112806 590454 113126 590486
rect 112806 590218 112848 590454
rect 113084 590218 113126 590454
rect 112806 590134 113126 590218
rect 112806 589898 112848 590134
rect 113084 589898 113126 590134
rect 112806 589866 113126 589898
rect 134875 590454 135195 590486
rect 134875 590218 134917 590454
rect 135153 590218 135195 590454
rect 134875 590134 135195 590218
rect 134875 589898 134917 590134
rect 135153 589898 135195 590134
rect 134875 589866 135195 589898
rect 140806 590454 141126 590486
rect 140806 590218 140848 590454
rect 141084 590218 141126 590454
rect 140806 590134 141126 590218
rect 140806 589898 140848 590134
rect 141084 589898 141126 590134
rect 140806 589866 141126 589898
rect 162875 590454 163195 590486
rect 162875 590218 162917 590454
rect 163153 590218 163195 590454
rect 162875 590134 163195 590218
rect 162875 589898 162917 590134
rect 163153 589898 163195 590134
rect 162875 589866 163195 589898
rect 168806 590454 169126 590486
rect 168806 590218 168848 590454
rect 169084 590218 169126 590454
rect 168806 590134 169126 590218
rect 168806 589898 168848 590134
rect 169084 589898 169126 590134
rect 168806 589866 169126 589898
rect 190875 590454 191195 590486
rect 190875 590218 190917 590454
rect 191153 590218 191195 590454
rect 190875 590134 191195 590218
rect 190875 589898 190917 590134
rect 191153 589898 191195 590134
rect 190875 589866 191195 589898
rect 196806 590454 197126 590486
rect 196806 590218 196848 590454
rect 197084 590218 197126 590454
rect 196806 590134 197126 590218
rect 196806 589898 196848 590134
rect 197084 589898 197126 590134
rect 196806 589866 197126 589898
rect 218875 590454 219195 590486
rect 218875 590218 218917 590454
rect 219153 590218 219195 590454
rect 218875 590134 219195 590218
rect 218875 589898 218917 590134
rect 219153 589898 219195 590134
rect 218875 589866 219195 589898
rect 224806 590454 225126 590486
rect 224806 590218 224848 590454
rect 225084 590218 225126 590454
rect 224806 590134 225126 590218
rect 224806 589898 224848 590134
rect 225084 589898 225126 590134
rect 224806 589866 225126 589898
rect 246875 590454 247195 590486
rect 246875 590218 246917 590454
rect 247153 590218 247195 590454
rect 246875 590134 247195 590218
rect 246875 589898 246917 590134
rect 247153 589898 247195 590134
rect 246875 589866 247195 589898
rect 252806 590454 253126 590486
rect 252806 590218 252848 590454
rect 253084 590218 253126 590454
rect 252806 590134 253126 590218
rect 252806 589898 252848 590134
rect 253084 589898 253126 590134
rect 252806 589866 253126 589898
rect 274875 590454 275195 590486
rect 274875 590218 274917 590454
rect 275153 590218 275195 590454
rect 274875 590134 275195 590218
rect 274875 589898 274917 590134
rect 275153 589898 275195 590134
rect 274875 589866 275195 589898
rect 280806 590454 281126 590486
rect 280806 590218 280848 590454
rect 281084 590218 281126 590454
rect 280806 590134 281126 590218
rect 280806 589898 280848 590134
rect 281084 589898 281126 590134
rect 280806 589866 281126 589898
rect 302875 590454 303195 590486
rect 302875 590218 302917 590454
rect 303153 590218 303195 590454
rect 302875 590134 303195 590218
rect 302875 589898 302917 590134
rect 303153 589898 303195 590134
rect 302875 589866 303195 589898
rect 308806 590454 309126 590486
rect 308806 590218 308848 590454
rect 309084 590218 309126 590454
rect 308806 590134 309126 590218
rect 308806 589898 308848 590134
rect 309084 589898 309126 590134
rect 308806 589866 309126 589898
rect 330875 590454 331195 590486
rect 330875 590218 330917 590454
rect 331153 590218 331195 590454
rect 330875 590134 331195 590218
rect 330875 589898 330917 590134
rect 331153 589898 331195 590134
rect 330875 589866 331195 589898
rect 336806 590454 337126 590486
rect 336806 590218 336848 590454
rect 337084 590218 337126 590454
rect 336806 590134 337126 590218
rect 336806 589898 336848 590134
rect 337084 589898 337126 590134
rect 336806 589866 337126 589898
rect 358875 590454 359195 590486
rect 358875 590218 358917 590454
rect 359153 590218 359195 590454
rect 358875 590134 359195 590218
rect 358875 589898 358917 590134
rect 359153 589898 359195 590134
rect 358875 589866 359195 589898
rect 364806 590454 365126 590486
rect 364806 590218 364848 590454
rect 365084 590218 365126 590454
rect 364806 590134 365126 590218
rect 364806 589898 364848 590134
rect 365084 589898 365126 590134
rect 364806 589866 365126 589898
rect 386875 590454 387195 590486
rect 386875 590218 386917 590454
rect 387153 590218 387195 590454
rect 386875 590134 387195 590218
rect 386875 589898 386917 590134
rect 387153 589898 387195 590134
rect 386875 589866 387195 589898
rect 392806 590454 393126 590486
rect 392806 590218 392848 590454
rect 393084 590218 393126 590454
rect 392806 590134 393126 590218
rect 392806 589898 392848 590134
rect 393084 589898 393126 590134
rect 392806 589866 393126 589898
rect 414875 590454 415195 590486
rect 414875 590218 414917 590454
rect 415153 590218 415195 590454
rect 414875 590134 415195 590218
rect 414875 589898 414917 590134
rect 415153 589898 415195 590134
rect 414875 589866 415195 589898
rect 420806 590454 421126 590486
rect 420806 590218 420848 590454
rect 421084 590218 421126 590454
rect 420806 590134 421126 590218
rect 420806 589898 420848 590134
rect 421084 589898 421126 590134
rect 420806 589866 421126 589898
rect 442875 590454 443195 590486
rect 442875 590218 442917 590454
rect 443153 590218 443195 590454
rect 442875 590134 443195 590218
rect 442875 589898 442917 590134
rect 443153 589898 443195 590134
rect 442875 589866 443195 589898
rect 448806 590454 449126 590486
rect 448806 590218 448848 590454
rect 449084 590218 449126 590454
rect 448806 590134 449126 590218
rect 448806 589898 448848 590134
rect 449084 589898 449126 590134
rect 448806 589866 449126 589898
rect 470875 590454 471195 590486
rect 470875 590218 470917 590454
rect 471153 590218 471195 590454
rect 470875 590134 471195 590218
rect 470875 589898 470917 590134
rect 471153 589898 471195 590134
rect 470875 589866 471195 589898
rect 476806 590454 477126 590486
rect 476806 590218 476848 590454
rect 477084 590218 477126 590454
rect 476806 590134 477126 590218
rect 476806 589898 476848 590134
rect 477084 589898 477126 590134
rect 476806 589866 477126 589898
rect 498875 590454 499195 590486
rect 498875 590218 498917 590454
rect 499153 590218 499195 590454
rect 498875 590134 499195 590218
rect 498875 589898 498917 590134
rect 499153 589898 499195 590134
rect 498875 589866 499195 589898
rect 504806 590454 505126 590486
rect 504806 590218 504848 590454
rect 505084 590218 505126 590454
rect 504806 590134 505126 590218
rect 504806 589898 504848 590134
rect 505084 589898 505126 590134
rect 504806 589866 505126 589898
rect 526875 590454 527195 590486
rect 526875 590218 526917 590454
rect 527153 590218 527195 590454
rect 526875 590134 527195 590218
rect 526875 589898 526917 590134
rect 527153 589898 527195 590134
rect 526875 589866 527195 589898
rect 532806 590454 533126 590486
rect 532806 590218 532848 590454
rect 533084 590218 533126 590454
rect 532806 590134 533126 590218
rect 532806 589898 532848 590134
rect 533084 589898 533126 590134
rect 532806 589866 533126 589898
rect 554875 590454 555195 590486
rect 554875 590218 554917 590454
rect 555153 590218 555195 590454
rect 554875 590134 555195 590218
rect 554875 589898 554917 590134
rect 555153 589898 555195 590134
rect 554875 589866 555195 589898
rect 560806 590454 561126 590486
rect 560806 590218 560848 590454
rect 561084 590218 561126 590454
rect 560806 590134 561126 590218
rect 560806 589898 560848 590134
rect 561084 589898 561126 590134
rect 560806 589866 561126 589898
rect -2006 566593 -1974 566829
rect -1738 566593 -1654 566829
rect -1418 566593 -1386 566829
rect -2006 566509 -1386 566593
rect -2006 566273 -1974 566509
rect -1738 566273 -1654 566509
rect -1418 566273 -1386 566509
rect -2006 539829 -1386 566273
rect 19910 566829 20230 566861
rect 19910 566593 19952 566829
rect 20188 566593 20230 566829
rect 19910 566509 20230 566593
rect 19910 566273 19952 566509
rect 20188 566273 20230 566509
rect 19910 566241 20230 566273
rect 25840 566829 26160 566861
rect 25840 566593 25882 566829
rect 26118 566593 26160 566829
rect 25840 566509 26160 566593
rect 25840 566273 25882 566509
rect 26118 566273 26160 566509
rect 25840 566241 26160 566273
rect 31771 566829 32091 566861
rect 31771 566593 31813 566829
rect 32049 566593 32091 566829
rect 31771 566509 32091 566593
rect 31771 566273 31813 566509
rect 32049 566273 32091 566509
rect 31771 566241 32091 566273
rect 47910 566829 48230 566861
rect 47910 566593 47952 566829
rect 48188 566593 48230 566829
rect 47910 566509 48230 566593
rect 47910 566273 47952 566509
rect 48188 566273 48230 566509
rect 47910 566241 48230 566273
rect 53840 566829 54160 566861
rect 53840 566593 53882 566829
rect 54118 566593 54160 566829
rect 53840 566509 54160 566593
rect 53840 566273 53882 566509
rect 54118 566273 54160 566509
rect 53840 566241 54160 566273
rect 59771 566829 60091 566861
rect 59771 566593 59813 566829
rect 60049 566593 60091 566829
rect 59771 566509 60091 566593
rect 59771 566273 59813 566509
rect 60049 566273 60091 566509
rect 59771 566241 60091 566273
rect 75910 566829 76230 566861
rect 75910 566593 75952 566829
rect 76188 566593 76230 566829
rect 75910 566509 76230 566593
rect 75910 566273 75952 566509
rect 76188 566273 76230 566509
rect 75910 566241 76230 566273
rect 81840 566829 82160 566861
rect 81840 566593 81882 566829
rect 82118 566593 82160 566829
rect 81840 566509 82160 566593
rect 81840 566273 81882 566509
rect 82118 566273 82160 566509
rect 81840 566241 82160 566273
rect 87771 566829 88091 566861
rect 87771 566593 87813 566829
rect 88049 566593 88091 566829
rect 87771 566509 88091 566593
rect 87771 566273 87813 566509
rect 88049 566273 88091 566509
rect 87771 566241 88091 566273
rect 103910 566829 104230 566861
rect 103910 566593 103952 566829
rect 104188 566593 104230 566829
rect 103910 566509 104230 566593
rect 103910 566273 103952 566509
rect 104188 566273 104230 566509
rect 103910 566241 104230 566273
rect 109840 566829 110160 566861
rect 109840 566593 109882 566829
rect 110118 566593 110160 566829
rect 109840 566509 110160 566593
rect 109840 566273 109882 566509
rect 110118 566273 110160 566509
rect 109840 566241 110160 566273
rect 115771 566829 116091 566861
rect 115771 566593 115813 566829
rect 116049 566593 116091 566829
rect 115771 566509 116091 566593
rect 115771 566273 115813 566509
rect 116049 566273 116091 566509
rect 115771 566241 116091 566273
rect 131910 566829 132230 566861
rect 131910 566593 131952 566829
rect 132188 566593 132230 566829
rect 131910 566509 132230 566593
rect 131910 566273 131952 566509
rect 132188 566273 132230 566509
rect 131910 566241 132230 566273
rect 137840 566829 138160 566861
rect 137840 566593 137882 566829
rect 138118 566593 138160 566829
rect 137840 566509 138160 566593
rect 137840 566273 137882 566509
rect 138118 566273 138160 566509
rect 137840 566241 138160 566273
rect 143771 566829 144091 566861
rect 143771 566593 143813 566829
rect 144049 566593 144091 566829
rect 143771 566509 144091 566593
rect 143771 566273 143813 566509
rect 144049 566273 144091 566509
rect 143771 566241 144091 566273
rect 159910 566829 160230 566861
rect 159910 566593 159952 566829
rect 160188 566593 160230 566829
rect 159910 566509 160230 566593
rect 159910 566273 159952 566509
rect 160188 566273 160230 566509
rect 159910 566241 160230 566273
rect 165840 566829 166160 566861
rect 165840 566593 165882 566829
rect 166118 566593 166160 566829
rect 165840 566509 166160 566593
rect 165840 566273 165882 566509
rect 166118 566273 166160 566509
rect 165840 566241 166160 566273
rect 171771 566829 172091 566861
rect 171771 566593 171813 566829
rect 172049 566593 172091 566829
rect 171771 566509 172091 566593
rect 171771 566273 171813 566509
rect 172049 566273 172091 566509
rect 171771 566241 172091 566273
rect 187910 566829 188230 566861
rect 187910 566593 187952 566829
rect 188188 566593 188230 566829
rect 187910 566509 188230 566593
rect 187910 566273 187952 566509
rect 188188 566273 188230 566509
rect 187910 566241 188230 566273
rect 193840 566829 194160 566861
rect 193840 566593 193882 566829
rect 194118 566593 194160 566829
rect 193840 566509 194160 566593
rect 193840 566273 193882 566509
rect 194118 566273 194160 566509
rect 193840 566241 194160 566273
rect 199771 566829 200091 566861
rect 199771 566593 199813 566829
rect 200049 566593 200091 566829
rect 199771 566509 200091 566593
rect 199771 566273 199813 566509
rect 200049 566273 200091 566509
rect 199771 566241 200091 566273
rect 215910 566829 216230 566861
rect 215910 566593 215952 566829
rect 216188 566593 216230 566829
rect 215910 566509 216230 566593
rect 215910 566273 215952 566509
rect 216188 566273 216230 566509
rect 215910 566241 216230 566273
rect 221840 566829 222160 566861
rect 221840 566593 221882 566829
rect 222118 566593 222160 566829
rect 221840 566509 222160 566593
rect 221840 566273 221882 566509
rect 222118 566273 222160 566509
rect 221840 566241 222160 566273
rect 227771 566829 228091 566861
rect 227771 566593 227813 566829
rect 228049 566593 228091 566829
rect 227771 566509 228091 566593
rect 227771 566273 227813 566509
rect 228049 566273 228091 566509
rect 227771 566241 228091 566273
rect 243910 566829 244230 566861
rect 243910 566593 243952 566829
rect 244188 566593 244230 566829
rect 243910 566509 244230 566593
rect 243910 566273 243952 566509
rect 244188 566273 244230 566509
rect 243910 566241 244230 566273
rect 249840 566829 250160 566861
rect 249840 566593 249882 566829
rect 250118 566593 250160 566829
rect 249840 566509 250160 566593
rect 249840 566273 249882 566509
rect 250118 566273 250160 566509
rect 249840 566241 250160 566273
rect 255771 566829 256091 566861
rect 255771 566593 255813 566829
rect 256049 566593 256091 566829
rect 255771 566509 256091 566593
rect 255771 566273 255813 566509
rect 256049 566273 256091 566509
rect 255771 566241 256091 566273
rect 271910 566829 272230 566861
rect 271910 566593 271952 566829
rect 272188 566593 272230 566829
rect 271910 566509 272230 566593
rect 271910 566273 271952 566509
rect 272188 566273 272230 566509
rect 271910 566241 272230 566273
rect 277840 566829 278160 566861
rect 277840 566593 277882 566829
rect 278118 566593 278160 566829
rect 277840 566509 278160 566593
rect 277840 566273 277882 566509
rect 278118 566273 278160 566509
rect 277840 566241 278160 566273
rect 283771 566829 284091 566861
rect 283771 566593 283813 566829
rect 284049 566593 284091 566829
rect 283771 566509 284091 566593
rect 283771 566273 283813 566509
rect 284049 566273 284091 566509
rect 283771 566241 284091 566273
rect 299910 566829 300230 566861
rect 299910 566593 299952 566829
rect 300188 566593 300230 566829
rect 299910 566509 300230 566593
rect 299910 566273 299952 566509
rect 300188 566273 300230 566509
rect 299910 566241 300230 566273
rect 305840 566829 306160 566861
rect 305840 566593 305882 566829
rect 306118 566593 306160 566829
rect 305840 566509 306160 566593
rect 305840 566273 305882 566509
rect 306118 566273 306160 566509
rect 305840 566241 306160 566273
rect 311771 566829 312091 566861
rect 311771 566593 311813 566829
rect 312049 566593 312091 566829
rect 311771 566509 312091 566593
rect 311771 566273 311813 566509
rect 312049 566273 312091 566509
rect 311771 566241 312091 566273
rect 327910 566829 328230 566861
rect 327910 566593 327952 566829
rect 328188 566593 328230 566829
rect 327910 566509 328230 566593
rect 327910 566273 327952 566509
rect 328188 566273 328230 566509
rect 327910 566241 328230 566273
rect 333840 566829 334160 566861
rect 333840 566593 333882 566829
rect 334118 566593 334160 566829
rect 333840 566509 334160 566593
rect 333840 566273 333882 566509
rect 334118 566273 334160 566509
rect 333840 566241 334160 566273
rect 339771 566829 340091 566861
rect 339771 566593 339813 566829
rect 340049 566593 340091 566829
rect 339771 566509 340091 566593
rect 339771 566273 339813 566509
rect 340049 566273 340091 566509
rect 339771 566241 340091 566273
rect 355910 566829 356230 566861
rect 355910 566593 355952 566829
rect 356188 566593 356230 566829
rect 355910 566509 356230 566593
rect 355910 566273 355952 566509
rect 356188 566273 356230 566509
rect 355910 566241 356230 566273
rect 361840 566829 362160 566861
rect 361840 566593 361882 566829
rect 362118 566593 362160 566829
rect 361840 566509 362160 566593
rect 361840 566273 361882 566509
rect 362118 566273 362160 566509
rect 361840 566241 362160 566273
rect 367771 566829 368091 566861
rect 367771 566593 367813 566829
rect 368049 566593 368091 566829
rect 367771 566509 368091 566593
rect 367771 566273 367813 566509
rect 368049 566273 368091 566509
rect 367771 566241 368091 566273
rect 383910 566829 384230 566861
rect 383910 566593 383952 566829
rect 384188 566593 384230 566829
rect 383910 566509 384230 566593
rect 383910 566273 383952 566509
rect 384188 566273 384230 566509
rect 383910 566241 384230 566273
rect 389840 566829 390160 566861
rect 389840 566593 389882 566829
rect 390118 566593 390160 566829
rect 389840 566509 390160 566593
rect 389840 566273 389882 566509
rect 390118 566273 390160 566509
rect 389840 566241 390160 566273
rect 395771 566829 396091 566861
rect 395771 566593 395813 566829
rect 396049 566593 396091 566829
rect 395771 566509 396091 566593
rect 395771 566273 395813 566509
rect 396049 566273 396091 566509
rect 395771 566241 396091 566273
rect 411910 566829 412230 566861
rect 411910 566593 411952 566829
rect 412188 566593 412230 566829
rect 411910 566509 412230 566593
rect 411910 566273 411952 566509
rect 412188 566273 412230 566509
rect 411910 566241 412230 566273
rect 417840 566829 418160 566861
rect 417840 566593 417882 566829
rect 418118 566593 418160 566829
rect 417840 566509 418160 566593
rect 417840 566273 417882 566509
rect 418118 566273 418160 566509
rect 417840 566241 418160 566273
rect 423771 566829 424091 566861
rect 423771 566593 423813 566829
rect 424049 566593 424091 566829
rect 423771 566509 424091 566593
rect 423771 566273 423813 566509
rect 424049 566273 424091 566509
rect 423771 566241 424091 566273
rect 439910 566829 440230 566861
rect 439910 566593 439952 566829
rect 440188 566593 440230 566829
rect 439910 566509 440230 566593
rect 439910 566273 439952 566509
rect 440188 566273 440230 566509
rect 439910 566241 440230 566273
rect 445840 566829 446160 566861
rect 445840 566593 445882 566829
rect 446118 566593 446160 566829
rect 445840 566509 446160 566593
rect 445840 566273 445882 566509
rect 446118 566273 446160 566509
rect 445840 566241 446160 566273
rect 451771 566829 452091 566861
rect 451771 566593 451813 566829
rect 452049 566593 452091 566829
rect 451771 566509 452091 566593
rect 451771 566273 451813 566509
rect 452049 566273 452091 566509
rect 451771 566241 452091 566273
rect 467910 566829 468230 566861
rect 467910 566593 467952 566829
rect 468188 566593 468230 566829
rect 467910 566509 468230 566593
rect 467910 566273 467952 566509
rect 468188 566273 468230 566509
rect 467910 566241 468230 566273
rect 473840 566829 474160 566861
rect 473840 566593 473882 566829
rect 474118 566593 474160 566829
rect 473840 566509 474160 566593
rect 473840 566273 473882 566509
rect 474118 566273 474160 566509
rect 473840 566241 474160 566273
rect 479771 566829 480091 566861
rect 479771 566593 479813 566829
rect 480049 566593 480091 566829
rect 479771 566509 480091 566593
rect 479771 566273 479813 566509
rect 480049 566273 480091 566509
rect 479771 566241 480091 566273
rect 495910 566829 496230 566861
rect 495910 566593 495952 566829
rect 496188 566593 496230 566829
rect 495910 566509 496230 566593
rect 495910 566273 495952 566509
rect 496188 566273 496230 566509
rect 495910 566241 496230 566273
rect 501840 566829 502160 566861
rect 501840 566593 501882 566829
rect 502118 566593 502160 566829
rect 501840 566509 502160 566593
rect 501840 566273 501882 566509
rect 502118 566273 502160 566509
rect 501840 566241 502160 566273
rect 507771 566829 508091 566861
rect 507771 566593 507813 566829
rect 508049 566593 508091 566829
rect 507771 566509 508091 566593
rect 507771 566273 507813 566509
rect 508049 566273 508091 566509
rect 507771 566241 508091 566273
rect 523910 566829 524230 566861
rect 523910 566593 523952 566829
rect 524188 566593 524230 566829
rect 523910 566509 524230 566593
rect 523910 566273 523952 566509
rect 524188 566273 524230 566509
rect 523910 566241 524230 566273
rect 529840 566829 530160 566861
rect 529840 566593 529882 566829
rect 530118 566593 530160 566829
rect 529840 566509 530160 566593
rect 529840 566273 529882 566509
rect 530118 566273 530160 566509
rect 529840 566241 530160 566273
rect 535771 566829 536091 566861
rect 535771 566593 535813 566829
rect 536049 566593 536091 566829
rect 535771 566509 536091 566593
rect 535771 566273 535813 566509
rect 536049 566273 536091 566509
rect 535771 566241 536091 566273
rect 551910 566829 552230 566861
rect 551910 566593 551952 566829
rect 552188 566593 552230 566829
rect 551910 566509 552230 566593
rect 551910 566273 551952 566509
rect 552188 566273 552230 566509
rect 551910 566241 552230 566273
rect 557840 566829 558160 566861
rect 557840 566593 557882 566829
rect 558118 566593 558160 566829
rect 557840 566509 558160 566593
rect 557840 566273 557882 566509
rect 558118 566273 558160 566509
rect 557840 566241 558160 566273
rect 563771 566829 564091 566861
rect 563771 566593 563813 566829
rect 564049 566593 564091 566829
rect 563771 566509 564091 566593
rect 563771 566273 563813 566509
rect 564049 566273 564091 566509
rect 563771 566241 564091 566273
rect 573494 566829 574114 593273
rect 573494 566593 573526 566829
rect 573762 566593 573846 566829
rect 574082 566593 574114 566829
rect 573494 566509 574114 566593
rect 573494 566273 573526 566509
rect 573762 566273 573846 566509
rect 574082 566273 574114 566509
rect 22874 563454 23194 563486
rect 22874 563218 22916 563454
rect 23152 563218 23194 563454
rect 22874 563134 23194 563218
rect 22874 562898 22916 563134
rect 23152 562898 23194 563134
rect 22874 562866 23194 562898
rect 28805 563454 29125 563486
rect 28805 563218 28847 563454
rect 29083 563218 29125 563454
rect 28805 563134 29125 563218
rect 28805 562898 28847 563134
rect 29083 562898 29125 563134
rect 28805 562866 29125 562898
rect 50874 563454 51194 563486
rect 50874 563218 50916 563454
rect 51152 563218 51194 563454
rect 50874 563134 51194 563218
rect 50874 562898 50916 563134
rect 51152 562898 51194 563134
rect 50874 562866 51194 562898
rect 56805 563454 57125 563486
rect 56805 563218 56847 563454
rect 57083 563218 57125 563454
rect 56805 563134 57125 563218
rect 56805 562898 56847 563134
rect 57083 562898 57125 563134
rect 56805 562866 57125 562898
rect 78874 563454 79194 563486
rect 78874 563218 78916 563454
rect 79152 563218 79194 563454
rect 78874 563134 79194 563218
rect 78874 562898 78916 563134
rect 79152 562898 79194 563134
rect 78874 562866 79194 562898
rect 84805 563454 85125 563486
rect 84805 563218 84847 563454
rect 85083 563218 85125 563454
rect 84805 563134 85125 563218
rect 84805 562898 84847 563134
rect 85083 562898 85125 563134
rect 84805 562866 85125 562898
rect 106874 563454 107194 563486
rect 106874 563218 106916 563454
rect 107152 563218 107194 563454
rect 106874 563134 107194 563218
rect 106874 562898 106916 563134
rect 107152 562898 107194 563134
rect 106874 562866 107194 562898
rect 112805 563454 113125 563486
rect 112805 563218 112847 563454
rect 113083 563218 113125 563454
rect 112805 563134 113125 563218
rect 112805 562898 112847 563134
rect 113083 562898 113125 563134
rect 112805 562866 113125 562898
rect 134874 563454 135194 563486
rect 134874 563218 134916 563454
rect 135152 563218 135194 563454
rect 134874 563134 135194 563218
rect 134874 562898 134916 563134
rect 135152 562898 135194 563134
rect 134874 562866 135194 562898
rect 140805 563454 141125 563486
rect 140805 563218 140847 563454
rect 141083 563218 141125 563454
rect 140805 563134 141125 563218
rect 140805 562898 140847 563134
rect 141083 562898 141125 563134
rect 140805 562866 141125 562898
rect 162874 563454 163194 563486
rect 162874 563218 162916 563454
rect 163152 563218 163194 563454
rect 162874 563134 163194 563218
rect 162874 562898 162916 563134
rect 163152 562898 163194 563134
rect 162874 562866 163194 562898
rect 168805 563454 169125 563486
rect 168805 563218 168847 563454
rect 169083 563218 169125 563454
rect 168805 563134 169125 563218
rect 168805 562898 168847 563134
rect 169083 562898 169125 563134
rect 168805 562866 169125 562898
rect 190874 563454 191194 563486
rect 190874 563218 190916 563454
rect 191152 563218 191194 563454
rect 190874 563134 191194 563218
rect 190874 562898 190916 563134
rect 191152 562898 191194 563134
rect 190874 562866 191194 562898
rect 196805 563454 197125 563486
rect 196805 563218 196847 563454
rect 197083 563218 197125 563454
rect 196805 563134 197125 563218
rect 196805 562898 196847 563134
rect 197083 562898 197125 563134
rect 196805 562866 197125 562898
rect 218874 563454 219194 563486
rect 218874 563218 218916 563454
rect 219152 563218 219194 563454
rect 218874 563134 219194 563218
rect 218874 562898 218916 563134
rect 219152 562898 219194 563134
rect 218874 562866 219194 562898
rect 224805 563454 225125 563486
rect 224805 563218 224847 563454
rect 225083 563218 225125 563454
rect 224805 563134 225125 563218
rect 224805 562898 224847 563134
rect 225083 562898 225125 563134
rect 224805 562866 225125 562898
rect 246874 563454 247194 563486
rect 246874 563218 246916 563454
rect 247152 563218 247194 563454
rect 246874 563134 247194 563218
rect 246874 562898 246916 563134
rect 247152 562898 247194 563134
rect 246874 562866 247194 562898
rect 252805 563454 253125 563486
rect 252805 563218 252847 563454
rect 253083 563218 253125 563454
rect 252805 563134 253125 563218
rect 252805 562898 252847 563134
rect 253083 562898 253125 563134
rect 252805 562866 253125 562898
rect 274874 563454 275194 563486
rect 274874 563218 274916 563454
rect 275152 563218 275194 563454
rect 274874 563134 275194 563218
rect 274874 562898 274916 563134
rect 275152 562898 275194 563134
rect 274874 562866 275194 562898
rect 280805 563454 281125 563486
rect 280805 563218 280847 563454
rect 281083 563218 281125 563454
rect 280805 563134 281125 563218
rect 280805 562898 280847 563134
rect 281083 562898 281125 563134
rect 280805 562866 281125 562898
rect 302874 563454 303194 563486
rect 302874 563218 302916 563454
rect 303152 563218 303194 563454
rect 302874 563134 303194 563218
rect 302874 562898 302916 563134
rect 303152 562898 303194 563134
rect 302874 562866 303194 562898
rect 308805 563454 309125 563486
rect 308805 563218 308847 563454
rect 309083 563218 309125 563454
rect 308805 563134 309125 563218
rect 308805 562898 308847 563134
rect 309083 562898 309125 563134
rect 308805 562866 309125 562898
rect 330874 563454 331194 563486
rect 330874 563218 330916 563454
rect 331152 563218 331194 563454
rect 330874 563134 331194 563218
rect 330874 562898 330916 563134
rect 331152 562898 331194 563134
rect 330874 562866 331194 562898
rect 336805 563454 337125 563486
rect 336805 563218 336847 563454
rect 337083 563218 337125 563454
rect 336805 563134 337125 563218
rect 336805 562898 336847 563134
rect 337083 562898 337125 563134
rect 336805 562866 337125 562898
rect 358874 563454 359194 563486
rect 358874 563218 358916 563454
rect 359152 563218 359194 563454
rect 358874 563134 359194 563218
rect 358874 562898 358916 563134
rect 359152 562898 359194 563134
rect 358874 562866 359194 562898
rect 364805 563454 365125 563486
rect 364805 563218 364847 563454
rect 365083 563218 365125 563454
rect 364805 563134 365125 563218
rect 364805 562898 364847 563134
rect 365083 562898 365125 563134
rect 364805 562866 365125 562898
rect 386874 563454 387194 563486
rect 386874 563218 386916 563454
rect 387152 563218 387194 563454
rect 386874 563134 387194 563218
rect 386874 562898 386916 563134
rect 387152 562898 387194 563134
rect 386874 562866 387194 562898
rect 392805 563454 393125 563486
rect 392805 563218 392847 563454
rect 393083 563218 393125 563454
rect 392805 563134 393125 563218
rect 392805 562898 392847 563134
rect 393083 562898 393125 563134
rect 392805 562866 393125 562898
rect 414874 563454 415194 563486
rect 414874 563218 414916 563454
rect 415152 563218 415194 563454
rect 414874 563134 415194 563218
rect 414874 562898 414916 563134
rect 415152 562898 415194 563134
rect 414874 562866 415194 562898
rect 420805 563454 421125 563486
rect 420805 563218 420847 563454
rect 421083 563218 421125 563454
rect 420805 563134 421125 563218
rect 420805 562898 420847 563134
rect 421083 562898 421125 563134
rect 420805 562866 421125 562898
rect 442874 563454 443194 563486
rect 442874 563218 442916 563454
rect 443152 563218 443194 563454
rect 442874 563134 443194 563218
rect 442874 562898 442916 563134
rect 443152 562898 443194 563134
rect 442874 562866 443194 562898
rect 448805 563454 449125 563486
rect 448805 563218 448847 563454
rect 449083 563218 449125 563454
rect 448805 563134 449125 563218
rect 448805 562898 448847 563134
rect 449083 562898 449125 563134
rect 448805 562866 449125 562898
rect 470874 563454 471194 563486
rect 470874 563218 470916 563454
rect 471152 563218 471194 563454
rect 470874 563134 471194 563218
rect 470874 562898 470916 563134
rect 471152 562898 471194 563134
rect 470874 562866 471194 562898
rect 476805 563454 477125 563486
rect 476805 563218 476847 563454
rect 477083 563218 477125 563454
rect 476805 563134 477125 563218
rect 476805 562898 476847 563134
rect 477083 562898 477125 563134
rect 476805 562866 477125 562898
rect 498874 563454 499194 563486
rect 498874 563218 498916 563454
rect 499152 563218 499194 563454
rect 498874 563134 499194 563218
rect 498874 562898 498916 563134
rect 499152 562898 499194 563134
rect 498874 562866 499194 562898
rect 504805 563454 505125 563486
rect 504805 563218 504847 563454
rect 505083 563218 505125 563454
rect 504805 563134 505125 563218
rect 504805 562898 504847 563134
rect 505083 562898 505125 563134
rect 504805 562866 505125 562898
rect 526874 563454 527194 563486
rect 526874 563218 526916 563454
rect 527152 563218 527194 563454
rect 526874 563134 527194 563218
rect 526874 562898 526916 563134
rect 527152 562898 527194 563134
rect 526874 562866 527194 562898
rect 532805 563454 533125 563486
rect 532805 563218 532847 563454
rect 533083 563218 533125 563454
rect 532805 563134 533125 563218
rect 532805 562898 532847 563134
rect 533083 562898 533125 563134
rect 532805 562866 533125 562898
rect 554874 563454 555194 563486
rect 554874 563218 554916 563454
rect 555152 563218 555194 563454
rect 554874 563134 555194 563218
rect 554874 562898 554916 563134
rect 555152 562898 555194 563134
rect 554874 562866 555194 562898
rect 560805 563454 561125 563486
rect 560805 563218 560847 563454
rect 561083 563218 561125 563454
rect 560805 563134 561125 563218
rect 560805 562898 560847 563134
rect 561083 562898 561125 563134
rect 560805 562866 561125 562898
rect -2006 539593 -1974 539829
rect -1738 539593 -1654 539829
rect -1418 539593 -1386 539829
rect -2006 539509 -1386 539593
rect -2006 539273 -1974 539509
rect -1738 539273 -1654 539509
rect -1418 539273 -1386 539509
rect -2006 512829 -1386 539273
rect 19909 539829 20229 539861
rect 19909 539593 19951 539829
rect 20187 539593 20229 539829
rect 19909 539509 20229 539593
rect 19909 539273 19951 539509
rect 20187 539273 20229 539509
rect 19909 539241 20229 539273
rect 25840 539829 26160 539861
rect 25840 539593 25882 539829
rect 26118 539593 26160 539829
rect 25840 539509 26160 539593
rect 25840 539273 25882 539509
rect 26118 539273 26160 539509
rect 25840 539241 26160 539273
rect 31770 539829 32090 539861
rect 31770 539593 31812 539829
rect 32048 539593 32090 539829
rect 31770 539509 32090 539593
rect 31770 539273 31812 539509
rect 32048 539273 32090 539509
rect 31770 539241 32090 539273
rect 47909 539829 48229 539861
rect 47909 539593 47951 539829
rect 48187 539593 48229 539829
rect 47909 539509 48229 539593
rect 47909 539273 47951 539509
rect 48187 539273 48229 539509
rect 47909 539241 48229 539273
rect 53840 539829 54160 539861
rect 53840 539593 53882 539829
rect 54118 539593 54160 539829
rect 53840 539509 54160 539593
rect 53840 539273 53882 539509
rect 54118 539273 54160 539509
rect 53840 539241 54160 539273
rect 59770 539829 60090 539861
rect 59770 539593 59812 539829
rect 60048 539593 60090 539829
rect 59770 539509 60090 539593
rect 59770 539273 59812 539509
rect 60048 539273 60090 539509
rect 59770 539241 60090 539273
rect 75909 539829 76229 539861
rect 75909 539593 75951 539829
rect 76187 539593 76229 539829
rect 75909 539509 76229 539593
rect 75909 539273 75951 539509
rect 76187 539273 76229 539509
rect 75909 539241 76229 539273
rect 81840 539829 82160 539861
rect 81840 539593 81882 539829
rect 82118 539593 82160 539829
rect 81840 539509 82160 539593
rect 81840 539273 81882 539509
rect 82118 539273 82160 539509
rect 81840 539241 82160 539273
rect 87770 539829 88090 539861
rect 87770 539593 87812 539829
rect 88048 539593 88090 539829
rect 87770 539509 88090 539593
rect 87770 539273 87812 539509
rect 88048 539273 88090 539509
rect 87770 539241 88090 539273
rect 103909 539829 104229 539861
rect 103909 539593 103951 539829
rect 104187 539593 104229 539829
rect 103909 539509 104229 539593
rect 103909 539273 103951 539509
rect 104187 539273 104229 539509
rect 103909 539241 104229 539273
rect 109840 539829 110160 539861
rect 109840 539593 109882 539829
rect 110118 539593 110160 539829
rect 109840 539509 110160 539593
rect 109840 539273 109882 539509
rect 110118 539273 110160 539509
rect 109840 539241 110160 539273
rect 115770 539829 116090 539861
rect 115770 539593 115812 539829
rect 116048 539593 116090 539829
rect 115770 539509 116090 539593
rect 115770 539273 115812 539509
rect 116048 539273 116090 539509
rect 115770 539241 116090 539273
rect 131909 539829 132229 539861
rect 131909 539593 131951 539829
rect 132187 539593 132229 539829
rect 131909 539509 132229 539593
rect 131909 539273 131951 539509
rect 132187 539273 132229 539509
rect 131909 539241 132229 539273
rect 137840 539829 138160 539861
rect 137840 539593 137882 539829
rect 138118 539593 138160 539829
rect 137840 539509 138160 539593
rect 137840 539273 137882 539509
rect 138118 539273 138160 539509
rect 137840 539241 138160 539273
rect 143770 539829 144090 539861
rect 143770 539593 143812 539829
rect 144048 539593 144090 539829
rect 143770 539509 144090 539593
rect 143770 539273 143812 539509
rect 144048 539273 144090 539509
rect 143770 539241 144090 539273
rect 159909 539829 160229 539861
rect 159909 539593 159951 539829
rect 160187 539593 160229 539829
rect 159909 539509 160229 539593
rect 159909 539273 159951 539509
rect 160187 539273 160229 539509
rect 159909 539241 160229 539273
rect 165840 539829 166160 539861
rect 165840 539593 165882 539829
rect 166118 539593 166160 539829
rect 165840 539509 166160 539593
rect 165840 539273 165882 539509
rect 166118 539273 166160 539509
rect 165840 539241 166160 539273
rect 171770 539829 172090 539861
rect 171770 539593 171812 539829
rect 172048 539593 172090 539829
rect 171770 539509 172090 539593
rect 171770 539273 171812 539509
rect 172048 539273 172090 539509
rect 171770 539241 172090 539273
rect 187909 539829 188229 539861
rect 187909 539593 187951 539829
rect 188187 539593 188229 539829
rect 187909 539509 188229 539593
rect 187909 539273 187951 539509
rect 188187 539273 188229 539509
rect 187909 539241 188229 539273
rect 193840 539829 194160 539861
rect 193840 539593 193882 539829
rect 194118 539593 194160 539829
rect 193840 539509 194160 539593
rect 193840 539273 193882 539509
rect 194118 539273 194160 539509
rect 193840 539241 194160 539273
rect 199770 539829 200090 539861
rect 199770 539593 199812 539829
rect 200048 539593 200090 539829
rect 199770 539509 200090 539593
rect 199770 539273 199812 539509
rect 200048 539273 200090 539509
rect 199770 539241 200090 539273
rect 215909 539829 216229 539861
rect 215909 539593 215951 539829
rect 216187 539593 216229 539829
rect 215909 539509 216229 539593
rect 215909 539273 215951 539509
rect 216187 539273 216229 539509
rect 215909 539241 216229 539273
rect 221840 539829 222160 539861
rect 221840 539593 221882 539829
rect 222118 539593 222160 539829
rect 221840 539509 222160 539593
rect 221840 539273 221882 539509
rect 222118 539273 222160 539509
rect 221840 539241 222160 539273
rect 227770 539829 228090 539861
rect 227770 539593 227812 539829
rect 228048 539593 228090 539829
rect 227770 539509 228090 539593
rect 227770 539273 227812 539509
rect 228048 539273 228090 539509
rect 227770 539241 228090 539273
rect 243909 539829 244229 539861
rect 243909 539593 243951 539829
rect 244187 539593 244229 539829
rect 243909 539509 244229 539593
rect 243909 539273 243951 539509
rect 244187 539273 244229 539509
rect 243909 539241 244229 539273
rect 249840 539829 250160 539861
rect 249840 539593 249882 539829
rect 250118 539593 250160 539829
rect 249840 539509 250160 539593
rect 249840 539273 249882 539509
rect 250118 539273 250160 539509
rect 249840 539241 250160 539273
rect 255770 539829 256090 539861
rect 255770 539593 255812 539829
rect 256048 539593 256090 539829
rect 255770 539509 256090 539593
rect 255770 539273 255812 539509
rect 256048 539273 256090 539509
rect 255770 539241 256090 539273
rect 271909 539829 272229 539861
rect 271909 539593 271951 539829
rect 272187 539593 272229 539829
rect 271909 539509 272229 539593
rect 271909 539273 271951 539509
rect 272187 539273 272229 539509
rect 271909 539241 272229 539273
rect 277840 539829 278160 539861
rect 277840 539593 277882 539829
rect 278118 539593 278160 539829
rect 277840 539509 278160 539593
rect 277840 539273 277882 539509
rect 278118 539273 278160 539509
rect 277840 539241 278160 539273
rect 283770 539829 284090 539861
rect 283770 539593 283812 539829
rect 284048 539593 284090 539829
rect 283770 539509 284090 539593
rect 283770 539273 283812 539509
rect 284048 539273 284090 539509
rect 283770 539241 284090 539273
rect 299909 539829 300229 539861
rect 299909 539593 299951 539829
rect 300187 539593 300229 539829
rect 299909 539509 300229 539593
rect 299909 539273 299951 539509
rect 300187 539273 300229 539509
rect 299909 539241 300229 539273
rect 305840 539829 306160 539861
rect 305840 539593 305882 539829
rect 306118 539593 306160 539829
rect 305840 539509 306160 539593
rect 305840 539273 305882 539509
rect 306118 539273 306160 539509
rect 305840 539241 306160 539273
rect 311770 539829 312090 539861
rect 311770 539593 311812 539829
rect 312048 539593 312090 539829
rect 311770 539509 312090 539593
rect 311770 539273 311812 539509
rect 312048 539273 312090 539509
rect 311770 539241 312090 539273
rect 327909 539829 328229 539861
rect 327909 539593 327951 539829
rect 328187 539593 328229 539829
rect 327909 539509 328229 539593
rect 327909 539273 327951 539509
rect 328187 539273 328229 539509
rect 327909 539241 328229 539273
rect 333840 539829 334160 539861
rect 333840 539593 333882 539829
rect 334118 539593 334160 539829
rect 333840 539509 334160 539593
rect 333840 539273 333882 539509
rect 334118 539273 334160 539509
rect 333840 539241 334160 539273
rect 339770 539829 340090 539861
rect 339770 539593 339812 539829
rect 340048 539593 340090 539829
rect 339770 539509 340090 539593
rect 339770 539273 339812 539509
rect 340048 539273 340090 539509
rect 339770 539241 340090 539273
rect 355909 539829 356229 539861
rect 355909 539593 355951 539829
rect 356187 539593 356229 539829
rect 355909 539509 356229 539593
rect 355909 539273 355951 539509
rect 356187 539273 356229 539509
rect 355909 539241 356229 539273
rect 361840 539829 362160 539861
rect 361840 539593 361882 539829
rect 362118 539593 362160 539829
rect 361840 539509 362160 539593
rect 361840 539273 361882 539509
rect 362118 539273 362160 539509
rect 361840 539241 362160 539273
rect 367770 539829 368090 539861
rect 367770 539593 367812 539829
rect 368048 539593 368090 539829
rect 367770 539509 368090 539593
rect 367770 539273 367812 539509
rect 368048 539273 368090 539509
rect 367770 539241 368090 539273
rect 383909 539829 384229 539861
rect 383909 539593 383951 539829
rect 384187 539593 384229 539829
rect 383909 539509 384229 539593
rect 383909 539273 383951 539509
rect 384187 539273 384229 539509
rect 383909 539241 384229 539273
rect 389840 539829 390160 539861
rect 389840 539593 389882 539829
rect 390118 539593 390160 539829
rect 389840 539509 390160 539593
rect 389840 539273 389882 539509
rect 390118 539273 390160 539509
rect 389840 539241 390160 539273
rect 395770 539829 396090 539861
rect 395770 539593 395812 539829
rect 396048 539593 396090 539829
rect 395770 539509 396090 539593
rect 395770 539273 395812 539509
rect 396048 539273 396090 539509
rect 395770 539241 396090 539273
rect 411909 539829 412229 539861
rect 411909 539593 411951 539829
rect 412187 539593 412229 539829
rect 411909 539509 412229 539593
rect 411909 539273 411951 539509
rect 412187 539273 412229 539509
rect 411909 539241 412229 539273
rect 417840 539829 418160 539861
rect 417840 539593 417882 539829
rect 418118 539593 418160 539829
rect 417840 539509 418160 539593
rect 417840 539273 417882 539509
rect 418118 539273 418160 539509
rect 417840 539241 418160 539273
rect 423770 539829 424090 539861
rect 423770 539593 423812 539829
rect 424048 539593 424090 539829
rect 423770 539509 424090 539593
rect 423770 539273 423812 539509
rect 424048 539273 424090 539509
rect 423770 539241 424090 539273
rect 439909 539829 440229 539861
rect 439909 539593 439951 539829
rect 440187 539593 440229 539829
rect 439909 539509 440229 539593
rect 439909 539273 439951 539509
rect 440187 539273 440229 539509
rect 439909 539241 440229 539273
rect 445840 539829 446160 539861
rect 445840 539593 445882 539829
rect 446118 539593 446160 539829
rect 445840 539509 446160 539593
rect 445840 539273 445882 539509
rect 446118 539273 446160 539509
rect 445840 539241 446160 539273
rect 451770 539829 452090 539861
rect 451770 539593 451812 539829
rect 452048 539593 452090 539829
rect 451770 539509 452090 539593
rect 451770 539273 451812 539509
rect 452048 539273 452090 539509
rect 451770 539241 452090 539273
rect 467909 539829 468229 539861
rect 467909 539593 467951 539829
rect 468187 539593 468229 539829
rect 467909 539509 468229 539593
rect 467909 539273 467951 539509
rect 468187 539273 468229 539509
rect 467909 539241 468229 539273
rect 473840 539829 474160 539861
rect 473840 539593 473882 539829
rect 474118 539593 474160 539829
rect 473840 539509 474160 539593
rect 473840 539273 473882 539509
rect 474118 539273 474160 539509
rect 473840 539241 474160 539273
rect 479770 539829 480090 539861
rect 479770 539593 479812 539829
rect 480048 539593 480090 539829
rect 479770 539509 480090 539593
rect 479770 539273 479812 539509
rect 480048 539273 480090 539509
rect 479770 539241 480090 539273
rect 495909 539829 496229 539861
rect 495909 539593 495951 539829
rect 496187 539593 496229 539829
rect 495909 539509 496229 539593
rect 495909 539273 495951 539509
rect 496187 539273 496229 539509
rect 495909 539241 496229 539273
rect 501840 539829 502160 539861
rect 501840 539593 501882 539829
rect 502118 539593 502160 539829
rect 501840 539509 502160 539593
rect 501840 539273 501882 539509
rect 502118 539273 502160 539509
rect 501840 539241 502160 539273
rect 507770 539829 508090 539861
rect 507770 539593 507812 539829
rect 508048 539593 508090 539829
rect 507770 539509 508090 539593
rect 507770 539273 507812 539509
rect 508048 539273 508090 539509
rect 507770 539241 508090 539273
rect 523909 539829 524229 539861
rect 523909 539593 523951 539829
rect 524187 539593 524229 539829
rect 523909 539509 524229 539593
rect 523909 539273 523951 539509
rect 524187 539273 524229 539509
rect 523909 539241 524229 539273
rect 529840 539829 530160 539861
rect 529840 539593 529882 539829
rect 530118 539593 530160 539829
rect 529840 539509 530160 539593
rect 529840 539273 529882 539509
rect 530118 539273 530160 539509
rect 529840 539241 530160 539273
rect 535770 539829 536090 539861
rect 535770 539593 535812 539829
rect 536048 539593 536090 539829
rect 535770 539509 536090 539593
rect 535770 539273 535812 539509
rect 536048 539273 536090 539509
rect 535770 539241 536090 539273
rect 551909 539829 552229 539861
rect 551909 539593 551951 539829
rect 552187 539593 552229 539829
rect 551909 539509 552229 539593
rect 551909 539273 551951 539509
rect 552187 539273 552229 539509
rect 551909 539241 552229 539273
rect 557840 539829 558160 539861
rect 557840 539593 557882 539829
rect 558118 539593 558160 539829
rect 557840 539509 558160 539593
rect 557840 539273 557882 539509
rect 558118 539273 558160 539509
rect 557840 539241 558160 539273
rect 563770 539829 564090 539861
rect 563770 539593 563812 539829
rect 564048 539593 564090 539829
rect 563770 539509 564090 539593
rect 563770 539273 563812 539509
rect 564048 539273 564090 539509
rect 563770 539241 564090 539273
rect 573494 539829 574114 566273
rect 573494 539593 573526 539829
rect 573762 539593 573846 539829
rect 574082 539593 574114 539829
rect 573494 539509 574114 539593
rect 573494 539273 573526 539509
rect 573762 539273 573846 539509
rect 574082 539273 574114 539509
rect 22875 536454 23195 536486
rect 22875 536218 22917 536454
rect 23153 536218 23195 536454
rect 22875 536134 23195 536218
rect 22875 535898 22917 536134
rect 23153 535898 23195 536134
rect 22875 535866 23195 535898
rect 28806 536454 29126 536486
rect 28806 536218 28848 536454
rect 29084 536218 29126 536454
rect 28806 536134 29126 536218
rect 28806 535898 28848 536134
rect 29084 535898 29126 536134
rect 28806 535866 29126 535898
rect 50875 536454 51195 536486
rect 50875 536218 50917 536454
rect 51153 536218 51195 536454
rect 50875 536134 51195 536218
rect 50875 535898 50917 536134
rect 51153 535898 51195 536134
rect 50875 535866 51195 535898
rect 56806 536454 57126 536486
rect 56806 536218 56848 536454
rect 57084 536218 57126 536454
rect 56806 536134 57126 536218
rect 56806 535898 56848 536134
rect 57084 535898 57126 536134
rect 56806 535866 57126 535898
rect 78875 536454 79195 536486
rect 78875 536218 78917 536454
rect 79153 536218 79195 536454
rect 78875 536134 79195 536218
rect 78875 535898 78917 536134
rect 79153 535898 79195 536134
rect 78875 535866 79195 535898
rect 84806 536454 85126 536486
rect 84806 536218 84848 536454
rect 85084 536218 85126 536454
rect 84806 536134 85126 536218
rect 84806 535898 84848 536134
rect 85084 535898 85126 536134
rect 84806 535866 85126 535898
rect 106875 536454 107195 536486
rect 106875 536218 106917 536454
rect 107153 536218 107195 536454
rect 106875 536134 107195 536218
rect 106875 535898 106917 536134
rect 107153 535898 107195 536134
rect 106875 535866 107195 535898
rect 112806 536454 113126 536486
rect 112806 536218 112848 536454
rect 113084 536218 113126 536454
rect 112806 536134 113126 536218
rect 112806 535898 112848 536134
rect 113084 535898 113126 536134
rect 112806 535866 113126 535898
rect 134875 536454 135195 536486
rect 134875 536218 134917 536454
rect 135153 536218 135195 536454
rect 134875 536134 135195 536218
rect 134875 535898 134917 536134
rect 135153 535898 135195 536134
rect 134875 535866 135195 535898
rect 140806 536454 141126 536486
rect 140806 536218 140848 536454
rect 141084 536218 141126 536454
rect 140806 536134 141126 536218
rect 140806 535898 140848 536134
rect 141084 535898 141126 536134
rect 140806 535866 141126 535898
rect 162875 536454 163195 536486
rect 162875 536218 162917 536454
rect 163153 536218 163195 536454
rect 162875 536134 163195 536218
rect 162875 535898 162917 536134
rect 163153 535898 163195 536134
rect 162875 535866 163195 535898
rect 168806 536454 169126 536486
rect 168806 536218 168848 536454
rect 169084 536218 169126 536454
rect 168806 536134 169126 536218
rect 168806 535898 168848 536134
rect 169084 535898 169126 536134
rect 168806 535866 169126 535898
rect 190875 536454 191195 536486
rect 190875 536218 190917 536454
rect 191153 536218 191195 536454
rect 190875 536134 191195 536218
rect 190875 535898 190917 536134
rect 191153 535898 191195 536134
rect 190875 535866 191195 535898
rect 196806 536454 197126 536486
rect 196806 536218 196848 536454
rect 197084 536218 197126 536454
rect 196806 536134 197126 536218
rect 196806 535898 196848 536134
rect 197084 535898 197126 536134
rect 196806 535866 197126 535898
rect 218875 536454 219195 536486
rect 218875 536218 218917 536454
rect 219153 536218 219195 536454
rect 218875 536134 219195 536218
rect 218875 535898 218917 536134
rect 219153 535898 219195 536134
rect 218875 535866 219195 535898
rect 224806 536454 225126 536486
rect 224806 536218 224848 536454
rect 225084 536218 225126 536454
rect 224806 536134 225126 536218
rect 224806 535898 224848 536134
rect 225084 535898 225126 536134
rect 224806 535866 225126 535898
rect 246875 536454 247195 536486
rect 246875 536218 246917 536454
rect 247153 536218 247195 536454
rect 246875 536134 247195 536218
rect 246875 535898 246917 536134
rect 247153 535898 247195 536134
rect 246875 535866 247195 535898
rect 252806 536454 253126 536486
rect 252806 536218 252848 536454
rect 253084 536218 253126 536454
rect 252806 536134 253126 536218
rect 252806 535898 252848 536134
rect 253084 535898 253126 536134
rect 252806 535866 253126 535898
rect 274875 536454 275195 536486
rect 274875 536218 274917 536454
rect 275153 536218 275195 536454
rect 274875 536134 275195 536218
rect 274875 535898 274917 536134
rect 275153 535898 275195 536134
rect 274875 535866 275195 535898
rect 280806 536454 281126 536486
rect 280806 536218 280848 536454
rect 281084 536218 281126 536454
rect 280806 536134 281126 536218
rect 280806 535898 280848 536134
rect 281084 535898 281126 536134
rect 280806 535866 281126 535898
rect 302875 536454 303195 536486
rect 302875 536218 302917 536454
rect 303153 536218 303195 536454
rect 302875 536134 303195 536218
rect 302875 535898 302917 536134
rect 303153 535898 303195 536134
rect 302875 535866 303195 535898
rect 308806 536454 309126 536486
rect 308806 536218 308848 536454
rect 309084 536218 309126 536454
rect 308806 536134 309126 536218
rect 308806 535898 308848 536134
rect 309084 535898 309126 536134
rect 308806 535866 309126 535898
rect 330875 536454 331195 536486
rect 330875 536218 330917 536454
rect 331153 536218 331195 536454
rect 330875 536134 331195 536218
rect 330875 535898 330917 536134
rect 331153 535898 331195 536134
rect 330875 535866 331195 535898
rect 336806 536454 337126 536486
rect 336806 536218 336848 536454
rect 337084 536218 337126 536454
rect 336806 536134 337126 536218
rect 336806 535898 336848 536134
rect 337084 535898 337126 536134
rect 336806 535866 337126 535898
rect 358875 536454 359195 536486
rect 358875 536218 358917 536454
rect 359153 536218 359195 536454
rect 358875 536134 359195 536218
rect 358875 535898 358917 536134
rect 359153 535898 359195 536134
rect 358875 535866 359195 535898
rect 364806 536454 365126 536486
rect 364806 536218 364848 536454
rect 365084 536218 365126 536454
rect 364806 536134 365126 536218
rect 364806 535898 364848 536134
rect 365084 535898 365126 536134
rect 364806 535866 365126 535898
rect 386875 536454 387195 536486
rect 386875 536218 386917 536454
rect 387153 536218 387195 536454
rect 386875 536134 387195 536218
rect 386875 535898 386917 536134
rect 387153 535898 387195 536134
rect 386875 535866 387195 535898
rect 392806 536454 393126 536486
rect 392806 536218 392848 536454
rect 393084 536218 393126 536454
rect 392806 536134 393126 536218
rect 392806 535898 392848 536134
rect 393084 535898 393126 536134
rect 392806 535866 393126 535898
rect 414875 536454 415195 536486
rect 414875 536218 414917 536454
rect 415153 536218 415195 536454
rect 414875 536134 415195 536218
rect 414875 535898 414917 536134
rect 415153 535898 415195 536134
rect 414875 535866 415195 535898
rect 420806 536454 421126 536486
rect 420806 536218 420848 536454
rect 421084 536218 421126 536454
rect 420806 536134 421126 536218
rect 420806 535898 420848 536134
rect 421084 535898 421126 536134
rect 420806 535866 421126 535898
rect 442875 536454 443195 536486
rect 442875 536218 442917 536454
rect 443153 536218 443195 536454
rect 442875 536134 443195 536218
rect 442875 535898 442917 536134
rect 443153 535898 443195 536134
rect 442875 535866 443195 535898
rect 448806 536454 449126 536486
rect 448806 536218 448848 536454
rect 449084 536218 449126 536454
rect 448806 536134 449126 536218
rect 448806 535898 448848 536134
rect 449084 535898 449126 536134
rect 448806 535866 449126 535898
rect 470875 536454 471195 536486
rect 470875 536218 470917 536454
rect 471153 536218 471195 536454
rect 470875 536134 471195 536218
rect 470875 535898 470917 536134
rect 471153 535898 471195 536134
rect 470875 535866 471195 535898
rect 476806 536454 477126 536486
rect 476806 536218 476848 536454
rect 477084 536218 477126 536454
rect 476806 536134 477126 536218
rect 476806 535898 476848 536134
rect 477084 535898 477126 536134
rect 476806 535866 477126 535898
rect 498875 536454 499195 536486
rect 498875 536218 498917 536454
rect 499153 536218 499195 536454
rect 498875 536134 499195 536218
rect 498875 535898 498917 536134
rect 499153 535898 499195 536134
rect 498875 535866 499195 535898
rect 504806 536454 505126 536486
rect 504806 536218 504848 536454
rect 505084 536218 505126 536454
rect 504806 536134 505126 536218
rect 504806 535898 504848 536134
rect 505084 535898 505126 536134
rect 504806 535866 505126 535898
rect 526875 536454 527195 536486
rect 526875 536218 526917 536454
rect 527153 536218 527195 536454
rect 526875 536134 527195 536218
rect 526875 535898 526917 536134
rect 527153 535898 527195 536134
rect 526875 535866 527195 535898
rect 532806 536454 533126 536486
rect 532806 536218 532848 536454
rect 533084 536218 533126 536454
rect 532806 536134 533126 536218
rect 532806 535898 532848 536134
rect 533084 535898 533126 536134
rect 532806 535866 533126 535898
rect 554875 536454 555195 536486
rect 554875 536218 554917 536454
rect 555153 536218 555195 536454
rect 554875 536134 555195 536218
rect 554875 535898 554917 536134
rect 555153 535898 555195 536134
rect 554875 535866 555195 535898
rect 560806 536454 561126 536486
rect 560806 536218 560848 536454
rect 561084 536218 561126 536454
rect 560806 536134 561126 536218
rect 560806 535898 560848 536134
rect 561084 535898 561126 536134
rect 560806 535866 561126 535898
rect -2006 512593 -1974 512829
rect -1738 512593 -1654 512829
rect -1418 512593 -1386 512829
rect -2006 512509 -1386 512593
rect -2006 512273 -1974 512509
rect -1738 512273 -1654 512509
rect -1418 512273 -1386 512509
rect -2006 485829 -1386 512273
rect 19910 512829 20230 512861
rect 19910 512593 19952 512829
rect 20188 512593 20230 512829
rect 19910 512509 20230 512593
rect 19910 512273 19952 512509
rect 20188 512273 20230 512509
rect 19910 512241 20230 512273
rect 25840 512829 26160 512861
rect 25840 512593 25882 512829
rect 26118 512593 26160 512829
rect 25840 512509 26160 512593
rect 25840 512273 25882 512509
rect 26118 512273 26160 512509
rect 25840 512241 26160 512273
rect 31771 512829 32091 512861
rect 31771 512593 31813 512829
rect 32049 512593 32091 512829
rect 31771 512509 32091 512593
rect 31771 512273 31813 512509
rect 32049 512273 32091 512509
rect 31771 512241 32091 512273
rect 47910 512829 48230 512861
rect 47910 512593 47952 512829
rect 48188 512593 48230 512829
rect 47910 512509 48230 512593
rect 47910 512273 47952 512509
rect 48188 512273 48230 512509
rect 47910 512241 48230 512273
rect 53840 512829 54160 512861
rect 53840 512593 53882 512829
rect 54118 512593 54160 512829
rect 53840 512509 54160 512593
rect 53840 512273 53882 512509
rect 54118 512273 54160 512509
rect 53840 512241 54160 512273
rect 59771 512829 60091 512861
rect 59771 512593 59813 512829
rect 60049 512593 60091 512829
rect 59771 512509 60091 512593
rect 59771 512273 59813 512509
rect 60049 512273 60091 512509
rect 59771 512241 60091 512273
rect 75910 512829 76230 512861
rect 75910 512593 75952 512829
rect 76188 512593 76230 512829
rect 75910 512509 76230 512593
rect 75910 512273 75952 512509
rect 76188 512273 76230 512509
rect 75910 512241 76230 512273
rect 81840 512829 82160 512861
rect 81840 512593 81882 512829
rect 82118 512593 82160 512829
rect 81840 512509 82160 512593
rect 81840 512273 81882 512509
rect 82118 512273 82160 512509
rect 81840 512241 82160 512273
rect 87771 512829 88091 512861
rect 87771 512593 87813 512829
rect 88049 512593 88091 512829
rect 87771 512509 88091 512593
rect 87771 512273 87813 512509
rect 88049 512273 88091 512509
rect 87771 512241 88091 512273
rect 103910 512829 104230 512861
rect 103910 512593 103952 512829
rect 104188 512593 104230 512829
rect 103910 512509 104230 512593
rect 103910 512273 103952 512509
rect 104188 512273 104230 512509
rect 103910 512241 104230 512273
rect 109840 512829 110160 512861
rect 109840 512593 109882 512829
rect 110118 512593 110160 512829
rect 109840 512509 110160 512593
rect 109840 512273 109882 512509
rect 110118 512273 110160 512509
rect 109840 512241 110160 512273
rect 115771 512829 116091 512861
rect 115771 512593 115813 512829
rect 116049 512593 116091 512829
rect 115771 512509 116091 512593
rect 115771 512273 115813 512509
rect 116049 512273 116091 512509
rect 115771 512241 116091 512273
rect 131910 512829 132230 512861
rect 131910 512593 131952 512829
rect 132188 512593 132230 512829
rect 131910 512509 132230 512593
rect 131910 512273 131952 512509
rect 132188 512273 132230 512509
rect 131910 512241 132230 512273
rect 137840 512829 138160 512861
rect 137840 512593 137882 512829
rect 138118 512593 138160 512829
rect 137840 512509 138160 512593
rect 137840 512273 137882 512509
rect 138118 512273 138160 512509
rect 137840 512241 138160 512273
rect 143771 512829 144091 512861
rect 143771 512593 143813 512829
rect 144049 512593 144091 512829
rect 143771 512509 144091 512593
rect 143771 512273 143813 512509
rect 144049 512273 144091 512509
rect 143771 512241 144091 512273
rect 159910 512829 160230 512861
rect 159910 512593 159952 512829
rect 160188 512593 160230 512829
rect 159910 512509 160230 512593
rect 159910 512273 159952 512509
rect 160188 512273 160230 512509
rect 159910 512241 160230 512273
rect 165840 512829 166160 512861
rect 165840 512593 165882 512829
rect 166118 512593 166160 512829
rect 165840 512509 166160 512593
rect 165840 512273 165882 512509
rect 166118 512273 166160 512509
rect 165840 512241 166160 512273
rect 171771 512829 172091 512861
rect 171771 512593 171813 512829
rect 172049 512593 172091 512829
rect 171771 512509 172091 512593
rect 171771 512273 171813 512509
rect 172049 512273 172091 512509
rect 171771 512241 172091 512273
rect 187910 512829 188230 512861
rect 187910 512593 187952 512829
rect 188188 512593 188230 512829
rect 187910 512509 188230 512593
rect 187910 512273 187952 512509
rect 188188 512273 188230 512509
rect 187910 512241 188230 512273
rect 193840 512829 194160 512861
rect 193840 512593 193882 512829
rect 194118 512593 194160 512829
rect 193840 512509 194160 512593
rect 193840 512273 193882 512509
rect 194118 512273 194160 512509
rect 193840 512241 194160 512273
rect 199771 512829 200091 512861
rect 199771 512593 199813 512829
rect 200049 512593 200091 512829
rect 199771 512509 200091 512593
rect 199771 512273 199813 512509
rect 200049 512273 200091 512509
rect 199771 512241 200091 512273
rect 215910 512829 216230 512861
rect 215910 512593 215952 512829
rect 216188 512593 216230 512829
rect 215910 512509 216230 512593
rect 215910 512273 215952 512509
rect 216188 512273 216230 512509
rect 215910 512241 216230 512273
rect 221840 512829 222160 512861
rect 221840 512593 221882 512829
rect 222118 512593 222160 512829
rect 221840 512509 222160 512593
rect 221840 512273 221882 512509
rect 222118 512273 222160 512509
rect 221840 512241 222160 512273
rect 227771 512829 228091 512861
rect 227771 512593 227813 512829
rect 228049 512593 228091 512829
rect 227771 512509 228091 512593
rect 227771 512273 227813 512509
rect 228049 512273 228091 512509
rect 227771 512241 228091 512273
rect 243910 512829 244230 512861
rect 243910 512593 243952 512829
rect 244188 512593 244230 512829
rect 243910 512509 244230 512593
rect 243910 512273 243952 512509
rect 244188 512273 244230 512509
rect 243910 512241 244230 512273
rect 249840 512829 250160 512861
rect 249840 512593 249882 512829
rect 250118 512593 250160 512829
rect 249840 512509 250160 512593
rect 249840 512273 249882 512509
rect 250118 512273 250160 512509
rect 249840 512241 250160 512273
rect 255771 512829 256091 512861
rect 255771 512593 255813 512829
rect 256049 512593 256091 512829
rect 255771 512509 256091 512593
rect 255771 512273 255813 512509
rect 256049 512273 256091 512509
rect 255771 512241 256091 512273
rect 271910 512829 272230 512861
rect 271910 512593 271952 512829
rect 272188 512593 272230 512829
rect 271910 512509 272230 512593
rect 271910 512273 271952 512509
rect 272188 512273 272230 512509
rect 271910 512241 272230 512273
rect 277840 512829 278160 512861
rect 277840 512593 277882 512829
rect 278118 512593 278160 512829
rect 277840 512509 278160 512593
rect 277840 512273 277882 512509
rect 278118 512273 278160 512509
rect 277840 512241 278160 512273
rect 283771 512829 284091 512861
rect 283771 512593 283813 512829
rect 284049 512593 284091 512829
rect 283771 512509 284091 512593
rect 283771 512273 283813 512509
rect 284049 512273 284091 512509
rect 283771 512241 284091 512273
rect 299910 512829 300230 512861
rect 299910 512593 299952 512829
rect 300188 512593 300230 512829
rect 299910 512509 300230 512593
rect 299910 512273 299952 512509
rect 300188 512273 300230 512509
rect 299910 512241 300230 512273
rect 305840 512829 306160 512861
rect 305840 512593 305882 512829
rect 306118 512593 306160 512829
rect 305840 512509 306160 512593
rect 305840 512273 305882 512509
rect 306118 512273 306160 512509
rect 305840 512241 306160 512273
rect 311771 512829 312091 512861
rect 311771 512593 311813 512829
rect 312049 512593 312091 512829
rect 311771 512509 312091 512593
rect 311771 512273 311813 512509
rect 312049 512273 312091 512509
rect 311771 512241 312091 512273
rect 327910 512829 328230 512861
rect 327910 512593 327952 512829
rect 328188 512593 328230 512829
rect 327910 512509 328230 512593
rect 327910 512273 327952 512509
rect 328188 512273 328230 512509
rect 327910 512241 328230 512273
rect 333840 512829 334160 512861
rect 333840 512593 333882 512829
rect 334118 512593 334160 512829
rect 333840 512509 334160 512593
rect 333840 512273 333882 512509
rect 334118 512273 334160 512509
rect 333840 512241 334160 512273
rect 339771 512829 340091 512861
rect 339771 512593 339813 512829
rect 340049 512593 340091 512829
rect 339771 512509 340091 512593
rect 339771 512273 339813 512509
rect 340049 512273 340091 512509
rect 339771 512241 340091 512273
rect 355910 512829 356230 512861
rect 355910 512593 355952 512829
rect 356188 512593 356230 512829
rect 355910 512509 356230 512593
rect 355910 512273 355952 512509
rect 356188 512273 356230 512509
rect 355910 512241 356230 512273
rect 361840 512829 362160 512861
rect 361840 512593 361882 512829
rect 362118 512593 362160 512829
rect 361840 512509 362160 512593
rect 361840 512273 361882 512509
rect 362118 512273 362160 512509
rect 361840 512241 362160 512273
rect 367771 512829 368091 512861
rect 367771 512593 367813 512829
rect 368049 512593 368091 512829
rect 367771 512509 368091 512593
rect 367771 512273 367813 512509
rect 368049 512273 368091 512509
rect 367771 512241 368091 512273
rect 383910 512829 384230 512861
rect 383910 512593 383952 512829
rect 384188 512593 384230 512829
rect 383910 512509 384230 512593
rect 383910 512273 383952 512509
rect 384188 512273 384230 512509
rect 383910 512241 384230 512273
rect 389840 512829 390160 512861
rect 389840 512593 389882 512829
rect 390118 512593 390160 512829
rect 389840 512509 390160 512593
rect 389840 512273 389882 512509
rect 390118 512273 390160 512509
rect 389840 512241 390160 512273
rect 395771 512829 396091 512861
rect 395771 512593 395813 512829
rect 396049 512593 396091 512829
rect 395771 512509 396091 512593
rect 395771 512273 395813 512509
rect 396049 512273 396091 512509
rect 395771 512241 396091 512273
rect 411910 512829 412230 512861
rect 411910 512593 411952 512829
rect 412188 512593 412230 512829
rect 411910 512509 412230 512593
rect 411910 512273 411952 512509
rect 412188 512273 412230 512509
rect 411910 512241 412230 512273
rect 417840 512829 418160 512861
rect 417840 512593 417882 512829
rect 418118 512593 418160 512829
rect 417840 512509 418160 512593
rect 417840 512273 417882 512509
rect 418118 512273 418160 512509
rect 417840 512241 418160 512273
rect 423771 512829 424091 512861
rect 423771 512593 423813 512829
rect 424049 512593 424091 512829
rect 423771 512509 424091 512593
rect 423771 512273 423813 512509
rect 424049 512273 424091 512509
rect 423771 512241 424091 512273
rect 439910 512829 440230 512861
rect 439910 512593 439952 512829
rect 440188 512593 440230 512829
rect 439910 512509 440230 512593
rect 439910 512273 439952 512509
rect 440188 512273 440230 512509
rect 439910 512241 440230 512273
rect 445840 512829 446160 512861
rect 445840 512593 445882 512829
rect 446118 512593 446160 512829
rect 445840 512509 446160 512593
rect 445840 512273 445882 512509
rect 446118 512273 446160 512509
rect 445840 512241 446160 512273
rect 451771 512829 452091 512861
rect 451771 512593 451813 512829
rect 452049 512593 452091 512829
rect 451771 512509 452091 512593
rect 451771 512273 451813 512509
rect 452049 512273 452091 512509
rect 451771 512241 452091 512273
rect 467910 512829 468230 512861
rect 467910 512593 467952 512829
rect 468188 512593 468230 512829
rect 467910 512509 468230 512593
rect 467910 512273 467952 512509
rect 468188 512273 468230 512509
rect 467910 512241 468230 512273
rect 473840 512829 474160 512861
rect 473840 512593 473882 512829
rect 474118 512593 474160 512829
rect 473840 512509 474160 512593
rect 473840 512273 473882 512509
rect 474118 512273 474160 512509
rect 473840 512241 474160 512273
rect 479771 512829 480091 512861
rect 479771 512593 479813 512829
rect 480049 512593 480091 512829
rect 479771 512509 480091 512593
rect 479771 512273 479813 512509
rect 480049 512273 480091 512509
rect 479771 512241 480091 512273
rect 495910 512829 496230 512861
rect 495910 512593 495952 512829
rect 496188 512593 496230 512829
rect 495910 512509 496230 512593
rect 495910 512273 495952 512509
rect 496188 512273 496230 512509
rect 495910 512241 496230 512273
rect 501840 512829 502160 512861
rect 501840 512593 501882 512829
rect 502118 512593 502160 512829
rect 501840 512509 502160 512593
rect 501840 512273 501882 512509
rect 502118 512273 502160 512509
rect 501840 512241 502160 512273
rect 507771 512829 508091 512861
rect 507771 512593 507813 512829
rect 508049 512593 508091 512829
rect 507771 512509 508091 512593
rect 507771 512273 507813 512509
rect 508049 512273 508091 512509
rect 507771 512241 508091 512273
rect 523910 512829 524230 512861
rect 523910 512593 523952 512829
rect 524188 512593 524230 512829
rect 523910 512509 524230 512593
rect 523910 512273 523952 512509
rect 524188 512273 524230 512509
rect 523910 512241 524230 512273
rect 529840 512829 530160 512861
rect 529840 512593 529882 512829
rect 530118 512593 530160 512829
rect 529840 512509 530160 512593
rect 529840 512273 529882 512509
rect 530118 512273 530160 512509
rect 529840 512241 530160 512273
rect 535771 512829 536091 512861
rect 535771 512593 535813 512829
rect 536049 512593 536091 512829
rect 535771 512509 536091 512593
rect 535771 512273 535813 512509
rect 536049 512273 536091 512509
rect 535771 512241 536091 512273
rect 551910 512829 552230 512861
rect 551910 512593 551952 512829
rect 552188 512593 552230 512829
rect 551910 512509 552230 512593
rect 551910 512273 551952 512509
rect 552188 512273 552230 512509
rect 551910 512241 552230 512273
rect 557840 512829 558160 512861
rect 557840 512593 557882 512829
rect 558118 512593 558160 512829
rect 557840 512509 558160 512593
rect 557840 512273 557882 512509
rect 558118 512273 558160 512509
rect 557840 512241 558160 512273
rect 563771 512829 564091 512861
rect 563771 512593 563813 512829
rect 564049 512593 564091 512829
rect 563771 512509 564091 512593
rect 563771 512273 563813 512509
rect 564049 512273 564091 512509
rect 563771 512241 564091 512273
rect 573494 512829 574114 539273
rect 573494 512593 573526 512829
rect 573762 512593 573846 512829
rect 574082 512593 574114 512829
rect 573494 512509 574114 512593
rect 573494 512273 573526 512509
rect 573762 512273 573846 512509
rect 574082 512273 574114 512509
rect 22874 509454 23194 509486
rect 22874 509218 22916 509454
rect 23152 509218 23194 509454
rect 22874 509134 23194 509218
rect 22874 508898 22916 509134
rect 23152 508898 23194 509134
rect 22874 508866 23194 508898
rect 28805 509454 29125 509486
rect 28805 509218 28847 509454
rect 29083 509218 29125 509454
rect 28805 509134 29125 509218
rect 28805 508898 28847 509134
rect 29083 508898 29125 509134
rect 28805 508866 29125 508898
rect 50874 509454 51194 509486
rect 50874 509218 50916 509454
rect 51152 509218 51194 509454
rect 50874 509134 51194 509218
rect 50874 508898 50916 509134
rect 51152 508898 51194 509134
rect 50874 508866 51194 508898
rect 56805 509454 57125 509486
rect 56805 509218 56847 509454
rect 57083 509218 57125 509454
rect 56805 509134 57125 509218
rect 56805 508898 56847 509134
rect 57083 508898 57125 509134
rect 56805 508866 57125 508898
rect 78874 509454 79194 509486
rect 78874 509218 78916 509454
rect 79152 509218 79194 509454
rect 78874 509134 79194 509218
rect 78874 508898 78916 509134
rect 79152 508898 79194 509134
rect 78874 508866 79194 508898
rect 84805 509454 85125 509486
rect 84805 509218 84847 509454
rect 85083 509218 85125 509454
rect 84805 509134 85125 509218
rect 84805 508898 84847 509134
rect 85083 508898 85125 509134
rect 84805 508866 85125 508898
rect 106874 509454 107194 509486
rect 106874 509218 106916 509454
rect 107152 509218 107194 509454
rect 106874 509134 107194 509218
rect 106874 508898 106916 509134
rect 107152 508898 107194 509134
rect 106874 508866 107194 508898
rect 112805 509454 113125 509486
rect 112805 509218 112847 509454
rect 113083 509218 113125 509454
rect 112805 509134 113125 509218
rect 112805 508898 112847 509134
rect 113083 508898 113125 509134
rect 112805 508866 113125 508898
rect 134874 509454 135194 509486
rect 134874 509218 134916 509454
rect 135152 509218 135194 509454
rect 134874 509134 135194 509218
rect 134874 508898 134916 509134
rect 135152 508898 135194 509134
rect 134874 508866 135194 508898
rect 140805 509454 141125 509486
rect 140805 509218 140847 509454
rect 141083 509218 141125 509454
rect 140805 509134 141125 509218
rect 140805 508898 140847 509134
rect 141083 508898 141125 509134
rect 140805 508866 141125 508898
rect 162874 509454 163194 509486
rect 162874 509218 162916 509454
rect 163152 509218 163194 509454
rect 162874 509134 163194 509218
rect 162874 508898 162916 509134
rect 163152 508898 163194 509134
rect 162874 508866 163194 508898
rect 168805 509454 169125 509486
rect 168805 509218 168847 509454
rect 169083 509218 169125 509454
rect 168805 509134 169125 509218
rect 168805 508898 168847 509134
rect 169083 508898 169125 509134
rect 168805 508866 169125 508898
rect 190874 509454 191194 509486
rect 190874 509218 190916 509454
rect 191152 509218 191194 509454
rect 190874 509134 191194 509218
rect 190874 508898 190916 509134
rect 191152 508898 191194 509134
rect 190874 508866 191194 508898
rect 196805 509454 197125 509486
rect 196805 509218 196847 509454
rect 197083 509218 197125 509454
rect 196805 509134 197125 509218
rect 196805 508898 196847 509134
rect 197083 508898 197125 509134
rect 196805 508866 197125 508898
rect 218874 509454 219194 509486
rect 218874 509218 218916 509454
rect 219152 509218 219194 509454
rect 218874 509134 219194 509218
rect 218874 508898 218916 509134
rect 219152 508898 219194 509134
rect 218874 508866 219194 508898
rect 224805 509454 225125 509486
rect 224805 509218 224847 509454
rect 225083 509218 225125 509454
rect 224805 509134 225125 509218
rect 224805 508898 224847 509134
rect 225083 508898 225125 509134
rect 224805 508866 225125 508898
rect 246874 509454 247194 509486
rect 246874 509218 246916 509454
rect 247152 509218 247194 509454
rect 246874 509134 247194 509218
rect 246874 508898 246916 509134
rect 247152 508898 247194 509134
rect 246874 508866 247194 508898
rect 252805 509454 253125 509486
rect 252805 509218 252847 509454
rect 253083 509218 253125 509454
rect 252805 509134 253125 509218
rect 252805 508898 252847 509134
rect 253083 508898 253125 509134
rect 252805 508866 253125 508898
rect 274874 509454 275194 509486
rect 274874 509218 274916 509454
rect 275152 509218 275194 509454
rect 274874 509134 275194 509218
rect 274874 508898 274916 509134
rect 275152 508898 275194 509134
rect 274874 508866 275194 508898
rect 280805 509454 281125 509486
rect 280805 509218 280847 509454
rect 281083 509218 281125 509454
rect 280805 509134 281125 509218
rect 280805 508898 280847 509134
rect 281083 508898 281125 509134
rect 280805 508866 281125 508898
rect 302874 509454 303194 509486
rect 302874 509218 302916 509454
rect 303152 509218 303194 509454
rect 302874 509134 303194 509218
rect 302874 508898 302916 509134
rect 303152 508898 303194 509134
rect 302874 508866 303194 508898
rect 308805 509454 309125 509486
rect 308805 509218 308847 509454
rect 309083 509218 309125 509454
rect 308805 509134 309125 509218
rect 308805 508898 308847 509134
rect 309083 508898 309125 509134
rect 308805 508866 309125 508898
rect 330874 509454 331194 509486
rect 330874 509218 330916 509454
rect 331152 509218 331194 509454
rect 330874 509134 331194 509218
rect 330874 508898 330916 509134
rect 331152 508898 331194 509134
rect 330874 508866 331194 508898
rect 336805 509454 337125 509486
rect 336805 509218 336847 509454
rect 337083 509218 337125 509454
rect 336805 509134 337125 509218
rect 336805 508898 336847 509134
rect 337083 508898 337125 509134
rect 336805 508866 337125 508898
rect 358874 509454 359194 509486
rect 358874 509218 358916 509454
rect 359152 509218 359194 509454
rect 358874 509134 359194 509218
rect 358874 508898 358916 509134
rect 359152 508898 359194 509134
rect 358874 508866 359194 508898
rect 364805 509454 365125 509486
rect 364805 509218 364847 509454
rect 365083 509218 365125 509454
rect 364805 509134 365125 509218
rect 364805 508898 364847 509134
rect 365083 508898 365125 509134
rect 364805 508866 365125 508898
rect 386874 509454 387194 509486
rect 386874 509218 386916 509454
rect 387152 509218 387194 509454
rect 386874 509134 387194 509218
rect 386874 508898 386916 509134
rect 387152 508898 387194 509134
rect 386874 508866 387194 508898
rect 392805 509454 393125 509486
rect 392805 509218 392847 509454
rect 393083 509218 393125 509454
rect 392805 509134 393125 509218
rect 392805 508898 392847 509134
rect 393083 508898 393125 509134
rect 392805 508866 393125 508898
rect 414874 509454 415194 509486
rect 414874 509218 414916 509454
rect 415152 509218 415194 509454
rect 414874 509134 415194 509218
rect 414874 508898 414916 509134
rect 415152 508898 415194 509134
rect 414874 508866 415194 508898
rect 420805 509454 421125 509486
rect 420805 509218 420847 509454
rect 421083 509218 421125 509454
rect 420805 509134 421125 509218
rect 420805 508898 420847 509134
rect 421083 508898 421125 509134
rect 420805 508866 421125 508898
rect 442874 509454 443194 509486
rect 442874 509218 442916 509454
rect 443152 509218 443194 509454
rect 442874 509134 443194 509218
rect 442874 508898 442916 509134
rect 443152 508898 443194 509134
rect 442874 508866 443194 508898
rect 448805 509454 449125 509486
rect 448805 509218 448847 509454
rect 449083 509218 449125 509454
rect 448805 509134 449125 509218
rect 448805 508898 448847 509134
rect 449083 508898 449125 509134
rect 448805 508866 449125 508898
rect 470874 509454 471194 509486
rect 470874 509218 470916 509454
rect 471152 509218 471194 509454
rect 470874 509134 471194 509218
rect 470874 508898 470916 509134
rect 471152 508898 471194 509134
rect 470874 508866 471194 508898
rect 476805 509454 477125 509486
rect 476805 509218 476847 509454
rect 477083 509218 477125 509454
rect 476805 509134 477125 509218
rect 476805 508898 476847 509134
rect 477083 508898 477125 509134
rect 476805 508866 477125 508898
rect 498874 509454 499194 509486
rect 498874 509218 498916 509454
rect 499152 509218 499194 509454
rect 498874 509134 499194 509218
rect 498874 508898 498916 509134
rect 499152 508898 499194 509134
rect 498874 508866 499194 508898
rect 504805 509454 505125 509486
rect 504805 509218 504847 509454
rect 505083 509218 505125 509454
rect 504805 509134 505125 509218
rect 504805 508898 504847 509134
rect 505083 508898 505125 509134
rect 504805 508866 505125 508898
rect 526874 509454 527194 509486
rect 526874 509218 526916 509454
rect 527152 509218 527194 509454
rect 526874 509134 527194 509218
rect 526874 508898 526916 509134
rect 527152 508898 527194 509134
rect 526874 508866 527194 508898
rect 532805 509454 533125 509486
rect 532805 509218 532847 509454
rect 533083 509218 533125 509454
rect 532805 509134 533125 509218
rect 532805 508898 532847 509134
rect 533083 508898 533125 509134
rect 532805 508866 533125 508898
rect 554874 509454 555194 509486
rect 554874 509218 554916 509454
rect 555152 509218 555194 509454
rect 554874 509134 555194 509218
rect 554874 508898 554916 509134
rect 555152 508898 555194 509134
rect 554874 508866 555194 508898
rect 560805 509454 561125 509486
rect 560805 509218 560847 509454
rect 561083 509218 561125 509454
rect 560805 509134 561125 509218
rect 560805 508898 560847 509134
rect 561083 508898 561125 509134
rect 560805 508866 561125 508898
rect -2006 485593 -1974 485829
rect -1738 485593 -1654 485829
rect -1418 485593 -1386 485829
rect -2006 485509 -1386 485593
rect -2006 485273 -1974 485509
rect -1738 485273 -1654 485509
rect -1418 485273 -1386 485509
rect -2006 458829 -1386 485273
rect 19909 485829 20229 485861
rect 19909 485593 19951 485829
rect 20187 485593 20229 485829
rect 19909 485509 20229 485593
rect 19909 485273 19951 485509
rect 20187 485273 20229 485509
rect 19909 485241 20229 485273
rect 25840 485829 26160 485861
rect 25840 485593 25882 485829
rect 26118 485593 26160 485829
rect 25840 485509 26160 485593
rect 25840 485273 25882 485509
rect 26118 485273 26160 485509
rect 25840 485241 26160 485273
rect 31770 485829 32090 485861
rect 31770 485593 31812 485829
rect 32048 485593 32090 485829
rect 31770 485509 32090 485593
rect 31770 485273 31812 485509
rect 32048 485273 32090 485509
rect 31770 485241 32090 485273
rect 47909 485829 48229 485861
rect 47909 485593 47951 485829
rect 48187 485593 48229 485829
rect 47909 485509 48229 485593
rect 47909 485273 47951 485509
rect 48187 485273 48229 485509
rect 47909 485241 48229 485273
rect 53840 485829 54160 485861
rect 53840 485593 53882 485829
rect 54118 485593 54160 485829
rect 53840 485509 54160 485593
rect 53840 485273 53882 485509
rect 54118 485273 54160 485509
rect 53840 485241 54160 485273
rect 59770 485829 60090 485861
rect 59770 485593 59812 485829
rect 60048 485593 60090 485829
rect 59770 485509 60090 485593
rect 59770 485273 59812 485509
rect 60048 485273 60090 485509
rect 59770 485241 60090 485273
rect 75909 485829 76229 485861
rect 75909 485593 75951 485829
rect 76187 485593 76229 485829
rect 75909 485509 76229 485593
rect 75909 485273 75951 485509
rect 76187 485273 76229 485509
rect 75909 485241 76229 485273
rect 81840 485829 82160 485861
rect 81840 485593 81882 485829
rect 82118 485593 82160 485829
rect 81840 485509 82160 485593
rect 81840 485273 81882 485509
rect 82118 485273 82160 485509
rect 81840 485241 82160 485273
rect 87770 485829 88090 485861
rect 87770 485593 87812 485829
rect 88048 485593 88090 485829
rect 87770 485509 88090 485593
rect 87770 485273 87812 485509
rect 88048 485273 88090 485509
rect 87770 485241 88090 485273
rect 103909 485829 104229 485861
rect 103909 485593 103951 485829
rect 104187 485593 104229 485829
rect 103909 485509 104229 485593
rect 103909 485273 103951 485509
rect 104187 485273 104229 485509
rect 103909 485241 104229 485273
rect 109840 485829 110160 485861
rect 109840 485593 109882 485829
rect 110118 485593 110160 485829
rect 109840 485509 110160 485593
rect 109840 485273 109882 485509
rect 110118 485273 110160 485509
rect 109840 485241 110160 485273
rect 115770 485829 116090 485861
rect 115770 485593 115812 485829
rect 116048 485593 116090 485829
rect 115770 485509 116090 485593
rect 115770 485273 115812 485509
rect 116048 485273 116090 485509
rect 115770 485241 116090 485273
rect 131909 485829 132229 485861
rect 131909 485593 131951 485829
rect 132187 485593 132229 485829
rect 131909 485509 132229 485593
rect 131909 485273 131951 485509
rect 132187 485273 132229 485509
rect 131909 485241 132229 485273
rect 137840 485829 138160 485861
rect 137840 485593 137882 485829
rect 138118 485593 138160 485829
rect 137840 485509 138160 485593
rect 137840 485273 137882 485509
rect 138118 485273 138160 485509
rect 137840 485241 138160 485273
rect 143770 485829 144090 485861
rect 143770 485593 143812 485829
rect 144048 485593 144090 485829
rect 143770 485509 144090 485593
rect 143770 485273 143812 485509
rect 144048 485273 144090 485509
rect 143770 485241 144090 485273
rect 159909 485829 160229 485861
rect 159909 485593 159951 485829
rect 160187 485593 160229 485829
rect 159909 485509 160229 485593
rect 159909 485273 159951 485509
rect 160187 485273 160229 485509
rect 159909 485241 160229 485273
rect 165840 485829 166160 485861
rect 165840 485593 165882 485829
rect 166118 485593 166160 485829
rect 165840 485509 166160 485593
rect 165840 485273 165882 485509
rect 166118 485273 166160 485509
rect 165840 485241 166160 485273
rect 171770 485829 172090 485861
rect 171770 485593 171812 485829
rect 172048 485593 172090 485829
rect 171770 485509 172090 485593
rect 171770 485273 171812 485509
rect 172048 485273 172090 485509
rect 171770 485241 172090 485273
rect 187909 485829 188229 485861
rect 187909 485593 187951 485829
rect 188187 485593 188229 485829
rect 187909 485509 188229 485593
rect 187909 485273 187951 485509
rect 188187 485273 188229 485509
rect 187909 485241 188229 485273
rect 193840 485829 194160 485861
rect 193840 485593 193882 485829
rect 194118 485593 194160 485829
rect 193840 485509 194160 485593
rect 193840 485273 193882 485509
rect 194118 485273 194160 485509
rect 193840 485241 194160 485273
rect 199770 485829 200090 485861
rect 199770 485593 199812 485829
rect 200048 485593 200090 485829
rect 199770 485509 200090 485593
rect 199770 485273 199812 485509
rect 200048 485273 200090 485509
rect 199770 485241 200090 485273
rect 215909 485829 216229 485861
rect 215909 485593 215951 485829
rect 216187 485593 216229 485829
rect 215909 485509 216229 485593
rect 215909 485273 215951 485509
rect 216187 485273 216229 485509
rect 215909 485241 216229 485273
rect 221840 485829 222160 485861
rect 221840 485593 221882 485829
rect 222118 485593 222160 485829
rect 221840 485509 222160 485593
rect 221840 485273 221882 485509
rect 222118 485273 222160 485509
rect 221840 485241 222160 485273
rect 227770 485829 228090 485861
rect 227770 485593 227812 485829
rect 228048 485593 228090 485829
rect 227770 485509 228090 485593
rect 227770 485273 227812 485509
rect 228048 485273 228090 485509
rect 227770 485241 228090 485273
rect 243909 485829 244229 485861
rect 243909 485593 243951 485829
rect 244187 485593 244229 485829
rect 243909 485509 244229 485593
rect 243909 485273 243951 485509
rect 244187 485273 244229 485509
rect 243909 485241 244229 485273
rect 249840 485829 250160 485861
rect 249840 485593 249882 485829
rect 250118 485593 250160 485829
rect 249840 485509 250160 485593
rect 249840 485273 249882 485509
rect 250118 485273 250160 485509
rect 249840 485241 250160 485273
rect 255770 485829 256090 485861
rect 255770 485593 255812 485829
rect 256048 485593 256090 485829
rect 255770 485509 256090 485593
rect 255770 485273 255812 485509
rect 256048 485273 256090 485509
rect 255770 485241 256090 485273
rect 271909 485829 272229 485861
rect 271909 485593 271951 485829
rect 272187 485593 272229 485829
rect 271909 485509 272229 485593
rect 271909 485273 271951 485509
rect 272187 485273 272229 485509
rect 271909 485241 272229 485273
rect 277840 485829 278160 485861
rect 277840 485593 277882 485829
rect 278118 485593 278160 485829
rect 277840 485509 278160 485593
rect 277840 485273 277882 485509
rect 278118 485273 278160 485509
rect 277840 485241 278160 485273
rect 283770 485829 284090 485861
rect 283770 485593 283812 485829
rect 284048 485593 284090 485829
rect 283770 485509 284090 485593
rect 283770 485273 283812 485509
rect 284048 485273 284090 485509
rect 283770 485241 284090 485273
rect 299909 485829 300229 485861
rect 299909 485593 299951 485829
rect 300187 485593 300229 485829
rect 299909 485509 300229 485593
rect 299909 485273 299951 485509
rect 300187 485273 300229 485509
rect 299909 485241 300229 485273
rect 305840 485829 306160 485861
rect 305840 485593 305882 485829
rect 306118 485593 306160 485829
rect 305840 485509 306160 485593
rect 305840 485273 305882 485509
rect 306118 485273 306160 485509
rect 305840 485241 306160 485273
rect 311770 485829 312090 485861
rect 311770 485593 311812 485829
rect 312048 485593 312090 485829
rect 311770 485509 312090 485593
rect 311770 485273 311812 485509
rect 312048 485273 312090 485509
rect 311770 485241 312090 485273
rect 327909 485829 328229 485861
rect 327909 485593 327951 485829
rect 328187 485593 328229 485829
rect 327909 485509 328229 485593
rect 327909 485273 327951 485509
rect 328187 485273 328229 485509
rect 327909 485241 328229 485273
rect 333840 485829 334160 485861
rect 333840 485593 333882 485829
rect 334118 485593 334160 485829
rect 333840 485509 334160 485593
rect 333840 485273 333882 485509
rect 334118 485273 334160 485509
rect 333840 485241 334160 485273
rect 339770 485829 340090 485861
rect 339770 485593 339812 485829
rect 340048 485593 340090 485829
rect 339770 485509 340090 485593
rect 339770 485273 339812 485509
rect 340048 485273 340090 485509
rect 339770 485241 340090 485273
rect 355909 485829 356229 485861
rect 355909 485593 355951 485829
rect 356187 485593 356229 485829
rect 355909 485509 356229 485593
rect 355909 485273 355951 485509
rect 356187 485273 356229 485509
rect 355909 485241 356229 485273
rect 361840 485829 362160 485861
rect 361840 485593 361882 485829
rect 362118 485593 362160 485829
rect 361840 485509 362160 485593
rect 361840 485273 361882 485509
rect 362118 485273 362160 485509
rect 361840 485241 362160 485273
rect 367770 485829 368090 485861
rect 367770 485593 367812 485829
rect 368048 485593 368090 485829
rect 367770 485509 368090 485593
rect 367770 485273 367812 485509
rect 368048 485273 368090 485509
rect 367770 485241 368090 485273
rect 383909 485829 384229 485861
rect 383909 485593 383951 485829
rect 384187 485593 384229 485829
rect 383909 485509 384229 485593
rect 383909 485273 383951 485509
rect 384187 485273 384229 485509
rect 383909 485241 384229 485273
rect 389840 485829 390160 485861
rect 389840 485593 389882 485829
rect 390118 485593 390160 485829
rect 389840 485509 390160 485593
rect 389840 485273 389882 485509
rect 390118 485273 390160 485509
rect 389840 485241 390160 485273
rect 395770 485829 396090 485861
rect 395770 485593 395812 485829
rect 396048 485593 396090 485829
rect 395770 485509 396090 485593
rect 395770 485273 395812 485509
rect 396048 485273 396090 485509
rect 395770 485241 396090 485273
rect 411909 485829 412229 485861
rect 411909 485593 411951 485829
rect 412187 485593 412229 485829
rect 411909 485509 412229 485593
rect 411909 485273 411951 485509
rect 412187 485273 412229 485509
rect 411909 485241 412229 485273
rect 417840 485829 418160 485861
rect 417840 485593 417882 485829
rect 418118 485593 418160 485829
rect 417840 485509 418160 485593
rect 417840 485273 417882 485509
rect 418118 485273 418160 485509
rect 417840 485241 418160 485273
rect 423770 485829 424090 485861
rect 423770 485593 423812 485829
rect 424048 485593 424090 485829
rect 423770 485509 424090 485593
rect 423770 485273 423812 485509
rect 424048 485273 424090 485509
rect 423770 485241 424090 485273
rect 439909 485829 440229 485861
rect 439909 485593 439951 485829
rect 440187 485593 440229 485829
rect 439909 485509 440229 485593
rect 439909 485273 439951 485509
rect 440187 485273 440229 485509
rect 439909 485241 440229 485273
rect 445840 485829 446160 485861
rect 445840 485593 445882 485829
rect 446118 485593 446160 485829
rect 445840 485509 446160 485593
rect 445840 485273 445882 485509
rect 446118 485273 446160 485509
rect 445840 485241 446160 485273
rect 451770 485829 452090 485861
rect 451770 485593 451812 485829
rect 452048 485593 452090 485829
rect 451770 485509 452090 485593
rect 451770 485273 451812 485509
rect 452048 485273 452090 485509
rect 451770 485241 452090 485273
rect 467909 485829 468229 485861
rect 467909 485593 467951 485829
rect 468187 485593 468229 485829
rect 467909 485509 468229 485593
rect 467909 485273 467951 485509
rect 468187 485273 468229 485509
rect 467909 485241 468229 485273
rect 473840 485829 474160 485861
rect 473840 485593 473882 485829
rect 474118 485593 474160 485829
rect 473840 485509 474160 485593
rect 473840 485273 473882 485509
rect 474118 485273 474160 485509
rect 473840 485241 474160 485273
rect 479770 485829 480090 485861
rect 479770 485593 479812 485829
rect 480048 485593 480090 485829
rect 479770 485509 480090 485593
rect 479770 485273 479812 485509
rect 480048 485273 480090 485509
rect 479770 485241 480090 485273
rect 495909 485829 496229 485861
rect 495909 485593 495951 485829
rect 496187 485593 496229 485829
rect 495909 485509 496229 485593
rect 495909 485273 495951 485509
rect 496187 485273 496229 485509
rect 495909 485241 496229 485273
rect 501840 485829 502160 485861
rect 501840 485593 501882 485829
rect 502118 485593 502160 485829
rect 501840 485509 502160 485593
rect 501840 485273 501882 485509
rect 502118 485273 502160 485509
rect 501840 485241 502160 485273
rect 507770 485829 508090 485861
rect 507770 485593 507812 485829
rect 508048 485593 508090 485829
rect 507770 485509 508090 485593
rect 507770 485273 507812 485509
rect 508048 485273 508090 485509
rect 507770 485241 508090 485273
rect 523909 485829 524229 485861
rect 523909 485593 523951 485829
rect 524187 485593 524229 485829
rect 523909 485509 524229 485593
rect 523909 485273 523951 485509
rect 524187 485273 524229 485509
rect 523909 485241 524229 485273
rect 529840 485829 530160 485861
rect 529840 485593 529882 485829
rect 530118 485593 530160 485829
rect 529840 485509 530160 485593
rect 529840 485273 529882 485509
rect 530118 485273 530160 485509
rect 529840 485241 530160 485273
rect 535770 485829 536090 485861
rect 535770 485593 535812 485829
rect 536048 485593 536090 485829
rect 535770 485509 536090 485593
rect 535770 485273 535812 485509
rect 536048 485273 536090 485509
rect 535770 485241 536090 485273
rect 551909 485829 552229 485861
rect 551909 485593 551951 485829
rect 552187 485593 552229 485829
rect 551909 485509 552229 485593
rect 551909 485273 551951 485509
rect 552187 485273 552229 485509
rect 551909 485241 552229 485273
rect 557840 485829 558160 485861
rect 557840 485593 557882 485829
rect 558118 485593 558160 485829
rect 557840 485509 558160 485593
rect 557840 485273 557882 485509
rect 558118 485273 558160 485509
rect 557840 485241 558160 485273
rect 563770 485829 564090 485861
rect 563770 485593 563812 485829
rect 564048 485593 564090 485829
rect 563770 485509 564090 485593
rect 563770 485273 563812 485509
rect 564048 485273 564090 485509
rect 563770 485241 564090 485273
rect 573494 485829 574114 512273
rect 573494 485593 573526 485829
rect 573762 485593 573846 485829
rect 574082 485593 574114 485829
rect 573494 485509 574114 485593
rect 573494 485273 573526 485509
rect 573762 485273 573846 485509
rect 574082 485273 574114 485509
rect 22875 482454 23195 482486
rect 22875 482218 22917 482454
rect 23153 482218 23195 482454
rect 22875 482134 23195 482218
rect 22875 481898 22917 482134
rect 23153 481898 23195 482134
rect 22875 481866 23195 481898
rect 28806 482454 29126 482486
rect 28806 482218 28848 482454
rect 29084 482218 29126 482454
rect 28806 482134 29126 482218
rect 28806 481898 28848 482134
rect 29084 481898 29126 482134
rect 28806 481866 29126 481898
rect 50875 482454 51195 482486
rect 50875 482218 50917 482454
rect 51153 482218 51195 482454
rect 50875 482134 51195 482218
rect 50875 481898 50917 482134
rect 51153 481898 51195 482134
rect 50875 481866 51195 481898
rect 56806 482454 57126 482486
rect 56806 482218 56848 482454
rect 57084 482218 57126 482454
rect 56806 482134 57126 482218
rect 56806 481898 56848 482134
rect 57084 481898 57126 482134
rect 56806 481866 57126 481898
rect 78875 482454 79195 482486
rect 78875 482218 78917 482454
rect 79153 482218 79195 482454
rect 78875 482134 79195 482218
rect 78875 481898 78917 482134
rect 79153 481898 79195 482134
rect 78875 481866 79195 481898
rect 84806 482454 85126 482486
rect 84806 482218 84848 482454
rect 85084 482218 85126 482454
rect 84806 482134 85126 482218
rect 84806 481898 84848 482134
rect 85084 481898 85126 482134
rect 84806 481866 85126 481898
rect 106875 482454 107195 482486
rect 106875 482218 106917 482454
rect 107153 482218 107195 482454
rect 106875 482134 107195 482218
rect 106875 481898 106917 482134
rect 107153 481898 107195 482134
rect 106875 481866 107195 481898
rect 112806 482454 113126 482486
rect 112806 482218 112848 482454
rect 113084 482218 113126 482454
rect 112806 482134 113126 482218
rect 112806 481898 112848 482134
rect 113084 481898 113126 482134
rect 112806 481866 113126 481898
rect 134875 482454 135195 482486
rect 134875 482218 134917 482454
rect 135153 482218 135195 482454
rect 134875 482134 135195 482218
rect 134875 481898 134917 482134
rect 135153 481898 135195 482134
rect 134875 481866 135195 481898
rect 140806 482454 141126 482486
rect 140806 482218 140848 482454
rect 141084 482218 141126 482454
rect 140806 482134 141126 482218
rect 140806 481898 140848 482134
rect 141084 481898 141126 482134
rect 140806 481866 141126 481898
rect 162875 482454 163195 482486
rect 162875 482218 162917 482454
rect 163153 482218 163195 482454
rect 162875 482134 163195 482218
rect 162875 481898 162917 482134
rect 163153 481898 163195 482134
rect 162875 481866 163195 481898
rect 168806 482454 169126 482486
rect 168806 482218 168848 482454
rect 169084 482218 169126 482454
rect 168806 482134 169126 482218
rect 168806 481898 168848 482134
rect 169084 481898 169126 482134
rect 168806 481866 169126 481898
rect 190875 482454 191195 482486
rect 190875 482218 190917 482454
rect 191153 482218 191195 482454
rect 190875 482134 191195 482218
rect 190875 481898 190917 482134
rect 191153 481898 191195 482134
rect 190875 481866 191195 481898
rect 196806 482454 197126 482486
rect 196806 482218 196848 482454
rect 197084 482218 197126 482454
rect 196806 482134 197126 482218
rect 196806 481898 196848 482134
rect 197084 481898 197126 482134
rect 196806 481866 197126 481898
rect 218875 482454 219195 482486
rect 218875 482218 218917 482454
rect 219153 482218 219195 482454
rect 218875 482134 219195 482218
rect 218875 481898 218917 482134
rect 219153 481898 219195 482134
rect 218875 481866 219195 481898
rect 224806 482454 225126 482486
rect 224806 482218 224848 482454
rect 225084 482218 225126 482454
rect 224806 482134 225126 482218
rect 224806 481898 224848 482134
rect 225084 481898 225126 482134
rect 224806 481866 225126 481898
rect 246875 482454 247195 482486
rect 246875 482218 246917 482454
rect 247153 482218 247195 482454
rect 246875 482134 247195 482218
rect 246875 481898 246917 482134
rect 247153 481898 247195 482134
rect 246875 481866 247195 481898
rect 252806 482454 253126 482486
rect 252806 482218 252848 482454
rect 253084 482218 253126 482454
rect 252806 482134 253126 482218
rect 252806 481898 252848 482134
rect 253084 481898 253126 482134
rect 252806 481866 253126 481898
rect 274875 482454 275195 482486
rect 274875 482218 274917 482454
rect 275153 482218 275195 482454
rect 274875 482134 275195 482218
rect 274875 481898 274917 482134
rect 275153 481898 275195 482134
rect 274875 481866 275195 481898
rect 280806 482454 281126 482486
rect 280806 482218 280848 482454
rect 281084 482218 281126 482454
rect 280806 482134 281126 482218
rect 280806 481898 280848 482134
rect 281084 481898 281126 482134
rect 280806 481866 281126 481898
rect 302875 482454 303195 482486
rect 302875 482218 302917 482454
rect 303153 482218 303195 482454
rect 302875 482134 303195 482218
rect 302875 481898 302917 482134
rect 303153 481898 303195 482134
rect 302875 481866 303195 481898
rect 308806 482454 309126 482486
rect 308806 482218 308848 482454
rect 309084 482218 309126 482454
rect 308806 482134 309126 482218
rect 308806 481898 308848 482134
rect 309084 481898 309126 482134
rect 308806 481866 309126 481898
rect 330875 482454 331195 482486
rect 330875 482218 330917 482454
rect 331153 482218 331195 482454
rect 330875 482134 331195 482218
rect 330875 481898 330917 482134
rect 331153 481898 331195 482134
rect 330875 481866 331195 481898
rect 336806 482454 337126 482486
rect 336806 482218 336848 482454
rect 337084 482218 337126 482454
rect 336806 482134 337126 482218
rect 336806 481898 336848 482134
rect 337084 481898 337126 482134
rect 336806 481866 337126 481898
rect 358875 482454 359195 482486
rect 358875 482218 358917 482454
rect 359153 482218 359195 482454
rect 358875 482134 359195 482218
rect 358875 481898 358917 482134
rect 359153 481898 359195 482134
rect 358875 481866 359195 481898
rect 364806 482454 365126 482486
rect 364806 482218 364848 482454
rect 365084 482218 365126 482454
rect 364806 482134 365126 482218
rect 364806 481898 364848 482134
rect 365084 481898 365126 482134
rect 364806 481866 365126 481898
rect 386875 482454 387195 482486
rect 386875 482218 386917 482454
rect 387153 482218 387195 482454
rect 386875 482134 387195 482218
rect 386875 481898 386917 482134
rect 387153 481898 387195 482134
rect 386875 481866 387195 481898
rect 392806 482454 393126 482486
rect 392806 482218 392848 482454
rect 393084 482218 393126 482454
rect 392806 482134 393126 482218
rect 392806 481898 392848 482134
rect 393084 481898 393126 482134
rect 392806 481866 393126 481898
rect 414875 482454 415195 482486
rect 414875 482218 414917 482454
rect 415153 482218 415195 482454
rect 414875 482134 415195 482218
rect 414875 481898 414917 482134
rect 415153 481898 415195 482134
rect 414875 481866 415195 481898
rect 420806 482454 421126 482486
rect 420806 482218 420848 482454
rect 421084 482218 421126 482454
rect 420806 482134 421126 482218
rect 420806 481898 420848 482134
rect 421084 481898 421126 482134
rect 420806 481866 421126 481898
rect 442875 482454 443195 482486
rect 442875 482218 442917 482454
rect 443153 482218 443195 482454
rect 442875 482134 443195 482218
rect 442875 481898 442917 482134
rect 443153 481898 443195 482134
rect 442875 481866 443195 481898
rect 448806 482454 449126 482486
rect 448806 482218 448848 482454
rect 449084 482218 449126 482454
rect 448806 482134 449126 482218
rect 448806 481898 448848 482134
rect 449084 481898 449126 482134
rect 448806 481866 449126 481898
rect 470875 482454 471195 482486
rect 470875 482218 470917 482454
rect 471153 482218 471195 482454
rect 470875 482134 471195 482218
rect 470875 481898 470917 482134
rect 471153 481898 471195 482134
rect 470875 481866 471195 481898
rect 476806 482454 477126 482486
rect 476806 482218 476848 482454
rect 477084 482218 477126 482454
rect 476806 482134 477126 482218
rect 476806 481898 476848 482134
rect 477084 481898 477126 482134
rect 476806 481866 477126 481898
rect 498875 482454 499195 482486
rect 498875 482218 498917 482454
rect 499153 482218 499195 482454
rect 498875 482134 499195 482218
rect 498875 481898 498917 482134
rect 499153 481898 499195 482134
rect 498875 481866 499195 481898
rect 504806 482454 505126 482486
rect 504806 482218 504848 482454
rect 505084 482218 505126 482454
rect 504806 482134 505126 482218
rect 504806 481898 504848 482134
rect 505084 481898 505126 482134
rect 504806 481866 505126 481898
rect 526875 482454 527195 482486
rect 526875 482218 526917 482454
rect 527153 482218 527195 482454
rect 526875 482134 527195 482218
rect 526875 481898 526917 482134
rect 527153 481898 527195 482134
rect 526875 481866 527195 481898
rect 532806 482454 533126 482486
rect 532806 482218 532848 482454
rect 533084 482218 533126 482454
rect 532806 482134 533126 482218
rect 532806 481898 532848 482134
rect 533084 481898 533126 482134
rect 532806 481866 533126 481898
rect 554875 482454 555195 482486
rect 554875 482218 554917 482454
rect 555153 482218 555195 482454
rect 554875 482134 555195 482218
rect 554875 481898 554917 482134
rect 555153 481898 555195 482134
rect 554875 481866 555195 481898
rect 560806 482454 561126 482486
rect 560806 482218 560848 482454
rect 561084 482218 561126 482454
rect 560806 482134 561126 482218
rect 560806 481898 560848 482134
rect 561084 481898 561126 482134
rect 560806 481866 561126 481898
rect -2006 458593 -1974 458829
rect -1738 458593 -1654 458829
rect -1418 458593 -1386 458829
rect -2006 458509 -1386 458593
rect -2006 458273 -1974 458509
rect -1738 458273 -1654 458509
rect -1418 458273 -1386 458509
rect -2006 431829 -1386 458273
rect 19910 458829 20230 458861
rect 19910 458593 19952 458829
rect 20188 458593 20230 458829
rect 19910 458509 20230 458593
rect 19910 458273 19952 458509
rect 20188 458273 20230 458509
rect 19910 458241 20230 458273
rect 25840 458829 26160 458861
rect 25840 458593 25882 458829
rect 26118 458593 26160 458829
rect 25840 458509 26160 458593
rect 25840 458273 25882 458509
rect 26118 458273 26160 458509
rect 25840 458241 26160 458273
rect 31771 458829 32091 458861
rect 31771 458593 31813 458829
rect 32049 458593 32091 458829
rect 31771 458509 32091 458593
rect 31771 458273 31813 458509
rect 32049 458273 32091 458509
rect 31771 458241 32091 458273
rect 47910 458829 48230 458861
rect 47910 458593 47952 458829
rect 48188 458593 48230 458829
rect 47910 458509 48230 458593
rect 47910 458273 47952 458509
rect 48188 458273 48230 458509
rect 47910 458241 48230 458273
rect 53840 458829 54160 458861
rect 53840 458593 53882 458829
rect 54118 458593 54160 458829
rect 53840 458509 54160 458593
rect 53840 458273 53882 458509
rect 54118 458273 54160 458509
rect 53840 458241 54160 458273
rect 59771 458829 60091 458861
rect 59771 458593 59813 458829
rect 60049 458593 60091 458829
rect 59771 458509 60091 458593
rect 59771 458273 59813 458509
rect 60049 458273 60091 458509
rect 59771 458241 60091 458273
rect 75910 458829 76230 458861
rect 75910 458593 75952 458829
rect 76188 458593 76230 458829
rect 75910 458509 76230 458593
rect 75910 458273 75952 458509
rect 76188 458273 76230 458509
rect 75910 458241 76230 458273
rect 81840 458829 82160 458861
rect 81840 458593 81882 458829
rect 82118 458593 82160 458829
rect 81840 458509 82160 458593
rect 81840 458273 81882 458509
rect 82118 458273 82160 458509
rect 81840 458241 82160 458273
rect 87771 458829 88091 458861
rect 87771 458593 87813 458829
rect 88049 458593 88091 458829
rect 87771 458509 88091 458593
rect 87771 458273 87813 458509
rect 88049 458273 88091 458509
rect 87771 458241 88091 458273
rect 103910 458829 104230 458861
rect 103910 458593 103952 458829
rect 104188 458593 104230 458829
rect 103910 458509 104230 458593
rect 103910 458273 103952 458509
rect 104188 458273 104230 458509
rect 103910 458241 104230 458273
rect 109840 458829 110160 458861
rect 109840 458593 109882 458829
rect 110118 458593 110160 458829
rect 109840 458509 110160 458593
rect 109840 458273 109882 458509
rect 110118 458273 110160 458509
rect 109840 458241 110160 458273
rect 115771 458829 116091 458861
rect 115771 458593 115813 458829
rect 116049 458593 116091 458829
rect 115771 458509 116091 458593
rect 115771 458273 115813 458509
rect 116049 458273 116091 458509
rect 115771 458241 116091 458273
rect 131910 458829 132230 458861
rect 131910 458593 131952 458829
rect 132188 458593 132230 458829
rect 131910 458509 132230 458593
rect 131910 458273 131952 458509
rect 132188 458273 132230 458509
rect 131910 458241 132230 458273
rect 137840 458829 138160 458861
rect 137840 458593 137882 458829
rect 138118 458593 138160 458829
rect 137840 458509 138160 458593
rect 137840 458273 137882 458509
rect 138118 458273 138160 458509
rect 137840 458241 138160 458273
rect 143771 458829 144091 458861
rect 143771 458593 143813 458829
rect 144049 458593 144091 458829
rect 143771 458509 144091 458593
rect 143771 458273 143813 458509
rect 144049 458273 144091 458509
rect 143771 458241 144091 458273
rect 159910 458829 160230 458861
rect 159910 458593 159952 458829
rect 160188 458593 160230 458829
rect 159910 458509 160230 458593
rect 159910 458273 159952 458509
rect 160188 458273 160230 458509
rect 159910 458241 160230 458273
rect 165840 458829 166160 458861
rect 165840 458593 165882 458829
rect 166118 458593 166160 458829
rect 165840 458509 166160 458593
rect 165840 458273 165882 458509
rect 166118 458273 166160 458509
rect 165840 458241 166160 458273
rect 171771 458829 172091 458861
rect 171771 458593 171813 458829
rect 172049 458593 172091 458829
rect 171771 458509 172091 458593
rect 171771 458273 171813 458509
rect 172049 458273 172091 458509
rect 171771 458241 172091 458273
rect 187910 458829 188230 458861
rect 187910 458593 187952 458829
rect 188188 458593 188230 458829
rect 187910 458509 188230 458593
rect 187910 458273 187952 458509
rect 188188 458273 188230 458509
rect 187910 458241 188230 458273
rect 193840 458829 194160 458861
rect 193840 458593 193882 458829
rect 194118 458593 194160 458829
rect 193840 458509 194160 458593
rect 193840 458273 193882 458509
rect 194118 458273 194160 458509
rect 193840 458241 194160 458273
rect 199771 458829 200091 458861
rect 199771 458593 199813 458829
rect 200049 458593 200091 458829
rect 199771 458509 200091 458593
rect 199771 458273 199813 458509
rect 200049 458273 200091 458509
rect 199771 458241 200091 458273
rect 215910 458829 216230 458861
rect 215910 458593 215952 458829
rect 216188 458593 216230 458829
rect 215910 458509 216230 458593
rect 215910 458273 215952 458509
rect 216188 458273 216230 458509
rect 215910 458241 216230 458273
rect 221840 458829 222160 458861
rect 221840 458593 221882 458829
rect 222118 458593 222160 458829
rect 221840 458509 222160 458593
rect 221840 458273 221882 458509
rect 222118 458273 222160 458509
rect 221840 458241 222160 458273
rect 227771 458829 228091 458861
rect 227771 458593 227813 458829
rect 228049 458593 228091 458829
rect 227771 458509 228091 458593
rect 227771 458273 227813 458509
rect 228049 458273 228091 458509
rect 227771 458241 228091 458273
rect 243910 458829 244230 458861
rect 243910 458593 243952 458829
rect 244188 458593 244230 458829
rect 243910 458509 244230 458593
rect 243910 458273 243952 458509
rect 244188 458273 244230 458509
rect 243910 458241 244230 458273
rect 249840 458829 250160 458861
rect 249840 458593 249882 458829
rect 250118 458593 250160 458829
rect 249840 458509 250160 458593
rect 249840 458273 249882 458509
rect 250118 458273 250160 458509
rect 249840 458241 250160 458273
rect 255771 458829 256091 458861
rect 255771 458593 255813 458829
rect 256049 458593 256091 458829
rect 255771 458509 256091 458593
rect 255771 458273 255813 458509
rect 256049 458273 256091 458509
rect 255771 458241 256091 458273
rect 271910 458829 272230 458861
rect 271910 458593 271952 458829
rect 272188 458593 272230 458829
rect 271910 458509 272230 458593
rect 271910 458273 271952 458509
rect 272188 458273 272230 458509
rect 271910 458241 272230 458273
rect 277840 458829 278160 458861
rect 277840 458593 277882 458829
rect 278118 458593 278160 458829
rect 277840 458509 278160 458593
rect 277840 458273 277882 458509
rect 278118 458273 278160 458509
rect 277840 458241 278160 458273
rect 283771 458829 284091 458861
rect 283771 458593 283813 458829
rect 284049 458593 284091 458829
rect 283771 458509 284091 458593
rect 283771 458273 283813 458509
rect 284049 458273 284091 458509
rect 283771 458241 284091 458273
rect 299910 458829 300230 458861
rect 299910 458593 299952 458829
rect 300188 458593 300230 458829
rect 299910 458509 300230 458593
rect 299910 458273 299952 458509
rect 300188 458273 300230 458509
rect 299910 458241 300230 458273
rect 305840 458829 306160 458861
rect 305840 458593 305882 458829
rect 306118 458593 306160 458829
rect 305840 458509 306160 458593
rect 305840 458273 305882 458509
rect 306118 458273 306160 458509
rect 305840 458241 306160 458273
rect 311771 458829 312091 458861
rect 311771 458593 311813 458829
rect 312049 458593 312091 458829
rect 311771 458509 312091 458593
rect 311771 458273 311813 458509
rect 312049 458273 312091 458509
rect 311771 458241 312091 458273
rect 327910 458829 328230 458861
rect 327910 458593 327952 458829
rect 328188 458593 328230 458829
rect 327910 458509 328230 458593
rect 327910 458273 327952 458509
rect 328188 458273 328230 458509
rect 327910 458241 328230 458273
rect 333840 458829 334160 458861
rect 333840 458593 333882 458829
rect 334118 458593 334160 458829
rect 333840 458509 334160 458593
rect 333840 458273 333882 458509
rect 334118 458273 334160 458509
rect 333840 458241 334160 458273
rect 339771 458829 340091 458861
rect 339771 458593 339813 458829
rect 340049 458593 340091 458829
rect 339771 458509 340091 458593
rect 339771 458273 339813 458509
rect 340049 458273 340091 458509
rect 339771 458241 340091 458273
rect 355910 458829 356230 458861
rect 355910 458593 355952 458829
rect 356188 458593 356230 458829
rect 355910 458509 356230 458593
rect 355910 458273 355952 458509
rect 356188 458273 356230 458509
rect 355910 458241 356230 458273
rect 361840 458829 362160 458861
rect 361840 458593 361882 458829
rect 362118 458593 362160 458829
rect 361840 458509 362160 458593
rect 361840 458273 361882 458509
rect 362118 458273 362160 458509
rect 361840 458241 362160 458273
rect 367771 458829 368091 458861
rect 367771 458593 367813 458829
rect 368049 458593 368091 458829
rect 367771 458509 368091 458593
rect 367771 458273 367813 458509
rect 368049 458273 368091 458509
rect 367771 458241 368091 458273
rect 383910 458829 384230 458861
rect 383910 458593 383952 458829
rect 384188 458593 384230 458829
rect 383910 458509 384230 458593
rect 383910 458273 383952 458509
rect 384188 458273 384230 458509
rect 383910 458241 384230 458273
rect 389840 458829 390160 458861
rect 389840 458593 389882 458829
rect 390118 458593 390160 458829
rect 389840 458509 390160 458593
rect 389840 458273 389882 458509
rect 390118 458273 390160 458509
rect 389840 458241 390160 458273
rect 395771 458829 396091 458861
rect 395771 458593 395813 458829
rect 396049 458593 396091 458829
rect 395771 458509 396091 458593
rect 395771 458273 395813 458509
rect 396049 458273 396091 458509
rect 395771 458241 396091 458273
rect 411910 458829 412230 458861
rect 411910 458593 411952 458829
rect 412188 458593 412230 458829
rect 411910 458509 412230 458593
rect 411910 458273 411952 458509
rect 412188 458273 412230 458509
rect 411910 458241 412230 458273
rect 417840 458829 418160 458861
rect 417840 458593 417882 458829
rect 418118 458593 418160 458829
rect 417840 458509 418160 458593
rect 417840 458273 417882 458509
rect 418118 458273 418160 458509
rect 417840 458241 418160 458273
rect 423771 458829 424091 458861
rect 423771 458593 423813 458829
rect 424049 458593 424091 458829
rect 423771 458509 424091 458593
rect 423771 458273 423813 458509
rect 424049 458273 424091 458509
rect 423771 458241 424091 458273
rect 439910 458829 440230 458861
rect 439910 458593 439952 458829
rect 440188 458593 440230 458829
rect 439910 458509 440230 458593
rect 439910 458273 439952 458509
rect 440188 458273 440230 458509
rect 439910 458241 440230 458273
rect 445840 458829 446160 458861
rect 445840 458593 445882 458829
rect 446118 458593 446160 458829
rect 445840 458509 446160 458593
rect 445840 458273 445882 458509
rect 446118 458273 446160 458509
rect 445840 458241 446160 458273
rect 451771 458829 452091 458861
rect 451771 458593 451813 458829
rect 452049 458593 452091 458829
rect 451771 458509 452091 458593
rect 451771 458273 451813 458509
rect 452049 458273 452091 458509
rect 451771 458241 452091 458273
rect 467910 458829 468230 458861
rect 467910 458593 467952 458829
rect 468188 458593 468230 458829
rect 467910 458509 468230 458593
rect 467910 458273 467952 458509
rect 468188 458273 468230 458509
rect 467910 458241 468230 458273
rect 473840 458829 474160 458861
rect 473840 458593 473882 458829
rect 474118 458593 474160 458829
rect 473840 458509 474160 458593
rect 473840 458273 473882 458509
rect 474118 458273 474160 458509
rect 473840 458241 474160 458273
rect 479771 458829 480091 458861
rect 479771 458593 479813 458829
rect 480049 458593 480091 458829
rect 479771 458509 480091 458593
rect 479771 458273 479813 458509
rect 480049 458273 480091 458509
rect 479771 458241 480091 458273
rect 495910 458829 496230 458861
rect 495910 458593 495952 458829
rect 496188 458593 496230 458829
rect 495910 458509 496230 458593
rect 495910 458273 495952 458509
rect 496188 458273 496230 458509
rect 495910 458241 496230 458273
rect 501840 458829 502160 458861
rect 501840 458593 501882 458829
rect 502118 458593 502160 458829
rect 501840 458509 502160 458593
rect 501840 458273 501882 458509
rect 502118 458273 502160 458509
rect 501840 458241 502160 458273
rect 507771 458829 508091 458861
rect 507771 458593 507813 458829
rect 508049 458593 508091 458829
rect 507771 458509 508091 458593
rect 507771 458273 507813 458509
rect 508049 458273 508091 458509
rect 507771 458241 508091 458273
rect 523910 458829 524230 458861
rect 523910 458593 523952 458829
rect 524188 458593 524230 458829
rect 523910 458509 524230 458593
rect 523910 458273 523952 458509
rect 524188 458273 524230 458509
rect 523910 458241 524230 458273
rect 529840 458829 530160 458861
rect 529840 458593 529882 458829
rect 530118 458593 530160 458829
rect 529840 458509 530160 458593
rect 529840 458273 529882 458509
rect 530118 458273 530160 458509
rect 529840 458241 530160 458273
rect 535771 458829 536091 458861
rect 535771 458593 535813 458829
rect 536049 458593 536091 458829
rect 535771 458509 536091 458593
rect 535771 458273 535813 458509
rect 536049 458273 536091 458509
rect 535771 458241 536091 458273
rect 551910 458829 552230 458861
rect 551910 458593 551952 458829
rect 552188 458593 552230 458829
rect 551910 458509 552230 458593
rect 551910 458273 551952 458509
rect 552188 458273 552230 458509
rect 551910 458241 552230 458273
rect 557840 458829 558160 458861
rect 557840 458593 557882 458829
rect 558118 458593 558160 458829
rect 557840 458509 558160 458593
rect 557840 458273 557882 458509
rect 558118 458273 558160 458509
rect 557840 458241 558160 458273
rect 563771 458829 564091 458861
rect 563771 458593 563813 458829
rect 564049 458593 564091 458829
rect 563771 458509 564091 458593
rect 563771 458273 563813 458509
rect 564049 458273 564091 458509
rect 563771 458241 564091 458273
rect 573494 458829 574114 485273
rect 573494 458593 573526 458829
rect 573762 458593 573846 458829
rect 574082 458593 574114 458829
rect 573494 458509 574114 458593
rect 573494 458273 573526 458509
rect 573762 458273 573846 458509
rect 574082 458273 574114 458509
rect 22874 455454 23194 455486
rect 22874 455218 22916 455454
rect 23152 455218 23194 455454
rect 22874 455134 23194 455218
rect 22874 454898 22916 455134
rect 23152 454898 23194 455134
rect 22874 454866 23194 454898
rect 28805 455454 29125 455486
rect 28805 455218 28847 455454
rect 29083 455218 29125 455454
rect 28805 455134 29125 455218
rect 28805 454898 28847 455134
rect 29083 454898 29125 455134
rect 28805 454866 29125 454898
rect 50874 455454 51194 455486
rect 50874 455218 50916 455454
rect 51152 455218 51194 455454
rect 50874 455134 51194 455218
rect 50874 454898 50916 455134
rect 51152 454898 51194 455134
rect 50874 454866 51194 454898
rect 56805 455454 57125 455486
rect 56805 455218 56847 455454
rect 57083 455218 57125 455454
rect 56805 455134 57125 455218
rect 56805 454898 56847 455134
rect 57083 454898 57125 455134
rect 56805 454866 57125 454898
rect 78874 455454 79194 455486
rect 78874 455218 78916 455454
rect 79152 455218 79194 455454
rect 78874 455134 79194 455218
rect 78874 454898 78916 455134
rect 79152 454898 79194 455134
rect 78874 454866 79194 454898
rect 84805 455454 85125 455486
rect 84805 455218 84847 455454
rect 85083 455218 85125 455454
rect 84805 455134 85125 455218
rect 84805 454898 84847 455134
rect 85083 454898 85125 455134
rect 84805 454866 85125 454898
rect 106874 455454 107194 455486
rect 106874 455218 106916 455454
rect 107152 455218 107194 455454
rect 106874 455134 107194 455218
rect 106874 454898 106916 455134
rect 107152 454898 107194 455134
rect 106874 454866 107194 454898
rect 112805 455454 113125 455486
rect 112805 455218 112847 455454
rect 113083 455218 113125 455454
rect 112805 455134 113125 455218
rect 112805 454898 112847 455134
rect 113083 454898 113125 455134
rect 112805 454866 113125 454898
rect 134874 455454 135194 455486
rect 134874 455218 134916 455454
rect 135152 455218 135194 455454
rect 134874 455134 135194 455218
rect 134874 454898 134916 455134
rect 135152 454898 135194 455134
rect 134874 454866 135194 454898
rect 140805 455454 141125 455486
rect 140805 455218 140847 455454
rect 141083 455218 141125 455454
rect 140805 455134 141125 455218
rect 140805 454898 140847 455134
rect 141083 454898 141125 455134
rect 140805 454866 141125 454898
rect 162874 455454 163194 455486
rect 162874 455218 162916 455454
rect 163152 455218 163194 455454
rect 162874 455134 163194 455218
rect 162874 454898 162916 455134
rect 163152 454898 163194 455134
rect 162874 454866 163194 454898
rect 168805 455454 169125 455486
rect 168805 455218 168847 455454
rect 169083 455218 169125 455454
rect 168805 455134 169125 455218
rect 168805 454898 168847 455134
rect 169083 454898 169125 455134
rect 168805 454866 169125 454898
rect 190874 455454 191194 455486
rect 190874 455218 190916 455454
rect 191152 455218 191194 455454
rect 190874 455134 191194 455218
rect 190874 454898 190916 455134
rect 191152 454898 191194 455134
rect 190874 454866 191194 454898
rect 196805 455454 197125 455486
rect 196805 455218 196847 455454
rect 197083 455218 197125 455454
rect 196805 455134 197125 455218
rect 196805 454898 196847 455134
rect 197083 454898 197125 455134
rect 196805 454866 197125 454898
rect 218874 455454 219194 455486
rect 218874 455218 218916 455454
rect 219152 455218 219194 455454
rect 218874 455134 219194 455218
rect 218874 454898 218916 455134
rect 219152 454898 219194 455134
rect 218874 454866 219194 454898
rect 224805 455454 225125 455486
rect 224805 455218 224847 455454
rect 225083 455218 225125 455454
rect 224805 455134 225125 455218
rect 224805 454898 224847 455134
rect 225083 454898 225125 455134
rect 224805 454866 225125 454898
rect 246874 455454 247194 455486
rect 246874 455218 246916 455454
rect 247152 455218 247194 455454
rect 246874 455134 247194 455218
rect 246874 454898 246916 455134
rect 247152 454898 247194 455134
rect 246874 454866 247194 454898
rect 252805 455454 253125 455486
rect 252805 455218 252847 455454
rect 253083 455218 253125 455454
rect 252805 455134 253125 455218
rect 252805 454898 252847 455134
rect 253083 454898 253125 455134
rect 252805 454866 253125 454898
rect 274874 455454 275194 455486
rect 274874 455218 274916 455454
rect 275152 455218 275194 455454
rect 274874 455134 275194 455218
rect 274874 454898 274916 455134
rect 275152 454898 275194 455134
rect 274874 454866 275194 454898
rect 280805 455454 281125 455486
rect 280805 455218 280847 455454
rect 281083 455218 281125 455454
rect 280805 455134 281125 455218
rect 280805 454898 280847 455134
rect 281083 454898 281125 455134
rect 280805 454866 281125 454898
rect 302874 455454 303194 455486
rect 302874 455218 302916 455454
rect 303152 455218 303194 455454
rect 302874 455134 303194 455218
rect 302874 454898 302916 455134
rect 303152 454898 303194 455134
rect 302874 454866 303194 454898
rect 308805 455454 309125 455486
rect 308805 455218 308847 455454
rect 309083 455218 309125 455454
rect 308805 455134 309125 455218
rect 308805 454898 308847 455134
rect 309083 454898 309125 455134
rect 308805 454866 309125 454898
rect 330874 455454 331194 455486
rect 330874 455218 330916 455454
rect 331152 455218 331194 455454
rect 330874 455134 331194 455218
rect 330874 454898 330916 455134
rect 331152 454898 331194 455134
rect 330874 454866 331194 454898
rect 336805 455454 337125 455486
rect 336805 455218 336847 455454
rect 337083 455218 337125 455454
rect 336805 455134 337125 455218
rect 336805 454898 336847 455134
rect 337083 454898 337125 455134
rect 336805 454866 337125 454898
rect 358874 455454 359194 455486
rect 358874 455218 358916 455454
rect 359152 455218 359194 455454
rect 358874 455134 359194 455218
rect 358874 454898 358916 455134
rect 359152 454898 359194 455134
rect 358874 454866 359194 454898
rect 364805 455454 365125 455486
rect 364805 455218 364847 455454
rect 365083 455218 365125 455454
rect 364805 455134 365125 455218
rect 364805 454898 364847 455134
rect 365083 454898 365125 455134
rect 364805 454866 365125 454898
rect 386874 455454 387194 455486
rect 386874 455218 386916 455454
rect 387152 455218 387194 455454
rect 386874 455134 387194 455218
rect 386874 454898 386916 455134
rect 387152 454898 387194 455134
rect 386874 454866 387194 454898
rect 392805 455454 393125 455486
rect 392805 455218 392847 455454
rect 393083 455218 393125 455454
rect 392805 455134 393125 455218
rect 392805 454898 392847 455134
rect 393083 454898 393125 455134
rect 392805 454866 393125 454898
rect 414874 455454 415194 455486
rect 414874 455218 414916 455454
rect 415152 455218 415194 455454
rect 414874 455134 415194 455218
rect 414874 454898 414916 455134
rect 415152 454898 415194 455134
rect 414874 454866 415194 454898
rect 420805 455454 421125 455486
rect 420805 455218 420847 455454
rect 421083 455218 421125 455454
rect 420805 455134 421125 455218
rect 420805 454898 420847 455134
rect 421083 454898 421125 455134
rect 420805 454866 421125 454898
rect 442874 455454 443194 455486
rect 442874 455218 442916 455454
rect 443152 455218 443194 455454
rect 442874 455134 443194 455218
rect 442874 454898 442916 455134
rect 443152 454898 443194 455134
rect 442874 454866 443194 454898
rect 448805 455454 449125 455486
rect 448805 455218 448847 455454
rect 449083 455218 449125 455454
rect 448805 455134 449125 455218
rect 448805 454898 448847 455134
rect 449083 454898 449125 455134
rect 448805 454866 449125 454898
rect 470874 455454 471194 455486
rect 470874 455218 470916 455454
rect 471152 455218 471194 455454
rect 470874 455134 471194 455218
rect 470874 454898 470916 455134
rect 471152 454898 471194 455134
rect 470874 454866 471194 454898
rect 476805 455454 477125 455486
rect 476805 455218 476847 455454
rect 477083 455218 477125 455454
rect 476805 455134 477125 455218
rect 476805 454898 476847 455134
rect 477083 454898 477125 455134
rect 476805 454866 477125 454898
rect 498874 455454 499194 455486
rect 498874 455218 498916 455454
rect 499152 455218 499194 455454
rect 498874 455134 499194 455218
rect 498874 454898 498916 455134
rect 499152 454898 499194 455134
rect 498874 454866 499194 454898
rect 504805 455454 505125 455486
rect 504805 455218 504847 455454
rect 505083 455218 505125 455454
rect 504805 455134 505125 455218
rect 504805 454898 504847 455134
rect 505083 454898 505125 455134
rect 504805 454866 505125 454898
rect 526874 455454 527194 455486
rect 526874 455218 526916 455454
rect 527152 455218 527194 455454
rect 526874 455134 527194 455218
rect 526874 454898 526916 455134
rect 527152 454898 527194 455134
rect 526874 454866 527194 454898
rect 532805 455454 533125 455486
rect 532805 455218 532847 455454
rect 533083 455218 533125 455454
rect 532805 455134 533125 455218
rect 532805 454898 532847 455134
rect 533083 454898 533125 455134
rect 532805 454866 533125 454898
rect 554874 455454 555194 455486
rect 554874 455218 554916 455454
rect 555152 455218 555194 455454
rect 554874 455134 555194 455218
rect 554874 454898 554916 455134
rect 555152 454898 555194 455134
rect 554874 454866 555194 454898
rect 560805 455454 561125 455486
rect 560805 455218 560847 455454
rect 561083 455218 561125 455454
rect 560805 455134 561125 455218
rect 560805 454898 560847 455134
rect 561083 454898 561125 455134
rect 560805 454866 561125 454898
rect -2006 431593 -1974 431829
rect -1738 431593 -1654 431829
rect -1418 431593 -1386 431829
rect -2006 431509 -1386 431593
rect -2006 431273 -1974 431509
rect -1738 431273 -1654 431509
rect -1418 431273 -1386 431509
rect -2006 404829 -1386 431273
rect 19909 431829 20229 431861
rect 19909 431593 19951 431829
rect 20187 431593 20229 431829
rect 19909 431509 20229 431593
rect 19909 431273 19951 431509
rect 20187 431273 20229 431509
rect 19909 431241 20229 431273
rect 25840 431829 26160 431861
rect 25840 431593 25882 431829
rect 26118 431593 26160 431829
rect 25840 431509 26160 431593
rect 25840 431273 25882 431509
rect 26118 431273 26160 431509
rect 25840 431241 26160 431273
rect 31770 431829 32090 431861
rect 31770 431593 31812 431829
rect 32048 431593 32090 431829
rect 31770 431509 32090 431593
rect 31770 431273 31812 431509
rect 32048 431273 32090 431509
rect 31770 431241 32090 431273
rect 47909 431829 48229 431861
rect 47909 431593 47951 431829
rect 48187 431593 48229 431829
rect 47909 431509 48229 431593
rect 47909 431273 47951 431509
rect 48187 431273 48229 431509
rect 47909 431241 48229 431273
rect 53840 431829 54160 431861
rect 53840 431593 53882 431829
rect 54118 431593 54160 431829
rect 53840 431509 54160 431593
rect 53840 431273 53882 431509
rect 54118 431273 54160 431509
rect 53840 431241 54160 431273
rect 59770 431829 60090 431861
rect 59770 431593 59812 431829
rect 60048 431593 60090 431829
rect 59770 431509 60090 431593
rect 59770 431273 59812 431509
rect 60048 431273 60090 431509
rect 59770 431241 60090 431273
rect 75909 431829 76229 431861
rect 75909 431593 75951 431829
rect 76187 431593 76229 431829
rect 75909 431509 76229 431593
rect 75909 431273 75951 431509
rect 76187 431273 76229 431509
rect 75909 431241 76229 431273
rect 81840 431829 82160 431861
rect 81840 431593 81882 431829
rect 82118 431593 82160 431829
rect 81840 431509 82160 431593
rect 81840 431273 81882 431509
rect 82118 431273 82160 431509
rect 81840 431241 82160 431273
rect 87770 431829 88090 431861
rect 87770 431593 87812 431829
rect 88048 431593 88090 431829
rect 87770 431509 88090 431593
rect 87770 431273 87812 431509
rect 88048 431273 88090 431509
rect 87770 431241 88090 431273
rect 103909 431829 104229 431861
rect 103909 431593 103951 431829
rect 104187 431593 104229 431829
rect 103909 431509 104229 431593
rect 103909 431273 103951 431509
rect 104187 431273 104229 431509
rect 103909 431241 104229 431273
rect 109840 431829 110160 431861
rect 109840 431593 109882 431829
rect 110118 431593 110160 431829
rect 109840 431509 110160 431593
rect 109840 431273 109882 431509
rect 110118 431273 110160 431509
rect 109840 431241 110160 431273
rect 115770 431829 116090 431861
rect 115770 431593 115812 431829
rect 116048 431593 116090 431829
rect 115770 431509 116090 431593
rect 115770 431273 115812 431509
rect 116048 431273 116090 431509
rect 115770 431241 116090 431273
rect 131909 431829 132229 431861
rect 131909 431593 131951 431829
rect 132187 431593 132229 431829
rect 131909 431509 132229 431593
rect 131909 431273 131951 431509
rect 132187 431273 132229 431509
rect 131909 431241 132229 431273
rect 137840 431829 138160 431861
rect 137840 431593 137882 431829
rect 138118 431593 138160 431829
rect 137840 431509 138160 431593
rect 137840 431273 137882 431509
rect 138118 431273 138160 431509
rect 137840 431241 138160 431273
rect 143770 431829 144090 431861
rect 143770 431593 143812 431829
rect 144048 431593 144090 431829
rect 143770 431509 144090 431593
rect 143770 431273 143812 431509
rect 144048 431273 144090 431509
rect 143770 431241 144090 431273
rect 159909 431829 160229 431861
rect 159909 431593 159951 431829
rect 160187 431593 160229 431829
rect 159909 431509 160229 431593
rect 159909 431273 159951 431509
rect 160187 431273 160229 431509
rect 159909 431241 160229 431273
rect 165840 431829 166160 431861
rect 165840 431593 165882 431829
rect 166118 431593 166160 431829
rect 165840 431509 166160 431593
rect 165840 431273 165882 431509
rect 166118 431273 166160 431509
rect 165840 431241 166160 431273
rect 171770 431829 172090 431861
rect 171770 431593 171812 431829
rect 172048 431593 172090 431829
rect 171770 431509 172090 431593
rect 171770 431273 171812 431509
rect 172048 431273 172090 431509
rect 171770 431241 172090 431273
rect 187909 431829 188229 431861
rect 187909 431593 187951 431829
rect 188187 431593 188229 431829
rect 187909 431509 188229 431593
rect 187909 431273 187951 431509
rect 188187 431273 188229 431509
rect 187909 431241 188229 431273
rect 193840 431829 194160 431861
rect 193840 431593 193882 431829
rect 194118 431593 194160 431829
rect 193840 431509 194160 431593
rect 193840 431273 193882 431509
rect 194118 431273 194160 431509
rect 193840 431241 194160 431273
rect 199770 431829 200090 431861
rect 199770 431593 199812 431829
rect 200048 431593 200090 431829
rect 199770 431509 200090 431593
rect 199770 431273 199812 431509
rect 200048 431273 200090 431509
rect 199770 431241 200090 431273
rect 215909 431829 216229 431861
rect 215909 431593 215951 431829
rect 216187 431593 216229 431829
rect 215909 431509 216229 431593
rect 215909 431273 215951 431509
rect 216187 431273 216229 431509
rect 215909 431241 216229 431273
rect 221840 431829 222160 431861
rect 221840 431593 221882 431829
rect 222118 431593 222160 431829
rect 221840 431509 222160 431593
rect 221840 431273 221882 431509
rect 222118 431273 222160 431509
rect 221840 431241 222160 431273
rect 227770 431829 228090 431861
rect 227770 431593 227812 431829
rect 228048 431593 228090 431829
rect 227770 431509 228090 431593
rect 227770 431273 227812 431509
rect 228048 431273 228090 431509
rect 227770 431241 228090 431273
rect 243909 431829 244229 431861
rect 243909 431593 243951 431829
rect 244187 431593 244229 431829
rect 243909 431509 244229 431593
rect 243909 431273 243951 431509
rect 244187 431273 244229 431509
rect 243909 431241 244229 431273
rect 249840 431829 250160 431861
rect 249840 431593 249882 431829
rect 250118 431593 250160 431829
rect 249840 431509 250160 431593
rect 249840 431273 249882 431509
rect 250118 431273 250160 431509
rect 249840 431241 250160 431273
rect 255770 431829 256090 431861
rect 255770 431593 255812 431829
rect 256048 431593 256090 431829
rect 255770 431509 256090 431593
rect 255770 431273 255812 431509
rect 256048 431273 256090 431509
rect 255770 431241 256090 431273
rect 271909 431829 272229 431861
rect 271909 431593 271951 431829
rect 272187 431593 272229 431829
rect 271909 431509 272229 431593
rect 271909 431273 271951 431509
rect 272187 431273 272229 431509
rect 271909 431241 272229 431273
rect 277840 431829 278160 431861
rect 277840 431593 277882 431829
rect 278118 431593 278160 431829
rect 277840 431509 278160 431593
rect 277840 431273 277882 431509
rect 278118 431273 278160 431509
rect 277840 431241 278160 431273
rect 283770 431829 284090 431861
rect 283770 431593 283812 431829
rect 284048 431593 284090 431829
rect 283770 431509 284090 431593
rect 283770 431273 283812 431509
rect 284048 431273 284090 431509
rect 283770 431241 284090 431273
rect 299909 431829 300229 431861
rect 299909 431593 299951 431829
rect 300187 431593 300229 431829
rect 299909 431509 300229 431593
rect 299909 431273 299951 431509
rect 300187 431273 300229 431509
rect 299909 431241 300229 431273
rect 305840 431829 306160 431861
rect 305840 431593 305882 431829
rect 306118 431593 306160 431829
rect 305840 431509 306160 431593
rect 305840 431273 305882 431509
rect 306118 431273 306160 431509
rect 305840 431241 306160 431273
rect 311770 431829 312090 431861
rect 311770 431593 311812 431829
rect 312048 431593 312090 431829
rect 311770 431509 312090 431593
rect 311770 431273 311812 431509
rect 312048 431273 312090 431509
rect 311770 431241 312090 431273
rect 327909 431829 328229 431861
rect 327909 431593 327951 431829
rect 328187 431593 328229 431829
rect 327909 431509 328229 431593
rect 327909 431273 327951 431509
rect 328187 431273 328229 431509
rect 327909 431241 328229 431273
rect 333840 431829 334160 431861
rect 333840 431593 333882 431829
rect 334118 431593 334160 431829
rect 333840 431509 334160 431593
rect 333840 431273 333882 431509
rect 334118 431273 334160 431509
rect 333840 431241 334160 431273
rect 339770 431829 340090 431861
rect 339770 431593 339812 431829
rect 340048 431593 340090 431829
rect 339770 431509 340090 431593
rect 339770 431273 339812 431509
rect 340048 431273 340090 431509
rect 339770 431241 340090 431273
rect 355909 431829 356229 431861
rect 355909 431593 355951 431829
rect 356187 431593 356229 431829
rect 355909 431509 356229 431593
rect 355909 431273 355951 431509
rect 356187 431273 356229 431509
rect 355909 431241 356229 431273
rect 361840 431829 362160 431861
rect 361840 431593 361882 431829
rect 362118 431593 362160 431829
rect 361840 431509 362160 431593
rect 361840 431273 361882 431509
rect 362118 431273 362160 431509
rect 361840 431241 362160 431273
rect 367770 431829 368090 431861
rect 367770 431593 367812 431829
rect 368048 431593 368090 431829
rect 367770 431509 368090 431593
rect 367770 431273 367812 431509
rect 368048 431273 368090 431509
rect 367770 431241 368090 431273
rect 383909 431829 384229 431861
rect 383909 431593 383951 431829
rect 384187 431593 384229 431829
rect 383909 431509 384229 431593
rect 383909 431273 383951 431509
rect 384187 431273 384229 431509
rect 383909 431241 384229 431273
rect 389840 431829 390160 431861
rect 389840 431593 389882 431829
rect 390118 431593 390160 431829
rect 389840 431509 390160 431593
rect 389840 431273 389882 431509
rect 390118 431273 390160 431509
rect 389840 431241 390160 431273
rect 395770 431829 396090 431861
rect 395770 431593 395812 431829
rect 396048 431593 396090 431829
rect 395770 431509 396090 431593
rect 395770 431273 395812 431509
rect 396048 431273 396090 431509
rect 395770 431241 396090 431273
rect 411909 431829 412229 431861
rect 411909 431593 411951 431829
rect 412187 431593 412229 431829
rect 411909 431509 412229 431593
rect 411909 431273 411951 431509
rect 412187 431273 412229 431509
rect 411909 431241 412229 431273
rect 417840 431829 418160 431861
rect 417840 431593 417882 431829
rect 418118 431593 418160 431829
rect 417840 431509 418160 431593
rect 417840 431273 417882 431509
rect 418118 431273 418160 431509
rect 417840 431241 418160 431273
rect 423770 431829 424090 431861
rect 423770 431593 423812 431829
rect 424048 431593 424090 431829
rect 423770 431509 424090 431593
rect 423770 431273 423812 431509
rect 424048 431273 424090 431509
rect 423770 431241 424090 431273
rect 439909 431829 440229 431861
rect 439909 431593 439951 431829
rect 440187 431593 440229 431829
rect 439909 431509 440229 431593
rect 439909 431273 439951 431509
rect 440187 431273 440229 431509
rect 439909 431241 440229 431273
rect 445840 431829 446160 431861
rect 445840 431593 445882 431829
rect 446118 431593 446160 431829
rect 445840 431509 446160 431593
rect 445840 431273 445882 431509
rect 446118 431273 446160 431509
rect 445840 431241 446160 431273
rect 451770 431829 452090 431861
rect 451770 431593 451812 431829
rect 452048 431593 452090 431829
rect 451770 431509 452090 431593
rect 451770 431273 451812 431509
rect 452048 431273 452090 431509
rect 451770 431241 452090 431273
rect 467909 431829 468229 431861
rect 467909 431593 467951 431829
rect 468187 431593 468229 431829
rect 467909 431509 468229 431593
rect 467909 431273 467951 431509
rect 468187 431273 468229 431509
rect 467909 431241 468229 431273
rect 473840 431829 474160 431861
rect 473840 431593 473882 431829
rect 474118 431593 474160 431829
rect 473840 431509 474160 431593
rect 473840 431273 473882 431509
rect 474118 431273 474160 431509
rect 473840 431241 474160 431273
rect 479770 431829 480090 431861
rect 479770 431593 479812 431829
rect 480048 431593 480090 431829
rect 479770 431509 480090 431593
rect 479770 431273 479812 431509
rect 480048 431273 480090 431509
rect 479770 431241 480090 431273
rect 495909 431829 496229 431861
rect 495909 431593 495951 431829
rect 496187 431593 496229 431829
rect 495909 431509 496229 431593
rect 495909 431273 495951 431509
rect 496187 431273 496229 431509
rect 495909 431241 496229 431273
rect 501840 431829 502160 431861
rect 501840 431593 501882 431829
rect 502118 431593 502160 431829
rect 501840 431509 502160 431593
rect 501840 431273 501882 431509
rect 502118 431273 502160 431509
rect 501840 431241 502160 431273
rect 507770 431829 508090 431861
rect 507770 431593 507812 431829
rect 508048 431593 508090 431829
rect 507770 431509 508090 431593
rect 507770 431273 507812 431509
rect 508048 431273 508090 431509
rect 507770 431241 508090 431273
rect 523909 431829 524229 431861
rect 523909 431593 523951 431829
rect 524187 431593 524229 431829
rect 523909 431509 524229 431593
rect 523909 431273 523951 431509
rect 524187 431273 524229 431509
rect 523909 431241 524229 431273
rect 529840 431829 530160 431861
rect 529840 431593 529882 431829
rect 530118 431593 530160 431829
rect 529840 431509 530160 431593
rect 529840 431273 529882 431509
rect 530118 431273 530160 431509
rect 529840 431241 530160 431273
rect 535770 431829 536090 431861
rect 535770 431593 535812 431829
rect 536048 431593 536090 431829
rect 535770 431509 536090 431593
rect 535770 431273 535812 431509
rect 536048 431273 536090 431509
rect 535770 431241 536090 431273
rect 551909 431829 552229 431861
rect 551909 431593 551951 431829
rect 552187 431593 552229 431829
rect 551909 431509 552229 431593
rect 551909 431273 551951 431509
rect 552187 431273 552229 431509
rect 551909 431241 552229 431273
rect 557840 431829 558160 431861
rect 557840 431593 557882 431829
rect 558118 431593 558160 431829
rect 557840 431509 558160 431593
rect 557840 431273 557882 431509
rect 558118 431273 558160 431509
rect 557840 431241 558160 431273
rect 563770 431829 564090 431861
rect 563770 431593 563812 431829
rect 564048 431593 564090 431829
rect 563770 431509 564090 431593
rect 563770 431273 563812 431509
rect 564048 431273 564090 431509
rect 563770 431241 564090 431273
rect 573494 431829 574114 458273
rect 573494 431593 573526 431829
rect 573762 431593 573846 431829
rect 574082 431593 574114 431829
rect 573494 431509 574114 431593
rect 573494 431273 573526 431509
rect 573762 431273 573846 431509
rect 574082 431273 574114 431509
rect 22875 428454 23195 428486
rect 22875 428218 22917 428454
rect 23153 428218 23195 428454
rect 22875 428134 23195 428218
rect 22875 427898 22917 428134
rect 23153 427898 23195 428134
rect 22875 427866 23195 427898
rect 28806 428454 29126 428486
rect 28806 428218 28848 428454
rect 29084 428218 29126 428454
rect 28806 428134 29126 428218
rect 28806 427898 28848 428134
rect 29084 427898 29126 428134
rect 28806 427866 29126 427898
rect 50875 428454 51195 428486
rect 50875 428218 50917 428454
rect 51153 428218 51195 428454
rect 50875 428134 51195 428218
rect 50875 427898 50917 428134
rect 51153 427898 51195 428134
rect 50875 427866 51195 427898
rect 56806 428454 57126 428486
rect 56806 428218 56848 428454
rect 57084 428218 57126 428454
rect 56806 428134 57126 428218
rect 56806 427898 56848 428134
rect 57084 427898 57126 428134
rect 56806 427866 57126 427898
rect 78875 428454 79195 428486
rect 78875 428218 78917 428454
rect 79153 428218 79195 428454
rect 78875 428134 79195 428218
rect 78875 427898 78917 428134
rect 79153 427898 79195 428134
rect 78875 427866 79195 427898
rect 84806 428454 85126 428486
rect 84806 428218 84848 428454
rect 85084 428218 85126 428454
rect 84806 428134 85126 428218
rect 84806 427898 84848 428134
rect 85084 427898 85126 428134
rect 84806 427866 85126 427898
rect 106875 428454 107195 428486
rect 106875 428218 106917 428454
rect 107153 428218 107195 428454
rect 106875 428134 107195 428218
rect 106875 427898 106917 428134
rect 107153 427898 107195 428134
rect 106875 427866 107195 427898
rect 112806 428454 113126 428486
rect 112806 428218 112848 428454
rect 113084 428218 113126 428454
rect 112806 428134 113126 428218
rect 112806 427898 112848 428134
rect 113084 427898 113126 428134
rect 112806 427866 113126 427898
rect 134875 428454 135195 428486
rect 134875 428218 134917 428454
rect 135153 428218 135195 428454
rect 134875 428134 135195 428218
rect 134875 427898 134917 428134
rect 135153 427898 135195 428134
rect 134875 427866 135195 427898
rect 140806 428454 141126 428486
rect 140806 428218 140848 428454
rect 141084 428218 141126 428454
rect 140806 428134 141126 428218
rect 140806 427898 140848 428134
rect 141084 427898 141126 428134
rect 140806 427866 141126 427898
rect 162875 428454 163195 428486
rect 162875 428218 162917 428454
rect 163153 428218 163195 428454
rect 162875 428134 163195 428218
rect 162875 427898 162917 428134
rect 163153 427898 163195 428134
rect 162875 427866 163195 427898
rect 168806 428454 169126 428486
rect 168806 428218 168848 428454
rect 169084 428218 169126 428454
rect 168806 428134 169126 428218
rect 168806 427898 168848 428134
rect 169084 427898 169126 428134
rect 168806 427866 169126 427898
rect 190875 428454 191195 428486
rect 190875 428218 190917 428454
rect 191153 428218 191195 428454
rect 190875 428134 191195 428218
rect 190875 427898 190917 428134
rect 191153 427898 191195 428134
rect 190875 427866 191195 427898
rect 196806 428454 197126 428486
rect 196806 428218 196848 428454
rect 197084 428218 197126 428454
rect 196806 428134 197126 428218
rect 196806 427898 196848 428134
rect 197084 427898 197126 428134
rect 196806 427866 197126 427898
rect 218875 428454 219195 428486
rect 218875 428218 218917 428454
rect 219153 428218 219195 428454
rect 218875 428134 219195 428218
rect 218875 427898 218917 428134
rect 219153 427898 219195 428134
rect 218875 427866 219195 427898
rect 224806 428454 225126 428486
rect 224806 428218 224848 428454
rect 225084 428218 225126 428454
rect 224806 428134 225126 428218
rect 224806 427898 224848 428134
rect 225084 427898 225126 428134
rect 224806 427866 225126 427898
rect 246875 428454 247195 428486
rect 246875 428218 246917 428454
rect 247153 428218 247195 428454
rect 246875 428134 247195 428218
rect 246875 427898 246917 428134
rect 247153 427898 247195 428134
rect 246875 427866 247195 427898
rect 252806 428454 253126 428486
rect 252806 428218 252848 428454
rect 253084 428218 253126 428454
rect 252806 428134 253126 428218
rect 252806 427898 252848 428134
rect 253084 427898 253126 428134
rect 252806 427866 253126 427898
rect 274875 428454 275195 428486
rect 274875 428218 274917 428454
rect 275153 428218 275195 428454
rect 274875 428134 275195 428218
rect 274875 427898 274917 428134
rect 275153 427898 275195 428134
rect 274875 427866 275195 427898
rect 280806 428454 281126 428486
rect 280806 428218 280848 428454
rect 281084 428218 281126 428454
rect 280806 428134 281126 428218
rect 280806 427898 280848 428134
rect 281084 427898 281126 428134
rect 280806 427866 281126 427898
rect 302875 428454 303195 428486
rect 302875 428218 302917 428454
rect 303153 428218 303195 428454
rect 302875 428134 303195 428218
rect 302875 427898 302917 428134
rect 303153 427898 303195 428134
rect 302875 427866 303195 427898
rect 308806 428454 309126 428486
rect 308806 428218 308848 428454
rect 309084 428218 309126 428454
rect 308806 428134 309126 428218
rect 308806 427898 308848 428134
rect 309084 427898 309126 428134
rect 308806 427866 309126 427898
rect 330875 428454 331195 428486
rect 330875 428218 330917 428454
rect 331153 428218 331195 428454
rect 330875 428134 331195 428218
rect 330875 427898 330917 428134
rect 331153 427898 331195 428134
rect 330875 427866 331195 427898
rect 336806 428454 337126 428486
rect 336806 428218 336848 428454
rect 337084 428218 337126 428454
rect 336806 428134 337126 428218
rect 336806 427898 336848 428134
rect 337084 427898 337126 428134
rect 336806 427866 337126 427898
rect 358875 428454 359195 428486
rect 358875 428218 358917 428454
rect 359153 428218 359195 428454
rect 358875 428134 359195 428218
rect 358875 427898 358917 428134
rect 359153 427898 359195 428134
rect 358875 427866 359195 427898
rect 364806 428454 365126 428486
rect 364806 428218 364848 428454
rect 365084 428218 365126 428454
rect 364806 428134 365126 428218
rect 364806 427898 364848 428134
rect 365084 427898 365126 428134
rect 364806 427866 365126 427898
rect 386875 428454 387195 428486
rect 386875 428218 386917 428454
rect 387153 428218 387195 428454
rect 386875 428134 387195 428218
rect 386875 427898 386917 428134
rect 387153 427898 387195 428134
rect 386875 427866 387195 427898
rect 392806 428454 393126 428486
rect 392806 428218 392848 428454
rect 393084 428218 393126 428454
rect 392806 428134 393126 428218
rect 392806 427898 392848 428134
rect 393084 427898 393126 428134
rect 392806 427866 393126 427898
rect 414875 428454 415195 428486
rect 414875 428218 414917 428454
rect 415153 428218 415195 428454
rect 414875 428134 415195 428218
rect 414875 427898 414917 428134
rect 415153 427898 415195 428134
rect 414875 427866 415195 427898
rect 420806 428454 421126 428486
rect 420806 428218 420848 428454
rect 421084 428218 421126 428454
rect 420806 428134 421126 428218
rect 420806 427898 420848 428134
rect 421084 427898 421126 428134
rect 420806 427866 421126 427898
rect 442875 428454 443195 428486
rect 442875 428218 442917 428454
rect 443153 428218 443195 428454
rect 442875 428134 443195 428218
rect 442875 427898 442917 428134
rect 443153 427898 443195 428134
rect 442875 427866 443195 427898
rect 448806 428454 449126 428486
rect 448806 428218 448848 428454
rect 449084 428218 449126 428454
rect 448806 428134 449126 428218
rect 448806 427898 448848 428134
rect 449084 427898 449126 428134
rect 448806 427866 449126 427898
rect 470875 428454 471195 428486
rect 470875 428218 470917 428454
rect 471153 428218 471195 428454
rect 470875 428134 471195 428218
rect 470875 427898 470917 428134
rect 471153 427898 471195 428134
rect 470875 427866 471195 427898
rect 476806 428454 477126 428486
rect 476806 428218 476848 428454
rect 477084 428218 477126 428454
rect 476806 428134 477126 428218
rect 476806 427898 476848 428134
rect 477084 427898 477126 428134
rect 476806 427866 477126 427898
rect 498875 428454 499195 428486
rect 498875 428218 498917 428454
rect 499153 428218 499195 428454
rect 498875 428134 499195 428218
rect 498875 427898 498917 428134
rect 499153 427898 499195 428134
rect 498875 427866 499195 427898
rect 504806 428454 505126 428486
rect 504806 428218 504848 428454
rect 505084 428218 505126 428454
rect 504806 428134 505126 428218
rect 504806 427898 504848 428134
rect 505084 427898 505126 428134
rect 504806 427866 505126 427898
rect 526875 428454 527195 428486
rect 526875 428218 526917 428454
rect 527153 428218 527195 428454
rect 526875 428134 527195 428218
rect 526875 427898 526917 428134
rect 527153 427898 527195 428134
rect 526875 427866 527195 427898
rect 532806 428454 533126 428486
rect 532806 428218 532848 428454
rect 533084 428218 533126 428454
rect 532806 428134 533126 428218
rect 532806 427898 532848 428134
rect 533084 427898 533126 428134
rect 532806 427866 533126 427898
rect 554875 428454 555195 428486
rect 554875 428218 554917 428454
rect 555153 428218 555195 428454
rect 554875 428134 555195 428218
rect 554875 427898 554917 428134
rect 555153 427898 555195 428134
rect 554875 427866 555195 427898
rect 560806 428454 561126 428486
rect 560806 428218 560848 428454
rect 561084 428218 561126 428454
rect 560806 428134 561126 428218
rect 560806 427898 560848 428134
rect 561084 427898 561126 428134
rect 560806 427866 561126 427898
rect -2006 404593 -1974 404829
rect -1738 404593 -1654 404829
rect -1418 404593 -1386 404829
rect -2006 404509 -1386 404593
rect -2006 404273 -1974 404509
rect -1738 404273 -1654 404509
rect -1418 404273 -1386 404509
rect -2006 377829 -1386 404273
rect 19910 404829 20230 404861
rect 19910 404593 19952 404829
rect 20188 404593 20230 404829
rect 19910 404509 20230 404593
rect 19910 404273 19952 404509
rect 20188 404273 20230 404509
rect 19910 404241 20230 404273
rect 25840 404829 26160 404861
rect 25840 404593 25882 404829
rect 26118 404593 26160 404829
rect 25840 404509 26160 404593
rect 25840 404273 25882 404509
rect 26118 404273 26160 404509
rect 25840 404241 26160 404273
rect 31771 404829 32091 404861
rect 31771 404593 31813 404829
rect 32049 404593 32091 404829
rect 31771 404509 32091 404593
rect 31771 404273 31813 404509
rect 32049 404273 32091 404509
rect 31771 404241 32091 404273
rect 47910 404829 48230 404861
rect 47910 404593 47952 404829
rect 48188 404593 48230 404829
rect 47910 404509 48230 404593
rect 47910 404273 47952 404509
rect 48188 404273 48230 404509
rect 47910 404241 48230 404273
rect 53840 404829 54160 404861
rect 53840 404593 53882 404829
rect 54118 404593 54160 404829
rect 53840 404509 54160 404593
rect 53840 404273 53882 404509
rect 54118 404273 54160 404509
rect 53840 404241 54160 404273
rect 59771 404829 60091 404861
rect 59771 404593 59813 404829
rect 60049 404593 60091 404829
rect 59771 404509 60091 404593
rect 59771 404273 59813 404509
rect 60049 404273 60091 404509
rect 59771 404241 60091 404273
rect 75910 404829 76230 404861
rect 75910 404593 75952 404829
rect 76188 404593 76230 404829
rect 75910 404509 76230 404593
rect 75910 404273 75952 404509
rect 76188 404273 76230 404509
rect 75910 404241 76230 404273
rect 81840 404829 82160 404861
rect 81840 404593 81882 404829
rect 82118 404593 82160 404829
rect 81840 404509 82160 404593
rect 81840 404273 81882 404509
rect 82118 404273 82160 404509
rect 81840 404241 82160 404273
rect 87771 404829 88091 404861
rect 87771 404593 87813 404829
rect 88049 404593 88091 404829
rect 87771 404509 88091 404593
rect 87771 404273 87813 404509
rect 88049 404273 88091 404509
rect 87771 404241 88091 404273
rect 103910 404829 104230 404861
rect 103910 404593 103952 404829
rect 104188 404593 104230 404829
rect 103910 404509 104230 404593
rect 103910 404273 103952 404509
rect 104188 404273 104230 404509
rect 103910 404241 104230 404273
rect 109840 404829 110160 404861
rect 109840 404593 109882 404829
rect 110118 404593 110160 404829
rect 109840 404509 110160 404593
rect 109840 404273 109882 404509
rect 110118 404273 110160 404509
rect 109840 404241 110160 404273
rect 115771 404829 116091 404861
rect 115771 404593 115813 404829
rect 116049 404593 116091 404829
rect 115771 404509 116091 404593
rect 115771 404273 115813 404509
rect 116049 404273 116091 404509
rect 115771 404241 116091 404273
rect 131910 404829 132230 404861
rect 131910 404593 131952 404829
rect 132188 404593 132230 404829
rect 131910 404509 132230 404593
rect 131910 404273 131952 404509
rect 132188 404273 132230 404509
rect 131910 404241 132230 404273
rect 137840 404829 138160 404861
rect 137840 404593 137882 404829
rect 138118 404593 138160 404829
rect 137840 404509 138160 404593
rect 137840 404273 137882 404509
rect 138118 404273 138160 404509
rect 137840 404241 138160 404273
rect 143771 404829 144091 404861
rect 143771 404593 143813 404829
rect 144049 404593 144091 404829
rect 143771 404509 144091 404593
rect 143771 404273 143813 404509
rect 144049 404273 144091 404509
rect 143771 404241 144091 404273
rect 159910 404829 160230 404861
rect 159910 404593 159952 404829
rect 160188 404593 160230 404829
rect 159910 404509 160230 404593
rect 159910 404273 159952 404509
rect 160188 404273 160230 404509
rect 159910 404241 160230 404273
rect 165840 404829 166160 404861
rect 165840 404593 165882 404829
rect 166118 404593 166160 404829
rect 165840 404509 166160 404593
rect 165840 404273 165882 404509
rect 166118 404273 166160 404509
rect 165840 404241 166160 404273
rect 171771 404829 172091 404861
rect 171771 404593 171813 404829
rect 172049 404593 172091 404829
rect 171771 404509 172091 404593
rect 171771 404273 171813 404509
rect 172049 404273 172091 404509
rect 171771 404241 172091 404273
rect 187910 404829 188230 404861
rect 187910 404593 187952 404829
rect 188188 404593 188230 404829
rect 187910 404509 188230 404593
rect 187910 404273 187952 404509
rect 188188 404273 188230 404509
rect 187910 404241 188230 404273
rect 193840 404829 194160 404861
rect 193840 404593 193882 404829
rect 194118 404593 194160 404829
rect 193840 404509 194160 404593
rect 193840 404273 193882 404509
rect 194118 404273 194160 404509
rect 193840 404241 194160 404273
rect 199771 404829 200091 404861
rect 199771 404593 199813 404829
rect 200049 404593 200091 404829
rect 199771 404509 200091 404593
rect 199771 404273 199813 404509
rect 200049 404273 200091 404509
rect 199771 404241 200091 404273
rect 215910 404829 216230 404861
rect 215910 404593 215952 404829
rect 216188 404593 216230 404829
rect 215910 404509 216230 404593
rect 215910 404273 215952 404509
rect 216188 404273 216230 404509
rect 215910 404241 216230 404273
rect 221840 404829 222160 404861
rect 221840 404593 221882 404829
rect 222118 404593 222160 404829
rect 221840 404509 222160 404593
rect 221840 404273 221882 404509
rect 222118 404273 222160 404509
rect 221840 404241 222160 404273
rect 227771 404829 228091 404861
rect 227771 404593 227813 404829
rect 228049 404593 228091 404829
rect 227771 404509 228091 404593
rect 227771 404273 227813 404509
rect 228049 404273 228091 404509
rect 227771 404241 228091 404273
rect 243910 404829 244230 404861
rect 243910 404593 243952 404829
rect 244188 404593 244230 404829
rect 243910 404509 244230 404593
rect 243910 404273 243952 404509
rect 244188 404273 244230 404509
rect 243910 404241 244230 404273
rect 249840 404829 250160 404861
rect 249840 404593 249882 404829
rect 250118 404593 250160 404829
rect 249840 404509 250160 404593
rect 249840 404273 249882 404509
rect 250118 404273 250160 404509
rect 249840 404241 250160 404273
rect 255771 404829 256091 404861
rect 255771 404593 255813 404829
rect 256049 404593 256091 404829
rect 255771 404509 256091 404593
rect 255771 404273 255813 404509
rect 256049 404273 256091 404509
rect 255771 404241 256091 404273
rect 271910 404829 272230 404861
rect 271910 404593 271952 404829
rect 272188 404593 272230 404829
rect 271910 404509 272230 404593
rect 271910 404273 271952 404509
rect 272188 404273 272230 404509
rect 271910 404241 272230 404273
rect 277840 404829 278160 404861
rect 277840 404593 277882 404829
rect 278118 404593 278160 404829
rect 277840 404509 278160 404593
rect 277840 404273 277882 404509
rect 278118 404273 278160 404509
rect 277840 404241 278160 404273
rect 283771 404829 284091 404861
rect 283771 404593 283813 404829
rect 284049 404593 284091 404829
rect 283771 404509 284091 404593
rect 283771 404273 283813 404509
rect 284049 404273 284091 404509
rect 283771 404241 284091 404273
rect 299910 404829 300230 404861
rect 299910 404593 299952 404829
rect 300188 404593 300230 404829
rect 299910 404509 300230 404593
rect 299910 404273 299952 404509
rect 300188 404273 300230 404509
rect 299910 404241 300230 404273
rect 305840 404829 306160 404861
rect 305840 404593 305882 404829
rect 306118 404593 306160 404829
rect 305840 404509 306160 404593
rect 305840 404273 305882 404509
rect 306118 404273 306160 404509
rect 305840 404241 306160 404273
rect 311771 404829 312091 404861
rect 311771 404593 311813 404829
rect 312049 404593 312091 404829
rect 311771 404509 312091 404593
rect 311771 404273 311813 404509
rect 312049 404273 312091 404509
rect 311771 404241 312091 404273
rect 327910 404829 328230 404861
rect 327910 404593 327952 404829
rect 328188 404593 328230 404829
rect 327910 404509 328230 404593
rect 327910 404273 327952 404509
rect 328188 404273 328230 404509
rect 327910 404241 328230 404273
rect 333840 404829 334160 404861
rect 333840 404593 333882 404829
rect 334118 404593 334160 404829
rect 333840 404509 334160 404593
rect 333840 404273 333882 404509
rect 334118 404273 334160 404509
rect 333840 404241 334160 404273
rect 339771 404829 340091 404861
rect 339771 404593 339813 404829
rect 340049 404593 340091 404829
rect 339771 404509 340091 404593
rect 339771 404273 339813 404509
rect 340049 404273 340091 404509
rect 339771 404241 340091 404273
rect 355910 404829 356230 404861
rect 355910 404593 355952 404829
rect 356188 404593 356230 404829
rect 355910 404509 356230 404593
rect 355910 404273 355952 404509
rect 356188 404273 356230 404509
rect 355910 404241 356230 404273
rect 361840 404829 362160 404861
rect 361840 404593 361882 404829
rect 362118 404593 362160 404829
rect 361840 404509 362160 404593
rect 361840 404273 361882 404509
rect 362118 404273 362160 404509
rect 361840 404241 362160 404273
rect 367771 404829 368091 404861
rect 367771 404593 367813 404829
rect 368049 404593 368091 404829
rect 367771 404509 368091 404593
rect 367771 404273 367813 404509
rect 368049 404273 368091 404509
rect 367771 404241 368091 404273
rect 383910 404829 384230 404861
rect 383910 404593 383952 404829
rect 384188 404593 384230 404829
rect 383910 404509 384230 404593
rect 383910 404273 383952 404509
rect 384188 404273 384230 404509
rect 383910 404241 384230 404273
rect 389840 404829 390160 404861
rect 389840 404593 389882 404829
rect 390118 404593 390160 404829
rect 389840 404509 390160 404593
rect 389840 404273 389882 404509
rect 390118 404273 390160 404509
rect 389840 404241 390160 404273
rect 395771 404829 396091 404861
rect 395771 404593 395813 404829
rect 396049 404593 396091 404829
rect 395771 404509 396091 404593
rect 395771 404273 395813 404509
rect 396049 404273 396091 404509
rect 395771 404241 396091 404273
rect 411910 404829 412230 404861
rect 411910 404593 411952 404829
rect 412188 404593 412230 404829
rect 411910 404509 412230 404593
rect 411910 404273 411952 404509
rect 412188 404273 412230 404509
rect 411910 404241 412230 404273
rect 417840 404829 418160 404861
rect 417840 404593 417882 404829
rect 418118 404593 418160 404829
rect 417840 404509 418160 404593
rect 417840 404273 417882 404509
rect 418118 404273 418160 404509
rect 417840 404241 418160 404273
rect 423771 404829 424091 404861
rect 423771 404593 423813 404829
rect 424049 404593 424091 404829
rect 423771 404509 424091 404593
rect 423771 404273 423813 404509
rect 424049 404273 424091 404509
rect 423771 404241 424091 404273
rect 439910 404829 440230 404861
rect 439910 404593 439952 404829
rect 440188 404593 440230 404829
rect 439910 404509 440230 404593
rect 439910 404273 439952 404509
rect 440188 404273 440230 404509
rect 439910 404241 440230 404273
rect 445840 404829 446160 404861
rect 445840 404593 445882 404829
rect 446118 404593 446160 404829
rect 445840 404509 446160 404593
rect 445840 404273 445882 404509
rect 446118 404273 446160 404509
rect 445840 404241 446160 404273
rect 451771 404829 452091 404861
rect 451771 404593 451813 404829
rect 452049 404593 452091 404829
rect 451771 404509 452091 404593
rect 451771 404273 451813 404509
rect 452049 404273 452091 404509
rect 451771 404241 452091 404273
rect 467910 404829 468230 404861
rect 467910 404593 467952 404829
rect 468188 404593 468230 404829
rect 467910 404509 468230 404593
rect 467910 404273 467952 404509
rect 468188 404273 468230 404509
rect 467910 404241 468230 404273
rect 473840 404829 474160 404861
rect 473840 404593 473882 404829
rect 474118 404593 474160 404829
rect 473840 404509 474160 404593
rect 473840 404273 473882 404509
rect 474118 404273 474160 404509
rect 473840 404241 474160 404273
rect 479771 404829 480091 404861
rect 479771 404593 479813 404829
rect 480049 404593 480091 404829
rect 479771 404509 480091 404593
rect 479771 404273 479813 404509
rect 480049 404273 480091 404509
rect 479771 404241 480091 404273
rect 495910 404829 496230 404861
rect 495910 404593 495952 404829
rect 496188 404593 496230 404829
rect 495910 404509 496230 404593
rect 495910 404273 495952 404509
rect 496188 404273 496230 404509
rect 495910 404241 496230 404273
rect 501840 404829 502160 404861
rect 501840 404593 501882 404829
rect 502118 404593 502160 404829
rect 501840 404509 502160 404593
rect 501840 404273 501882 404509
rect 502118 404273 502160 404509
rect 501840 404241 502160 404273
rect 507771 404829 508091 404861
rect 507771 404593 507813 404829
rect 508049 404593 508091 404829
rect 507771 404509 508091 404593
rect 507771 404273 507813 404509
rect 508049 404273 508091 404509
rect 507771 404241 508091 404273
rect 523910 404829 524230 404861
rect 523910 404593 523952 404829
rect 524188 404593 524230 404829
rect 523910 404509 524230 404593
rect 523910 404273 523952 404509
rect 524188 404273 524230 404509
rect 523910 404241 524230 404273
rect 529840 404829 530160 404861
rect 529840 404593 529882 404829
rect 530118 404593 530160 404829
rect 529840 404509 530160 404593
rect 529840 404273 529882 404509
rect 530118 404273 530160 404509
rect 529840 404241 530160 404273
rect 535771 404829 536091 404861
rect 535771 404593 535813 404829
rect 536049 404593 536091 404829
rect 535771 404509 536091 404593
rect 535771 404273 535813 404509
rect 536049 404273 536091 404509
rect 535771 404241 536091 404273
rect 551910 404829 552230 404861
rect 551910 404593 551952 404829
rect 552188 404593 552230 404829
rect 551910 404509 552230 404593
rect 551910 404273 551952 404509
rect 552188 404273 552230 404509
rect 551910 404241 552230 404273
rect 557840 404829 558160 404861
rect 557840 404593 557882 404829
rect 558118 404593 558160 404829
rect 557840 404509 558160 404593
rect 557840 404273 557882 404509
rect 558118 404273 558160 404509
rect 557840 404241 558160 404273
rect 563771 404829 564091 404861
rect 563771 404593 563813 404829
rect 564049 404593 564091 404829
rect 563771 404509 564091 404593
rect 563771 404273 563813 404509
rect 564049 404273 564091 404509
rect 563771 404241 564091 404273
rect 573494 404829 574114 431273
rect 573494 404593 573526 404829
rect 573762 404593 573846 404829
rect 574082 404593 574114 404829
rect 573494 404509 574114 404593
rect 573494 404273 573526 404509
rect 573762 404273 573846 404509
rect 574082 404273 574114 404509
rect 22874 401454 23194 401486
rect 22874 401218 22916 401454
rect 23152 401218 23194 401454
rect 22874 401134 23194 401218
rect 22874 400898 22916 401134
rect 23152 400898 23194 401134
rect 22874 400866 23194 400898
rect 28805 401454 29125 401486
rect 28805 401218 28847 401454
rect 29083 401218 29125 401454
rect 28805 401134 29125 401218
rect 28805 400898 28847 401134
rect 29083 400898 29125 401134
rect 28805 400866 29125 400898
rect 50874 401454 51194 401486
rect 50874 401218 50916 401454
rect 51152 401218 51194 401454
rect 50874 401134 51194 401218
rect 50874 400898 50916 401134
rect 51152 400898 51194 401134
rect 50874 400866 51194 400898
rect 56805 401454 57125 401486
rect 56805 401218 56847 401454
rect 57083 401218 57125 401454
rect 56805 401134 57125 401218
rect 56805 400898 56847 401134
rect 57083 400898 57125 401134
rect 56805 400866 57125 400898
rect 78874 401454 79194 401486
rect 78874 401218 78916 401454
rect 79152 401218 79194 401454
rect 78874 401134 79194 401218
rect 78874 400898 78916 401134
rect 79152 400898 79194 401134
rect 78874 400866 79194 400898
rect 84805 401454 85125 401486
rect 84805 401218 84847 401454
rect 85083 401218 85125 401454
rect 84805 401134 85125 401218
rect 84805 400898 84847 401134
rect 85083 400898 85125 401134
rect 84805 400866 85125 400898
rect 106874 401454 107194 401486
rect 106874 401218 106916 401454
rect 107152 401218 107194 401454
rect 106874 401134 107194 401218
rect 106874 400898 106916 401134
rect 107152 400898 107194 401134
rect 106874 400866 107194 400898
rect 112805 401454 113125 401486
rect 112805 401218 112847 401454
rect 113083 401218 113125 401454
rect 112805 401134 113125 401218
rect 112805 400898 112847 401134
rect 113083 400898 113125 401134
rect 112805 400866 113125 400898
rect 134874 401454 135194 401486
rect 134874 401218 134916 401454
rect 135152 401218 135194 401454
rect 134874 401134 135194 401218
rect 134874 400898 134916 401134
rect 135152 400898 135194 401134
rect 134874 400866 135194 400898
rect 140805 401454 141125 401486
rect 140805 401218 140847 401454
rect 141083 401218 141125 401454
rect 140805 401134 141125 401218
rect 140805 400898 140847 401134
rect 141083 400898 141125 401134
rect 140805 400866 141125 400898
rect 162874 401454 163194 401486
rect 162874 401218 162916 401454
rect 163152 401218 163194 401454
rect 162874 401134 163194 401218
rect 162874 400898 162916 401134
rect 163152 400898 163194 401134
rect 162874 400866 163194 400898
rect 168805 401454 169125 401486
rect 168805 401218 168847 401454
rect 169083 401218 169125 401454
rect 168805 401134 169125 401218
rect 168805 400898 168847 401134
rect 169083 400898 169125 401134
rect 168805 400866 169125 400898
rect 190874 401454 191194 401486
rect 190874 401218 190916 401454
rect 191152 401218 191194 401454
rect 190874 401134 191194 401218
rect 190874 400898 190916 401134
rect 191152 400898 191194 401134
rect 190874 400866 191194 400898
rect 196805 401454 197125 401486
rect 196805 401218 196847 401454
rect 197083 401218 197125 401454
rect 196805 401134 197125 401218
rect 196805 400898 196847 401134
rect 197083 400898 197125 401134
rect 196805 400866 197125 400898
rect 218874 401454 219194 401486
rect 218874 401218 218916 401454
rect 219152 401218 219194 401454
rect 218874 401134 219194 401218
rect 218874 400898 218916 401134
rect 219152 400898 219194 401134
rect 218874 400866 219194 400898
rect 224805 401454 225125 401486
rect 224805 401218 224847 401454
rect 225083 401218 225125 401454
rect 224805 401134 225125 401218
rect 224805 400898 224847 401134
rect 225083 400898 225125 401134
rect 224805 400866 225125 400898
rect 246874 401454 247194 401486
rect 246874 401218 246916 401454
rect 247152 401218 247194 401454
rect 246874 401134 247194 401218
rect 246874 400898 246916 401134
rect 247152 400898 247194 401134
rect 246874 400866 247194 400898
rect 252805 401454 253125 401486
rect 252805 401218 252847 401454
rect 253083 401218 253125 401454
rect 252805 401134 253125 401218
rect 252805 400898 252847 401134
rect 253083 400898 253125 401134
rect 252805 400866 253125 400898
rect 274874 401454 275194 401486
rect 274874 401218 274916 401454
rect 275152 401218 275194 401454
rect 274874 401134 275194 401218
rect 274874 400898 274916 401134
rect 275152 400898 275194 401134
rect 274874 400866 275194 400898
rect 280805 401454 281125 401486
rect 280805 401218 280847 401454
rect 281083 401218 281125 401454
rect 280805 401134 281125 401218
rect 280805 400898 280847 401134
rect 281083 400898 281125 401134
rect 280805 400866 281125 400898
rect 302874 401454 303194 401486
rect 302874 401218 302916 401454
rect 303152 401218 303194 401454
rect 302874 401134 303194 401218
rect 302874 400898 302916 401134
rect 303152 400898 303194 401134
rect 302874 400866 303194 400898
rect 308805 401454 309125 401486
rect 308805 401218 308847 401454
rect 309083 401218 309125 401454
rect 308805 401134 309125 401218
rect 308805 400898 308847 401134
rect 309083 400898 309125 401134
rect 308805 400866 309125 400898
rect 330874 401454 331194 401486
rect 330874 401218 330916 401454
rect 331152 401218 331194 401454
rect 330874 401134 331194 401218
rect 330874 400898 330916 401134
rect 331152 400898 331194 401134
rect 330874 400866 331194 400898
rect 336805 401454 337125 401486
rect 336805 401218 336847 401454
rect 337083 401218 337125 401454
rect 336805 401134 337125 401218
rect 336805 400898 336847 401134
rect 337083 400898 337125 401134
rect 336805 400866 337125 400898
rect 358874 401454 359194 401486
rect 358874 401218 358916 401454
rect 359152 401218 359194 401454
rect 358874 401134 359194 401218
rect 358874 400898 358916 401134
rect 359152 400898 359194 401134
rect 358874 400866 359194 400898
rect 364805 401454 365125 401486
rect 364805 401218 364847 401454
rect 365083 401218 365125 401454
rect 364805 401134 365125 401218
rect 364805 400898 364847 401134
rect 365083 400898 365125 401134
rect 364805 400866 365125 400898
rect 386874 401454 387194 401486
rect 386874 401218 386916 401454
rect 387152 401218 387194 401454
rect 386874 401134 387194 401218
rect 386874 400898 386916 401134
rect 387152 400898 387194 401134
rect 386874 400866 387194 400898
rect 392805 401454 393125 401486
rect 392805 401218 392847 401454
rect 393083 401218 393125 401454
rect 392805 401134 393125 401218
rect 392805 400898 392847 401134
rect 393083 400898 393125 401134
rect 392805 400866 393125 400898
rect 414874 401454 415194 401486
rect 414874 401218 414916 401454
rect 415152 401218 415194 401454
rect 414874 401134 415194 401218
rect 414874 400898 414916 401134
rect 415152 400898 415194 401134
rect 414874 400866 415194 400898
rect 420805 401454 421125 401486
rect 420805 401218 420847 401454
rect 421083 401218 421125 401454
rect 420805 401134 421125 401218
rect 420805 400898 420847 401134
rect 421083 400898 421125 401134
rect 420805 400866 421125 400898
rect 442874 401454 443194 401486
rect 442874 401218 442916 401454
rect 443152 401218 443194 401454
rect 442874 401134 443194 401218
rect 442874 400898 442916 401134
rect 443152 400898 443194 401134
rect 442874 400866 443194 400898
rect 448805 401454 449125 401486
rect 448805 401218 448847 401454
rect 449083 401218 449125 401454
rect 448805 401134 449125 401218
rect 448805 400898 448847 401134
rect 449083 400898 449125 401134
rect 448805 400866 449125 400898
rect 470874 401454 471194 401486
rect 470874 401218 470916 401454
rect 471152 401218 471194 401454
rect 470874 401134 471194 401218
rect 470874 400898 470916 401134
rect 471152 400898 471194 401134
rect 470874 400866 471194 400898
rect 476805 401454 477125 401486
rect 476805 401218 476847 401454
rect 477083 401218 477125 401454
rect 476805 401134 477125 401218
rect 476805 400898 476847 401134
rect 477083 400898 477125 401134
rect 476805 400866 477125 400898
rect 498874 401454 499194 401486
rect 498874 401218 498916 401454
rect 499152 401218 499194 401454
rect 498874 401134 499194 401218
rect 498874 400898 498916 401134
rect 499152 400898 499194 401134
rect 498874 400866 499194 400898
rect 504805 401454 505125 401486
rect 504805 401218 504847 401454
rect 505083 401218 505125 401454
rect 504805 401134 505125 401218
rect 504805 400898 504847 401134
rect 505083 400898 505125 401134
rect 504805 400866 505125 400898
rect 526874 401454 527194 401486
rect 526874 401218 526916 401454
rect 527152 401218 527194 401454
rect 526874 401134 527194 401218
rect 526874 400898 526916 401134
rect 527152 400898 527194 401134
rect 526874 400866 527194 400898
rect 532805 401454 533125 401486
rect 532805 401218 532847 401454
rect 533083 401218 533125 401454
rect 532805 401134 533125 401218
rect 532805 400898 532847 401134
rect 533083 400898 533125 401134
rect 532805 400866 533125 400898
rect 554874 401454 555194 401486
rect 554874 401218 554916 401454
rect 555152 401218 555194 401454
rect 554874 401134 555194 401218
rect 554874 400898 554916 401134
rect 555152 400898 555194 401134
rect 554874 400866 555194 400898
rect 560805 401454 561125 401486
rect 560805 401218 560847 401454
rect 561083 401218 561125 401454
rect 560805 401134 561125 401218
rect 560805 400898 560847 401134
rect 561083 400898 561125 401134
rect 560805 400866 561125 400898
rect -2006 377593 -1974 377829
rect -1738 377593 -1654 377829
rect -1418 377593 -1386 377829
rect -2006 377509 -1386 377593
rect -2006 377273 -1974 377509
rect -1738 377273 -1654 377509
rect -1418 377273 -1386 377509
rect -2006 350829 -1386 377273
rect 19909 377829 20229 377861
rect 19909 377593 19951 377829
rect 20187 377593 20229 377829
rect 19909 377509 20229 377593
rect 19909 377273 19951 377509
rect 20187 377273 20229 377509
rect 19909 377241 20229 377273
rect 25840 377829 26160 377861
rect 25840 377593 25882 377829
rect 26118 377593 26160 377829
rect 25840 377509 26160 377593
rect 25840 377273 25882 377509
rect 26118 377273 26160 377509
rect 25840 377241 26160 377273
rect 31770 377829 32090 377861
rect 31770 377593 31812 377829
rect 32048 377593 32090 377829
rect 31770 377509 32090 377593
rect 31770 377273 31812 377509
rect 32048 377273 32090 377509
rect 31770 377241 32090 377273
rect 47909 377829 48229 377861
rect 47909 377593 47951 377829
rect 48187 377593 48229 377829
rect 47909 377509 48229 377593
rect 47909 377273 47951 377509
rect 48187 377273 48229 377509
rect 47909 377241 48229 377273
rect 53840 377829 54160 377861
rect 53840 377593 53882 377829
rect 54118 377593 54160 377829
rect 53840 377509 54160 377593
rect 53840 377273 53882 377509
rect 54118 377273 54160 377509
rect 53840 377241 54160 377273
rect 59770 377829 60090 377861
rect 59770 377593 59812 377829
rect 60048 377593 60090 377829
rect 59770 377509 60090 377593
rect 59770 377273 59812 377509
rect 60048 377273 60090 377509
rect 59770 377241 60090 377273
rect 75909 377829 76229 377861
rect 75909 377593 75951 377829
rect 76187 377593 76229 377829
rect 75909 377509 76229 377593
rect 75909 377273 75951 377509
rect 76187 377273 76229 377509
rect 75909 377241 76229 377273
rect 81840 377829 82160 377861
rect 81840 377593 81882 377829
rect 82118 377593 82160 377829
rect 81840 377509 82160 377593
rect 81840 377273 81882 377509
rect 82118 377273 82160 377509
rect 81840 377241 82160 377273
rect 87770 377829 88090 377861
rect 87770 377593 87812 377829
rect 88048 377593 88090 377829
rect 87770 377509 88090 377593
rect 87770 377273 87812 377509
rect 88048 377273 88090 377509
rect 87770 377241 88090 377273
rect 103909 377829 104229 377861
rect 103909 377593 103951 377829
rect 104187 377593 104229 377829
rect 103909 377509 104229 377593
rect 103909 377273 103951 377509
rect 104187 377273 104229 377509
rect 103909 377241 104229 377273
rect 109840 377829 110160 377861
rect 109840 377593 109882 377829
rect 110118 377593 110160 377829
rect 109840 377509 110160 377593
rect 109840 377273 109882 377509
rect 110118 377273 110160 377509
rect 109840 377241 110160 377273
rect 115770 377829 116090 377861
rect 115770 377593 115812 377829
rect 116048 377593 116090 377829
rect 115770 377509 116090 377593
rect 115770 377273 115812 377509
rect 116048 377273 116090 377509
rect 115770 377241 116090 377273
rect 131909 377829 132229 377861
rect 131909 377593 131951 377829
rect 132187 377593 132229 377829
rect 131909 377509 132229 377593
rect 131909 377273 131951 377509
rect 132187 377273 132229 377509
rect 131909 377241 132229 377273
rect 137840 377829 138160 377861
rect 137840 377593 137882 377829
rect 138118 377593 138160 377829
rect 137840 377509 138160 377593
rect 137840 377273 137882 377509
rect 138118 377273 138160 377509
rect 137840 377241 138160 377273
rect 143770 377829 144090 377861
rect 143770 377593 143812 377829
rect 144048 377593 144090 377829
rect 143770 377509 144090 377593
rect 143770 377273 143812 377509
rect 144048 377273 144090 377509
rect 143770 377241 144090 377273
rect 159909 377829 160229 377861
rect 159909 377593 159951 377829
rect 160187 377593 160229 377829
rect 159909 377509 160229 377593
rect 159909 377273 159951 377509
rect 160187 377273 160229 377509
rect 159909 377241 160229 377273
rect 165840 377829 166160 377861
rect 165840 377593 165882 377829
rect 166118 377593 166160 377829
rect 165840 377509 166160 377593
rect 165840 377273 165882 377509
rect 166118 377273 166160 377509
rect 165840 377241 166160 377273
rect 171770 377829 172090 377861
rect 171770 377593 171812 377829
rect 172048 377593 172090 377829
rect 171770 377509 172090 377593
rect 171770 377273 171812 377509
rect 172048 377273 172090 377509
rect 171770 377241 172090 377273
rect 187909 377829 188229 377861
rect 187909 377593 187951 377829
rect 188187 377593 188229 377829
rect 187909 377509 188229 377593
rect 187909 377273 187951 377509
rect 188187 377273 188229 377509
rect 187909 377241 188229 377273
rect 193840 377829 194160 377861
rect 193840 377593 193882 377829
rect 194118 377593 194160 377829
rect 193840 377509 194160 377593
rect 193840 377273 193882 377509
rect 194118 377273 194160 377509
rect 193840 377241 194160 377273
rect 199770 377829 200090 377861
rect 199770 377593 199812 377829
rect 200048 377593 200090 377829
rect 199770 377509 200090 377593
rect 199770 377273 199812 377509
rect 200048 377273 200090 377509
rect 199770 377241 200090 377273
rect 215909 377829 216229 377861
rect 215909 377593 215951 377829
rect 216187 377593 216229 377829
rect 215909 377509 216229 377593
rect 215909 377273 215951 377509
rect 216187 377273 216229 377509
rect 215909 377241 216229 377273
rect 221840 377829 222160 377861
rect 221840 377593 221882 377829
rect 222118 377593 222160 377829
rect 221840 377509 222160 377593
rect 221840 377273 221882 377509
rect 222118 377273 222160 377509
rect 221840 377241 222160 377273
rect 227770 377829 228090 377861
rect 227770 377593 227812 377829
rect 228048 377593 228090 377829
rect 227770 377509 228090 377593
rect 227770 377273 227812 377509
rect 228048 377273 228090 377509
rect 227770 377241 228090 377273
rect 243909 377829 244229 377861
rect 243909 377593 243951 377829
rect 244187 377593 244229 377829
rect 243909 377509 244229 377593
rect 243909 377273 243951 377509
rect 244187 377273 244229 377509
rect 243909 377241 244229 377273
rect 249840 377829 250160 377861
rect 249840 377593 249882 377829
rect 250118 377593 250160 377829
rect 249840 377509 250160 377593
rect 249840 377273 249882 377509
rect 250118 377273 250160 377509
rect 249840 377241 250160 377273
rect 255770 377829 256090 377861
rect 255770 377593 255812 377829
rect 256048 377593 256090 377829
rect 255770 377509 256090 377593
rect 255770 377273 255812 377509
rect 256048 377273 256090 377509
rect 255770 377241 256090 377273
rect 271909 377829 272229 377861
rect 271909 377593 271951 377829
rect 272187 377593 272229 377829
rect 271909 377509 272229 377593
rect 271909 377273 271951 377509
rect 272187 377273 272229 377509
rect 271909 377241 272229 377273
rect 277840 377829 278160 377861
rect 277840 377593 277882 377829
rect 278118 377593 278160 377829
rect 277840 377509 278160 377593
rect 277840 377273 277882 377509
rect 278118 377273 278160 377509
rect 277840 377241 278160 377273
rect 283770 377829 284090 377861
rect 283770 377593 283812 377829
rect 284048 377593 284090 377829
rect 283770 377509 284090 377593
rect 283770 377273 283812 377509
rect 284048 377273 284090 377509
rect 283770 377241 284090 377273
rect 299909 377829 300229 377861
rect 299909 377593 299951 377829
rect 300187 377593 300229 377829
rect 299909 377509 300229 377593
rect 299909 377273 299951 377509
rect 300187 377273 300229 377509
rect 299909 377241 300229 377273
rect 305840 377829 306160 377861
rect 305840 377593 305882 377829
rect 306118 377593 306160 377829
rect 305840 377509 306160 377593
rect 305840 377273 305882 377509
rect 306118 377273 306160 377509
rect 305840 377241 306160 377273
rect 311770 377829 312090 377861
rect 311770 377593 311812 377829
rect 312048 377593 312090 377829
rect 311770 377509 312090 377593
rect 311770 377273 311812 377509
rect 312048 377273 312090 377509
rect 311770 377241 312090 377273
rect 327909 377829 328229 377861
rect 327909 377593 327951 377829
rect 328187 377593 328229 377829
rect 327909 377509 328229 377593
rect 327909 377273 327951 377509
rect 328187 377273 328229 377509
rect 327909 377241 328229 377273
rect 333840 377829 334160 377861
rect 333840 377593 333882 377829
rect 334118 377593 334160 377829
rect 333840 377509 334160 377593
rect 333840 377273 333882 377509
rect 334118 377273 334160 377509
rect 333840 377241 334160 377273
rect 339770 377829 340090 377861
rect 339770 377593 339812 377829
rect 340048 377593 340090 377829
rect 339770 377509 340090 377593
rect 339770 377273 339812 377509
rect 340048 377273 340090 377509
rect 339770 377241 340090 377273
rect 355909 377829 356229 377861
rect 355909 377593 355951 377829
rect 356187 377593 356229 377829
rect 355909 377509 356229 377593
rect 355909 377273 355951 377509
rect 356187 377273 356229 377509
rect 355909 377241 356229 377273
rect 361840 377829 362160 377861
rect 361840 377593 361882 377829
rect 362118 377593 362160 377829
rect 361840 377509 362160 377593
rect 361840 377273 361882 377509
rect 362118 377273 362160 377509
rect 361840 377241 362160 377273
rect 367770 377829 368090 377861
rect 367770 377593 367812 377829
rect 368048 377593 368090 377829
rect 367770 377509 368090 377593
rect 367770 377273 367812 377509
rect 368048 377273 368090 377509
rect 367770 377241 368090 377273
rect 383909 377829 384229 377861
rect 383909 377593 383951 377829
rect 384187 377593 384229 377829
rect 383909 377509 384229 377593
rect 383909 377273 383951 377509
rect 384187 377273 384229 377509
rect 383909 377241 384229 377273
rect 389840 377829 390160 377861
rect 389840 377593 389882 377829
rect 390118 377593 390160 377829
rect 389840 377509 390160 377593
rect 389840 377273 389882 377509
rect 390118 377273 390160 377509
rect 389840 377241 390160 377273
rect 395770 377829 396090 377861
rect 395770 377593 395812 377829
rect 396048 377593 396090 377829
rect 395770 377509 396090 377593
rect 395770 377273 395812 377509
rect 396048 377273 396090 377509
rect 395770 377241 396090 377273
rect 411909 377829 412229 377861
rect 411909 377593 411951 377829
rect 412187 377593 412229 377829
rect 411909 377509 412229 377593
rect 411909 377273 411951 377509
rect 412187 377273 412229 377509
rect 411909 377241 412229 377273
rect 417840 377829 418160 377861
rect 417840 377593 417882 377829
rect 418118 377593 418160 377829
rect 417840 377509 418160 377593
rect 417840 377273 417882 377509
rect 418118 377273 418160 377509
rect 417840 377241 418160 377273
rect 423770 377829 424090 377861
rect 423770 377593 423812 377829
rect 424048 377593 424090 377829
rect 423770 377509 424090 377593
rect 423770 377273 423812 377509
rect 424048 377273 424090 377509
rect 423770 377241 424090 377273
rect 439909 377829 440229 377861
rect 439909 377593 439951 377829
rect 440187 377593 440229 377829
rect 439909 377509 440229 377593
rect 439909 377273 439951 377509
rect 440187 377273 440229 377509
rect 439909 377241 440229 377273
rect 445840 377829 446160 377861
rect 445840 377593 445882 377829
rect 446118 377593 446160 377829
rect 445840 377509 446160 377593
rect 445840 377273 445882 377509
rect 446118 377273 446160 377509
rect 445840 377241 446160 377273
rect 451770 377829 452090 377861
rect 451770 377593 451812 377829
rect 452048 377593 452090 377829
rect 451770 377509 452090 377593
rect 451770 377273 451812 377509
rect 452048 377273 452090 377509
rect 451770 377241 452090 377273
rect 467909 377829 468229 377861
rect 467909 377593 467951 377829
rect 468187 377593 468229 377829
rect 467909 377509 468229 377593
rect 467909 377273 467951 377509
rect 468187 377273 468229 377509
rect 467909 377241 468229 377273
rect 473840 377829 474160 377861
rect 473840 377593 473882 377829
rect 474118 377593 474160 377829
rect 473840 377509 474160 377593
rect 473840 377273 473882 377509
rect 474118 377273 474160 377509
rect 473840 377241 474160 377273
rect 479770 377829 480090 377861
rect 479770 377593 479812 377829
rect 480048 377593 480090 377829
rect 479770 377509 480090 377593
rect 479770 377273 479812 377509
rect 480048 377273 480090 377509
rect 479770 377241 480090 377273
rect 495909 377829 496229 377861
rect 495909 377593 495951 377829
rect 496187 377593 496229 377829
rect 495909 377509 496229 377593
rect 495909 377273 495951 377509
rect 496187 377273 496229 377509
rect 495909 377241 496229 377273
rect 501840 377829 502160 377861
rect 501840 377593 501882 377829
rect 502118 377593 502160 377829
rect 501840 377509 502160 377593
rect 501840 377273 501882 377509
rect 502118 377273 502160 377509
rect 501840 377241 502160 377273
rect 507770 377829 508090 377861
rect 507770 377593 507812 377829
rect 508048 377593 508090 377829
rect 507770 377509 508090 377593
rect 507770 377273 507812 377509
rect 508048 377273 508090 377509
rect 507770 377241 508090 377273
rect 523909 377829 524229 377861
rect 523909 377593 523951 377829
rect 524187 377593 524229 377829
rect 523909 377509 524229 377593
rect 523909 377273 523951 377509
rect 524187 377273 524229 377509
rect 523909 377241 524229 377273
rect 529840 377829 530160 377861
rect 529840 377593 529882 377829
rect 530118 377593 530160 377829
rect 529840 377509 530160 377593
rect 529840 377273 529882 377509
rect 530118 377273 530160 377509
rect 529840 377241 530160 377273
rect 535770 377829 536090 377861
rect 535770 377593 535812 377829
rect 536048 377593 536090 377829
rect 535770 377509 536090 377593
rect 535770 377273 535812 377509
rect 536048 377273 536090 377509
rect 535770 377241 536090 377273
rect 551909 377829 552229 377861
rect 551909 377593 551951 377829
rect 552187 377593 552229 377829
rect 551909 377509 552229 377593
rect 551909 377273 551951 377509
rect 552187 377273 552229 377509
rect 551909 377241 552229 377273
rect 557840 377829 558160 377861
rect 557840 377593 557882 377829
rect 558118 377593 558160 377829
rect 557840 377509 558160 377593
rect 557840 377273 557882 377509
rect 558118 377273 558160 377509
rect 557840 377241 558160 377273
rect 563770 377829 564090 377861
rect 563770 377593 563812 377829
rect 564048 377593 564090 377829
rect 563770 377509 564090 377593
rect 563770 377273 563812 377509
rect 564048 377273 564090 377509
rect 563770 377241 564090 377273
rect 573494 377829 574114 404273
rect 573494 377593 573526 377829
rect 573762 377593 573846 377829
rect 574082 377593 574114 377829
rect 573494 377509 574114 377593
rect 573494 377273 573526 377509
rect 573762 377273 573846 377509
rect 574082 377273 574114 377509
rect 22875 374454 23195 374486
rect 22875 374218 22917 374454
rect 23153 374218 23195 374454
rect 22875 374134 23195 374218
rect 22875 373898 22917 374134
rect 23153 373898 23195 374134
rect 22875 373866 23195 373898
rect 28806 374454 29126 374486
rect 28806 374218 28848 374454
rect 29084 374218 29126 374454
rect 28806 374134 29126 374218
rect 28806 373898 28848 374134
rect 29084 373898 29126 374134
rect 28806 373866 29126 373898
rect 50875 374454 51195 374486
rect 50875 374218 50917 374454
rect 51153 374218 51195 374454
rect 50875 374134 51195 374218
rect 50875 373898 50917 374134
rect 51153 373898 51195 374134
rect 50875 373866 51195 373898
rect 56806 374454 57126 374486
rect 56806 374218 56848 374454
rect 57084 374218 57126 374454
rect 56806 374134 57126 374218
rect 56806 373898 56848 374134
rect 57084 373898 57126 374134
rect 56806 373866 57126 373898
rect 78875 374454 79195 374486
rect 78875 374218 78917 374454
rect 79153 374218 79195 374454
rect 78875 374134 79195 374218
rect 78875 373898 78917 374134
rect 79153 373898 79195 374134
rect 78875 373866 79195 373898
rect 84806 374454 85126 374486
rect 84806 374218 84848 374454
rect 85084 374218 85126 374454
rect 84806 374134 85126 374218
rect 84806 373898 84848 374134
rect 85084 373898 85126 374134
rect 84806 373866 85126 373898
rect 106875 374454 107195 374486
rect 106875 374218 106917 374454
rect 107153 374218 107195 374454
rect 106875 374134 107195 374218
rect 106875 373898 106917 374134
rect 107153 373898 107195 374134
rect 106875 373866 107195 373898
rect 112806 374454 113126 374486
rect 112806 374218 112848 374454
rect 113084 374218 113126 374454
rect 112806 374134 113126 374218
rect 112806 373898 112848 374134
rect 113084 373898 113126 374134
rect 112806 373866 113126 373898
rect 134875 374454 135195 374486
rect 134875 374218 134917 374454
rect 135153 374218 135195 374454
rect 134875 374134 135195 374218
rect 134875 373898 134917 374134
rect 135153 373898 135195 374134
rect 134875 373866 135195 373898
rect 140806 374454 141126 374486
rect 140806 374218 140848 374454
rect 141084 374218 141126 374454
rect 140806 374134 141126 374218
rect 140806 373898 140848 374134
rect 141084 373898 141126 374134
rect 140806 373866 141126 373898
rect 162875 374454 163195 374486
rect 162875 374218 162917 374454
rect 163153 374218 163195 374454
rect 162875 374134 163195 374218
rect 162875 373898 162917 374134
rect 163153 373898 163195 374134
rect 162875 373866 163195 373898
rect 168806 374454 169126 374486
rect 168806 374218 168848 374454
rect 169084 374218 169126 374454
rect 168806 374134 169126 374218
rect 168806 373898 168848 374134
rect 169084 373898 169126 374134
rect 168806 373866 169126 373898
rect 190875 374454 191195 374486
rect 190875 374218 190917 374454
rect 191153 374218 191195 374454
rect 190875 374134 191195 374218
rect 190875 373898 190917 374134
rect 191153 373898 191195 374134
rect 190875 373866 191195 373898
rect 196806 374454 197126 374486
rect 196806 374218 196848 374454
rect 197084 374218 197126 374454
rect 196806 374134 197126 374218
rect 196806 373898 196848 374134
rect 197084 373898 197126 374134
rect 196806 373866 197126 373898
rect 218875 374454 219195 374486
rect 218875 374218 218917 374454
rect 219153 374218 219195 374454
rect 218875 374134 219195 374218
rect 218875 373898 218917 374134
rect 219153 373898 219195 374134
rect 218875 373866 219195 373898
rect 224806 374454 225126 374486
rect 224806 374218 224848 374454
rect 225084 374218 225126 374454
rect 224806 374134 225126 374218
rect 224806 373898 224848 374134
rect 225084 373898 225126 374134
rect 224806 373866 225126 373898
rect 246875 374454 247195 374486
rect 246875 374218 246917 374454
rect 247153 374218 247195 374454
rect 246875 374134 247195 374218
rect 246875 373898 246917 374134
rect 247153 373898 247195 374134
rect 246875 373866 247195 373898
rect 252806 374454 253126 374486
rect 252806 374218 252848 374454
rect 253084 374218 253126 374454
rect 252806 374134 253126 374218
rect 252806 373898 252848 374134
rect 253084 373898 253126 374134
rect 252806 373866 253126 373898
rect 274875 374454 275195 374486
rect 274875 374218 274917 374454
rect 275153 374218 275195 374454
rect 274875 374134 275195 374218
rect 274875 373898 274917 374134
rect 275153 373898 275195 374134
rect 274875 373866 275195 373898
rect 280806 374454 281126 374486
rect 280806 374218 280848 374454
rect 281084 374218 281126 374454
rect 280806 374134 281126 374218
rect 280806 373898 280848 374134
rect 281084 373898 281126 374134
rect 280806 373866 281126 373898
rect 302875 374454 303195 374486
rect 302875 374218 302917 374454
rect 303153 374218 303195 374454
rect 302875 374134 303195 374218
rect 302875 373898 302917 374134
rect 303153 373898 303195 374134
rect 302875 373866 303195 373898
rect 308806 374454 309126 374486
rect 308806 374218 308848 374454
rect 309084 374218 309126 374454
rect 308806 374134 309126 374218
rect 308806 373898 308848 374134
rect 309084 373898 309126 374134
rect 308806 373866 309126 373898
rect 330875 374454 331195 374486
rect 330875 374218 330917 374454
rect 331153 374218 331195 374454
rect 330875 374134 331195 374218
rect 330875 373898 330917 374134
rect 331153 373898 331195 374134
rect 330875 373866 331195 373898
rect 336806 374454 337126 374486
rect 336806 374218 336848 374454
rect 337084 374218 337126 374454
rect 336806 374134 337126 374218
rect 336806 373898 336848 374134
rect 337084 373898 337126 374134
rect 336806 373866 337126 373898
rect 358875 374454 359195 374486
rect 358875 374218 358917 374454
rect 359153 374218 359195 374454
rect 358875 374134 359195 374218
rect 358875 373898 358917 374134
rect 359153 373898 359195 374134
rect 358875 373866 359195 373898
rect 364806 374454 365126 374486
rect 364806 374218 364848 374454
rect 365084 374218 365126 374454
rect 364806 374134 365126 374218
rect 364806 373898 364848 374134
rect 365084 373898 365126 374134
rect 364806 373866 365126 373898
rect 386875 374454 387195 374486
rect 386875 374218 386917 374454
rect 387153 374218 387195 374454
rect 386875 374134 387195 374218
rect 386875 373898 386917 374134
rect 387153 373898 387195 374134
rect 386875 373866 387195 373898
rect 392806 374454 393126 374486
rect 392806 374218 392848 374454
rect 393084 374218 393126 374454
rect 392806 374134 393126 374218
rect 392806 373898 392848 374134
rect 393084 373898 393126 374134
rect 392806 373866 393126 373898
rect 414875 374454 415195 374486
rect 414875 374218 414917 374454
rect 415153 374218 415195 374454
rect 414875 374134 415195 374218
rect 414875 373898 414917 374134
rect 415153 373898 415195 374134
rect 414875 373866 415195 373898
rect 420806 374454 421126 374486
rect 420806 374218 420848 374454
rect 421084 374218 421126 374454
rect 420806 374134 421126 374218
rect 420806 373898 420848 374134
rect 421084 373898 421126 374134
rect 420806 373866 421126 373898
rect 442875 374454 443195 374486
rect 442875 374218 442917 374454
rect 443153 374218 443195 374454
rect 442875 374134 443195 374218
rect 442875 373898 442917 374134
rect 443153 373898 443195 374134
rect 442875 373866 443195 373898
rect 448806 374454 449126 374486
rect 448806 374218 448848 374454
rect 449084 374218 449126 374454
rect 448806 374134 449126 374218
rect 448806 373898 448848 374134
rect 449084 373898 449126 374134
rect 448806 373866 449126 373898
rect 470875 374454 471195 374486
rect 470875 374218 470917 374454
rect 471153 374218 471195 374454
rect 470875 374134 471195 374218
rect 470875 373898 470917 374134
rect 471153 373898 471195 374134
rect 470875 373866 471195 373898
rect 476806 374454 477126 374486
rect 476806 374218 476848 374454
rect 477084 374218 477126 374454
rect 476806 374134 477126 374218
rect 476806 373898 476848 374134
rect 477084 373898 477126 374134
rect 476806 373866 477126 373898
rect 498875 374454 499195 374486
rect 498875 374218 498917 374454
rect 499153 374218 499195 374454
rect 498875 374134 499195 374218
rect 498875 373898 498917 374134
rect 499153 373898 499195 374134
rect 498875 373866 499195 373898
rect 504806 374454 505126 374486
rect 504806 374218 504848 374454
rect 505084 374218 505126 374454
rect 504806 374134 505126 374218
rect 504806 373898 504848 374134
rect 505084 373898 505126 374134
rect 504806 373866 505126 373898
rect 526875 374454 527195 374486
rect 526875 374218 526917 374454
rect 527153 374218 527195 374454
rect 526875 374134 527195 374218
rect 526875 373898 526917 374134
rect 527153 373898 527195 374134
rect 526875 373866 527195 373898
rect 532806 374454 533126 374486
rect 532806 374218 532848 374454
rect 533084 374218 533126 374454
rect 532806 374134 533126 374218
rect 532806 373898 532848 374134
rect 533084 373898 533126 374134
rect 532806 373866 533126 373898
rect 554875 374454 555195 374486
rect 554875 374218 554917 374454
rect 555153 374218 555195 374454
rect 554875 374134 555195 374218
rect 554875 373898 554917 374134
rect 555153 373898 555195 374134
rect 554875 373866 555195 373898
rect 560806 374454 561126 374486
rect 560806 374218 560848 374454
rect 561084 374218 561126 374454
rect 560806 374134 561126 374218
rect 560806 373898 560848 374134
rect 561084 373898 561126 374134
rect 560806 373866 561126 373898
rect -2006 350593 -1974 350829
rect -1738 350593 -1654 350829
rect -1418 350593 -1386 350829
rect -2006 350509 -1386 350593
rect -2006 350273 -1974 350509
rect -1738 350273 -1654 350509
rect -1418 350273 -1386 350509
rect -2006 323829 -1386 350273
rect 19910 350829 20230 350861
rect 19910 350593 19952 350829
rect 20188 350593 20230 350829
rect 19910 350509 20230 350593
rect 19910 350273 19952 350509
rect 20188 350273 20230 350509
rect 19910 350241 20230 350273
rect 25840 350829 26160 350861
rect 25840 350593 25882 350829
rect 26118 350593 26160 350829
rect 25840 350509 26160 350593
rect 25840 350273 25882 350509
rect 26118 350273 26160 350509
rect 25840 350241 26160 350273
rect 31771 350829 32091 350861
rect 31771 350593 31813 350829
rect 32049 350593 32091 350829
rect 31771 350509 32091 350593
rect 31771 350273 31813 350509
rect 32049 350273 32091 350509
rect 31771 350241 32091 350273
rect 47910 350829 48230 350861
rect 47910 350593 47952 350829
rect 48188 350593 48230 350829
rect 47910 350509 48230 350593
rect 47910 350273 47952 350509
rect 48188 350273 48230 350509
rect 47910 350241 48230 350273
rect 53840 350829 54160 350861
rect 53840 350593 53882 350829
rect 54118 350593 54160 350829
rect 53840 350509 54160 350593
rect 53840 350273 53882 350509
rect 54118 350273 54160 350509
rect 53840 350241 54160 350273
rect 59771 350829 60091 350861
rect 59771 350593 59813 350829
rect 60049 350593 60091 350829
rect 59771 350509 60091 350593
rect 59771 350273 59813 350509
rect 60049 350273 60091 350509
rect 59771 350241 60091 350273
rect 75910 350829 76230 350861
rect 75910 350593 75952 350829
rect 76188 350593 76230 350829
rect 75910 350509 76230 350593
rect 75910 350273 75952 350509
rect 76188 350273 76230 350509
rect 75910 350241 76230 350273
rect 81840 350829 82160 350861
rect 81840 350593 81882 350829
rect 82118 350593 82160 350829
rect 81840 350509 82160 350593
rect 81840 350273 81882 350509
rect 82118 350273 82160 350509
rect 81840 350241 82160 350273
rect 87771 350829 88091 350861
rect 87771 350593 87813 350829
rect 88049 350593 88091 350829
rect 87771 350509 88091 350593
rect 87771 350273 87813 350509
rect 88049 350273 88091 350509
rect 87771 350241 88091 350273
rect 103910 350829 104230 350861
rect 103910 350593 103952 350829
rect 104188 350593 104230 350829
rect 103910 350509 104230 350593
rect 103910 350273 103952 350509
rect 104188 350273 104230 350509
rect 103910 350241 104230 350273
rect 109840 350829 110160 350861
rect 109840 350593 109882 350829
rect 110118 350593 110160 350829
rect 109840 350509 110160 350593
rect 109840 350273 109882 350509
rect 110118 350273 110160 350509
rect 109840 350241 110160 350273
rect 115771 350829 116091 350861
rect 115771 350593 115813 350829
rect 116049 350593 116091 350829
rect 115771 350509 116091 350593
rect 115771 350273 115813 350509
rect 116049 350273 116091 350509
rect 115771 350241 116091 350273
rect 131910 350829 132230 350861
rect 131910 350593 131952 350829
rect 132188 350593 132230 350829
rect 131910 350509 132230 350593
rect 131910 350273 131952 350509
rect 132188 350273 132230 350509
rect 131910 350241 132230 350273
rect 137840 350829 138160 350861
rect 137840 350593 137882 350829
rect 138118 350593 138160 350829
rect 137840 350509 138160 350593
rect 137840 350273 137882 350509
rect 138118 350273 138160 350509
rect 137840 350241 138160 350273
rect 143771 350829 144091 350861
rect 143771 350593 143813 350829
rect 144049 350593 144091 350829
rect 143771 350509 144091 350593
rect 143771 350273 143813 350509
rect 144049 350273 144091 350509
rect 143771 350241 144091 350273
rect 159910 350829 160230 350861
rect 159910 350593 159952 350829
rect 160188 350593 160230 350829
rect 159910 350509 160230 350593
rect 159910 350273 159952 350509
rect 160188 350273 160230 350509
rect 159910 350241 160230 350273
rect 165840 350829 166160 350861
rect 165840 350593 165882 350829
rect 166118 350593 166160 350829
rect 165840 350509 166160 350593
rect 165840 350273 165882 350509
rect 166118 350273 166160 350509
rect 165840 350241 166160 350273
rect 171771 350829 172091 350861
rect 171771 350593 171813 350829
rect 172049 350593 172091 350829
rect 171771 350509 172091 350593
rect 171771 350273 171813 350509
rect 172049 350273 172091 350509
rect 171771 350241 172091 350273
rect 187910 350829 188230 350861
rect 187910 350593 187952 350829
rect 188188 350593 188230 350829
rect 187910 350509 188230 350593
rect 187910 350273 187952 350509
rect 188188 350273 188230 350509
rect 187910 350241 188230 350273
rect 193840 350829 194160 350861
rect 193840 350593 193882 350829
rect 194118 350593 194160 350829
rect 193840 350509 194160 350593
rect 193840 350273 193882 350509
rect 194118 350273 194160 350509
rect 193840 350241 194160 350273
rect 199771 350829 200091 350861
rect 199771 350593 199813 350829
rect 200049 350593 200091 350829
rect 199771 350509 200091 350593
rect 199771 350273 199813 350509
rect 200049 350273 200091 350509
rect 199771 350241 200091 350273
rect 215910 350829 216230 350861
rect 215910 350593 215952 350829
rect 216188 350593 216230 350829
rect 215910 350509 216230 350593
rect 215910 350273 215952 350509
rect 216188 350273 216230 350509
rect 215910 350241 216230 350273
rect 221840 350829 222160 350861
rect 221840 350593 221882 350829
rect 222118 350593 222160 350829
rect 221840 350509 222160 350593
rect 221840 350273 221882 350509
rect 222118 350273 222160 350509
rect 221840 350241 222160 350273
rect 227771 350829 228091 350861
rect 227771 350593 227813 350829
rect 228049 350593 228091 350829
rect 227771 350509 228091 350593
rect 227771 350273 227813 350509
rect 228049 350273 228091 350509
rect 227771 350241 228091 350273
rect 243910 350829 244230 350861
rect 243910 350593 243952 350829
rect 244188 350593 244230 350829
rect 243910 350509 244230 350593
rect 243910 350273 243952 350509
rect 244188 350273 244230 350509
rect 243910 350241 244230 350273
rect 249840 350829 250160 350861
rect 249840 350593 249882 350829
rect 250118 350593 250160 350829
rect 249840 350509 250160 350593
rect 249840 350273 249882 350509
rect 250118 350273 250160 350509
rect 249840 350241 250160 350273
rect 255771 350829 256091 350861
rect 255771 350593 255813 350829
rect 256049 350593 256091 350829
rect 255771 350509 256091 350593
rect 255771 350273 255813 350509
rect 256049 350273 256091 350509
rect 255771 350241 256091 350273
rect 271910 350829 272230 350861
rect 271910 350593 271952 350829
rect 272188 350593 272230 350829
rect 271910 350509 272230 350593
rect 271910 350273 271952 350509
rect 272188 350273 272230 350509
rect 271910 350241 272230 350273
rect 277840 350829 278160 350861
rect 277840 350593 277882 350829
rect 278118 350593 278160 350829
rect 277840 350509 278160 350593
rect 277840 350273 277882 350509
rect 278118 350273 278160 350509
rect 277840 350241 278160 350273
rect 283771 350829 284091 350861
rect 283771 350593 283813 350829
rect 284049 350593 284091 350829
rect 283771 350509 284091 350593
rect 283771 350273 283813 350509
rect 284049 350273 284091 350509
rect 283771 350241 284091 350273
rect 299910 350829 300230 350861
rect 299910 350593 299952 350829
rect 300188 350593 300230 350829
rect 299910 350509 300230 350593
rect 299910 350273 299952 350509
rect 300188 350273 300230 350509
rect 299910 350241 300230 350273
rect 305840 350829 306160 350861
rect 305840 350593 305882 350829
rect 306118 350593 306160 350829
rect 305840 350509 306160 350593
rect 305840 350273 305882 350509
rect 306118 350273 306160 350509
rect 305840 350241 306160 350273
rect 311771 350829 312091 350861
rect 311771 350593 311813 350829
rect 312049 350593 312091 350829
rect 311771 350509 312091 350593
rect 311771 350273 311813 350509
rect 312049 350273 312091 350509
rect 311771 350241 312091 350273
rect 327910 350829 328230 350861
rect 327910 350593 327952 350829
rect 328188 350593 328230 350829
rect 327910 350509 328230 350593
rect 327910 350273 327952 350509
rect 328188 350273 328230 350509
rect 327910 350241 328230 350273
rect 333840 350829 334160 350861
rect 333840 350593 333882 350829
rect 334118 350593 334160 350829
rect 333840 350509 334160 350593
rect 333840 350273 333882 350509
rect 334118 350273 334160 350509
rect 333840 350241 334160 350273
rect 339771 350829 340091 350861
rect 339771 350593 339813 350829
rect 340049 350593 340091 350829
rect 339771 350509 340091 350593
rect 339771 350273 339813 350509
rect 340049 350273 340091 350509
rect 339771 350241 340091 350273
rect 355910 350829 356230 350861
rect 355910 350593 355952 350829
rect 356188 350593 356230 350829
rect 355910 350509 356230 350593
rect 355910 350273 355952 350509
rect 356188 350273 356230 350509
rect 355910 350241 356230 350273
rect 361840 350829 362160 350861
rect 361840 350593 361882 350829
rect 362118 350593 362160 350829
rect 361840 350509 362160 350593
rect 361840 350273 361882 350509
rect 362118 350273 362160 350509
rect 361840 350241 362160 350273
rect 367771 350829 368091 350861
rect 367771 350593 367813 350829
rect 368049 350593 368091 350829
rect 367771 350509 368091 350593
rect 367771 350273 367813 350509
rect 368049 350273 368091 350509
rect 367771 350241 368091 350273
rect 383910 350829 384230 350861
rect 383910 350593 383952 350829
rect 384188 350593 384230 350829
rect 383910 350509 384230 350593
rect 383910 350273 383952 350509
rect 384188 350273 384230 350509
rect 383910 350241 384230 350273
rect 389840 350829 390160 350861
rect 389840 350593 389882 350829
rect 390118 350593 390160 350829
rect 389840 350509 390160 350593
rect 389840 350273 389882 350509
rect 390118 350273 390160 350509
rect 389840 350241 390160 350273
rect 395771 350829 396091 350861
rect 395771 350593 395813 350829
rect 396049 350593 396091 350829
rect 395771 350509 396091 350593
rect 395771 350273 395813 350509
rect 396049 350273 396091 350509
rect 395771 350241 396091 350273
rect 411910 350829 412230 350861
rect 411910 350593 411952 350829
rect 412188 350593 412230 350829
rect 411910 350509 412230 350593
rect 411910 350273 411952 350509
rect 412188 350273 412230 350509
rect 411910 350241 412230 350273
rect 417840 350829 418160 350861
rect 417840 350593 417882 350829
rect 418118 350593 418160 350829
rect 417840 350509 418160 350593
rect 417840 350273 417882 350509
rect 418118 350273 418160 350509
rect 417840 350241 418160 350273
rect 423771 350829 424091 350861
rect 423771 350593 423813 350829
rect 424049 350593 424091 350829
rect 423771 350509 424091 350593
rect 423771 350273 423813 350509
rect 424049 350273 424091 350509
rect 423771 350241 424091 350273
rect 439910 350829 440230 350861
rect 439910 350593 439952 350829
rect 440188 350593 440230 350829
rect 439910 350509 440230 350593
rect 439910 350273 439952 350509
rect 440188 350273 440230 350509
rect 439910 350241 440230 350273
rect 445840 350829 446160 350861
rect 445840 350593 445882 350829
rect 446118 350593 446160 350829
rect 445840 350509 446160 350593
rect 445840 350273 445882 350509
rect 446118 350273 446160 350509
rect 445840 350241 446160 350273
rect 451771 350829 452091 350861
rect 451771 350593 451813 350829
rect 452049 350593 452091 350829
rect 451771 350509 452091 350593
rect 451771 350273 451813 350509
rect 452049 350273 452091 350509
rect 451771 350241 452091 350273
rect 467910 350829 468230 350861
rect 467910 350593 467952 350829
rect 468188 350593 468230 350829
rect 467910 350509 468230 350593
rect 467910 350273 467952 350509
rect 468188 350273 468230 350509
rect 467910 350241 468230 350273
rect 473840 350829 474160 350861
rect 473840 350593 473882 350829
rect 474118 350593 474160 350829
rect 473840 350509 474160 350593
rect 473840 350273 473882 350509
rect 474118 350273 474160 350509
rect 473840 350241 474160 350273
rect 479771 350829 480091 350861
rect 479771 350593 479813 350829
rect 480049 350593 480091 350829
rect 479771 350509 480091 350593
rect 479771 350273 479813 350509
rect 480049 350273 480091 350509
rect 479771 350241 480091 350273
rect 495910 350829 496230 350861
rect 495910 350593 495952 350829
rect 496188 350593 496230 350829
rect 495910 350509 496230 350593
rect 495910 350273 495952 350509
rect 496188 350273 496230 350509
rect 495910 350241 496230 350273
rect 501840 350829 502160 350861
rect 501840 350593 501882 350829
rect 502118 350593 502160 350829
rect 501840 350509 502160 350593
rect 501840 350273 501882 350509
rect 502118 350273 502160 350509
rect 501840 350241 502160 350273
rect 507771 350829 508091 350861
rect 507771 350593 507813 350829
rect 508049 350593 508091 350829
rect 507771 350509 508091 350593
rect 507771 350273 507813 350509
rect 508049 350273 508091 350509
rect 507771 350241 508091 350273
rect 523910 350829 524230 350861
rect 523910 350593 523952 350829
rect 524188 350593 524230 350829
rect 523910 350509 524230 350593
rect 523910 350273 523952 350509
rect 524188 350273 524230 350509
rect 523910 350241 524230 350273
rect 529840 350829 530160 350861
rect 529840 350593 529882 350829
rect 530118 350593 530160 350829
rect 529840 350509 530160 350593
rect 529840 350273 529882 350509
rect 530118 350273 530160 350509
rect 529840 350241 530160 350273
rect 535771 350829 536091 350861
rect 535771 350593 535813 350829
rect 536049 350593 536091 350829
rect 535771 350509 536091 350593
rect 535771 350273 535813 350509
rect 536049 350273 536091 350509
rect 535771 350241 536091 350273
rect 551910 350829 552230 350861
rect 551910 350593 551952 350829
rect 552188 350593 552230 350829
rect 551910 350509 552230 350593
rect 551910 350273 551952 350509
rect 552188 350273 552230 350509
rect 551910 350241 552230 350273
rect 557840 350829 558160 350861
rect 557840 350593 557882 350829
rect 558118 350593 558160 350829
rect 557840 350509 558160 350593
rect 557840 350273 557882 350509
rect 558118 350273 558160 350509
rect 557840 350241 558160 350273
rect 563771 350829 564091 350861
rect 563771 350593 563813 350829
rect 564049 350593 564091 350829
rect 563771 350509 564091 350593
rect 563771 350273 563813 350509
rect 564049 350273 564091 350509
rect 563771 350241 564091 350273
rect 573494 350829 574114 377273
rect 573494 350593 573526 350829
rect 573762 350593 573846 350829
rect 574082 350593 574114 350829
rect 573494 350509 574114 350593
rect 573494 350273 573526 350509
rect 573762 350273 573846 350509
rect 574082 350273 574114 350509
rect 22874 347454 23194 347486
rect 22874 347218 22916 347454
rect 23152 347218 23194 347454
rect 22874 347134 23194 347218
rect 22874 346898 22916 347134
rect 23152 346898 23194 347134
rect 22874 346866 23194 346898
rect 28805 347454 29125 347486
rect 28805 347218 28847 347454
rect 29083 347218 29125 347454
rect 28805 347134 29125 347218
rect 28805 346898 28847 347134
rect 29083 346898 29125 347134
rect 28805 346866 29125 346898
rect 50874 347454 51194 347486
rect 50874 347218 50916 347454
rect 51152 347218 51194 347454
rect 50874 347134 51194 347218
rect 50874 346898 50916 347134
rect 51152 346898 51194 347134
rect 50874 346866 51194 346898
rect 56805 347454 57125 347486
rect 56805 347218 56847 347454
rect 57083 347218 57125 347454
rect 56805 347134 57125 347218
rect 56805 346898 56847 347134
rect 57083 346898 57125 347134
rect 56805 346866 57125 346898
rect 78874 347454 79194 347486
rect 78874 347218 78916 347454
rect 79152 347218 79194 347454
rect 78874 347134 79194 347218
rect 78874 346898 78916 347134
rect 79152 346898 79194 347134
rect 78874 346866 79194 346898
rect 84805 347454 85125 347486
rect 84805 347218 84847 347454
rect 85083 347218 85125 347454
rect 84805 347134 85125 347218
rect 84805 346898 84847 347134
rect 85083 346898 85125 347134
rect 84805 346866 85125 346898
rect 106874 347454 107194 347486
rect 106874 347218 106916 347454
rect 107152 347218 107194 347454
rect 106874 347134 107194 347218
rect 106874 346898 106916 347134
rect 107152 346898 107194 347134
rect 106874 346866 107194 346898
rect 112805 347454 113125 347486
rect 112805 347218 112847 347454
rect 113083 347218 113125 347454
rect 112805 347134 113125 347218
rect 112805 346898 112847 347134
rect 113083 346898 113125 347134
rect 112805 346866 113125 346898
rect 134874 347454 135194 347486
rect 134874 347218 134916 347454
rect 135152 347218 135194 347454
rect 134874 347134 135194 347218
rect 134874 346898 134916 347134
rect 135152 346898 135194 347134
rect 134874 346866 135194 346898
rect 140805 347454 141125 347486
rect 140805 347218 140847 347454
rect 141083 347218 141125 347454
rect 140805 347134 141125 347218
rect 140805 346898 140847 347134
rect 141083 346898 141125 347134
rect 140805 346866 141125 346898
rect 162874 347454 163194 347486
rect 162874 347218 162916 347454
rect 163152 347218 163194 347454
rect 162874 347134 163194 347218
rect 162874 346898 162916 347134
rect 163152 346898 163194 347134
rect 162874 346866 163194 346898
rect 168805 347454 169125 347486
rect 168805 347218 168847 347454
rect 169083 347218 169125 347454
rect 168805 347134 169125 347218
rect 168805 346898 168847 347134
rect 169083 346898 169125 347134
rect 168805 346866 169125 346898
rect 190874 347454 191194 347486
rect 190874 347218 190916 347454
rect 191152 347218 191194 347454
rect 190874 347134 191194 347218
rect 190874 346898 190916 347134
rect 191152 346898 191194 347134
rect 190874 346866 191194 346898
rect 196805 347454 197125 347486
rect 196805 347218 196847 347454
rect 197083 347218 197125 347454
rect 196805 347134 197125 347218
rect 196805 346898 196847 347134
rect 197083 346898 197125 347134
rect 196805 346866 197125 346898
rect 218874 347454 219194 347486
rect 218874 347218 218916 347454
rect 219152 347218 219194 347454
rect 218874 347134 219194 347218
rect 218874 346898 218916 347134
rect 219152 346898 219194 347134
rect 218874 346866 219194 346898
rect 224805 347454 225125 347486
rect 224805 347218 224847 347454
rect 225083 347218 225125 347454
rect 224805 347134 225125 347218
rect 224805 346898 224847 347134
rect 225083 346898 225125 347134
rect 224805 346866 225125 346898
rect 246874 347454 247194 347486
rect 246874 347218 246916 347454
rect 247152 347218 247194 347454
rect 246874 347134 247194 347218
rect 246874 346898 246916 347134
rect 247152 346898 247194 347134
rect 246874 346866 247194 346898
rect 252805 347454 253125 347486
rect 252805 347218 252847 347454
rect 253083 347218 253125 347454
rect 252805 347134 253125 347218
rect 252805 346898 252847 347134
rect 253083 346898 253125 347134
rect 252805 346866 253125 346898
rect 274874 347454 275194 347486
rect 274874 347218 274916 347454
rect 275152 347218 275194 347454
rect 274874 347134 275194 347218
rect 274874 346898 274916 347134
rect 275152 346898 275194 347134
rect 274874 346866 275194 346898
rect 280805 347454 281125 347486
rect 280805 347218 280847 347454
rect 281083 347218 281125 347454
rect 280805 347134 281125 347218
rect 280805 346898 280847 347134
rect 281083 346898 281125 347134
rect 280805 346866 281125 346898
rect 302874 347454 303194 347486
rect 302874 347218 302916 347454
rect 303152 347218 303194 347454
rect 302874 347134 303194 347218
rect 302874 346898 302916 347134
rect 303152 346898 303194 347134
rect 302874 346866 303194 346898
rect 308805 347454 309125 347486
rect 308805 347218 308847 347454
rect 309083 347218 309125 347454
rect 308805 347134 309125 347218
rect 308805 346898 308847 347134
rect 309083 346898 309125 347134
rect 308805 346866 309125 346898
rect 330874 347454 331194 347486
rect 330874 347218 330916 347454
rect 331152 347218 331194 347454
rect 330874 347134 331194 347218
rect 330874 346898 330916 347134
rect 331152 346898 331194 347134
rect 330874 346866 331194 346898
rect 336805 347454 337125 347486
rect 336805 347218 336847 347454
rect 337083 347218 337125 347454
rect 336805 347134 337125 347218
rect 336805 346898 336847 347134
rect 337083 346898 337125 347134
rect 336805 346866 337125 346898
rect 358874 347454 359194 347486
rect 358874 347218 358916 347454
rect 359152 347218 359194 347454
rect 358874 347134 359194 347218
rect 358874 346898 358916 347134
rect 359152 346898 359194 347134
rect 358874 346866 359194 346898
rect 364805 347454 365125 347486
rect 364805 347218 364847 347454
rect 365083 347218 365125 347454
rect 364805 347134 365125 347218
rect 364805 346898 364847 347134
rect 365083 346898 365125 347134
rect 364805 346866 365125 346898
rect 386874 347454 387194 347486
rect 386874 347218 386916 347454
rect 387152 347218 387194 347454
rect 386874 347134 387194 347218
rect 386874 346898 386916 347134
rect 387152 346898 387194 347134
rect 386874 346866 387194 346898
rect 392805 347454 393125 347486
rect 392805 347218 392847 347454
rect 393083 347218 393125 347454
rect 392805 347134 393125 347218
rect 392805 346898 392847 347134
rect 393083 346898 393125 347134
rect 392805 346866 393125 346898
rect 414874 347454 415194 347486
rect 414874 347218 414916 347454
rect 415152 347218 415194 347454
rect 414874 347134 415194 347218
rect 414874 346898 414916 347134
rect 415152 346898 415194 347134
rect 414874 346866 415194 346898
rect 420805 347454 421125 347486
rect 420805 347218 420847 347454
rect 421083 347218 421125 347454
rect 420805 347134 421125 347218
rect 420805 346898 420847 347134
rect 421083 346898 421125 347134
rect 420805 346866 421125 346898
rect 442874 347454 443194 347486
rect 442874 347218 442916 347454
rect 443152 347218 443194 347454
rect 442874 347134 443194 347218
rect 442874 346898 442916 347134
rect 443152 346898 443194 347134
rect 442874 346866 443194 346898
rect 448805 347454 449125 347486
rect 448805 347218 448847 347454
rect 449083 347218 449125 347454
rect 448805 347134 449125 347218
rect 448805 346898 448847 347134
rect 449083 346898 449125 347134
rect 448805 346866 449125 346898
rect 470874 347454 471194 347486
rect 470874 347218 470916 347454
rect 471152 347218 471194 347454
rect 470874 347134 471194 347218
rect 470874 346898 470916 347134
rect 471152 346898 471194 347134
rect 470874 346866 471194 346898
rect 476805 347454 477125 347486
rect 476805 347218 476847 347454
rect 477083 347218 477125 347454
rect 476805 347134 477125 347218
rect 476805 346898 476847 347134
rect 477083 346898 477125 347134
rect 476805 346866 477125 346898
rect 498874 347454 499194 347486
rect 498874 347218 498916 347454
rect 499152 347218 499194 347454
rect 498874 347134 499194 347218
rect 498874 346898 498916 347134
rect 499152 346898 499194 347134
rect 498874 346866 499194 346898
rect 504805 347454 505125 347486
rect 504805 347218 504847 347454
rect 505083 347218 505125 347454
rect 504805 347134 505125 347218
rect 504805 346898 504847 347134
rect 505083 346898 505125 347134
rect 504805 346866 505125 346898
rect 526874 347454 527194 347486
rect 526874 347218 526916 347454
rect 527152 347218 527194 347454
rect 526874 347134 527194 347218
rect 526874 346898 526916 347134
rect 527152 346898 527194 347134
rect 526874 346866 527194 346898
rect 532805 347454 533125 347486
rect 532805 347218 532847 347454
rect 533083 347218 533125 347454
rect 532805 347134 533125 347218
rect 532805 346898 532847 347134
rect 533083 346898 533125 347134
rect 532805 346866 533125 346898
rect 554874 347454 555194 347486
rect 554874 347218 554916 347454
rect 555152 347218 555194 347454
rect 554874 347134 555194 347218
rect 554874 346898 554916 347134
rect 555152 346898 555194 347134
rect 554874 346866 555194 346898
rect 560805 347454 561125 347486
rect 560805 347218 560847 347454
rect 561083 347218 561125 347454
rect 560805 347134 561125 347218
rect 560805 346898 560847 347134
rect 561083 346898 561125 347134
rect 560805 346866 561125 346898
rect -2006 323593 -1974 323829
rect -1738 323593 -1654 323829
rect -1418 323593 -1386 323829
rect -2006 323509 -1386 323593
rect -2006 323273 -1974 323509
rect -1738 323273 -1654 323509
rect -1418 323273 -1386 323509
rect -2006 296829 -1386 323273
rect 19909 323829 20229 323861
rect 19909 323593 19951 323829
rect 20187 323593 20229 323829
rect 19909 323509 20229 323593
rect 19909 323273 19951 323509
rect 20187 323273 20229 323509
rect 19909 323241 20229 323273
rect 25840 323829 26160 323861
rect 25840 323593 25882 323829
rect 26118 323593 26160 323829
rect 25840 323509 26160 323593
rect 25840 323273 25882 323509
rect 26118 323273 26160 323509
rect 25840 323241 26160 323273
rect 31770 323829 32090 323861
rect 31770 323593 31812 323829
rect 32048 323593 32090 323829
rect 31770 323509 32090 323593
rect 31770 323273 31812 323509
rect 32048 323273 32090 323509
rect 31770 323241 32090 323273
rect 47909 323829 48229 323861
rect 47909 323593 47951 323829
rect 48187 323593 48229 323829
rect 47909 323509 48229 323593
rect 47909 323273 47951 323509
rect 48187 323273 48229 323509
rect 47909 323241 48229 323273
rect 53840 323829 54160 323861
rect 53840 323593 53882 323829
rect 54118 323593 54160 323829
rect 53840 323509 54160 323593
rect 53840 323273 53882 323509
rect 54118 323273 54160 323509
rect 53840 323241 54160 323273
rect 59770 323829 60090 323861
rect 59770 323593 59812 323829
rect 60048 323593 60090 323829
rect 59770 323509 60090 323593
rect 59770 323273 59812 323509
rect 60048 323273 60090 323509
rect 59770 323241 60090 323273
rect 75909 323829 76229 323861
rect 75909 323593 75951 323829
rect 76187 323593 76229 323829
rect 75909 323509 76229 323593
rect 75909 323273 75951 323509
rect 76187 323273 76229 323509
rect 75909 323241 76229 323273
rect 81840 323829 82160 323861
rect 81840 323593 81882 323829
rect 82118 323593 82160 323829
rect 81840 323509 82160 323593
rect 81840 323273 81882 323509
rect 82118 323273 82160 323509
rect 81840 323241 82160 323273
rect 87770 323829 88090 323861
rect 87770 323593 87812 323829
rect 88048 323593 88090 323829
rect 87770 323509 88090 323593
rect 87770 323273 87812 323509
rect 88048 323273 88090 323509
rect 87770 323241 88090 323273
rect 103909 323829 104229 323861
rect 103909 323593 103951 323829
rect 104187 323593 104229 323829
rect 103909 323509 104229 323593
rect 103909 323273 103951 323509
rect 104187 323273 104229 323509
rect 103909 323241 104229 323273
rect 109840 323829 110160 323861
rect 109840 323593 109882 323829
rect 110118 323593 110160 323829
rect 109840 323509 110160 323593
rect 109840 323273 109882 323509
rect 110118 323273 110160 323509
rect 109840 323241 110160 323273
rect 115770 323829 116090 323861
rect 115770 323593 115812 323829
rect 116048 323593 116090 323829
rect 115770 323509 116090 323593
rect 115770 323273 115812 323509
rect 116048 323273 116090 323509
rect 115770 323241 116090 323273
rect 131909 323829 132229 323861
rect 131909 323593 131951 323829
rect 132187 323593 132229 323829
rect 131909 323509 132229 323593
rect 131909 323273 131951 323509
rect 132187 323273 132229 323509
rect 131909 323241 132229 323273
rect 137840 323829 138160 323861
rect 137840 323593 137882 323829
rect 138118 323593 138160 323829
rect 137840 323509 138160 323593
rect 137840 323273 137882 323509
rect 138118 323273 138160 323509
rect 137840 323241 138160 323273
rect 143770 323829 144090 323861
rect 143770 323593 143812 323829
rect 144048 323593 144090 323829
rect 143770 323509 144090 323593
rect 143770 323273 143812 323509
rect 144048 323273 144090 323509
rect 143770 323241 144090 323273
rect 159909 323829 160229 323861
rect 159909 323593 159951 323829
rect 160187 323593 160229 323829
rect 159909 323509 160229 323593
rect 159909 323273 159951 323509
rect 160187 323273 160229 323509
rect 159909 323241 160229 323273
rect 165840 323829 166160 323861
rect 165840 323593 165882 323829
rect 166118 323593 166160 323829
rect 165840 323509 166160 323593
rect 165840 323273 165882 323509
rect 166118 323273 166160 323509
rect 165840 323241 166160 323273
rect 171770 323829 172090 323861
rect 171770 323593 171812 323829
rect 172048 323593 172090 323829
rect 171770 323509 172090 323593
rect 171770 323273 171812 323509
rect 172048 323273 172090 323509
rect 171770 323241 172090 323273
rect 187909 323829 188229 323861
rect 187909 323593 187951 323829
rect 188187 323593 188229 323829
rect 187909 323509 188229 323593
rect 187909 323273 187951 323509
rect 188187 323273 188229 323509
rect 187909 323241 188229 323273
rect 193840 323829 194160 323861
rect 193840 323593 193882 323829
rect 194118 323593 194160 323829
rect 193840 323509 194160 323593
rect 193840 323273 193882 323509
rect 194118 323273 194160 323509
rect 193840 323241 194160 323273
rect 199770 323829 200090 323861
rect 199770 323593 199812 323829
rect 200048 323593 200090 323829
rect 199770 323509 200090 323593
rect 199770 323273 199812 323509
rect 200048 323273 200090 323509
rect 199770 323241 200090 323273
rect 215909 323829 216229 323861
rect 215909 323593 215951 323829
rect 216187 323593 216229 323829
rect 215909 323509 216229 323593
rect 215909 323273 215951 323509
rect 216187 323273 216229 323509
rect 215909 323241 216229 323273
rect 221840 323829 222160 323861
rect 221840 323593 221882 323829
rect 222118 323593 222160 323829
rect 221840 323509 222160 323593
rect 221840 323273 221882 323509
rect 222118 323273 222160 323509
rect 221840 323241 222160 323273
rect 227770 323829 228090 323861
rect 227770 323593 227812 323829
rect 228048 323593 228090 323829
rect 227770 323509 228090 323593
rect 227770 323273 227812 323509
rect 228048 323273 228090 323509
rect 227770 323241 228090 323273
rect 243909 323829 244229 323861
rect 243909 323593 243951 323829
rect 244187 323593 244229 323829
rect 243909 323509 244229 323593
rect 243909 323273 243951 323509
rect 244187 323273 244229 323509
rect 243909 323241 244229 323273
rect 249840 323829 250160 323861
rect 249840 323593 249882 323829
rect 250118 323593 250160 323829
rect 249840 323509 250160 323593
rect 249840 323273 249882 323509
rect 250118 323273 250160 323509
rect 249840 323241 250160 323273
rect 255770 323829 256090 323861
rect 255770 323593 255812 323829
rect 256048 323593 256090 323829
rect 255770 323509 256090 323593
rect 255770 323273 255812 323509
rect 256048 323273 256090 323509
rect 255770 323241 256090 323273
rect 271909 323829 272229 323861
rect 271909 323593 271951 323829
rect 272187 323593 272229 323829
rect 271909 323509 272229 323593
rect 271909 323273 271951 323509
rect 272187 323273 272229 323509
rect 271909 323241 272229 323273
rect 277840 323829 278160 323861
rect 277840 323593 277882 323829
rect 278118 323593 278160 323829
rect 277840 323509 278160 323593
rect 277840 323273 277882 323509
rect 278118 323273 278160 323509
rect 277840 323241 278160 323273
rect 283770 323829 284090 323861
rect 283770 323593 283812 323829
rect 284048 323593 284090 323829
rect 283770 323509 284090 323593
rect 283770 323273 283812 323509
rect 284048 323273 284090 323509
rect 283770 323241 284090 323273
rect 299909 323829 300229 323861
rect 299909 323593 299951 323829
rect 300187 323593 300229 323829
rect 299909 323509 300229 323593
rect 299909 323273 299951 323509
rect 300187 323273 300229 323509
rect 299909 323241 300229 323273
rect 305840 323829 306160 323861
rect 305840 323593 305882 323829
rect 306118 323593 306160 323829
rect 305840 323509 306160 323593
rect 305840 323273 305882 323509
rect 306118 323273 306160 323509
rect 305840 323241 306160 323273
rect 311770 323829 312090 323861
rect 311770 323593 311812 323829
rect 312048 323593 312090 323829
rect 311770 323509 312090 323593
rect 311770 323273 311812 323509
rect 312048 323273 312090 323509
rect 311770 323241 312090 323273
rect 327909 323829 328229 323861
rect 327909 323593 327951 323829
rect 328187 323593 328229 323829
rect 327909 323509 328229 323593
rect 327909 323273 327951 323509
rect 328187 323273 328229 323509
rect 327909 323241 328229 323273
rect 333840 323829 334160 323861
rect 333840 323593 333882 323829
rect 334118 323593 334160 323829
rect 333840 323509 334160 323593
rect 333840 323273 333882 323509
rect 334118 323273 334160 323509
rect 333840 323241 334160 323273
rect 339770 323829 340090 323861
rect 339770 323593 339812 323829
rect 340048 323593 340090 323829
rect 339770 323509 340090 323593
rect 339770 323273 339812 323509
rect 340048 323273 340090 323509
rect 339770 323241 340090 323273
rect 355909 323829 356229 323861
rect 355909 323593 355951 323829
rect 356187 323593 356229 323829
rect 355909 323509 356229 323593
rect 355909 323273 355951 323509
rect 356187 323273 356229 323509
rect 355909 323241 356229 323273
rect 361840 323829 362160 323861
rect 361840 323593 361882 323829
rect 362118 323593 362160 323829
rect 361840 323509 362160 323593
rect 361840 323273 361882 323509
rect 362118 323273 362160 323509
rect 361840 323241 362160 323273
rect 367770 323829 368090 323861
rect 367770 323593 367812 323829
rect 368048 323593 368090 323829
rect 367770 323509 368090 323593
rect 367770 323273 367812 323509
rect 368048 323273 368090 323509
rect 367770 323241 368090 323273
rect 383909 323829 384229 323861
rect 383909 323593 383951 323829
rect 384187 323593 384229 323829
rect 383909 323509 384229 323593
rect 383909 323273 383951 323509
rect 384187 323273 384229 323509
rect 383909 323241 384229 323273
rect 389840 323829 390160 323861
rect 389840 323593 389882 323829
rect 390118 323593 390160 323829
rect 389840 323509 390160 323593
rect 389840 323273 389882 323509
rect 390118 323273 390160 323509
rect 389840 323241 390160 323273
rect 395770 323829 396090 323861
rect 395770 323593 395812 323829
rect 396048 323593 396090 323829
rect 395770 323509 396090 323593
rect 395770 323273 395812 323509
rect 396048 323273 396090 323509
rect 395770 323241 396090 323273
rect 411909 323829 412229 323861
rect 411909 323593 411951 323829
rect 412187 323593 412229 323829
rect 411909 323509 412229 323593
rect 411909 323273 411951 323509
rect 412187 323273 412229 323509
rect 411909 323241 412229 323273
rect 417840 323829 418160 323861
rect 417840 323593 417882 323829
rect 418118 323593 418160 323829
rect 417840 323509 418160 323593
rect 417840 323273 417882 323509
rect 418118 323273 418160 323509
rect 417840 323241 418160 323273
rect 423770 323829 424090 323861
rect 423770 323593 423812 323829
rect 424048 323593 424090 323829
rect 423770 323509 424090 323593
rect 423770 323273 423812 323509
rect 424048 323273 424090 323509
rect 423770 323241 424090 323273
rect 439909 323829 440229 323861
rect 439909 323593 439951 323829
rect 440187 323593 440229 323829
rect 439909 323509 440229 323593
rect 439909 323273 439951 323509
rect 440187 323273 440229 323509
rect 439909 323241 440229 323273
rect 445840 323829 446160 323861
rect 445840 323593 445882 323829
rect 446118 323593 446160 323829
rect 445840 323509 446160 323593
rect 445840 323273 445882 323509
rect 446118 323273 446160 323509
rect 445840 323241 446160 323273
rect 451770 323829 452090 323861
rect 451770 323593 451812 323829
rect 452048 323593 452090 323829
rect 451770 323509 452090 323593
rect 451770 323273 451812 323509
rect 452048 323273 452090 323509
rect 451770 323241 452090 323273
rect 467909 323829 468229 323861
rect 467909 323593 467951 323829
rect 468187 323593 468229 323829
rect 467909 323509 468229 323593
rect 467909 323273 467951 323509
rect 468187 323273 468229 323509
rect 467909 323241 468229 323273
rect 473840 323829 474160 323861
rect 473840 323593 473882 323829
rect 474118 323593 474160 323829
rect 473840 323509 474160 323593
rect 473840 323273 473882 323509
rect 474118 323273 474160 323509
rect 473840 323241 474160 323273
rect 479770 323829 480090 323861
rect 479770 323593 479812 323829
rect 480048 323593 480090 323829
rect 479770 323509 480090 323593
rect 479770 323273 479812 323509
rect 480048 323273 480090 323509
rect 479770 323241 480090 323273
rect 495909 323829 496229 323861
rect 495909 323593 495951 323829
rect 496187 323593 496229 323829
rect 495909 323509 496229 323593
rect 495909 323273 495951 323509
rect 496187 323273 496229 323509
rect 495909 323241 496229 323273
rect 501840 323829 502160 323861
rect 501840 323593 501882 323829
rect 502118 323593 502160 323829
rect 501840 323509 502160 323593
rect 501840 323273 501882 323509
rect 502118 323273 502160 323509
rect 501840 323241 502160 323273
rect 507770 323829 508090 323861
rect 507770 323593 507812 323829
rect 508048 323593 508090 323829
rect 507770 323509 508090 323593
rect 507770 323273 507812 323509
rect 508048 323273 508090 323509
rect 507770 323241 508090 323273
rect 523909 323829 524229 323861
rect 523909 323593 523951 323829
rect 524187 323593 524229 323829
rect 523909 323509 524229 323593
rect 523909 323273 523951 323509
rect 524187 323273 524229 323509
rect 523909 323241 524229 323273
rect 529840 323829 530160 323861
rect 529840 323593 529882 323829
rect 530118 323593 530160 323829
rect 529840 323509 530160 323593
rect 529840 323273 529882 323509
rect 530118 323273 530160 323509
rect 529840 323241 530160 323273
rect 535770 323829 536090 323861
rect 535770 323593 535812 323829
rect 536048 323593 536090 323829
rect 535770 323509 536090 323593
rect 535770 323273 535812 323509
rect 536048 323273 536090 323509
rect 535770 323241 536090 323273
rect 551909 323829 552229 323861
rect 551909 323593 551951 323829
rect 552187 323593 552229 323829
rect 551909 323509 552229 323593
rect 551909 323273 551951 323509
rect 552187 323273 552229 323509
rect 551909 323241 552229 323273
rect 557840 323829 558160 323861
rect 557840 323593 557882 323829
rect 558118 323593 558160 323829
rect 557840 323509 558160 323593
rect 557840 323273 557882 323509
rect 558118 323273 558160 323509
rect 557840 323241 558160 323273
rect 563770 323829 564090 323861
rect 563770 323593 563812 323829
rect 564048 323593 564090 323829
rect 563770 323509 564090 323593
rect 563770 323273 563812 323509
rect 564048 323273 564090 323509
rect 563770 323241 564090 323273
rect 573494 323829 574114 350273
rect 573494 323593 573526 323829
rect 573762 323593 573846 323829
rect 574082 323593 574114 323829
rect 573494 323509 574114 323593
rect 573494 323273 573526 323509
rect 573762 323273 573846 323509
rect 574082 323273 574114 323509
rect 22875 320454 23195 320486
rect 22875 320218 22917 320454
rect 23153 320218 23195 320454
rect 22875 320134 23195 320218
rect 22875 319898 22917 320134
rect 23153 319898 23195 320134
rect 22875 319866 23195 319898
rect 28806 320454 29126 320486
rect 28806 320218 28848 320454
rect 29084 320218 29126 320454
rect 28806 320134 29126 320218
rect 28806 319898 28848 320134
rect 29084 319898 29126 320134
rect 28806 319866 29126 319898
rect 50875 320454 51195 320486
rect 50875 320218 50917 320454
rect 51153 320218 51195 320454
rect 50875 320134 51195 320218
rect 50875 319898 50917 320134
rect 51153 319898 51195 320134
rect 50875 319866 51195 319898
rect 56806 320454 57126 320486
rect 56806 320218 56848 320454
rect 57084 320218 57126 320454
rect 56806 320134 57126 320218
rect 56806 319898 56848 320134
rect 57084 319898 57126 320134
rect 56806 319866 57126 319898
rect 78875 320454 79195 320486
rect 78875 320218 78917 320454
rect 79153 320218 79195 320454
rect 78875 320134 79195 320218
rect 78875 319898 78917 320134
rect 79153 319898 79195 320134
rect 78875 319866 79195 319898
rect 84806 320454 85126 320486
rect 84806 320218 84848 320454
rect 85084 320218 85126 320454
rect 84806 320134 85126 320218
rect 84806 319898 84848 320134
rect 85084 319898 85126 320134
rect 84806 319866 85126 319898
rect 106875 320454 107195 320486
rect 106875 320218 106917 320454
rect 107153 320218 107195 320454
rect 106875 320134 107195 320218
rect 106875 319898 106917 320134
rect 107153 319898 107195 320134
rect 106875 319866 107195 319898
rect 112806 320454 113126 320486
rect 112806 320218 112848 320454
rect 113084 320218 113126 320454
rect 112806 320134 113126 320218
rect 112806 319898 112848 320134
rect 113084 319898 113126 320134
rect 112806 319866 113126 319898
rect 134875 320454 135195 320486
rect 134875 320218 134917 320454
rect 135153 320218 135195 320454
rect 134875 320134 135195 320218
rect 134875 319898 134917 320134
rect 135153 319898 135195 320134
rect 134875 319866 135195 319898
rect 140806 320454 141126 320486
rect 140806 320218 140848 320454
rect 141084 320218 141126 320454
rect 140806 320134 141126 320218
rect 140806 319898 140848 320134
rect 141084 319898 141126 320134
rect 140806 319866 141126 319898
rect 162875 320454 163195 320486
rect 162875 320218 162917 320454
rect 163153 320218 163195 320454
rect 162875 320134 163195 320218
rect 162875 319898 162917 320134
rect 163153 319898 163195 320134
rect 162875 319866 163195 319898
rect 168806 320454 169126 320486
rect 168806 320218 168848 320454
rect 169084 320218 169126 320454
rect 168806 320134 169126 320218
rect 168806 319898 168848 320134
rect 169084 319898 169126 320134
rect 168806 319866 169126 319898
rect 190875 320454 191195 320486
rect 190875 320218 190917 320454
rect 191153 320218 191195 320454
rect 190875 320134 191195 320218
rect 190875 319898 190917 320134
rect 191153 319898 191195 320134
rect 190875 319866 191195 319898
rect 196806 320454 197126 320486
rect 196806 320218 196848 320454
rect 197084 320218 197126 320454
rect 196806 320134 197126 320218
rect 196806 319898 196848 320134
rect 197084 319898 197126 320134
rect 196806 319866 197126 319898
rect 218875 320454 219195 320486
rect 218875 320218 218917 320454
rect 219153 320218 219195 320454
rect 218875 320134 219195 320218
rect 218875 319898 218917 320134
rect 219153 319898 219195 320134
rect 218875 319866 219195 319898
rect 224806 320454 225126 320486
rect 224806 320218 224848 320454
rect 225084 320218 225126 320454
rect 224806 320134 225126 320218
rect 224806 319898 224848 320134
rect 225084 319898 225126 320134
rect 224806 319866 225126 319898
rect 246875 320454 247195 320486
rect 246875 320218 246917 320454
rect 247153 320218 247195 320454
rect 246875 320134 247195 320218
rect 246875 319898 246917 320134
rect 247153 319898 247195 320134
rect 246875 319866 247195 319898
rect 252806 320454 253126 320486
rect 252806 320218 252848 320454
rect 253084 320218 253126 320454
rect 252806 320134 253126 320218
rect 252806 319898 252848 320134
rect 253084 319898 253126 320134
rect 252806 319866 253126 319898
rect 274875 320454 275195 320486
rect 274875 320218 274917 320454
rect 275153 320218 275195 320454
rect 274875 320134 275195 320218
rect 274875 319898 274917 320134
rect 275153 319898 275195 320134
rect 274875 319866 275195 319898
rect 280806 320454 281126 320486
rect 280806 320218 280848 320454
rect 281084 320218 281126 320454
rect 280806 320134 281126 320218
rect 280806 319898 280848 320134
rect 281084 319898 281126 320134
rect 280806 319866 281126 319898
rect 302875 320454 303195 320486
rect 302875 320218 302917 320454
rect 303153 320218 303195 320454
rect 302875 320134 303195 320218
rect 302875 319898 302917 320134
rect 303153 319898 303195 320134
rect 302875 319866 303195 319898
rect 308806 320454 309126 320486
rect 308806 320218 308848 320454
rect 309084 320218 309126 320454
rect 308806 320134 309126 320218
rect 308806 319898 308848 320134
rect 309084 319898 309126 320134
rect 308806 319866 309126 319898
rect 330875 320454 331195 320486
rect 330875 320218 330917 320454
rect 331153 320218 331195 320454
rect 330875 320134 331195 320218
rect 330875 319898 330917 320134
rect 331153 319898 331195 320134
rect 330875 319866 331195 319898
rect 336806 320454 337126 320486
rect 336806 320218 336848 320454
rect 337084 320218 337126 320454
rect 336806 320134 337126 320218
rect 336806 319898 336848 320134
rect 337084 319898 337126 320134
rect 336806 319866 337126 319898
rect 358875 320454 359195 320486
rect 358875 320218 358917 320454
rect 359153 320218 359195 320454
rect 358875 320134 359195 320218
rect 358875 319898 358917 320134
rect 359153 319898 359195 320134
rect 358875 319866 359195 319898
rect 364806 320454 365126 320486
rect 364806 320218 364848 320454
rect 365084 320218 365126 320454
rect 364806 320134 365126 320218
rect 364806 319898 364848 320134
rect 365084 319898 365126 320134
rect 364806 319866 365126 319898
rect 386875 320454 387195 320486
rect 386875 320218 386917 320454
rect 387153 320218 387195 320454
rect 386875 320134 387195 320218
rect 386875 319898 386917 320134
rect 387153 319898 387195 320134
rect 386875 319866 387195 319898
rect 392806 320454 393126 320486
rect 392806 320218 392848 320454
rect 393084 320218 393126 320454
rect 392806 320134 393126 320218
rect 392806 319898 392848 320134
rect 393084 319898 393126 320134
rect 392806 319866 393126 319898
rect 414875 320454 415195 320486
rect 414875 320218 414917 320454
rect 415153 320218 415195 320454
rect 414875 320134 415195 320218
rect 414875 319898 414917 320134
rect 415153 319898 415195 320134
rect 414875 319866 415195 319898
rect 420806 320454 421126 320486
rect 420806 320218 420848 320454
rect 421084 320218 421126 320454
rect 420806 320134 421126 320218
rect 420806 319898 420848 320134
rect 421084 319898 421126 320134
rect 420806 319866 421126 319898
rect 442875 320454 443195 320486
rect 442875 320218 442917 320454
rect 443153 320218 443195 320454
rect 442875 320134 443195 320218
rect 442875 319898 442917 320134
rect 443153 319898 443195 320134
rect 442875 319866 443195 319898
rect 448806 320454 449126 320486
rect 448806 320218 448848 320454
rect 449084 320218 449126 320454
rect 448806 320134 449126 320218
rect 448806 319898 448848 320134
rect 449084 319898 449126 320134
rect 448806 319866 449126 319898
rect 470875 320454 471195 320486
rect 470875 320218 470917 320454
rect 471153 320218 471195 320454
rect 470875 320134 471195 320218
rect 470875 319898 470917 320134
rect 471153 319898 471195 320134
rect 470875 319866 471195 319898
rect 476806 320454 477126 320486
rect 476806 320218 476848 320454
rect 477084 320218 477126 320454
rect 476806 320134 477126 320218
rect 476806 319898 476848 320134
rect 477084 319898 477126 320134
rect 476806 319866 477126 319898
rect 498875 320454 499195 320486
rect 498875 320218 498917 320454
rect 499153 320218 499195 320454
rect 498875 320134 499195 320218
rect 498875 319898 498917 320134
rect 499153 319898 499195 320134
rect 498875 319866 499195 319898
rect 504806 320454 505126 320486
rect 504806 320218 504848 320454
rect 505084 320218 505126 320454
rect 504806 320134 505126 320218
rect 504806 319898 504848 320134
rect 505084 319898 505126 320134
rect 504806 319866 505126 319898
rect 526875 320454 527195 320486
rect 526875 320218 526917 320454
rect 527153 320218 527195 320454
rect 526875 320134 527195 320218
rect 526875 319898 526917 320134
rect 527153 319898 527195 320134
rect 526875 319866 527195 319898
rect 532806 320454 533126 320486
rect 532806 320218 532848 320454
rect 533084 320218 533126 320454
rect 532806 320134 533126 320218
rect 532806 319898 532848 320134
rect 533084 319898 533126 320134
rect 532806 319866 533126 319898
rect 554875 320454 555195 320486
rect 554875 320218 554917 320454
rect 555153 320218 555195 320454
rect 554875 320134 555195 320218
rect 554875 319898 554917 320134
rect 555153 319898 555195 320134
rect 554875 319866 555195 319898
rect 560806 320454 561126 320486
rect 560806 320218 560848 320454
rect 561084 320218 561126 320454
rect 560806 320134 561126 320218
rect 560806 319898 560848 320134
rect 561084 319898 561126 320134
rect 560806 319866 561126 319898
rect -2006 296593 -1974 296829
rect -1738 296593 -1654 296829
rect -1418 296593 -1386 296829
rect -2006 296509 -1386 296593
rect -2006 296273 -1974 296509
rect -1738 296273 -1654 296509
rect -1418 296273 -1386 296509
rect -2006 269829 -1386 296273
rect 19910 296829 20230 296861
rect 19910 296593 19952 296829
rect 20188 296593 20230 296829
rect 19910 296509 20230 296593
rect 19910 296273 19952 296509
rect 20188 296273 20230 296509
rect 19910 296241 20230 296273
rect 25840 296829 26160 296861
rect 25840 296593 25882 296829
rect 26118 296593 26160 296829
rect 25840 296509 26160 296593
rect 25840 296273 25882 296509
rect 26118 296273 26160 296509
rect 25840 296241 26160 296273
rect 31771 296829 32091 296861
rect 31771 296593 31813 296829
rect 32049 296593 32091 296829
rect 31771 296509 32091 296593
rect 31771 296273 31813 296509
rect 32049 296273 32091 296509
rect 31771 296241 32091 296273
rect 47910 296829 48230 296861
rect 47910 296593 47952 296829
rect 48188 296593 48230 296829
rect 47910 296509 48230 296593
rect 47910 296273 47952 296509
rect 48188 296273 48230 296509
rect 47910 296241 48230 296273
rect 53840 296829 54160 296861
rect 53840 296593 53882 296829
rect 54118 296593 54160 296829
rect 53840 296509 54160 296593
rect 53840 296273 53882 296509
rect 54118 296273 54160 296509
rect 53840 296241 54160 296273
rect 59771 296829 60091 296861
rect 59771 296593 59813 296829
rect 60049 296593 60091 296829
rect 59771 296509 60091 296593
rect 59771 296273 59813 296509
rect 60049 296273 60091 296509
rect 59771 296241 60091 296273
rect 75910 296829 76230 296861
rect 75910 296593 75952 296829
rect 76188 296593 76230 296829
rect 75910 296509 76230 296593
rect 75910 296273 75952 296509
rect 76188 296273 76230 296509
rect 75910 296241 76230 296273
rect 81840 296829 82160 296861
rect 81840 296593 81882 296829
rect 82118 296593 82160 296829
rect 81840 296509 82160 296593
rect 81840 296273 81882 296509
rect 82118 296273 82160 296509
rect 81840 296241 82160 296273
rect 87771 296829 88091 296861
rect 87771 296593 87813 296829
rect 88049 296593 88091 296829
rect 87771 296509 88091 296593
rect 87771 296273 87813 296509
rect 88049 296273 88091 296509
rect 87771 296241 88091 296273
rect 103910 296829 104230 296861
rect 103910 296593 103952 296829
rect 104188 296593 104230 296829
rect 103910 296509 104230 296593
rect 103910 296273 103952 296509
rect 104188 296273 104230 296509
rect 103910 296241 104230 296273
rect 109840 296829 110160 296861
rect 109840 296593 109882 296829
rect 110118 296593 110160 296829
rect 109840 296509 110160 296593
rect 109840 296273 109882 296509
rect 110118 296273 110160 296509
rect 109840 296241 110160 296273
rect 115771 296829 116091 296861
rect 115771 296593 115813 296829
rect 116049 296593 116091 296829
rect 115771 296509 116091 296593
rect 115771 296273 115813 296509
rect 116049 296273 116091 296509
rect 115771 296241 116091 296273
rect 131910 296829 132230 296861
rect 131910 296593 131952 296829
rect 132188 296593 132230 296829
rect 131910 296509 132230 296593
rect 131910 296273 131952 296509
rect 132188 296273 132230 296509
rect 131910 296241 132230 296273
rect 137840 296829 138160 296861
rect 137840 296593 137882 296829
rect 138118 296593 138160 296829
rect 137840 296509 138160 296593
rect 137840 296273 137882 296509
rect 138118 296273 138160 296509
rect 137840 296241 138160 296273
rect 143771 296829 144091 296861
rect 143771 296593 143813 296829
rect 144049 296593 144091 296829
rect 143771 296509 144091 296593
rect 143771 296273 143813 296509
rect 144049 296273 144091 296509
rect 143771 296241 144091 296273
rect 159910 296829 160230 296861
rect 159910 296593 159952 296829
rect 160188 296593 160230 296829
rect 159910 296509 160230 296593
rect 159910 296273 159952 296509
rect 160188 296273 160230 296509
rect 159910 296241 160230 296273
rect 165840 296829 166160 296861
rect 165840 296593 165882 296829
rect 166118 296593 166160 296829
rect 165840 296509 166160 296593
rect 165840 296273 165882 296509
rect 166118 296273 166160 296509
rect 165840 296241 166160 296273
rect 171771 296829 172091 296861
rect 171771 296593 171813 296829
rect 172049 296593 172091 296829
rect 171771 296509 172091 296593
rect 171771 296273 171813 296509
rect 172049 296273 172091 296509
rect 171771 296241 172091 296273
rect 187910 296829 188230 296861
rect 187910 296593 187952 296829
rect 188188 296593 188230 296829
rect 187910 296509 188230 296593
rect 187910 296273 187952 296509
rect 188188 296273 188230 296509
rect 187910 296241 188230 296273
rect 193840 296829 194160 296861
rect 193840 296593 193882 296829
rect 194118 296593 194160 296829
rect 193840 296509 194160 296593
rect 193840 296273 193882 296509
rect 194118 296273 194160 296509
rect 193840 296241 194160 296273
rect 199771 296829 200091 296861
rect 199771 296593 199813 296829
rect 200049 296593 200091 296829
rect 199771 296509 200091 296593
rect 199771 296273 199813 296509
rect 200049 296273 200091 296509
rect 199771 296241 200091 296273
rect 215910 296829 216230 296861
rect 215910 296593 215952 296829
rect 216188 296593 216230 296829
rect 215910 296509 216230 296593
rect 215910 296273 215952 296509
rect 216188 296273 216230 296509
rect 215910 296241 216230 296273
rect 221840 296829 222160 296861
rect 221840 296593 221882 296829
rect 222118 296593 222160 296829
rect 221840 296509 222160 296593
rect 221840 296273 221882 296509
rect 222118 296273 222160 296509
rect 221840 296241 222160 296273
rect 227771 296829 228091 296861
rect 227771 296593 227813 296829
rect 228049 296593 228091 296829
rect 227771 296509 228091 296593
rect 227771 296273 227813 296509
rect 228049 296273 228091 296509
rect 227771 296241 228091 296273
rect 243910 296829 244230 296861
rect 243910 296593 243952 296829
rect 244188 296593 244230 296829
rect 243910 296509 244230 296593
rect 243910 296273 243952 296509
rect 244188 296273 244230 296509
rect 243910 296241 244230 296273
rect 249840 296829 250160 296861
rect 249840 296593 249882 296829
rect 250118 296593 250160 296829
rect 249840 296509 250160 296593
rect 249840 296273 249882 296509
rect 250118 296273 250160 296509
rect 249840 296241 250160 296273
rect 255771 296829 256091 296861
rect 255771 296593 255813 296829
rect 256049 296593 256091 296829
rect 255771 296509 256091 296593
rect 255771 296273 255813 296509
rect 256049 296273 256091 296509
rect 255771 296241 256091 296273
rect 271910 296829 272230 296861
rect 271910 296593 271952 296829
rect 272188 296593 272230 296829
rect 271910 296509 272230 296593
rect 271910 296273 271952 296509
rect 272188 296273 272230 296509
rect 271910 296241 272230 296273
rect 277840 296829 278160 296861
rect 277840 296593 277882 296829
rect 278118 296593 278160 296829
rect 277840 296509 278160 296593
rect 277840 296273 277882 296509
rect 278118 296273 278160 296509
rect 277840 296241 278160 296273
rect 283771 296829 284091 296861
rect 283771 296593 283813 296829
rect 284049 296593 284091 296829
rect 283771 296509 284091 296593
rect 283771 296273 283813 296509
rect 284049 296273 284091 296509
rect 283771 296241 284091 296273
rect 299910 296829 300230 296861
rect 299910 296593 299952 296829
rect 300188 296593 300230 296829
rect 299910 296509 300230 296593
rect 299910 296273 299952 296509
rect 300188 296273 300230 296509
rect 299910 296241 300230 296273
rect 305840 296829 306160 296861
rect 305840 296593 305882 296829
rect 306118 296593 306160 296829
rect 305840 296509 306160 296593
rect 305840 296273 305882 296509
rect 306118 296273 306160 296509
rect 305840 296241 306160 296273
rect 311771 296829 312091 296861
rect 311771 296593 311813 296829
rect 312049 296593 312091 296829
rect 311771 296509 312091 296593
rect 311771 296273 311813 296509
rect 312049 296273 312091 296509
rect 311771 296241 312091 296273
rect 327910 296829 328230 296861
rect 327910 296593 327952 296829
rect 328188 296593 328230 296829
rect 327910 296509 328230 296593
rect 327910 296273 327952 296509
rect 328188 296273 328230 296509
rect 327910 296241 328230 296273
rect 333840 296829 334160 296861
rect 333840 296593 333882 296829
rect 334118 296593 334160 296829
rect 333840 296509 334160 296593
rect 333840 296273 333882 296509
rect 334118 296273 334160 296509
rect 333840 296241 334160 296273
rect 339771 296829 340091 296861
rect 339771 296593 339813 296829
rect 340049 296593 340091 296829
rect 339771 296509 340091 296593
rect 339771 296273 339813 296509
rect 340049 296273 340091 296509
rect 339771 296241 340091 296273
rect 355910 296829 356230 296861
rect 355910 296593 355952 296829
rect 356188 296593 356230 296829
rect 355910 296509 356230 296593
rect 355910 296273 355952 296509
rect 356188 296273 356230 296509
rect 355910 296241 356230 296273
rect 361840 296829 362160 296861
rect 361840 296593 361882 296829
rect 362118 296593 362160 296829
rect 361840 296509 362160 296593
rect 361840 296273 361882 296509
rect 362118 296273 362160 296509
rect 361840 296241 362160 296273
rect 367771 296829 368091 296861
rect 367771 296593 367813 296829
rect 368049 296593 368091 296829
rect 367771 296509 368091 296593
rect 367771 296273 367813 296509
rect 368049 296273 368091 296509
rect 367771 296241 368091 296273
rect 383910 296829 384230 296861
rect 383910 296593 383952 296829
rect 384188 296593 384230 296829
rect 383910 296509 384230 296593
rect 383910 296273 383952 296509
rect 384188 296273 384230 296509
rect 383910 296241 384230 296273
rect 389840 296829 390160 296861
rect 389840 296593 389882 296829
rect 390118 296593 390160 296829
rect 389840 296509 390160 296593
rect 389840 296273 389882 296509
rect 390118 296273 390160 296509
rect 389840 296241 390160 296273
rect 395771 296829 396091 296861
rect 395771 296593 395813 296829
rect 396049 296593 396091 296829
rect 395771 296509 396091 296593
rect 395771 296273 395813 296509
rect 396049 296273 396091 296509
rect 395771 296241 396091 296273
rect 411910 296829 412230 296861
rect 411910 296593 411952 296829
rect 412188 296593 412230 296829
rect 411910 296509 412230 296593
rect 411910 296273 411952 296509
rect 412188 296273 412230 296509
rect 411910 296241 412230 296273
rect 417840 296829 418160 296861
rect 417840 296593 417882 296829
rect 418118 296593 418160 296829
rect 417840 296509 418160 296593
rect 417840 296273 417882 296509
rect 418118 296273 418160 296509
rect 417840 296241 418160 296273
rect 423771 296829 424091 296861
rect 423771 296593 423813 296829
rect 424049 296593 424091 296829
rect 423771 296509 424091 296593
rect 423771 296273 423813 296509
rect 424049 296273 424091 296509
rect 423771 296241 424091 296273
rect 439910 296829 440230 296861
rect 439910 296593 439952 296829
rect 440188 296593 440230 296829
rect 439910 296509 440230 296593
rect 439910 296273 439952 296509
rect 440188 296273 440230 296509
rect 439910 296241 440230 296273
rect 445840 296829 446160 296861
rect 445840 296593 445882 296829
rect 446118 296593 446160 296829
rect 445840 296509 446160 296593
rect 445840 296273 445882 296509
rect 446118 296273 446160 296509
rect 445840 296241 446160 296273
rect 451771 296829 452091 296861
rect 451771 296593 451813 296829
rect 452049 296593 452091 296829
rect 451771 296509 452091 296593
rect 451771 296273 451813 296509
rect 452049 296273 452091 296509
rect 451771 296241 452091 296273
rect 467910 296829 468230 296861
rect 467910 296593 467952 296829
rect 468188 296593 468230 296829
rect 467910 296509 468230 296593
rect 467910 296273 467952 296509
rect 468188 296273 468230 296509
rect 467910 296241 468230 296273
rect 473840 296829 474160 296861
rect 473840 296593 473882 296829
rect 474118 296593 474160 296829
rect 473840 296509 474160 296593
rect 473840 296273 473882 296509
rect 474118 296273 474160 296509
rect 473840 296241 474160 296273
rect 479771 296829 480091 296861
rect 479771 296593 479813 296829
rect 480049 296593 480091 296829
rect 479771 296509 480091 296593
rect 479771 296273 479813 296509
rect 480049 296273 480091 296509
rect 479771 296241 480091 296273
rect 495910 296829 496230 296861
rect 495910 296593 495952 296829
rect 496188 296593 496230 296829
rect 495910 296509 496230 296593
rect 495910 296273 495952 296509
rect 496188 296273 496230 296509
rect 495910 296241 496230 296273
rect 501840 296829 502160 296861
rect 501840 296593 501882 296829
rect 502118 296593 502160 296829
rect 501840 296509 502160 296593
rect 501840 296273 501882 296509
rect 502118 296273 502160 296509
rect 501840 296241 502160 296273
rect 507771 296829 508091 296861
rect 507771 296593 507813 296829
rect 508049 296593 508091 296829
rect 507771 296509 508091 296593
rect 507771 296273 507813 296509
rect 508049 296273 508091 296509
rect 507771 296241 508091 296273
rect 523910 296829 524230 296861
rect 523910 296593 523952 296829
rect 524188 296593 524230 296829
rect 523910 296509 524230 296593
rect 523910 296273 523952 296509
rect 524188 296273 524230 296509
rect 523910 296241 524230 296273
rect 529840 296829 530160 296861
rect 529840 296593 529882 296829
rect 530118 296593 530160 296829
rect 529840 296509 530160 296593
rect 529840 296273 529882 296509
rect 530118 296273 530160 296509
rect 529840 296241 530160 296273
rect 535771 296829 536091 296861
rect 535771 296593 535813 296829
rect 536049 296593 536091 296829
rect 535771 296509 536091 296593
rect 535771 296273 535813 296509
rect 536049 296273 536091 296509
rect 535771 296241 536091 296273
rect 551910 296829 552230 296861
rect 551910 296593 551952 296829
rect 552188 296593 552230 296829
rect 551910 296509 552230 296593
rect 551910 296273 551952 296509
rect 552188 296273 552230 296509
rect 551910 296241 552230 296273
rect 557840 296829 558160 296861
rect 557840 296593 557882 296829
rect 558118 296593 558160 296829
rect 557840 296509 558160 296593
rect 557840 296273 557882 296509
rect 558118 296273 558160 296509
rect 557840 296241 558160 296273
rect 563771 296829 564091 296861
rect 563771 296593 563813 296829
rect 564049 296593 564091 296829
rect 563771 296509 564091 296593
rect 563771 296273 563813 296509
rect 564049 296273 564091 296509
rect 563771 296241 564091 296273
rect 573494 296829 574114 323273
rect 573494 296593 573526 296829
rect 573762 296593 573846 296829
rect 574082 296593 574114 296829
rect 573494 296509 574114 296593
rect 573494 296273 573526 296509
rect 573762 296273 573846 296509
rect 574082 296273 574114 296509
rect 22874 293454 23194 293486
rect 22874 293218 22916 293454
rect 23152 293218 23194 293454
rect 22874 293134 23194 293218
rect 22874 292898 22916 293134
rect 23152 292898 23194 293134
rect 22874 292866 23194 292898
rect 28805 293454 29125 293486
rect 28805 293218 28847 293454
rect 29083 293218 29125 293454
rect 28805 293134 29125 293218
rect 28805 292898 28847 293134
rect 29083 292898 29125 293134
rect 28805 292866 29125 292898
rect 50874 293454 51194 293486
rect 50874 293218 50916 293454
rect 51152 293218 51194 293454
rect 50874 293134 51194 293218
rect 50874 292898 50916 293134
rect 51152 292898 51194 293134
rect 50874 292866 51194 292898
rect 56805 293454 57125 293486
rect 56805 293218 56847 293454
rect 57083 293218 57125 293454
rect 56805 293134 57125 293218
rect 56805 292898 56847 293134
rect 57083 292898 57125 293134
rect 56805 292866 57125 292898
rect 78874 293454 79194 293486
rect 78874 293218 78916 293454
rect 79152 293218 79194 293454
rect 78874 293134 79194 293218
rect 78874 292898 78916 293134
rect 79152 292898 79194 293134
rect 78874 292866 79194 292898
rect 84805 293454 85125 293486
rect 84805 293218 84847 293454
rect 85083 293218 85125 293454
rect 84805 293134 85125 293218
rect 84805 292898 84847 293134
rect 85083 292898 85125 293134
rect 84805 292866 85125 292898
rect 106874 293454 107194 293486
rect 106874 293218 106916 293454
rect 107152 293218 107194 293454
rect 106874 293134 107194 293218
rect 106874 292898 106916 293134
rect 107152 292898 107194 293134
rect 106874 292866 107194 292898
rect 112805 293454 113125 293486
rect 112805 293218 112847 293454
rect 113083 293218 113125 293454
rect 112805 293134 113125 293218
rect 112805 292898 112847 293134
rect 113083 292898 113125 293134
rect 112805 292866 113125 292898
rect 134874 293454 135194 293486
rect 134874 293218 134916 293454
rect 135152 293218 135194 293454
rect 134874 293134 135194 293218
rect 134874 292898 134916 293134
rect 135152 292898 135194 293134
rect 134874 292866 135194 292898
rect 140805 293454 141125 293486
rect 140805 293218 140847 293454
rect 141083 293218 141125 293454
rect 140805 293134 141125 293218
rect 140805 292898 140847 293134
rect 141083 292898 141125 293134
rect 140805 292866 141125 292898
rect 162874 293454 163194 293486
rect 162874 293218 162916 293454
rect 163152 293218 163194 293454
rect 162874 293134 163194 293218
rect 162874 292898 162916 293134
rect 163152 292898 163194 293134
rect 162874 292866 163194 292898
rect 168805 293454 169125 293486
rect 168805 293218 168847 293454
rect 169083 293218 169125 293454
rect 168805 293134 169125 293218
rect 168805 292898 168847 293134
rect 169083 292898 169125 293134
rect 168805 292866 169125 292898
rect 190874 293454 191194 293486
rect 190874 293218 190916 293454
rect 191152 293218 191194 293454
rect 190874 293134 191194 293218
rect 190874 292898 190916 293134
rect 191152 292898 191194 293134
rect 190874 292866 191194 292898
rect 196805 293454 197125 293486
rect 196805 293218 196847 293454
rect 197083 293218 197125 293454
rect 196805 293134 197125 293218
rect 196805 292898 196847 293134
rect 197083 292898 197125 293134
rect 196805 292866 197125 292898
rect 218874 293454 219194 293486
rect 218874 293218 218916 293454
rect 219152 293218 219194 293454
rect 218874 293134 219194 293218
rect 218874 292898 218916 293134
rect 219152 292898 219194 293134
rect 218874 292866 219194 292898
rect 224805 293454 225125 293486
rect 224805 293218 224847 293454
rect 225083 293218 225125 293454
rect 224805 293134 225125 293218
rect 224805 292898 224847 293134
rect 225083 292898 225125 293134
rect 224805 292866 225125 292898
rect 246874 293454 247194 293486
rect 246874 293218 246916 293454
rect 247152 293218 247194 293454
rect 246874 293134 247194 293218
rect 246874 292898 246916 293134
rect 247152 292898 247194 293134
rect 246874 292866 247194 292898
rect 252805 293454 253125 293486
rect 252805 293218 252847 293454
rect 253083 293218 253125 293454
rect 252805 293134 253125 293218
rect 252805 292898 252847 293134
rect 253083 292898 253125 293134
rect 252805 292866 253125 292898
rect 274874 293454 275194 293486
rect 274874 293218 274916 293454
rect 275152 293218 275194 293454
rect 274874 293134 275194 293218
rect 274874 292898 274916 293134
rect 275152 292898 275194 293134
rect 274874 292866 275194 292898
rect 280805 293454 281125 293486
rect 280805 293218 280847 293454
rect 281083 293218 281125 293454
rect 280805 293134 281125 293218
rect 280805 292898 280847 293134
rect 281083 292898 281125 293134
rect 280805 292866 281125 292898
rect 302874 293454 303194 293486
rect 302874 293218 302916 293454
rect 303152 293218 303194 293454
rect 302874 293134 303194 293218
rect 302874 292898 302916 293134
rect 303152 292898 303194 293134
rect 302874 292866 303194 292898
rect 308805 293454 309125 293486
rect 308805 293218 308847 293454
rect 309083 293218 309125 293454
rect 308805 293134 309125 293218
rect 308805 292898 308847 293134
rect 309083 292898 309125 293134
rect 308805 292866 309125 292898
rect 330874 293454 331194 293486
rect 330874 293218 330916 293454
rect 331152 293218 331194 293454
rect 330874 293134 331194 293218
rect 330874 292898 330916 293134
rect 331152 292898 331194 293134
rect 330874 292866 331194 292898
rect 336805 293454 337125 293486
rect 336805 293218 336847 293454
rect 337083 293218 337125 293454
rect 336805 293134 337125 293218
rect 336805 292898 336847 293134
rect 337083 292898 337125 293134
rect 336805 292866 337125 292898
rect 358874 293454 359194 293486
rect 358874 293218 358916 293454
rect 359152 293218 359194 293454
rect 358874 293134 359194 293218
rect 358874 292898 358916 293134
rect 359152 292898 359194 293134
rect 358874 292866 359194 292898
rect 364805 293454 365125 293486
rect 364805 293218 364847 293454
rect 365083 293218 365125 293454
rect 364805 293134 365125 293218
rect 364805 292898 364847 293134
rect 365083 292898 365125 293134
rect 364805 292866 365125 292898
rect 386874 293454 387194 293486
rect 386874 293218 386916 293454
rect 387152 293218 387194 293454
rect 386874 293134 387194 293218
rect 386874 292898 386916 293134
rect 387152 292898 387194 293134
rect 386874 292866 387194 292898
rect 392805 293454 393125 293486
rect 392805 293218 392847 293454
rect 393083 293218 393125 293454
rect 392805 293134 393125 293218
rect 392805 292898 392847 293134
rect 393083 292898 393125 293134
rect 392805 292866 393125 292898
rect 414874 293454 415194 293486
rect 414874 293218 414916 293454
rect 415152 293218 415194 293454
rect 414874 293134 415194 293218
rect 414874 292898 414916 293134
rect 415152 292898 415194 293134
rect 414874 292866 415194 292898
rect 420805 293454 421125 293486
rect 420805 293218 420847 293454
rect 421083 293218 421125 293454
rect 420805 293134 421125 293218
rect 420805 292898 420847 293134
rect 421083 292898 421125 293134
rect 420805 292866 421125 292898
rect 442874 293454 443194 293486
rect 442874 293218 442916 293454
rect 443152 293218 443194 293454
rect 442874 293134 443194 293218
rect 442874 292898 442916 293134
rect 443152 292898 443194 293134
rect 442874 292866 443194 292898
rect 448805 293454 449125 293486
rect 448805 293218 448847 293454
rect 449083 293218 449125 293454
rect 448805 293134 449125 293218
rect 448805 292898 448847 293134
rect 449083 292898 449125 293134
rect 448805 292866 449125 292898
rect 470874 293454 471194 293486
rect 470874 293218 470916 293454
rect 471152 293218 471194 293454
rect 470874 293134 471194 293218
rect 470874 292898 470916 293134
rect 471152 292898 471194 293134
rect 470874 292866 471194 292898
rect 476805 293454 477125 293486
rect 476805 293218 476847 293454
rect 477083 293218 477125 293454
rect 476805 293134 477125 293218
rect 476805 292898 476847 293134
rect 477083 292898 477125 293134
rect 476805 292866 477125 292898
rect 498874 293454 499194 293486
rect 498874 293218 498916 293454
rect 499152 293218 499194 293454
rect 498874 293134 499194 293218
rect 498874 292898 498916 293134
rect 499152 292898 499194 293134
rect 498874 292866 499194 292898
rect 504805 293454 505125 293486
rect 504805 293218 504847 293454
rect 505083 293218 505125 293454
rect 504805 293134 505125 293218
rect 504805 292898 504847 293134
rect 505083 292898 505125 293134
rect 504805 292866 505125 292898
rect 526874 293454 527194 293486
rect 526874 293218 526916 293454
rect 527152 293218 527194 293454
rect 526874 293134 527194 293218
rect 526874 292898 526916 293134
rect 527152 292898 527194 293134
rect 526874 292866 527194 292898
rect 532805 293454 533125 293486
rect 532805 293218 532847 293454
rect 533083 293218 533125 293454
rect 532805 293134 533125 293218
rect 532805 292898 532847 293134
rect 533083 292898 533125 293134
rect 532805 292866 533125 292898
rect 554874 293454 555194 293486
rect 554874 293218 554916 293454
rect 555152 293218 555194 293454
rect 554874 293134 555194 293218
rect 554874 292898 554916 293134
rect 555152 292898 555194 293134
rect 554874 292866 555194 292898
rect 560805 293454 561125 293486
rect 560805 293218 560847 293454
rect 561083 293218 561125 293454
rect 560805 293134 561125 293218
rect 560805 292898 560847 293134
rect 561083 292898 561125 293134
rect 560805 292866 561125 292898
rect -2006 269593 -1974 269829
rect -1738 269593 -1654 269829
rect -1418 269593 -1386 269829
rect -2006 269509 -1386 269593
rect -2006 269273 -1974 269509
rect -1738 269273 -1654 269509
rect -1418 269273 -1386 269509
rect -2006 242829 -1386 269273
rect 19909 269829 20229 269861
rect 19909 269593 19951 269829
rect 20187 269593 20229 269829
rect 19909 269509 20229 269593
rect 19909 269273 19951 269509
rect 20187 269273 20229 269509
rect 19909 269241 20229 269273
rect 25840 269829 26160 269861
rect 25840 269593 25882 269829
rect 26118 269593 26160 269829
rect 25840 269509 26160 269593
rect 25840 269273 25882 269509
rect 26118 269273 26160 269509
rect 25840 269241 26160 269273
rect 31770 269829 32090 269861
rect 31770 269593 31812 269829
rect 32048 269593 32090 269829
rect 31770 269509 32090 269593
rect 31770 269273 31812 269509
rect 32048 269273 32090 269509
rect 31770 269241 32090 269273
rect 47909 269829 48229 269861
rect 47909 269593 47951 269829
rect 48187 269593 48229 269829
rect 47909 269509 48229 269593
rect 47909 269273 47951 269509
rect 48187 269273 48229 269509
rect 47909 269241 48229 269273
rect 53840 269829 54160 269861
rect 53840 269593 53882 269829
rect 54118 269593 54160 269829
rect 53840 269509 54160 269593
rect 53840 269273 53882 269509
rect 54118 269273 54160 269509
rect 53840 269241 54160 269273
rect 59770 269829 60090 269861
rect 59770 269593 59812 269829
rect 60048 269593 60090 269829
rect 59770 269509 60090 269593
rect 59770 269273 59812 269509
rect 60048 269273 60090 269509
rect 59770 269241 60090 269273
rect 75909 269829 76229 269861
rect 75909 269593 75951 269829
rect 76187 269593 76229 269829
rect 75909 269509 76229 269593
rect 75909 269273 75951 269509
rect 76187 269273 76229 269509
rect 75909 269241 76229 269273
rect 81840 269829 82160 269861
rect 81840 269593 81882 269829
rect 82118 269593 82160 269829
rect 81840 269509 82160 269593
rect 81840 269273 81882 269509
rect 82118 269273 82160 269509
rect 81840 269241 82160 269273
rect 87770 269829 88090 269861
rect 87770 269593 87812 269829
rect 88048 269593 88090 269829
rect 87770 269509 88090 269593
rect 87770 269273 87812 269509
rect 88048 269273 88090 269509
rect 87770 269241 88090 269273
rect 103909 269829 104229 269861
rect 103909 269593 103951 269829
rect 104187 269593 104229 269829
rect 103909 269509 104229 269593
rect 103909 269273 103951 269509
rect 104187 269273 104229 269509
rect 103909 269241 104229 269273
rect 109840 269829 110160 269861
rect 109840 269593 109882 269829
rect 110118 269593 110160 269829
rect 109840 269509 110160 269593
rect 109840 269273 109882 269509
rect 110118 269273 110160 269509
rect 109840 269241 110160 269273
rect 115770 269829 116090 269861
rect 115770 269593 115812 269829
rect 116048 269593 116090 269829
rect 115770 269509 116090 269593
rect 115770 269273 115812 269509
rect 116048 269273 116090 269509
rect 115770 269241 116090 269273
rect 131909 269829 132229 269861
rect 131909 269593 131951 269829
rect 132187 269593 132229 269829
rect 131909 269509 132229 269593
rect 131909 269273 131951 269509
rect 132187 269273 132229 269509
rect 131909 269241 132229 269273
rect 137840 269829 138160 269861
rect 137840 269593 137882 269829
rect 138118 269593 138160 269829
rect 137840 269509 138160 269593
rect 137840 269273 137882 269509
rect 138118 269273 138160 269509
rect 137840 269241 138160 269273
rect 143770 269829 144090 269861
rect 143770 269593 143812 269829
rect 144048 269593 144090 269829
rect 143770 269509 144090 269593
rect 143770 269273 143812 269509
rect 144048 269273 144090 269509
rect 143770 269241 144090 269273
rect 159909 269829 160229 269861
rect 159909 269593 159951 269829
rect 160187 269593 160229 269829
rect 159909 269509 160229 269593
rect 159909 269273 159951 269509
rect 160187 269273 160229 269509
rect 159909 269241 160229 269273
rect 165840 269829 166160 269861
rect 165840 269593 165882 269829
rect 166118 269593 166160 269829
rect 165840 269509 166160 269593
rect 165840 269273 165882 269509
rect 166118 269273 166160 269509
rect 165840 269241 166160 269273
rect 171770 269829 172090 269861
rect 171770 269593 171812 269829
rect 172048 269593 172090 269829
rect 171770 269509 172090 269593
rect 171770 269273 171812 269509
rect 172048 269273 172090 269509
rect 171770 269241 172090 269273
rect 187909 269829 188229 269861
rect 187909 269593 187951 269829
rect 188187 269593 188229 269829
rect 187909 269509 188229 269593
rect 187909 269273 187951 269509
rect 188187 269273 188229 269509
rect 187909 269241 188229 269273
rect 193840 269829 194160 269861
rect 193840 269593 193882 269829
rect 194118 269593 194160 269829
rect 193840 269509 194160 269593
rect 193840 269273 193882 269509
rect 194118 269273 194160 269509
rect 193840 269241 194160 269273
rect 199770 269829 200090 269861
rect 199770 269593 199812 269829
rect 200048 269593 200090 269829
rect 199770 269509 200090 269593
rect 199770 269273 199812 269509
rect 200048 269273 200090 269509
rect 199770 269241 200090 269273
rect 215909 269829 216229 269861
rect 215909 269593 215951 269829
rect 216187 269593 216229 269829
rect 215909 269509 216229 269593
rect 215909 269273 215951 269509
rect 216187 269273 216229 269509
rect 215909 269241 216229 269273
rect 221840 269829 222160 269861
rect 221840 269593 221882 269829
rect 222118 269593 222160 269829
rect 221840 269509 222160 269593
rect 221840 269273 221882 269509
rect 222118 269273 222160 269509
rect 221840 269241 222160 269273
rect 227770 269829 228090 269861
rect 227770 269593 227812 269829
rect 228048 269593 228090 269829
rect 227770 269509 228090 269593
rect 227770 269273 227812 269509
rect 228048 269273 228090 269509
rect 227770 269241 228090 269273
rect 243909 269829 244229 269861
rect 243909 269593 243951 269829
rect 244187 269593 244229 269829
rect 243909 269509 244229 269593
rect 243909 269273 243951 269509
rect 244187 269273 244229 269509
rect 243909 269241 244229 269273
rect 249840 269829 250160 269861
rect 249840 269593 249882 269829
rect 250118 269593 250160 269829
rect 249840 269509 250160 269593
rect 249840 269273 249882 269509
rect 250118 269273 250160 269509
rect 249840 269241 250160 269273
rect 255770 269829 256090 269861
rect 255770 269593 255812 269829
rect 256048 269593 256090 269829
rect 255770 269509 256090 269593
rect 255770 269273 255812 269509
rect 256048 269273 256090 269509
rect 255770 269241 256090 269273
rect 271909 269829 272229 269861
rect 271909 269593 271951 269829
rect 272187 269593 272229 269829
rect 271909 269509 272229 269593
rect 271909 269273 271951 269509
rect 272187 269273 272229 269509
rect 271909 269241 272229 269273
rect 277840 269829 278160 269861
rect 277840 269593 277882 269829
rect 278118 269593 278160 269829
rect 277840 269509 278160 269593
rect 277840 269273 277882 269509
rect 278118 269273 278160 269509
rect 277840 269241 278160 269273
rect 283770 269829 284090 269861
rect 283770 269593 283812 269829
rect 284048 269593 284090 269829
rect 283770 269509 284090 269593
rect 283770 269273 283812 269509
rect 284048 269273 284090 269509
rect 283770 269241 284090 269273
rect 299909 269829 300229 269861
rect 299909 269593 299951 269829
rect 300187 269593 300229 269829
rect 299909 269509 300229 269593
rect 299909 269273 299951 269509
rect 300187 269273 300229 269509
rect 299909 269241 300229 269273
rect 305840 269829 306160 269861
rect 305840 269593 305882 269829
rect 306118 269593 306160 269829
rect 305840 269509 306160 269593
rect 305840 269273 305882 269509
rect 306118 269273 306160 269509
rect 305840 269241 306160 269273
rect 311770 269829 312090 269861
rect 311770 269593 311812 269829
rect 312048 269593 312090 269829
rect 311770 269509 312090 269593
rect 311770 269273 311812 269509
rect 312048 269273 312090 269509
rect 311770 269241 312090 269273
rect 327909 269829 328229 269861
rect 327909 269593 327951 269829
rect 328187 269593 328229 269829
rect 327909 269509 328229 269593
rect 327909 269273 327951 269509
rect 328187 269273 328229 269509
rect 327909 269241 328229 269273
rect 333840 269829 334160 269861
rect 333840 269593 333882 269829
rect 334118 269593 334160 269829
rect 333840 269509 334160 269593
rect 333840 269273 333882 269509
rect 334118 269273 334160 269509
rect 333840 269241 334160 269273
rect 339770 269829 340090 269861
rect 339770 269593 339812 269829
rect 340048 269593 340090 269829
rect 339770 269509 340090 269593
rect 339770 269273 339812 269509
rect 340048 269273 340090 269509
rect 339770 269241 340090 269273
rect 355909 269829 356229 269861
rect 355909 269593 355951 269829
rect 356187 269593 356229 269829
rect 355909 269509 356229 269593
rect 355909 269273 355951 269509
rect 356187 269273 356229 269509
rect 355909 269241 356229 269273
rect 361840 269829 362160 269861
rect 361840 269593 361882 269829
rect 362118 269593 362160 269829
rect 361840 269509 362160 269593
rect 361840 269273 361882 269509
rect 362118 269273 362160 269509
rect 361840 269241 362160 269273
rect 367770 269829 368090 269861
rect 367770 269593 367812 269829
rect 368048 269593 368090 269829
rect 367770 269509 368090 269593
rect 367770 269273 367812 269509
rect 368048 269273 368090 269509
rect 367770 269241 368090 269273
rect 383909 269829 384229 269861
rect 383909 269593 383951 269829
rect 384187 269593 384229 269829
rect 383909 269509 384229 269593
rect 383909 269273 383951 269509
rect 384187 269273 384229 269509
rect 383909 269241 384229 269273
rect 389840 269829 390160 269861
rect 389840 269593 389882 269829
rect 390118 269593 390160 269829
rect 389840 269509 390160 269593
rect 389840 269273 389882 269509
rect 390118 269273 390160 269509
rect 389840 269241 390160 269273
rect 395770 269829 396090 269861
rect 395770 269593 395812 269829
rect 396048 269593 396090 269829
rect 395770 269509 396090 269593
rect 395770 269273 395812 269509
rect 396048 269273 396090 269509
rect 395770 269241 396090 269273
rect 411909 269829 412229 269861
rect 411909 269593 411951 269829
rect 412187 269593 412229 269829
rect 411909 269509 412229 269593
rect 411909 269273 411951 269509
rect 412187 269273 412229 269509
rect 411909 269241 412229 269273
rect 417840 269829 418160 269861
rect 417840 269593 417882 269829
rect 418118 269593 418160 269829
rect 417840 269509 418160 269593
rect 417840 269273 417882 269509
rect 418118 269273 418160 269509
rect 417840 269241 418160 269273
rect 423770 269829 424090 269861
rect 423770 269593 423812 269829
rect 424048 269593 424090 269829
rect 423770 269509 424090 269593
rect 423770 269273 423812 269509
rect 424048 269273 424090 269509
rect 423770 269241 424090 269273
rect 439909 269829 440229 269861
rect 439909 269593 439951 269829
rect 440187 269593 440229 269829
rect 439909 269509 440229 269593
rect 439909 269273 439951 269509
rect 440187 269273 440229 269509
rect 439909 269241 440229 269273
rect 445840 269829 446160 269861
rect 445840 269593 445882 269829
rect 446118 269593 446160 269829
rect 445840 269509 446160 269593
rect 445840 269273 445882 269509
rect 446118 269273 446160 269509
rect 445840 269241 446160 269273
rect 451770 269829 452090 269861
rect 451770 269593 451812 269829
rect 452048 269593 452090 269829
rect 451770 269509 452090 269593
rect 451770 269273 451812 269509
rect 452048 269273 452090 269509
rect 451770 269241 452090 269273
rect 467909 269829 468229 269861
rect 467909 269593 467951 269829
rect 468187 269593 468229 269829
rect 467909 269509 468229 269593
rect 467909 269273 467951 269509
rect 468187 269273 468229 269509
rect 467909 269241 468229 269273
rect 473840 269829 474160 269861
rect 473840 269593 473882 269829
rect 474118 269593 474160 269829
rect 473840 269509 474160 269593
rect 473840 269273 473882 269509
rect 474118 269273 474160 269509
rect 473840 269241 474160 269273
rect 479770 269829 480090 269861
rect 479770 269593 479812 269829
rect 480048 269593 480090 269829
rect 479770 269509 480090 269593
rect 479770 269273 479812 269509
rect 480048 269273 480090 269509
rect 479770 269241 480090 269273
rect 495909 269829 496229 269861
rect 495909 269593 495951 269829
rect 496187 269593 496229 269829
rect 495909 269509 496229 269593
rect 495909 269273 495951 269509
rect 496187 269273 496229 269509
rect 495909 269241 496229 269273
rect 501840 269829 502160 269861
rect 501840 269593 501882 269829
rect 502118 269593 502160 269829
rect 501840 269509 502160 269593
rect 501840 269273 501882 269509
rect 502118 269273 502160 269509
rect 501840 269241 502160 269273
rect 507770 269829 508090 269861
rect 507770 269593 507812 269829
rect 508048 269593 508090 269829
rect 507770 269509 508090 269593
rect 507770 269273 507812 269509
rect 508048 269273 508090 269509
rect 507770 269241 508090 269273
rect 523909 269829 524229 269861
rect 523909 269593 523951 269829
rect 524187 269593 524229 269829
rect 523909 269509 524229 269593
rect 523909 269273 523951 269509
rect 524187 269273 524229 269509
rect 523909 269241 524229 269273
rect 529840 269829 530160 269861
rect 529840 269593 529882 269829
rect 530118 269593 530160 269829
rect 529840 269509 530160 269593
rect 529840 269273 529882 269509
rect 530118 269273 530160 269509
rect 529840 269241 530160 269273
rect 535770 269829 536090 269861
rect 535770 269593 535812 269829
rect 536048 269593 536090 269829
rect 535770 269509 536090 269593
rect 535770 269273 535812 269509
rect 536048 269273 536090 269509
rect 535770 269241 536090 269273
rect 551909 269829 552229 269861
rect 551909 269593 551951 269829
rect 552187 269593 552229 269829
rect 551909 269509 552229 269593
rect 551909 269273 551951 269509
rect 552187 269273 552229 269509
rect 551909 269241 552229 269273
rect 557840 269829 558160 269861
rect 557840 269593 557882 269829
rect 558118 269593 558160 269829
rect 557840 269509 558160 269593
rect 557840 269273 557882 269509
rect 558118 269273 558160 269509
rect 557840 269241 558160 269273
rect 563770 269829 564090 269861
rect 563770 269593 563812 269829
rect 564048 269593 564090 269829
rect 563770 269509 564090 269593
rect 563770 269273 563812 269509
rect 564048 269273 564090 269509
rect 563770 269241 564090 269273
rect 573494 269829 574114 296273
rect 573494 269593 573526 269829
rect 573762 269593 573846 269829
rect 574082 269593 574114 269829
rect 573494 269509 574114 269593
rect 573494 269273 573526 269509
rect 573762 269273 573846 269509
rect 574082 269273 574114 269509
rect 22875 266454 23195 266486
rect 22875 266218 22917 266454
rect 23153 266218 23195 266454
rect 22875 266134 23195 266218
rect 22875 265898 22917 266134
rect 23153 265898 23195 266134
rect 22875 265866 23195 265898
rect 28806 266454 29126 266486
rect 28806 266218 28848 266454
rect 29084 266218 29126 266454
rect 28806 266134 29126 266218
rect 28806 265898 28848 266134
rect 29084 265898 29126 266134
rect 28806 265866 29126 265898
rect 50875 266454 51195 266486
rect 50875 266218 50917 266454
rect 51153 266218 51195 266454
rect 50875 266134 51195 266218
rect 50875 265898 50917 266134
rect 51153 265898 51195 266134
rect 50875 265866 51195 265898
rect 56806 266454 57126 266486
rect 56806 266218 56848 266454
rect 57084 266218 57126 266454
rect 56806 266134 57126 266218
rect 56806 265898 56848 266134
rect 57084 265898 57126 266134
rect 56806 265866 57126 265898
rect 78875 266454 79195 266486
rect 78875 266218 78917 266454
rect 79153 266218 79195 266454
rect 78875 266134 79195 266218
rect 78875 265898 78917 266134
rect 79153 265898 79195 266134
rect 78875 265866 79195 265898
rect 84806 266454 85126 266486
rect 84806 266218 84848 266454
rect 85084 266218 85126 266454
rect 84806 266134 85126 266218
rect 84806 265898 84848 266134
rect 85084 265898 85126 266134
rect 84806 265866 85126 265898
rect 106875 266454 107195 266486
rect 106875 266218 106917 266454
rect 107153 266218 107195 266454
rect 106875 266134 107195 266218
rect 106875 265898 106917 266134
rect 107153 265898 107195 266134
rect 106875 265866 107195 265898
rect 112806 266454 113126 266486
rect 112806 266218 112848 266454
rect 113084 266218 113126 266454
rect 112806 266134 113126 266218
rect 112806 265898 112848 266134
rect 113084 265898 113126 266134
rect 112806 265866 113126 265898
rect 134875 266454 135195 266486
rect 134875 266218 134917 266454
rect 135153 266218 135195 266454
rect 134875 266134 135195 266218
rect 134875 265898 134917 266134
rect 135153 265898 135195 266134
rect 134875 265866 135195 265898
rect 140806 266454 141126 266486
rect 140806 266218 140848 266454
rect 141084 266218 141126 266454
rect 140806 266134 141126 266218
rect 140806 265898 140848 266134
rect 141084 265898 141126 266134
rect 140806 265866 141126 265898
rect 162875 266454 163195 266486
rect 162875 266218 162917 266454
rect 163153 266218 163195 266454
rect 162875 266134 163195 266218
rect 162875 265898 162917 266134
rect 163153 265898 163195 266134
rect 162875 265866 163195 265898
rect 168806 266454 169126 266486
rect 168806 266218 168848 266454
rect 169084 266218 169126 266454
rect 168806 266134 169126 266218
rect 168806 265898 168848 266134
rect 169084 265898 169126 266134
rect 168806 265866 169126 265898
rect 190875 266454 191195 266486
rect 190875 266218 190917 266454
rect 191153 266218 191195 266454
rect 190875 266134 191195 266218
rect 190875 265898 190917 266134
rect 191153 265898 191195 266134
rect 190875 265866 191195 265898
rect 196806 266454 197126 266486
rect 196806 266218 196848 266454
rect 197084 266218 197126 266454
rect 196806 266134 197126 266218
rect 196806 265898 196848 266134
rect 197084 265898 197126 266134
rect 196806 265866 197126 265898
rect 218875 266454 219195 266486
rect 218875 266218 218917 266454
rect 219153 266218 219195 266454
rect 218875 266134 219195 266218
rect 218875 265898 218917 266134
rect 219153 265898 219195 266134
rect 218875 265866 219195 265898
rect 224806 266454 225126 266486
rect 224806 266218 224848 266454
rect 225084 266218 225126 266454
rect 224806 266134 225126 266218
rect 224806 265898 224848 266134
rect 225084 265898 225126 266134
rect 224806 265866 225126 265898
rect 246875 266454 247195 266486
rect 246875 266218 246917 266454
rect 247153 266218 247195 266454
rect 246875 266134 247195 266218
rect 246875 265898 246917 266134
rect 247153 265898 247195 266134
rect 246875 265866 247195 265898
rect 252806 266454 253126 266486
rect 252806 266218 252848 266454
rect 253084 266218 253126 266454
rect 252806 266134 253126 266218
rect 252806 265898 252848 266134
rect 253084 265898 253126 266134
rect 252806 265866 253126 265898
rect 274875 266454 275195 266486
rect 274875 266218 274917 266454
rect 275153 266218 275195 266454
rect 274875 266134 275195 266218
rect 274875 265898 274917 266134
rect 275153 265898 275195 266134
rect 274875 265866 275195 265898
rect 280806 266454 281126 266486
rect 280806 266218 280848 266454
rect 281084 266218 281126 266454
rect 280806 266134 281126 266218
rect 280806 265898 280848 266134
rect 281084 265898 281126 266134
rect 280806 265866 281126 265898
rect 302875 266454 303195 266486
rect 302875 266218 302917 266454
rect 303153 266218 303195 266454
rect 302875 266134 303195 266218
rect 302875 265898 302917 266134
rect 303153 265898 303195 266134
rect 302875 265866 303195 265898
rect 308806 266454 309126 266486
rect 308806 266218 308848 266454
rect 309084 266218 309126 266454
rect 308806 266134 309126 266218
rect 308806 265898 308848 266134
rect 309084 265898 309126 266134
rect 308806 265866 309126 265898
rect 330875 266454 331195 266486
rect 330875 266218 330917 266454
rect 331153 266218 331195 266454
rect 330875 266134 331195 266218
rect 330875 265898 330917 266134
rect 331153 265898 331195 266134
rect 330875 265866 331195 265898
rect 336806 266454 337126 266486
rect 336806 266218 336848 266454
rect 337084 266218 337126 266454
rect 336806 266134 337126 266218
rect 336806 265898 336848 266134
rect 337084 265898 337126 266134
rect 336806 265866 337126 265898
rect 358875 266454 359195 266486
rect 358875 266218 358917 266454
rect 359153 266218 359195 266454
rect 358875 266134 359195 266218
rect 358875 265898 358917 266134
rect 359153 265898 359195 266134
rect 358875 265866 359195 265898
rect 364806 266454 365126 266486
rect 364806 266218 364848 266454
rect 365084 266218 365126 266454
rect 364806 266134 365126 266218
rect 364806 265898 364848 266134
rect 365084 265898 365126 266134
rect 364806 265866 365126 265898
rect 386875 266454 387195 266486
rect 386875 266218 386917 266454
rect 387153 266218 387195 266454
rect 386875 266134 387195 266218
rect 386875 265898 386917 266134
rect 387153 265898 387195 266134
rect 386875 265866 387195 265898
rect 392806 266454 393126 266486
rect 392806 266218 392848 266454
rect 393084 266218 393126 266454
rect 392806 266134 393126 266218
rect 392806 265898 392848 266134
rect 393084 265898 393126 266134
rect 392806 265866 393126 265898
rect 414875 266454 415195 266486
rect 414875 266218 414917 266454
rect 415153 266218 415195 266454
rect 414875 266134 415195 266218
rect 414875 265898 414917 266134
rect 415153 265898 415195 266134
rect 414875 265866 415195 265898
rect 420806 266454 421126 266486
rect 420806 266218 420848 266454
rect 421084 266218 421126 266454
rect 420806 266134 421126 266218
rect 420806 265898 420848 266134
rect 421084 265898 421126 266134
rect 420806 265866 421126 265898
rect 442875 266454 443195 266486
rect 442875 266218 442917 266454
rect 443153 266218 443195 266454
rect 442875 266134 443195 266218
rect 442875 265898 442917 266134
rect 443153 265898 443195 266134
rect 442875 265866 443195 265898
rect 448806 266454 449126 266486
rect 448806 266218 448848 266454
rect 449084 266218 449126 266454
rect 448806 266134 449126 266218
rect 448806 265898 448848 266134
rect 449084 265898 449126 266134
rect 448806 265866 449126 265898
rect 470875 266454 471195 266486
rect 470875 266218 470917 266454
rect 471153 266218 471195 266454
rect 470875 266134 471195 266218
rect 470875 265898 470917 266134
rect 471153 265898 471195 266134
rect 470875 265866 471195 265898
rect 476806 266454 477126 266486
rect 476806 266218 476848 266454
rect 477084 266218 477126 266454
rect 476806 266134 477126 266218
rect 476806 265898 476848 266134
rect 477084 265898 477126 266134
rect 476806 265866 477126 265898
rect 498875 266454 499195 266486
rect 498875 266218 498917 266454
rect 499153 266218 499195 266454
rect 498875 266134 499195 266218
rect 498875 265898 498917 266134
rect 499153 265898 499195 266134
rect 498875 265866 499195 265898
rect 504806 266454 505126 266486
rect 504806 266218 504848 266454
rect 505084 266218 505126 266454
rect 504806 266134 505126 266218
rect 504806 265898 504848 266134
rect 505084 265898 505126 266134
rect 504806 265866 505126 265898
rect 526875 266454 527195 266486
rect 526875 266218 526917 266454
rect 527153 266218 527195 266454
rect 526875 266134 527195 266218
rect 526875 265898 526917 266134
rect 527153 265898 527195 266134
rect 526875 265866 527195 265898
rect 532806 266454 533126 266486
rect 532806 266218 532848 266454
rect 533084 266218 533126 266454
rect 532806 266134 533126 266218
rect 532806 265898 532848 266134
rect 533084 265898 533126 266134
rect 532806 265866 533126 265898
rect 554875 266454 555195 266486
rect 554875 266218 554917 266454
rect 555153 266218 555195 266454
rect 554875 266134 555195 266218
rect 554875 265898 554917 266134
rect 555153 265898 555195 266134
rect 554875 265866 555195 265898
rect 560806 266454 561126 266486
rect 560806 266218 560848 266454
rect 561084 266218 561126 266454
rect 560806 266134 561126 266218
rect 560806 265898 560848 266134
rect 561084 265898 561126 266134
rect 560806 265866 561126 265898
rect -2006 242593 -1974 242829
rect -1738 242593 -1654 242829
rect -1418 242593 -1386 242829
rect -2006 242509 -1386 242593
rect -2006 242273 -1974 242509
rect -1738 242273 -1654 242509
rect -1418 242273 -1386 242509
rect -2006 215829 -1386 242273
rect 19910 242829 20230 242861
rect 19910 242593 19952 242829
rect 20188 242593 20230 242829
rect 19910 242509 20230 242593
rect 19910 242273 19952 242509
rect 20188 242273 20230 242509
rect 19910 242241 20230 242273
rect 25840 242829 26160 242861
rect 25840 242593 25882 242829
rect 26118 242593 26160 242829
rect 25840 242509 26160 242593
rect 25840 242273 25882 242509
rect 26118 242273 26160 242509
rect 25840 242241 26160 242273
rect 31771 242829 32091 242861
rect 31771 242593 31813 242829
rect 32049 242593 32091 242829
rect 31771 242509 32091 242593
rect 31771 242273 31813 242509
rect 32049 242273 32091 242509
rect 31771 242241 32091 242273
rect 47910 242829 48230 242861
rect 47910 242593 47952 242829
rect 48188 242593 48230 242829
rect 47910 242509 48230 242593
rect 47910 242273 47952 242509
rect 48188 242273 48230 242509
rect 47910 242241 48230 242273
rect 53840 242829 54160 242861
rect 53840 242593 53882 242829
rect 54118 242593 54160 242829
rect 53840 242509 54160 242593
rect 53840 242273 53882 242509
rect 54118 242273 54160 242509
rect 53840 242241 54160 242273
rect 59771 242829 60091 242861
rect 59771 242593 59813 242829
rect 60049 242593 60091 242829
rect 59771 242509 60091 242593
rect 59771 242273 59813 242509
rect 60049 242273 60091 242509
rect 59771 242241 60091 242273
rect 75910 242829 76230 242861
rect 75910 242593 75952 242829
rect 76188 242593 76230 242829
rect 75910 242509 76230 242593
rect 75910 242273 75952 242509
rect 76188 242273 76230 242509
rect 75910 242241 76230 242273
rect 81840 242829 82160 242861
rect 81840 242593 81882 242829
rect 82118 242593 82160 242829
rect 81840 242509 82160 242593
rect 81840 242273 81882 242509
rect 82118 242273 82160 242509
rect 81840 242241 82160 242273
rect 87771 242829 88091 242861
rect 87771 242593 87813 242829
rect 88049 242593 88091 242829
rect 87771 242509 88091 242593
rect 87771 242273 87813 242509
rect 88049 242273 88091 242509
rect 87771 242241 88091 242273
rect 103910 242829 104230 242861
rect 103910 242593 103952 242829
rect 104188 242593 104230 242829
rect 103910 242509 104230 242593
rect 103910 242273 103952 242509
rect 104188 242273 104230 242509
rect 103910 242241 104230 242273
rect 109840 242829 110160 242861
rect 109840 242593 109882 242829
rect 110118 242593 110160 242829
rect 109840 242509 110160 242593
rect 109840 242273 109882 242509
rect 110118 242273 110160 242509
rect 109840 242241 110160 242273
rect 115771 242829 116091 242861
rect 115771 242593 115813 242829
rect 116049 242593 116091 242829
rect 115771 242509 116091 242593
rect 115771 242273 115813 242509
rect 116049 242273 116091 242509
rect 115771 242241 116091 242273
rect 131910 242829 132230 242861
rect 131910 242593 131952 242829
rect 132188 242593 132230 242829
rect 131910 242509 132230 242593
rect 131910 242273 131952 242509
rect 132188 242273 132230 242509
rect 131910 242241 132230 242273
rect 137840 242829 138160 242861
rect 137840 242593 137882 242829
rect 138118 242593 138160 242829
rect 137840 242509 138160 242593
rect 137840 242273 137882 242509
rect 138118 242273 138160 242509
rect 137840 242241 138160 242273
rect 143771 242829 144091 242861
rect 143771 242593 143813 242829
rect 144049 242593 144091 242829
rect 143771 242509 144091 242593
rect 143771 242273 143813 242509
rect 144049 242273 144091 242509
rect 143771 242241 144091 242273
rect 159910 242829 160230 242861
rect 159910 242593 159952 242829
rect 160188 242593 160230 242829
rect 159910 242509 160230 242593
rect 159910 242273 159952 242509
rect 160188 242273 160230 242509
rect 159910 242241 160230 242273
rect 165840 242829 166160 242861
rect 165840 242593 165882 242829
rect 166118 242593 166160 242829
rect 165840 242509 166160 242593
rect 165840 242273 165882 242509
rect 166118 242273 166160 242509
rect 165840 242241 166160 242273
rect 171771 242829 172091 242861
rect 171771 242593 171813 242829
rect 172049 242593 172091 242829
rect 171771 242509 172091 242593
rect 171771 242273 171813 242509
rect 172049 242273 172091 242509
rect 171771 242241 172091 242273
rect 187910 242829 188230 242861
rect 187910 242593 187952 242829
rect 188188 242593 188230 242829
rect 187910 242509 188230 242593
rect 187910 242273 187952 242509
rect 188188 242273 188230 242509
rect 187910 242241 188230 242273
rect 193840 242829 194160 242861
rect 193840 242593 193882 242829
rect 194118 242593 194160 242829
rect 193840 242509 194160 242593
rect 193840 242273 193882 242509
rect 194118 242273 194160 242509
rect 193840 242241 194160 242273
rect 199771 242829 200091 242861
rect 199771 242593 199813 242829
rect 200049 242593 200091 242829
rect 199771 242509 200091 242593
rect 199771 242273 199813 242509
rect 200049 242273 200091 242509
rect 199771 242241 200091 242273
rect 215910 242829 216230 242861
rect 215910 242593 215952 242829
rect 216188 242593 216230 242829
rect 215910 242509 216230 242593
rect 215910 242273 215952 242509
rect 216188 242273 216230 242509
rect 215910 242241 216230 242273
rect 221840 242829 222160 242861
rect 221840 242593 221882 242829
rect 222118 242593 222160 242829
rect 221840 242509 222160 242593
rect 221840 242273 221882 242509
rect 222118 242273 222160 242509
rect 221840 242241 222160 242273
rect 227771 242829 228091 242861
rect 227771 242593 227813 242829
rect 228049 242593 228091 242829
rect 227771 242509 228091 242593
rect 227771 242273 227813 242509
rect 228049 242273 228091 242509
rect 227771 242241 228091 242273
rect 243910 242829 244230 242861
rect 243910 242593 243952 242829
rect 244188 242593 244230 242829
rect 243910 242509 244230 242593
rect 243910 242273 243952 242509
rect 244188 242273 244230 242509
rect 243910 242241 244230 242273
rect 249840 242829 250160 242861
rect 249840 242593 249882 242829
rect 250118 242593 250160 242829
rect 249840 242509 250160 242593
rect 249840 242273 249882 242509
rect 250118 242273 250160 242509
rect 249840 242241 250160 242273
rect 255771 242829 256091 242861
rect 255771 242593 255813 242829
rect 256049 242593 256091 242829
rect 255771 242509 256091 242593
rect 255771 242273 255813 242509
rect 256049 242273 256091 242509
rect 255771 242241 256091 242273
rect 271910 242829 272230 242861
rect 271910 242593 271952 242829
rect 272188 242593 272230 242829
rect 271910 242509 272230 242593
rect 271910 242273 271952 242509
rect 272188 242273 272230 242509
rect 271910 242241 272230 242273
rect 277840 242829 278160 242861
rect 277840 242593 277882 242829
rect 278118 242593 278160 242829
rect 277840 242509 278160 242593
rect 277840 242273 277882 242509
rect 278118 242273 278160 242509
rect 277840 242241 278160 242273
rect 283771 242829 284091 242861
rect 283771 242593 283813 242829
rect 284049 242593 284091 242829
rect 283771 242509 284091 242593
rect 283771 242273 283813 242509
rect 284049 242273 284091 242509
rect 283771 242241 284091 242273
rect 299910 242829 300230 242861
rect 299910 242593 299952 242829
rect 300188 242593 300230 242829
rect 299910 242509 300230 242593
rect 299910 242273 299952 242509
rect 300188 242273 300230 242509
rect 299910 242241 300230 242273
rect 305840 242829 306160 242861
rect 305840 242593 305882 242829
rect 306118 242593 306160 242829
rect 305840 242509 306160 242593
rect 305840 242273 305882 242509
rect 306118 242273 306160 242509
rect 305840 242241 306160 242273
rect 311771 242829 312091 242861
rect 311771 242593 311813 242829
rect 312049 242593 312091 242829
rect 311771 242509 312091 242593
rect 311771 242273 311813 242509
rect 312049 242273 312091 242509
rect 311771 242241 312091 242273
rect 327910 242829 328230 242861
rect 327910 242593 327952 242829
rect 328188 242593 328230 242829
rect 327910 242509 328230 242593
rect 327910 242273 327952 242509
rect 328188 242273 328230 242509
rect 327910 242241 328230 242273
rect 333840 242829 334160 242861
rect 333840 242593 333882 242829
rect 334118 242593 334160 242829
rect 333840 242509 334160 242593
rect 333840 242273 333882 242509
rect 334118 242273 334160 242509
rect 333840 242241 334160 242273
rect 339771 242829 340091 242861
rect 339771 242593 339813 242829
rect 340049 242593 340091 242829
rect 339771 242509 340091 242593
rect 339771 242273 339813 242509
rect 340049 242273 340091 242509
rect 339771 242241 340091 242273
rect 355910 242829 356230 242861
rect 355910 242593 355952 242829
rect 356188 242593 356230 242829
rect 355910 242509 356230 242593
rect 355910 242273 355952 242509
rect 356188 242273 356230 242509
rect 355910 242241 356230 242273
rect 361840 242829 362160 242861
rect 361840 242593 361882 242829
rect 362118 242593 362160 242829
rect 361840 242509 362160 242593
rect 361840 242273 361882 242509
rect 362118 242273 362160 242509
rect 361840 242241 362160 242273
rect 367771 242829 368091 242861
rect 367771 242593 367813 242829
rect 368049 242593 368091 242829
rect 367771 242509 368091 242593
rect 367771 242273 367813 242509
rect 368049 242273 368091 242509
rect 367771 242241 368091 242273
rect 383910 242829 384230 242861
rect 383910 242593 383952 242829
rect 384188 242593 384230 242829
rect 383910 242509 384230 242593
rect 383910 242273 383952 242509
rect 384188 242273 384230 242509
rect 383910 242241 384230 242273
rect 389840 242829 390160 242861
rect 389840 242593 389882 242829
rect 390118 242593 390160 242829
rect 389840 242509 390160 242593
rect 389840 242273 389882 242509
rect 390118 242273 390160 242509
rect 389840 242241 390160 242273
rect 395771 242829 396091 242861
rect 395771 242593 395813 242829
rect 396049 242593 396091 242829
rect 395771 242509 396091 242593
rect 395771 242273 395813 242509
rect 396049 242273 396091 242509
rect 395771 242241 396091 242273
rect 411910 242829 412230 242861
rect 411910 242593 411952 242829
rect 412188 242593 412230 242829
rect 411910 242509 412230 242593
rect 411910 242273 411952 242509
rect 412188 242273 412230 242509
rect 411910 242241 412230 242273
rect 417840 242829 418160 242861
rect 417840 242593 417882 242829
rect 418118 242593 418160 242829
rect 417840 242509 418160 242593
rect 417840 242273 417882 242509
rect 418118 242273 418160 242509
rect 417840 242241 418160 242273
rect 423771 242829 424091 242861
rect 423771 242593 423813 242829
rect 424049 242593 424091 242829
rect 423771 242509 424091 242593
rect 423771 242273 423813 242509
rect 424049 242273 424091 242509
rect 423771 242241 424091 242273
rect 439910 242829 440230 242861
rect 439910 242593 439952 242829
rect 440188 242593 440230 242829
rect 439910 242509 440230 242593
rect 439910 242273 439952 242509
rect 440188 242273 440230 242509
rect 439910 242241 440230 242273
rect 445840 242829 446160 242861
rect 445840 242593 445882 242829
rect 446118 242593 446160 242829
rect 445840 242509 446160 242593
rect 445840 242273 445882 242509
rect 446118 242273 446160 242509
rect 445840 242241 446160 242273
rect 451771 242829 452091 242861
rect 451771 242593 451813 242829
rect 452049 242593 452091 242829
rect 451771 242509 452091 242593
rect 451771 242273 451813 242509
rect 452049 242273 452091 242509
rect 451771 242241 452091 242273
rect 467910 242829 468230 242861
rect 467910 242593 467952 242829
rect 468188 242593 468230 242829
rect 467910 242509 468230 242593
rect 467910 242273 467952 242509
rect 468188 242273 468230 242509
rect 467910 242241 468230 242273
rect 473840 242829 474160 242861
rect 473840 242593 473882 242829
rect 474118 242593 474160 242829
rect 473840 242509 474160 242593
rect 473840 242273 473882 242509
rect 474118 242273 474160 242509
rect 473840 242241 474160 242273
rect 479771 242829 480091 242861
rect 479771 242593 479813 242829
rect 480049 242593 480091 242829
rect 479771 242509 480091 242593
rect 479771 242273 479813 242509
rect 480049 242273 480091 242509
rect 479771 242241 480091 242273
rect 495910 242829 496230 242861
rect 495910 242593 495952 242829
rect 496188 242593 496230 242829
rect 495910 242509 496230 242593
rect 495910 242273 495952 242509
rect 496188 242273 496230 242509
rect 495910 242241 496230 242273
rect 501840 242829 502160 242861
rect 501840 242593 501882 242829
rect 502118 242593 502160 242829
rect 501840 242509 502160 242593
rect 501840 242273 501882 242509
rect 502118 242273 502160 242509
rect 501840 242241 502160 242273
rect 507771 242829 508091 242861
rect 507771 242593 507813 242829
rect 508049 242593 508091 242829
rect 507771 242509 508091 242593
rect 507771 242273 507813 242509
rect 508049 242273 508091 242509
rect 507771 242241 508091 242273
rect 523910 242829 524230 242861
rect 523910 242593 523952 242829
rect 524188 242593 524230 242829
rect 523910 242509 524230 242593
rect 523910 242273 523952 242509
rect 524188 242273 524230 242509
rect 523910 242241 524230 242273
rect 529840 242829 530160 242861
rect 529840 242593 529882 242829
rect 530118 242593 530160 242829
rect 529840 242509 530160 242593
rect 529840 242273 529882 242509
rect 530118 242273 530160 242509
rect 529840 242241 530160 242273
rect 535771 242829 536091 242861
rect 535771 242593 535813 242829
rect 536049 242593 536091 242829
rect 535771 242509 536091 242593
rect 535771 242273 535813 242509
rect 536049 242273 536091 242509
rect 535771 242241 536091 242273
rect 551910 242829 552230 242861
rect 551910 242593 551952 242829
rect 552188 242593 552230 242829
rect 551910 242509 552230 242593
rect 551910 242273 551952 242509
rect 552188 242273 552230 242509
rect 551910 242241 552230 242273
rect 557840 242829 558160 242861
rect 557840 242593 557882 242829
rect 558118 242593 558160 242829
rect 557840 242509 558160 242593
rect 557840 242273 557882 242509
rect 558118 242273 558160 242509
rect 557840 242241 558160 242273
rect 563771 242829 564091 242861
rect 563771 242593 563813 242829
rect 564049 242593 564091 242829
rect 563771 242509 564091 242593
rect 563771 242273 563813 242509
rect 564049 242273 564091 242509
rect 563771 242241 564091 242273
rect 573494 242829 574114 269273
rect 573494 242593 573526 242829
rect 573762 242593 573846 242829
rect 574082 242593 574114 242829
rect 573494 242509 574114 242593
rect 573494 242273 573526 242509
rect 573762 242273 573846 242509
rect 574082 242273 574114 242509
rect 22874 239454 23194 239486
rect 22874 239218 22916 239454
rect 23152 239218 23194 239454
rect 22874 239134 23194 239218
rect 22874 238898 22916 239134
rect 23152 238898 23194 239134
rect 22874 238866 23194 238898
rect 28805 239454 29125 239486
rect 28805 239218 28847 239454
rect 29083 239218 29125 239454
rect 28805 239134 29125 239218
rect 28805 238898 28847 239134
rect 29083 238898 29125 239134
rect 28805 238866 29125 238898
rect 50874 239454 51194 239486
rect 50874 239218 50916 239454
rect 51152 239218 51194 239454
rect 50874 239134 51194 239218
rect 50874 238898 50916 239134
rect 51152 238898 51194 239134
rect 50874 238866 51194 238898
rect 56805 239454 57125 239486
rect 56805 239218 56847 239454
rect 57083 239218 57125 239454
rect 56805 239134 57125 239218
rect 56805 238898 56847 239134
rect 57083 238898 57125 239134
rect 56805 238866 57125 238898
rect 78874 239454 79194 239486
rect 78874 239218 78916 239454
rect 79152 239218 79194 239454
rect 78874 239134 79194 239218
rect 78874 238898 78916 239134
rect 79152 238898 79194 239134
rect 78874 238866 79194 238898
rect 84805 239454 85125 239486
rect 84805 239218 84847 239454
rect 85083 239218 85125 239454
rect 84805 239134 85125 239218
rect 84805 238898 84847 239134
rect 85083 238898 85125 239134
rect 84805 238866 85125 238898
rect 106874 239454 107194 239486
rect 106874 239218 106916 239454
rect 107152 239218 107194 239454
rect 106874 239134 107194 239218
rect 106874 238898 106916 239134
rect 107152 238898 107194 239134
rect 106874 238866 107194 238898
rect 112805 239454 113125 239486
rect 112805 239218 112847 239454
rect 113083 239218 113125 239454
rect 112805 239134 113125 239218
rect 112805 238898 112847 239134
rect 113083 238898 113125 239134
rect 112805 238866 113125 238898
rect 134874 239454 135194 239486
rect 134874 239218 134916 239454
rect 135152 239218 135194 239454
rect 134874 239134 135194 239218
rect 134874 238898 134916 239134
rect 135152 238898 135194 239134
rect 134874 238866 135194 238898
rect 140805 239454 141125 239486
rect 140805 239218 140847 239454
rect 141083 239218 141125 239454
rect 140805 239134 141125 239218
rect 140805 238898 140847 239134
rect 141083 238898 141125 239134
rect 140805 238866 141125 238898
rect 162874 239454 163194 239486
rect 162874 239218 162916 239454
rect 163152 239218 163194 239454
rect 162874 239134 163194 239218
rect 162874 238898 162916 239134
rect 163152 238898 163194 239134
rect 162874 238866 163194 238898
rect 168805 239454 169125 239486
rect 168805 239218 168847 239454
rect 169083 239218 169125 239454
rect 168805 239134 169125 239218
rect 168805 238898 168847 239134
rect 169083 238898 169125 239134
rect 168805 238866 169125 238898
rect 190874 239454 191194 239486
rect 190874 239218 190916 239454
rect 191152 239218 191194 239454
rect 190874 239134 191194 239218
rect 190874 238898 190916 239134
rect 191152 238898 191194 239134
rect 190874 238866 191194 238898
rect 196805 239454 197125 239486
rect 196805 239218 196847 239454
rect 197083 239218 197125 239454
rect 196805 239134 197125 239218
rect 196805 238898 196847 239134
rect 197083 238898 197125 239134
rect 196805 238866 197125 238898
rect 218874 239454 219194 239486
rect 218874 239218 218916 239454
rect 219152 239218 219194 239454
rect 218874 239134 219194 239218
rect 218874 238898 218916 239134
rect 219152 238898 219194 239134
rect 218874 238866 219194 238898
rect 224805 239454 225125 239486
rect 224805 239218 224847 239454
rect 225083 239218 225125 239454
rect 224805 239134 225125 239218
rect 224805 238898 224847 239134
rect 225083 238898 225125 239134
rect 224805 238866 225125 238898
rect 246874 239454 247194 239486
rect 246874 239218 246916 239454
rect 247152 239218 247194 239454
rect 246874 239134 247194 239218
rect 246874 238898 246916 239134
rect 247152 238898 247194 239134
rect 246874 238866 247194 238898
rect 252805 239454 253125 239486
rect 252805 239218 252847 239454
rect 253083 239218 253125 239454
rect 252805 239134 253125 239218
rect 252805 238898 252847 239134
rect 253083 238898 253125 239134
rect 252805 238866 253125 238898
rect 274874 239454 275194 239486
rect 274874 239218 274916 239454
rect 275152 239218 275194 239454
rect 274874 239134 275194 239218
rect 274874 238898 274916 239134
rect 275152 238898 275194 239134
rect 274874 238866 275194 238898
rect 280805 239454 281125 239486
rect 280805 239218 280847 239454
rect 281083 239218 281125 239454
rect 280805 239134 281125 239218
rect 280805 238898 280847 239134
rect 281083 238898 281125 239134
rect 280805 238866 281125 238898
rect 302874 239454 303194 239486
rect 302874 239218 302916 239454
rect 303152 239218 303194 239454
rect 302874 239134 303194 239218
rect 302874 238898 302916 239134
rect 303152 238898 303194 239134
rect 302874 238866 303194 238898
rect 308805 239454 309125 239486
rect 308805 239218 308847 239454
rect 309083 239218 309125 239454
rect 308805 239134 309125 239218
rect 308805 238898 308847 239134
rect 309083 238898 309125 239134
rect 308805 238866 309125 238898
rect 330874 239454 331194 239486
rect 330874 239218 330916 239454
rect 331152 239218 331194 239454
rect 330874 239134 331194 239218
rect 330874 238898 330916 239134
rect 331152 238898 331194 239134
rect 330874 238866 331194 238898
rect 336805 239454 337125 239486
rect 336805 239218 336847 239454
rect 337083 239218 337125 239454
rect 336805 239134 337125 239218
rect 336805 238898 336847 239134
rect 337083 238898 337125 239134
rect 336805 238866 337125 238898
rect 358874 239454 359194 239486
rect 358874 239218 358916 239454
rect 359152 239218 359194 239454
rect 358874 239134 359194 239218
rect 358874 238898 358916 239134
rect 359152 238898 359194 239134
rect 358874 238866 359194 238898
rect 364805 239454 365125 239486
rect 364805 239218 364847 239454
rect 365083 239218 365125 239454
rect 364805 239134 365125 239218
rect 364805 238898 364847 239134
rect 365083 238898 365125 239134
rect 364805 238866 365125 238898
rect 386874 239454 387194 239486
rect 386874 239218 386916 239454
rect 387152 239218 387194 239454
rect 386874 239134 387194 239218
rect 386874 238898 386916 239134
rect 387152 238898 387194 239134
rect 386874 238866 387194 238898
rect 392805 239454 393125 239486
rect 392805 239218 392847 239454
rect 393083 239218 393125 239454
rect 392805 239134 393125 239218
rect 392805 238898 392847 239134
rect 393083 238898 393125 239134
rect 392805 238866 393125 238898
rect 414874 239454 415194 239486
rect 414874 239218 414916 239454
rect 415152 239218 415194 239454
rect 414874 239134 415194 239218
rect 414874 238898 414916 239134
rect 415152 238898 415194 239134
rect 414874 238866 415194 238898
rect 420805 239454 421125 239486
rect 420805 239218 420847 239454
rect 421083 239218 421125 239454
rect 420805 239134 421125 239218
rect 420805 238898 420847 239134
rect 421083 238898 421125 239134
rect 420805 238866 421125 238898
rect 442874 239454 443194 239486
rect 442874 239218 442916 239454
rect 443152 239218 443194 239454
rect 442874 239134 443194 239218
rect 442874 238898 442916 239134
rect 443152 238898 443194 239134
rect 442874 238866 443194 238898
rect 448805 239454 449125 239486
rect 448805 239218 448847 239454
rect 449083 239218 449125 239454
rect 448805 239134 449125 239218
rect 448805 238898 448847 239134
rect 449083 238898 449125 239134
rect 448805 238866 449125 238898
rect 470874 239454 471194 239486
rect 470874 239218 470916 239454
rect 471152 239218 471194 239454
rect 470874 239134 471194 239218
rect 470874 238898 470916 239134
rect 471152 238898 471194 239134
rect 470874 238866 471194 238898
rect 476805 239454 477125 239486
rect 476805 239218 476847 239454
rect 477083 239218 477125 239454
rect 476805 239134 477125 239218
rect 476805 238898 476847 239134
rect 477083 238898 477125 239134
rect 476805 238866 477125 238898
rect 498874 239454 499194 239486
rect 498874 239218 498916 239454
rect 499152 239218 499194 239454
rect 498874 239134 499194 239218
rect 498874 238898 498916 239134
rect 499152 238898 499194 239134
rect 498874 238866 499194 238898
rect 504805 239454 505125 239486
rect 504805 239218 504847 239454
rect 505083 239218 505125 239454
rect 504805 239134 505125 239218
rect 504805 238898 504847 239134
rect 505083 238898 505125 239134
rect 504805 238866 505125 238898
rect 526874 239454 527194 239486
rect 526874 239218 526916 239454
rect 527152 239218 527194 239454
rect 526874 239134 527194 239218
rect 526874 238898 526916 239134
rect 527152 238898 527194 239134
rect 526874 238866 527194 238898
rect 532805 239454 533125 239486
rect 532805 239218 532847 239454
rect 533083 239218 533125 239454
rect 532805 239134 533125 239218
rect 532805 238898 532847 239134
rect 533083 238898 533125 239134
rect 532805 238866 533125 238898
rect 554874 239454 555194 239486
rect 554874 239218 554916 239454
rect 555152 239218 555194 239454
rect 554874 239134 555194 239218
rect 554874 238898 554916 239134
rect 555152 238898 555194 239134
rect 554874 238866 555194 238898
rect 560805 239454 561125 239486
rect 560805 239218 560847 239454
rect 561083 239218 561125 239454
rect 560805 239134 561125 239218
rect 560805 238898 560847 239134
rect 561083 238898 561125 239134
rect 560805 238866 561125 238898
rect -2006 215593 -1974 215829
rect -1738 215593 -1654 215829
rect -1418 215593 -1386 215829
rect -2006 215509 -1386 215593
rect -2006 215273 -1974 215509
rect -1738 215273 -1654 215509
rect -1418 215273 -1386 215509
rect -2006 188829 -1386 215273
rect 19909 215829 20229 215861
rect 19909 215593 19951 215829
rect 20187 215593 20229 215829
rect 19909 215509 20229 215593
rect 19909 215273 19951 215509
rect 20187 215273 20229 215509
rect 19909 215241 20229 215273
rect 25840 215829 26160 215861
rect 25840 215593 25882 215829
rect 26118 215593 26160 215829
rect 25840 215509 26160 215593
rect 25840 215273 25882 215509
rect 26118 215273 26160 215509
rect 25840 215241 26160 215273
rect 31770 215829 32090 215861
rect 31770 215593 31812 215829
rect 32048 215593 32090 215829
rect 31770 215509 32090 215593
rect 31770 215273 31812 215509
rect 32048 215273 32090 215509
rect 31770 215241 32090 215273
rect 47909 215829 48229 215861
rect 47909 215593 47951 215829
rect 48187 215593 48229 215829
rect 47909 215509 48229 215593
rect 47909 215273 47951 215509
rect 48187 215273 48229 215509
rect 47909 215241 48229 215273
rect 53840 215829 54160 215861
rect 53840 215593 53882 215829
rect 54118 215593 54160 215829
rect 53840 215509 54160 215593
rect 53840 215273 53882 215509
rect 54118 215273 54160 215509
rect 53840 215241 54160 215273
rect 59770 215829 60090 215861
rect 59770 215593 59812 215829
rect 60048 215593 60090 215829
rect 59770 215509 60090 215593
rect 59770 215273 59812 215509
rect 60048 215273 60090 215509
rect 59770 215241 60090 215273
rect 75909 215829 76229 215861
rect 75909 215593 75951 215829
rect 76187 215593 76229 215829
rect 75909 215509 76229 215593
rect 75909 215273 75951 215509
rect 76187 215273 76229 215509
rect 75909 215241 76229 215273
rect 81840 215829 82160 215861
rect 81840 215593 81882 215829
rect 82118 215593 82160 215829
rect 81840 215509 82160 215593
rect 81840 215273 81882 215509
rect 82118 215273 82160 215509
rect 81840 215241 82160 215273
rect 87770 215829 88090 215861
rect 87770 215593 87812 215829
rect 88048 215593 88090 215829
rect 87770 215509 88090 215593
rect 87770 215273 87812 215509
rect 88048 215273 88090 215509
rect 87770 215241 88090 215273
rect 103909 215829 104229 215861
rect 103909 215593 103951 215829
rect 104187 215593 104229 215829
rect 103909 215509 104229 215593
rect 103909 215273 103951 215509
rect 104187 215273 104229 215509
rect 103909 215241 104229 215273
rect 109840 215829 110160 215861
rect 109840 215593 109882 215829
rect 110118 215593 110160 215829
rect 109840 215509 110160 215593
rect 109840 215273 109882 215509
rect 110118 215273 110160 215509
rect 109840 215241 110160 215273
rect 115770 215829 116090 215861
rect 115770 215593 115812 215829
rect 116048 215593 116090 215829
rect 115770 215509 116090 215593
rect 115770 215273 115812 215509
rect 116048 215273 116090 215509
rect 115770 215241 116090 215273
rect 131909 215829 132229 215861
rect 131909 215593 131951 215829
rect 132187 215593 132229 215829
rect 131909 215509 132229 215593
rect 131909 215273 131951 215509
rect 132187 215273 132229 215509
rect 131909 215241 132229 215273
rect 137840 215829 138160 215861
rect 137840 215593 137882 215829
rect 138118 215593 138160 215829
rect 137840 215509 138160 215593
rect 137840 215273 137882 215509
rect 138118 215273 138160 215509
rect 137840 215241 138160 215273
rect 143770 215829 144090 215861
rect 143770 215593 143812 215829
rect 144048 215593 144090 215829
rect 143770 215509 144090 215593
rect 143770 215273 143812 215509
rect 144048 215273 144090 215509
rect 143770 215241 144090 215273
rect 159909 215829 160229 215861
rect 159909 215593 159951 215829
rect 160187 215593 160229 215829
rect 159909 215509 160229 215593
rect 159909 215273 159951 215509
rect 160187 215273 160229 215509
rect 159909 215241 160229 215273
rect 165840 215829 166160 215861
rect 165840 215593 165882 215829
rect 166118 215593 166160 215829
rect 165840 215509 166160 215593
rect 165840 215273 165882 215509
rect 166118 215273 166160 215509
rect 165840 215241 166160 215273
rect 171770 215829 172090 215861
rect 171770 215593 171812 215829
rect 172048 215593 172090 215829
rect 171770 215509 172090 215593
rect 171770 215273 171812 215509
rect 172048 215273 172090 215509
rect 171770 215241 172090 215273
rect 187909 215829 188229 215861
rect 187909 215593 187951 215829
rect 188187 215593 188229 215829
rect 187909 215509 188229 215593
rect 187909 215273 187951 215509
rect 188187 215273 188229 215509
rect 187909 215241 188229 215273
rect 193840 215829 194160 215861
rect 193840 215593 193882 215829
rect 194118 215593 194160 215829
rect 193840 215509 194160 215593
rect 193840 215273 193882 215509
rect 194118 215273 194160 215509
rect 193840 215241 194160 215273
rect 199770 215829 200090 215861
rect 199770 215593 199812 215829
rect 200048 215593 200090 215829
rect 199770 215509 200090 215593
rect 199770 215273 199812 215509
rect 200048 215273 200090 215509
rect 199770 215241 200090 215273
rect 215909 215829 216229 215861
rect 215909 215593 215951 215829
rect 216187 215593 216229 215829
rect 215909 215509 216229 215593
rect 215909 215273 215951 215509
rect 216187 215273 216229 215509
rect 215909 215241 216229 215273
rect 221840 215829 222160 215861
rect 221840 215593 221882 215829
rect 222118 215593 222160 215829
rect 221840 215509 222160 215593
rect 221840 215273 221882 215509
rect 222118 215273 222160 215509
rect 221840 215241 222160 215273
rect 227770 215829 228090 215861
rect 227770 215593 227812 215829
rect 228048 215593 228090 215829
rect 227770 215509 228090 215593
rect 227770 215273 227812 215509
rect 228048 215273 228090 215509
rect 227770 215241 228090 215273
rect 243909 215829 244229 215861
rect 243909 215593 243951 215829
rect 244187 215593 244229 215829
rect 243909 215509 244229 215593
rect 243909 215273 243951 215509
rect 244187 215273 244229 215509
rect 243909 215241 244229 215273
rect 249840 215829 250160 215861
rect 249840 215593 249882 215829
rect 250118 215593 250160 215829
rect 249840 215509 250160 215593
rect 249840 215273 249882 215509
rect 250118 215273 250160 215509
rect 249840 215241 250160 215273
rect 255770 215829 256090 215861
rect 255770 215593 255812 215829
rect 256048 215593 256090 215829
rect 255770 215509 256090 215593
rect 255770 215273 255812 215509
rect 256048 215273 256090 215509
rect 255770 215241 256090 215273
rect 271909 215829 272229 215861
rect 271909 215593 271951 215829
rect 272187 215593 272229 215829
rect 271909 215509 272229 215593
rect 271909 215273 271951 215509
rect 272187 215273 272229 215509
rect 271909 215241 272229 215273
rect 277840 215829 278160 215861
rect 277840 215593 277882 215829
rect 278118 215593 278160 215829
rect 277840 215509 278160 215593
rect 277840 215273 277882 215509
rect 278118 215273 278160 215509
rect 277840 215241 278160 215273
rect 283770 215829 284090 215861
rect 283770 215593 283812 215829
rect 284048 215593 284090 215829
rect 283770 215509 284090 215593
rect 283770 215273 283812 215509
rect 284048 215273 284090 215509
rect 283770 215241 284090 215273
rect 299909 215829 300229 215861
rect 299909 215593 299951 215829
rect 300187 215593 300229 215829
rect 299909 215509 300229 215593
rect 299909 215273 299951 215509
rect 300187 215273 300229 215509
rect 299909 215241 300229 215273
rect 305840 215829 306160 215861
rect 305840 215593 305882 215829
rect 306118 215593 306160 215829
rect 305840 215509 306160 215593
rect 305840 215273 305882 215509
rect 306118 215273 306160 215509
rect 305840 215241 306160 215273
rect 311770 215829 312090 215861
rect 311770 215593 311812 215829
rect 312048 215593 312090 215829
rect 311770 215509 312090 215593
rect 311770 215273 311812 215509
rect 312048 215273 312090 215509
rect 311770 215241 312090 215273
rect 327909 215829 328229 215861
rect 327909 215593 327951 215829
rect 328187 215593 328229 215829
rect 327909 215509 328229 215593
rect 327909 215273 327951 215509
rect 328187 215273 328229 215509
rect 327909 215241 328229 215273
rect 333840 215829 334160 215861
rect 333840 215593 333882 215829
rect 334118 215593 334160 215829
rect 333840 215509 334160 215593
rect 333840 215273 333882 215509
rect 334118 215273 334160 215509
rect 333840 215241 334160 215273
rect 339770 215829 340090 215861
rect 339770 215593 339812 215829
rect 340048 215593 340090 215829
rect 339770 215509 340090 215593
rect 339770 215273 339812 215509
rect 340048 215273 340090 215509
rect 339770 215241 340090 215273
rect 355909 215829 356229 215861
rect 355909 215593 355951 215829
rect 356187 215593 356229 215829
rect 355909 215509 356229 215593
rect 355909 215273 355951 215509
rect 356187 215273 356229 215509
rect 355909 215241 356229 215273
rect 361840 215829 362160 215861
rect 361840 215593 361882 215829
rect 362118 215593 362160 215829
rect 361840 215509 362160 215593
rect 361840 215273 361882 215509
rect 362118 215273 362160 215509
rect 361840 215241 362160 215273
rect 367770 215829 368090 215861
rect 367770 215593 367812 215829
rect 368048 215593 368090 215829
rect 367770 215509 368090 215593
rect 367770 215273 367812 215509
rect 368048 215273 368090 215509
rect 367770 215241 368090 215273
rect 383909 215829 384229 215861
rect 383909 215593 383951 215829
rect 384187 215593 384229 215829
rect 383909 215509 384229 215593
rect 383909 215273 383951 215509
rect 384187 215273 384229 215509
rect 383909 215241 384229 215273
rect 389840 215829 390160 215861
rect 389840 215593 389882 215829
rect 390118 215593 390160 215829
rect 389840 215509 390160 215593
rect 389840 215273 389882 215509
rect 390118 215273 390160 215509
rect 389840 215241 390160 215273
rect 395770 215829 396090 215861
rect 395770 215593 395812 215829
rect 396048 215593 396090 215829
rect 395770 215509 396090 215593
rect 395770 215273 395812 215509
rect 396048 215273 396090 215509
rect 395770 215241 396090 215273
rect 411909 215829 412229 215861
rect 411909 215593 411951 215829
rect 412187 215593 412229 215829
rect 411909 215509 412229 215593
rect 411909 215273 411951 215509
rect 412187 215273 412229 215509
rect 411909 215241 412229 215273
rect 417840 215829 418160 215861
rect 417840 215593 417882 215829
rect 418118 215593 418160 215829
rect 417840 215509 418160 215593
rect 417840 215273 417882 215509
rect 418118 215273 418160 215509
rect 417840 215241 418160 215273
rect 423770 215829 424090 215861
rect 423770 215593 423812 215829
rect 424048 215593 424090 215829
rect 423770 215509 424090 215593
rect 423770 215273 423812 215509
rect 424048 215273 424090 215509
rect 423770 215241 424090 215273
rect 439909 215829 440229 215861
rect 439909 215593 439951 215829
rect 440187 215593 440229 215829
rect 439909 215509 440229 215593
rect 439909 215273 439951 215509
rect 440187 215273 440229 215509
rect 439909 215241 440229 215273
rect 445840 215829 446160 215861
rect 445840 215593 445882 215829
rect 446118 215593 446160 215829
rect 445840 215509 446160 215593
rect 445840 215273 445882 215509
rect 446118 215273 446160 215509
rect 445840 215241 446160 215273
rect 451770 215829 452090 215861
rect 451770 215593 451812 215829
rect 452048 215593 452090 215829
rect 451770 215509 452090 215593
rect 451770 215273 451812 215509
rect 452048 215273 452090 215509
rect 451770 215241 452090 215273
rect 467909 215829 468229 215861
rect 467909 215593 467951 215829
rect 468187 215593 468229 215829
rect 467909 215509 468229 215593
rect 467909 215273 467951 215509
rect 468187 215273 468229 215509
rect 467909 215241 468229 215273
rect 473840 215829 474160 215861
rect 473840 215593 473882 215829
rect 474118 215593 474160 215829
rect 473840 215509 474160 215593
rect 473840 215273 473882 215509
rect 474118 215273 474160 215509
rect 473840 215241 474160 215273
rect 479770 215829 480090 215861
rect 479770 215593 479812 215829
rect 480048 215593 480090 215829
rect 479770 215509 480090 215593
rect 479770 215273 479812 215509
rect 480048 215273 480090 215509
rect 479770 215241 480090 215273
rect 495909 215829 496229 215861
rect 495909 215593 495951 215829
rect 496187 215593 496229 215829
rect 495909 215509 496229 215593
rect 495909 215273 495951 215509
rect 496187 215273 496229 215509
rect 495909 215241 496229 215273
rect 501840 215829 502160 215861
rect 501840 215593 501882 215829
rect 502118 215593 502160 215829
rect 501840 215509 502160 215593
rect 501840 215273 501882 215509
rect 502118 215273 502160 215509
rect 501840 215241 502160 215273
rect 507770 215829 508090 215861
rect 507770 215593 507812 215829
rect 508048 215593 508090 215829
rect 507770 215509 508090 215593
rect 507770 215273 507812 215509
rect 508048 215273 508090 215509
rect 507770 215241 508090 215273
rect 523909 215829 524229 215861
rect 523909 215593 523951 215829
rect 524187 215593 524229 215829
rect 523909 215509 524229 215593
rect 523909 215273 523951 215509
rect 524187 215273 524229 215509
rect 523909 215241 524229 215273
rect 529840 215829 530160 215861
rect 529840 215593 529882 215829
rect 530118 215593 530160 215829
rect 529840 215509 530160 215593
rect 529840 215273 529882 215509
rect 530118 215273 530160 215509
rect 529840 215241 530160 215273
rect 535770 215829 536090 215861
rect 535770 215593 535812 215829
rect 536048 215593 536090 215829
rect 535770 215509 536090 215593
rect 535770 215273 535812 215509
rect 536048 215273 536090 215509
rect 535770 215241 536090 215273
rect 551909 215829 552229 215861
rect 551909 215593 551951 215829
rect 552187 215593 552229 215829
rect 551909 215509 552229 215593
rect 551909 215273 551951 215509
rect 552187 215273 552229 215509
rect 551909 215241 552229 215273
rect 557840 215829 558160 215861
rect 557840 215593 557882 215829
rect 558118 215593 558160 215829
rect 557840 215509 558160 215593
rect 557840 215273 557882 215509
rect 558118 215273 558160 215509
rect 557840 215241 558160 215273
rect 563770 215829 564090 215861
rect 563770 215593 563812 215829
rect 564048 215593 564090 215829
rect 563770 215509 564090 215593
rect 563770 215273 563812 215509
rect 564048 215273 564090 215509
rect 563770 215241 564090 215273
rect 573494 215829 574114 242273
rect 573494 215593 573526 215829
rect 573762 215593 573846 215829
rect 574082 215593 574114 215829
rect 573494 215509 574114 215593
rect 573494 215273 573526 215509
rect 573762 215273 573846 215509
rect 574082 215273 574114 215509
rect 22875 212454 23195 212486
rect 22875 212218 22917 212454
rect 23153 212218 23195 212454
rect 22875 212134 23195 212218
rect 22875 211898 22917 212134
rect 23153 211898 23195 212134
rect 22875 211866 23195 211898
rect 28806 212454 29126 212486
rect 28806 212218 28848 212454
rect 29084 212218 29126 212454
rect 28806 212134 29126 212218
rect 28806 211898 28848 212134
rect 29084 211898 29126 212134
rect 28806 211866 29126 211898
rect 50875 212454 51195 212486
rect 50875 212218 50917 212454
rect 51153 212218 51195 212454
rect 50875 212134 51195 212218
rect 50875 211898 50917 212134
rect 51153 211898 51195 212134
rect 50875 211866 51195 211898
rect 56806 212454 57126 212486
rect 56806 212218 56848 212454
rect 57084 212218 57126 212454
rect 56806 212134 57126 212218
rect 56806 211898 56848 212134
rect 57084 211898 57126 212134
rect 56806 211866 57126 211898
rect 78875 212454 79195 212486
rect 78875 212218 78917 212454
rect 79153 212218 79195 212454
rect 78875 212134 79195 212218
rect 78875 211898 78917 212134
rect 79153 211898 79195 212134
rect 78875 211866 79195 211898
rect 84806 212454 85126 212486
rect 84806 212218 84848 212454
rect 85084 212218 85126 212454
rect 84806 212134 85126 212218
rect 84806 211898 84848 212134
rect 85084 211898 85126 212134
rect 84806 211866 85126 211898
rect 106875 212454 107195 212486
rect 106875 212218 106917 212454
rect 107153 212218 107195 212454
rect 106875 212134 107195 212218
rect 106875 211898 106917 212134
rect 107153 211898 107195 212134
rect 106875 211866 107195 211898
rect 112806 212454 113126 212486
rect 112806 212218 112848 212454
rect 113084 212218 113126 212454
rect 112806 212134 113126 212218
rect 112806 211898 112848 212134
rect 113084 211898 113126 212134
rect 112806 211866 113126 211898
rect 134875 212454 135195 212486
rect 134875 212218 134917 212454
rect 135153 212218 135195 212454
rect 134875 212134 135195 212218
rect 134875 211898 134917 212134
rect 135153 211898 135195 212134
rect 134875 211866 135195 211898
rect 140806 212454 141126 212486
rect 140806 212218 140848 212454
rect 141084 212218 141126 212454
rect 140806 212134 141126 212218
rect 140806 211898 140848 212134
rect 141084 211898 141126 212134
rect 140806 211866 141126 211898
rect 162875 212454 163195 212486
rect 162875 212218 162917 212454
rect 163153 212218 163195 212454
rect 162875 212134 163195 212218
rect 162875 211898 162917 212134
rect 163153 211898 163195 212134
rect 162875 211866 163195 211898
rect 168806 212454 169126 212486
rect 168806 212218 168848 212454
rect 169084 212218 169126 212454
rect 168806 212134 169126 212218
rect 168806 211898 168848 212134
rect 169084 211898 169126 212134
rect 168806 211866 169126 211898
rect 190875 212454 191195 212486
rect 190875 212218 190917 212454
rect 191153 212218 191195 212454
rect 190875 212134 191195 212218
rect 190875 211898 190917 212134
rect 191153 211898 191195 212134
rect 190875 211866 191195 211898
rect 196806 212454 197126 212486
rect 196806 212218 196848 212454
rect 197084 212218 197126 212454
rect 196806 212134 197126 212218
rect 196806 211898 196848 212134
rect 197084 211898 197126 212134
rect 196806 211866 197126 211898
rect 218875 212454 219195 212486
rect 218875 212218 218917 212454
rect 219153 212218 219195 212454
rect 218875 212134 219195 212218
rect 218875 211898 218917 212134
rect 219153 211898 219195 212134
rect 218875 211866 219195 211898
rect 224806 212454 225126 212486
rect 224806 212218 224848 212454
rect 225084 212218 225126 212454
rect 224806 212134 225126 212218
rect 224806 211898 224848 212134
rect 225084 211898 225126 212134
rect 224806 211866 225126 211898
rect 246875 212454 247195 212486
rect 246875 212218 246917 212454
rect 247153 212218 247195 212454
rect 246875 212134 247195 212218
rect 246875 211898 246917 212134
rect 247153 211898 247195 212134
rect 246875 211866 247195 211898
rect 252806 212454 253126 212486
rect 252806 212218 252848 212454
rect 253084 212218 253126 212454
rect 252806 212134 253126 212218
rect 252806 211898 252848 212134
rect 253084 211898 253126 212134
rect 252806 211866 253126 211898
rect 274875 212454 275195 212486
rect 274875 212218 274917 212454
rect 275153 212218 275195 212454
rect 274875 212134 275195 212218
rect 274875 211898 274917 212134
rect 275153 211898 275195 212134
rect 274875 211866 275195 211898
rect 280806 212454 281126 212486
rect 280806 212218 280848 212454
rect 281084 212218 281126 212454
rect 280806 212134 281126 212218
rect 280806 211898 280848 212134
rect 281084 211898 281126 212134
rect 280806 211866 281126 211898
rect 302875 212454 303195 212486
rect 302875 212218 302917 212454
rect 303153 212218 303195 212454
rect 302875 212134 303195 212218
rect 302875 211898 302917 212134
rect 303153 211898 303195 212134
rect 302875 211866 303195 211898
rect 308806 212454 309126 212486
rect 308806 212218 308848 212454
rect 309084 212218 309126 212454
rect 308806 212134 309126 212218
rect 308806 211898 308848 212134
rect 309084 211898 309126 212134
rect 308806 211866 309126 211898
rect 330875 212454 331195 212486
rect 330875 212218 330917 212454
rect 331153 212218 331195 212454
rect 330875 212134 331195 212218
rect 330875 211898 330917 212134
rect 331153 211898 331195 212134
rect 330875 211866 331195 211898
rect 336806 212454 337126 212486
rect 336806 212218 336848 212454
rect 337084 212218 337126 212454
rect 336806 212134 337126 212218
rect 336806 211898 336848 212134
rect 337084 211898 337126 212134
rect 336806 211866 337126 211898
rect 358875 212454 359195 212486
rect 358875 212218 358917 212454
rect 359153 212218 359195 212454
rect 358875 212134 359195 212218
rect 358875 211898 358917 212134
rect 359153 211898 359195 212134
rect 358875 211866 359195 211898
rect 364806 212454 365126 212486
rect 364806 212218 364848 212454
rect 365084 212218 365126 212454
rect 364806 212134 365126 212218
rect 364806 211898 364848 212134
rect 365084 211898 365126 212134
rect 364806 211866 365126 211898
rect 386875 212454 387195 212486
rect 386875 212218 386917 212454
rect 387153 212218 387195 212454
rect 386875 212134 387195 212218
rect 386875 211898 386917 212134
rect 387153 211898 387195 212134
rect 386875 211866 387195 211898
rect 392806 212454 393126 212486
rect 392806 212218 392848 212454
rect 393084 212218 393126 212454
rect 392806 212134 393126 212218
rect 392806 211898 392848 212134
rect 393084 211898 393126 212134
rect 392806 211866 393126 211898
rect 414875 212454 415195 212486
rect 414875 212218 414917 212454
rect 415153 212218 415195 212454
rect 414875 212134 415195 212218
rect 414875 211898 414917 212134
rect 415153 211898 415195 212134
rect 414875 211866 415195 211898
rect 420806 212454 421126 212486
rect 420806 212218 420848 212454
rect 421084 212218 421126 212454
rect 420806 212134 421126 212218
rect 420806 211898 420848 212134
rect 421084 211898 421126 212134
rect 420806 211866 421126 211898
rect 442875 212454 443195 212486
rect 442875 212218 442917 212454
rect 443153 212218 443195 212454
rect 442875 212134 443195 212218
rect 442875 211898 442917 212134
rect 443153 211898 443195 212134
rect 442875 211866 443195 211898
rect 448806 212454 449126 212486
rect 448806 212218 448848 212454
rect 449084 212218 449126 212454
rect 448806 212134 449126 212218
rect 448806 211898 448848 212134
rect 449084 211898 449126 212134
rect 448806 211866 449126 211898
rect 470875 212454 471195 212486
rect 470875 212218 470917 212454
rect 471153 212218 471195 212454
rect 470875 212134 471195 212218
rect 470875 211898 470917 212134
rect 471153 211898 471195 212134
rect 470875 211866 471195 211898
rect 476806 212454 477126 212486
rect 476806 212218 476848 212454
rect 477084 212218 477126 212454
rect 476806 212134 477126 212218
rect 476806 211898 476848 212134
rect 477084 211898 477126 212134
rect 476806 211866 477126 211898
rect 498875 212454 499195 212486
rect 498875 212218 498917 212454
rect 499153 212218 499195 212454
rect 498875 212134 499195 212218
rect 498875 211898 498917 212134
rect 499153 211898 499195 212134
rect 498875 211866 499195 211898
rect 504806 212454 505126 212486
rect 504806 212218 504848 212454
rect 505084 212218 505126 212454
rect 504806 212134 505126 212218
rect 504806 211898 504848 212134
rect 505084 211898 505126 212134
rect 504806 211866 505126 211898
rect 526875 212454 527195 212486
rect 526875 212218 526917 212454
rect 527153 212218 527195 212454
rect 526875 212134 527195 212218
rect 526875 211898 526917 212134
rect 527153 211898 527195 212134
rect 526875 211866 527195 211898
rect 532806 212454 533126 212486
rect 532806 212218 532848 212454
rect 533084 212218 533126 212454
rect 532806 212134 533126 212218
rect 532806 211898 532848 212134
rect 533084 211898 533126 212134
rect 532806 211866 533126 211898
rect 554875 212454 555195 212486
rect 554875 212218 554917 212454
rect 555153 212218 555195 212454
rect 554875 212134 555195 212218
rect 554875 211898 554917 212134
rect 555153 211898 555195 212134
rect 554875 211866 555195 211898
rect 560806 212454 561126 212486
rect 560806 212218 560848 212454
rect 561084 212218 561126 212454
rect 560806 212134 561126 212218
rect 560806 211898 560848 212134
rect 561084 211898 561126 212134
rect 560806 211866 561126 211898
rect -2006 188593 -1974 188829
rect -1738 188593 -1654 188829
rect -1418 188593 -1386 188829
rect -2006 188509 -1386 188593
rect -2006 188273 -1974 188509
rect -1738 188273 -1654 188509
rect -1418 188273 -1386 188509
rect -2006 161829 -1386 188273
rect 19910 188829 20230 188861
rect 19910 188593 19952 188829
rect 20188 188593 20230 188829
rect 19910 188509 20230 188593
rect 19910 188273 19952 188509
rect 20188 188273 20230 188509
rect 19910 188241 20230 188273
rect 25840 188829 26160 188861
rect 25840 188593 25882 188829
rect 26118 188593 26160 188829
rect 25840 188509 26160 188593
rect 25840 188273 25882 188509
rect 26118 188273 26160 188509
rect 25840 188241 26160 188273
rect 31771 188829 32091 188861
rect 31771 188593 31813 188829
rect 32049 188593 32091 188829
rect 31771 188509 32091 188593
rect 31771 188273 31813 188509
rect 32049 188273 32091 188509
rect 31771 188241 32091 188273
rect 47910 188829 48230 188861
rect 47910 188593 47952 188829
rect 48188 188593 48230 188829
rect 47910 188509 48230 188593
rect 47910 188273 47952 188509
rect 48188 188273 48230 188509
rect 47910 188241 48230 188273
rect 53840 188829 54160 188861
rect 53840 188593 53882 188829
rect 54118 188593 54160 188829
rect 53840 188509 54160 188593
rect 53840 188273 53882 188509
rect 54118 188273 54160 188509
rect 53840 188241 54160 188273
rect 59771 188829 60091 188861
rect 59771 188593 59813 188829
rect 60049 188593 60091 188829
rect 59771 188509 60091 188593
rect 59771 188273 59813 188509
rect 60049 188273 60091 188509
rect 59771 188241 60091 188273
rect 75910 188829 76230 188861
rect 75910 188593 75952 188829
rect 76188 188593 76230 188829
rect 75910 188509 76230 188593
rect 75910 188273 75952 188509
rect 76188 188273 76230 188509
rect 75910 188241 76230 188273
rect 81840 188829 82160 188861
rect 81840 188593 81882 188829
rect 82118 188593 82160 188829
rect 81840 188509 82160 188593
rect 81840 188273 81882 188509
rect 82118 188273 82160 188509
rect 81840 188241 82160 188273
rect 87771 188829 88091 188861
rect 87771 188593 87813 188829
rect 88049 188593 88091 188829
rect 87771 188509 88091 188593
rect 87771 188273 87813 188509
rect 88049 188273 88091 188509
rect 87771 188241 88091 188273
rect 103910 188829 104230 188861
rect 103910 188593 103952 188829
rect 104188 188593 104230 188829
rect 103910 188509 104230 188593
rect 103910 188273 103952 188509
rect 104188 188273 104230 188509
rect 103910 188241 104230 188273
rect 109840 188829 110160 188861
rect 109840 188593 109882 188829
rect 110118 188593 110160 188829
rect 109840 188509 110160 188593
rect 109840 188273 109882 188509
rect 110118 188273 110160 188509
rect 109840 188241 110160 188273
rect 115771 188829 116091 188861
rect 115771 188593 115813 188829
rect 116049 188593 116091 188829
rect 115771 188509 116091 188593
rect 115771 188273 115813 188509
rect 116049 188273 116091 188509
rect 115771 188241 116091 188273
rect 131910 188829 132230 188861
rect 131910 188593 131952 188829
rect 132188 188593 132230 188829
rect 131910 188509 132230 188593
rect 131910 188273 131952 188509
rect 132188 188273 132230 188509
rect 131910 188241 132230 188273
rect 137840 188829 138160 188861
rect 137840 188593 137882 188829
rect 138118 188593 138160 188829
rect 137840 188509 138160 188593
rect 137840 188273 137882 188509
rect 138118 188273 138160 188509
rect 137840 188241 138160 188273
rect 143771 188829 144091 188861
rect 143771 188593 143813 188829
rect 144049 188593 144091 188829
rect 143771 188509 144091 188593
rect 143771 188273 143813 188509
rect 144049 188273 144091 188509
rect 143771 188241 144091 188273
rect 159910 188829 160230 188861
rect 159910 188593 159952 188829
rect 160188 188593 160230 188829
rect 159910 188509 160230 188593
rect 159910 188273 159952 188509
rect 160188 188273 160230 188509
rect 159910 188241 160230 188273
rect 165840 188829 166160 188861
rect 165840 188593 165882 188829
rect 166118 188593 166160 188829
rect 165840 188509 166160 188593
rect 165840 188273 165882 188509
rect 166118 188273 166160 188509
rect 165840 188241 166160 188273
rect 171771 188829 172091 188861
rect 171771 188593 171813 188829
rect 172049 188593 172091 188829
rect 171771 188509 172091 188593
rect 171771 188273 171813 188509
rect 172049 188273 172091 188509
rect 171771 188241 172091 188273
rect 187910 188829 188230 188861
rect 187910 188593 187952 188829
rect 188188 188593 188230 188829
rect 187910 188509 188230 188593
rect 187910 188273 187952 188509
rect 188188 188273 188230 188509
rect 187910 188241 188230 188273
rect 193840 188829 194160 188861
rect 193840 188593 193882 188829
rect 194118 188593 194160 188829
rect 193840 188509 194160 188593
rect 193840 188273 193882 188509
rect 194118 188273 194160 188509
rect 193840 188241 194160 188273
rect 199771 188829 200091 188861
rect 199771 188593 199813 188829
rect 200049 188593 200091 188829
rect 199771 188509 200091 188593
rect 199771 188273 199813 188509
rect 200049 188273 200091 188509
rect 199771 188241 200091 188273
rect 215910 188829 216230 188861
rect 215910 188593 215952 188829
rect 216188 188593 216230 188829
rect 215910 188509 216230 188593
rect 215910 188273 215952 188509
rect 216188 188273 216230 188509
rect 215910 188241 216230 188273
rect 221840 188829 222160 188861
rect 221840 188593 221882 188829
rect 222118 188593 222160 188829
rect 221840 188509 222160 188593
rect 221840 188273 221882 188509
rect 222118 188273 222160 188509
rect 221840 188241 222160 188273
rect 227771 188829 228091 188861
rect 227771 188593 227813 188829
rect 228049 188593 228091 188829
rect 227771 188509 228091 188593
rect 227771 188273 227813 188509
rect 228049 188273 228091 188509
rect 227771 188241 228091 188273
rect 243910 188829 244230 188861
rect 243910 188593 243952 188829
rect 244188 188593 244230 188829
rect 243910 188509 244230 188593
rect 243910 188273 243952 188509
rect 244188 188273 244230 188509
rect 243910 188241 244230 188273
rect 249840 188829 250160 188861
rect 249840 188593 249882 188829
rect 250118 188593 250160 188829
rect 249840 188509 250160 188593
rect 249840 188273 249882 188509
rect 250118 188273 250160 188509
rect 249840 188241 250160 188273
rect 255771 188829 256091 188861
rect 255771 188593 255813 188829
rect 256049 188593 256091 188829
rect 255771 188509 256091 188593
rect 255771 188273 255813 188509
rect 256049 188273 256091 188509
rect 255771 188241 256091 188273
rect 271910 188829 272230 188861
rect 271910 188593 271952 188829
rect 272188 188593 272230 188829
rect 271910 188509 272230 188593
rect 271910 188273 271952 188509
rect 272188 188273 272230 188509
rect 271910 188241 272230 188273
rect 277840 188829 278160 188861
rect 277840 188593 277882 188829
rect 278118 188593 278160 188829
rect 277840 188509 278160 188593
rect 277840 188273 277882 188509
rect 278118 188273 278160 188509
rect 277840 188241 278160 188273
rect 283771 188829 284091 188861
rect 283771 188593 283813 188829
rect 284049 188593 284091 188829
rect 283771 188509 284091 188593
rect 283771 188273 283813 188509
rect 284049 188273 284091 188509
rect 283771 188241 284091 188273
rect 299910 188829 300230 188861
rect 299910 188593 299952 188829
rect 300188 188593 300230 188829
rect 299910 188509 300230 188593
rect 299910 188273 299952 188509
rect 300188 188273 300230 188509
rect 299910 188241 300230 188273
rect 305840 188829 306160 188861
rect 305840 188593 305882 188829
rect 306118 188593 306160 188829
rect 305840 188509 306160 188593
rect 305840 188273 305882 188509
rect 306118 188273 306160 188509
rect 305840 188241 306160 188273
rect 311771 188829 312091 188861
rect 311771 188593 311813 188829
rect 312049 188593 312091 188829
rect 311771 188509 312091 188593
rect 311771 188273 311813 188509
rect 312049 188273 312091 188509
rect 311771 188241 312091 188273
rect 327910 188829 328230 188861
rect 327910 188593 327952 188829
rect 328188 188593 328230 188829
rect 327910 188509 328230 188593
rect 327910 188273 327952 188509
rect 328188 188273 328230 188509
rect 327910 188241 328230 188273
rect 333840 188829 334160 188861
rect 333840 188593 333882 188829
rect 334118 188593 334160 188829
rect 333840 188509 334160 188593
rect 333840 188273 333882 188509
rect 334118 188273 334160 188509
rect 333840 188241 334160 188273
rect 339771 188829 340091 188861
rect 339771 188593 339813 188829
rect 340049 188593 340091 188829
rect 339771 188509 340091 188593
rect 339771 188273 339813 188509
rect 340049 188273 340091 188509
rect 339771 188241 340091 188273
rect 355910 188829 356230 188861
rect 355910 188593 355952 188829
rect 356188 188593 356230 188829
rect 355910 188509 356230 188593
rect 355910 188273 355952 188509
rect 356188 188273 356230 188509
rect 355910 188241 356230 188273
rect 361840 188829 362160 188861
rect 361840 188593 361882 188829
rect 362118 188593 362160 188829
rect 361840 188509 362160 188593
rect 361840 188273 361882 188509
rect 362118 188273 362160 188509
rect 361840 188241 362160 188273
rect 367771 188829 368091 188861
rect 367771 188593 367813 188829
rect 368049 188593 368091 188829
rect 367771 188509 368091 188593
rect 367771 188273 367813 188509
rect 368049 188273 368091 188509
rect 367771 188241 368091 188273
rect 383910 188829 384230 188861
rect 383910 188593 383952 188829
rect 384188 188593 384230 188829
rect 383910 188509 384230 188593
rect 383910 188273 383952 188509
rect 384188 188273 384230 188509
rect 383910 188241 384230 188273
rect 389840 188829 390160 188861
rect 389840 188593 389882 188829
rect 390118 188593 390160 188829
rect 389840 188509 390160 188593
rect 389840 188273 389882 188509
rect 390118 188273 390160 188509
rect 389840 188241 390160 188273
rect 395771 188829 396091 188861
rect 395771 188593 395813 188829
rect 396049 188593 396091 188829
rect 395771 188509 396091 188593
rect 395771 188273 395813 188509
rect 396049 188273 396091 188509
rect 395771 188241 396091 188273
rect 411910 188829 412230 188861
rect 411910 188593 411952 188829
rect 412188 188593 412230 188829
rect 411910 188509 412230 188593
rect 411910 188273 411952 188509
rect 412188 188273 412230 188509
rect 411910 188241 412230 188273
rect 417840 188829 418160 188861
rect 417840 188593 417882 188829
rect 418118 188593 418160 188829
rect 417840 188509 418160 188593
rect 417840 188273 417882 188509
rect 418118 188273 418160 188509
rect 417840 188241 418160 188273
rect 423771 188829 424091 188861
rect 423771 188593 423813 188829
rect 424049 188593 424091 188829
rect 423771 188509 424091 188593
rect 423771 188273 423813 188509
rect 424049 188273 424091 188509
rect 423771 188241 424091 188273
rect 439910 188829 440230 188861
rect 439910 188593 439952 188829
rect 440188 188593 440230 188829
rect 439910 188509 440230 188593
rect 439910 188273 439952 188509
rect 440188 188273 440230 188509
rect 439910 188241 440230 188273
rect 445840 188829 446160 188861
rect 445840 188593 445882 188829
rect 446118 188593 446160 188829
rect 445840 188509 446160 188593
rect 445840 188273 445882 188509
rect 446118 188273 446160 188509
rect 445840 188241 446160 188273
rect 451771 188829 452091 188861
rect 451771 188593 451813 188829
rect 452049 188593 452091 188829
rect 451771 188509 452091 188593
rect 451771 188273 451813 188509
rect 452049 188273 452091 188509
rect 451771 188241 452091 188273
rect 467910 188829 468230 188861
rect 467910 188593 467952 188829
rect 468188 188593 468230 188829
rect 467910 188509 468230 188593
rect 467910 188273 467952 188509
rect 468188 188273 468230 188509
rect 467910 188241 468230 188273
rect 473840 188829 474160 188861
rect 473840 188593 473882 188829
rect 474118 188593 474160 188829
rect 473840 188509 474160 188593
rect 473840 188273 473882 188509
rect 474118 188273 474160 188509
rect 473840 188241 474160 188273
rect 479771 188829 480091 188861
rect 479771 188593 479813 188829
rect 480049 188593 480091 188829
rect 479771 188509 480091 188593
rect 479771 188273 479813 188509
rect 480049 188273 480091 188509
rect 479771 188241 480091 188273
rect 495910 188829 496230 188861
rect 495910 188593 495952 188829
rect 496188 188593 496230 188829
rect 495910 188509 496230 188593
rect 495910 188273 495952 188509
rect 496188 188273 496230 188509
rect 495910 188241 496230 188273
rect 501840 188829 502160 188861
rect 501840 188593 501882 188829
rect 502118 188593 502160 188829
rect 501840 188509 502160 188593
rect 501840 188273 501882 188509
rect 502118 188273 502160 188509
rect 501840 188241 502160 188273
rect 507771 188829 508091 188861
rect 507771 188593 507813 188829
rect 508049 188593 508091 188829
rect 507771 188509 508091 188593
rect 507771 188273 507813 188509
rect 508049 188273 508091 188509
rect 507771 188241 508091 188273
rect 523910 188829 524230 188861
rect 523910 188593 523952 188829
rect 524188 188593 524230 188829
rect 523910 188509 524230 188593
rect 523910 188273 523952 188509
rect 524188 188273 524230 188509
rect 523910 188241 524230 188273
rect 529840 188829 530160 188861
rect 529840 188593 529882 188829
rect 530118 188593 530160 188829
rect 529840 188509 530160 188593
rect 529840 188273 529882 188509
rect 530118 188273 530160 188509
rect 529840 188241 530160 188273
rect 535771 188829 536091 188861
rect 535771 188593 535813 188829
rect 536049 188593 536091 188829
rect 535771 188509 536091 188593
rect 535771 188273 535813 188509
rect 536049 188273 536091 188509
rect 535771 188241 536091 188273
rect 551910 188829 552230 188861
rect 551910 188593 551952 188829
rect 552188 188593 552230 188829
rect 551910 188509 552230 188593
rect 551910 188273 551952 188509
rect 552188 188273 552230 188509
rect 551910 188241 552230 188273
rect 557840 188829 558160 188861
rect 557840 188593 557882 188829
rect 558118 188593 558160 188829
rect 557840 188509 558160 188593
rect 557840 188273 557882 188509
rect 558118 188273 558160 188509
rect 557840 188241 558160 188273
rect 563771 188829 564091 188861
rect 563771 188593 563813 188829
rect 564049 188593 564091 188829
rect 563771 188509 564091 188593
rect 563771 188273 563813 188509
rect 564049 188273 564091 188509
rect 563771 188241 564091 188273
rect 573494 188829 574114 215273
rect 573494 188593 573526 188829
rect 573762 188593 573846 188829
rect 574082 188593 574114 188829
rect 573494 188509 574114 188593
rect 573494 188273 573526 188509
rect 573762 188273 573846 188509
rect 574082 188273 574114 188509
rect 22874 185454 23194 185486
rect 22874 185218 22916 185454
rect 23152 185218 23194 185454
rect 22874 185134 23194 185218
rect 22874 184898 22916 185134
rect 23152 184898 23194 185134
rect 22874 184866 23194 184898
rect 28805 185454 29125 185486
rect 28805 185218 28847 185454
rect 29083 185218 29125 185454
rect 28805 185134 29125 185218
rect 28805 184898 28847 185134
rect 29083 184898 29125 185134
rect 28805 184866 29125 184898
rect 50874 185454 51194 185486
rect 50874 185218 50916 185454
rect 51152 185218 51194 185454
rect 50874 185134 51194 185218
rect 50874 184898 50916 185134
rect 51152 184898 51194 185134
rect 50874 184866 51194 184898
rect 56805 185454 57125 185486
rect 56805 185218 56847 185454
rect 57083 185218 57125 185454
rect 56805 185134 57125 185218
rect 56805 184898 56847 185134
rect 57083 184898 57125 185134
rect 56805 184866 57125 184898
rect 78874 185454 79194 185486
rect 78874 185218 78916 185454
rect 79152 185218 79194 185454
rect 78874 185134 79194 185218
rect 78874 184898 78916 185134
rect 79152 184898 79194 185134
rect 78874 184866 79194 184898
rect 84805 185454 85125 185486
rect 84805 185218 84847 185454
rect 85083 185218 85125 185454
rect 84805 185134 85125 185218
rect 84805 184898 84847 185134
rect 85083 184898 85125 185134
rect 84805 184866 85125 184898
rect 106874 185454 107194 185486
rect 106874 185218 106916 185454
rect 107152 185218 107194 185454
rect 106874 185134 107194 185218
rect 106874 184898 106916 185134
rect 107152 184898 107194 185134
rect 106874 184866 107194 184898
rect 112805 185454 113125 185486
rect 112805 185218 112847 185454
rect 113083 185218 113125 185454
rect 112805 185134 113125 185218
rect 112805 184898 112847 185134
rect 113083 184898 113125 185134
rect 112805 184866 113125 184898
rect 134874 185454 135194 185486
rect 134874 185218 134916 185454
rect 135152 185218 135194 185454
rect 134874 185134 135194 185218
rect 134874 184898 134916 185134
rect 135152 184898 135194 185134
rect 134874 184866 135194 184898
rect 140805 185454 141125 185486
rect 140805 185218 140847 185454
rect 141083 185218 141125 185454
rect 140805 185134 141125 185218
rect 140805 184898 140847 185134
rect 141083 184898 141125 185134
rect 140805 184866 141125 184898
rect 162874 185454 163194 185486
rect 162874 185218 162916 185454
rect 163152 185218 163194 185454
rect 162874 185134 163194 185218
rect 162874 184898 162916 185134
rect 163152 184898 163194 185134
rect 162874 184866 163194 184898
rect 168805 185454 169125 185486
rect 168805 185218 168847 185454
rect 169083 185218 169125 185454
rect 168805 185134 169125 185218
rect 168805 184898 168847 185134
rect 169083 184898 169125 185134
rect 168805 184866 169125 184898
rect 190874 185454 191194 185486
rect 190874 185218 190916 185454
rect 191152 185218 191194 185454
rect 190874 185134 191194 185218
rect 190874 184898 190916 185134
rect 191152 184898 191194 185134
rect 190874 184866 191194 184898
rect 196805 185454 197125 185486
rect 196805 185218 196847 185454
rect 197083 185218 197125 185454
rect 196805 185134 197125 185218
rect 196805 184898 196847 185134
rect 197083 184898 197125 185134
rect 196805 184866 197125 184898
rect 218874 185454 219194 185486
rect 218874 185218 218916 185454
rect 219152 185218 219194 185454
rect 218874 185134 219194 185218
rect 218874 184898 218916 185134
rect 219152 184898 219194 185134
rect 218874 184866 219194 184898
rect 224805 185454 225125 185486
rect 224805 185218 224847 185454
rect 225083 185218 225125 185454
rect 224805 185134 225125 185218
rect 224805 184898 224847 185134
rect 225083 184898 225125 185134
rect 224805 184866 225125 184898
rect 246874 185454 247194 185486
rect 246874 185218 246916 185454
rect 247152 185218 247194 185454
rect 246874 185134 247194 185218
rect 246874 184898 246916 185134
rect 247152 184898 247194 185134
rect 246874 184866 247194 184898
rect 252805 185454 253125 185486
rect 252805 185218 252847 185454
rect 253083 185218 253125 185454
rect 252805 185134 253125 185218
rect 252805 184898 252847 185134
rect 253083 184898 253125 185134
rect 252805 184866 253125 184898
rect 274874 185454 275194 185486
rect 274874 185218 274916 185454
rect 275152 185218 275194 185454
rect 274874 185134 275194 185218
rect 274874 184898 274916 185134
rect 275152 184898 275194 185134
rect 274874 184866 275194 184898
rect 280805 185454 281125 185486
rect 280805 185218 280847 185454
rect 281083 185218 281125 185454
rect 280805 185134 281125 185218
rect 280805 184898 280847 185134
rect 281083 184898 281125 185134
rect 280805 184866 281125 184898
rect 302874 185454 303194 185486
rect 302874 185218 302916 185454
rect 303152 185218 303194 185454
rect 302874 185134 303194 185218
rect 302874 184898 302916 185134
rect 303152 184898 303194 185134
rect 302874 184866 303194 184898
rect 308805 185454 309125 185486
rect 308805 185218 308847 185454
rect 309083 185218 309125 185454
rect 308805 185134 309125 185218
rect 308805 184898 308847 185134
rect 309083 184898 309125 185134
rect 308805 184866 309125 184898
rect 330874 185454 331194 185486
rect 330874 185218 330916 185454
rect 331152 185218 331194 185454
rect 330874 185134 331194 185218
rect 330874 184898 330916 185134
rect 331152 184898 331194 185134
rect 330874 184866 331194 184898
rect 336805 185454 337125 185486
rect 336805 185218 336847 185454
rect 337083 185218 337125 185454
rect 336805 185134 337125 185218
rect 336805 184898 336847 185134
rect 337083 184898 337125 185134
rect 336805 184866 337125 184898
rect 358874 185454 359194 185486
rect 358874 185218 358916 185454
rect 359152 185218 359194 185454
rect 358874 185134 359194 185218
rect 358874 184898 358916 185134
rect 359152 184898 359194 185134
rect 358874 184866 359194 184898
rect 364805 185454 365125 185486
rect 364805 185218 364847 185454
rect 365083 185218 365125 185454
rect 364805 185134 365125 185218
rect 364805 184898 364847 185134
rect 365083 184898 365125 185134
rect 364805 184866 365125 184898
rect 386874 185454 387194 185486
rect 386874 185218 386916 185454
rect 387152 185218 387194 185454
rect 386874 185134 387194 185218
rect 386874 184898 386916 185134
rect 387152 184898 387194 185134
rect 386874 184866 387194 184898
rect 392805 185454 393125 185486
rect 392805 185218 392847 185454
rect 393083 185218 393125 185454
rect 392805 185134 393125 185218
rect 392805 184898 392847 185134
rect 393083 184898 393125 185134
rect 392805 184866 393125 184898
rect 414874 185454 415194 185486
rect 414874 185218 414916 185454
rect 415152 185218 415194 185454
rect 414874 185134 415194 185218
rect 414874 184898 414916 185134
rect 415152 184898 415194 185134
rect 414874 184866 415194 184898
rect 420805 185454 421125 185486
rect 420805 185218 420847 185454
rect 421083 185218 421125 185454
rect 420805 185134 421125 185218
rect 420805 184898 420847 185134
rect 421083 184898 421125 185134
rect 420805 184866 421125 184898
rect 442874 185454 443194 185486
rect 442874 185218 442916 185454
rect 443152 185218 443194 185454
rect 442874 185134 443194 185218
rect 442874 184898 442916 185134
rect 443152 184898 443194 185134
rect 442874 184866 443194 184898
rect 448805 185454 449125 185486
rect 448805 185218 448847 185454
rect 449083 185218 449125 185454
rect 448805 185134 449125 185218
rect 448805 184898 448847 185134
rect 449083 184898 449125 185134
rect 448805 184866 449125 184898
rect 470874 185454 471194 185486
rect 470874 185218 470916 185454
rect 471152 185218 471194 185454
rect 470874 185134 471194 185218
rect 470874 184898 470916 185134
rect 471152 184898 471194 185134
rect 470874 184866 471194 184898
rect 476805 185454 477125 185486
rect 476805 185218 476847 185454
rect 477083 185218 477125 185454
rect 476805 185134 477125 185218
rect 476805 184898 476847 185134
rect 477083 184898 477125 185134
rect 476805 184866 477125 184898
rect 498874 185454 499194 185486
rect 498874 185218 498916 185454
rect 499152 185218 499194 185454
rect 498874 185134 499194 185218
rect 498874 184898 498916 185134
rect 499152 184898 499194 185134
rect 498874 184866 499194 184898
rect 504805 185454 505125 185486
rect 504805 185218 504847 185454
rect 505083 185218 505125 185454
rect 504805 185134 505125 185218
rect 504805 184898 504847 185134
rect 505083 184898 505125 185134
rect 504805 184866 505125 184898
rect 526874 185454 527194 185486
rect 526874 185218 526916 185454
rect 527152 185218 527194 185454
rect 526874 185134 527194 185218
rect 526874 184898 526916 185134
rect 527152 184898 527194 185134
rect 526874 184866 527194 184898
rect 532805 185454 533125 185486
rect 532805 185218 532847 185454
rect 533083 185218 533125 185454
rect 532805 185134 533125 185218
rect 532805 184898 532847 185134
rect 533083 184898 533125 185134
rect 532805 184866 533125 184898
rect 554874 185454 555194 185486
rect 554874 185218 554916 185454
rect 555152 185218 555194 185454
rect 554874 185134 555194 185218
rect 554874 184898 554916 185134
rect 555152 184898 555194 185134
rect 554874 184866 555194 184898
rect 560805 185454 561125 185486
rect 560805 185218 560847 185454
rect 561083 185218 561125 185454
rect 560805 185134 561125 185218
rect 560805 184898 560847 185134
rect 561083 184898 561125 185134
rect 560805 184866 561125 184898
rect -2006 161593 -1974 161829
rect -1738 161593 -1654 161829
rect -1418 161593 -1386 161829
rect -2006 161509 -1386 161593
rect -2006 161273 -1974 161509
rect -1738 161273 -1654 161509
rect -1418 161273 -1386 161509
rect -2006 134829 -1386 161273
rect 19909 161829 20229 161861
rect 19909 161593 19951 161829
rect 20187 161593 20229 161829
rect 19909 161509 20229 161593
rect 19909 161273 19951 161509
rect 20187 161273 20229 161509
rect 19909 161241 20229 161273
rect 25840 161829 26160 161861
rect 25840 161593 25882 161829
rect 26118 161593 26160 161829
rect 25840 161509 26160 161593
rect 25840 161273 25882 161509
rect 26118 161273 26160 161509
rect 25840 161241 26160 161273
rect 31770 161829 32090 161861
rect 31770 161593 31812 161829
rect 32048 161593 32090 161829
rect 31770 161509 32090 161593
rect 31770 161273 31812 161509
rect 32048 161273 32090 161509
rect 31770 161241 32090 161273
rect 47909 161829 48229 161861
rect 47909 161593 47951 161829
rect 48187 161593 48229 161829
rect 47909 161509 48229 161593
rect 47909 161273 47951 161509
rect 48187 161273 48229 161509
rect 47909 161241 48229 161273
rect 53840 161829 54160 161861
rect 53840 161593 53882 161829
rect 54118 161593 54160 161829
rect 53840 161509 54160 161593
rect 53840 161273 53882 161509
rect 54118 161273 54160 161509
rect 53840 161241 54160 161273
rect 59770 161829 60090 161861
rect 59770 161593 59812 161829
rect 60048 161593 60090 161829
rect 59770 161509 60090 161593
rect 59770 161273 59812 161509
rect 60048 161273 60090 161509
rect 59770 161241 60090 161273
rect 75909 161829 76229 161861
rect 75909 161593 75951 161829
rect 76187 161593 76229 161829
rect 75909 161509 76229 161593
rect 75909 161273 75951 161509
rect 76187 161273 76229 161509
rect 75909 161241 76229 161273
rect 81840 161829 82160 161861
rect 81840 161593 81882 161829
rect 82118 161593 82160 161829
rect 81840 161509 82160 161593
rect 81840 161273 81882 161509
rect 82118 161273 82160 161509
rect 81840 161241 82160 161273
rect 87770 161829 88090 161861
rect 87770 161593 87812 161829
rect 88048 161593 88090 161829
rect 87770 161509 88090 161593
rect 87770 161273 87812 161509
rect 88048 161273 88090 161509
rect 87770 161241 88090 161273
rect 103909 161829 104229 161861
rect 103909 161593 103951 161829
rect 104187 161593 104229 161829
rect 103909 161509 104229 161593
rect 103909 161273 103951 161509
rect 104187 161273 104229 161509
rect 103909 161241 104229 161273
rect 109840 161829 110160 161861
rect 109840 161593 109882 161829
rect 110118 161593 110160 161829
rect 109840 161509 110160 161593
rect 109840 161273 109882 161509
rect 110118 161273 110160 161509
rect 109840 161241 110160 161273
rect 115770 161829 116090 161861
rect 115770 161593 115812 161829
rect 116048 161593 116090 161829
rect 115770 161509 116090 161593
rect 115770 161273 115812 161509
rect 116048 161273 116090 161509
rect 115770 161241 116090 161273
rect 131909 161829 132229 161861
rect 131909 161593 131951 161829
rect 132187 161593 132229 161829
rect 131909 161509 132229 161593
rect 131909 161273 131951 161509
rect 132187 161273 132229 161509
rect 131909 161241 132229 161273
rect 137840 161829 138160 161861
rect 137840 161593 137882 161829
rect 138118 161593 138160 161829
rect 137840 161509 138160 161593
rect 137840 161273 137882 161509
rect 138118 161273 138160 161509
rect 137840 161241 138160 161273
rect 143770 161829 144090 161861
rect 143770 161593 143812 161829
rect 144048 161593 144090 161829
rect 143770 161509 144090 161593
rect 143770 161273 143812 161509
rect 144048 161273 144090 161509
rect 143770 161241 144090 161273
rect 159909 161829 160229 161861
rect 159909 161593 159951 161829
rect 160187 161593 160229 161829
rect 159909 161509 160229 161593
rect 159909 161273 159951 161509
rect 160187 161273 160229 161509
rect 159909 161241 160229 161273
rect 165840 161829 166160 161861
rect 165840 161593 165882 161829
rect 166118 161593 166160 161829
rect 165840 161509 166160 161593
rect 165840 161273 165882 161509
rect 166118 161273 166160 161509
rect 165840 161241 166160 161273
rect 171770 161829 172090 161861
rect 171770 161593 171812 161829
rect 172048 161593 172090 161829
rect 171770 161509 172090 161593
rect 171770 161273 171812 161509
rect 172048 161273 172090 161509
rect 171770 161241 172090 161273
rect 187909 161829 188229 161861
rect 187909 161593 187951 161829
rect 188187 161593 188229 161829
rect 187909 161509 188229 161593
rect 187909 161273 187951 161509
rect 188187 161273 188229 161509
rect 187909 161241 188229 161273
rect 193840 161829 194160 161861
rect 193840 161593 193882 161829
rect 194118 161593 194160 161829
rect 193840 161509 194160 161593
rect 193840 161273 193882 161509
rect 194118 161273 194160 161509
rect 193840 161241 194160 161273
rect 199770 161829 200090 161861
rect 199770 161593 199812 161829
rect 200048 161593 200090 161829
rect 199770 161509 200090 161593
rect 199770 161273 199812 161509
rect 200048 161273 200090 161509
rect 199770 161241 200090 161273
rect 215909 161829 216229 161861
rect 215909 161593 215951 161829
rect 216187 161593 216229 161829
rect 215909 161509 216229 161593
rect 215909 161273 215951 161509
rect 216187 161273 216229 161509
rect 215909 161241 216229 161273
rect 221840 161829 222160 161861
rect 221840 161593 221882 161829
rect 222118 161593 222160 161829
rect 221840 161509 222160 161593
rect 221840 161273 221882 161509
rect 222118 161273 222160 161509
rect 221840 161241 222160 161273
rect 227770 161829 228090 161861
rect 227770 161593 227812 161829
rect 228048 161593 228090 161829
rect 227770 161509 228090 161593
rect 227770 161273 227812 161509
rect 228048 161273 228090 161509
rect 227770 161241 228090 161273
rect 243909 161829 244229 161861
rect 243909 161593 243951 161829
rect 244187 161593 244229 161829
rect 243909 161509 244229 161593
rect 243909 161273 243951 161509
rect 244187 161273 244229 161509
rect 243909 161241 244229 161273
rect 249840 161829 250160 161861
rect 249840 161593 249882 161829
rect 250118 161593 250160 161829
rect 249840 161509 250160 161593
rect 249840 161273 249882 161509
rect 250118 161273 250160 161509
rect 249840 161241 250160 161273
rect 255770 161829 256090 161861
rect 255770 161593 255812 161829
rect 256048 161593 256090 161829
rect 255770 161509 256090 161593
rect 255770 161273 255812 161509
rect 256048 161273 256090 161509
rect 255770 161241 256090 161273
rect 271909 161829 272229 161861
rect 271909 161593 271951 161829
rect 272187 161593 272229 161829
rect 271909 161509 272229 161593
rect 271909 161273 271951 161509
rect 272187 161273 272229 161509
rect 271909 161241 272229 161273
rect 277840 161829 278160 161861
rect 277840 161593 277882 161829
rect 278118 161593 278160 161829
rect 277840 161509 278160 161593
rect 277840 161273 277882 161509
rect 278118 161273 278160 161509
rect 277840 161241 278160 161273
rect 283770 161829 284090 161861
rect 283770 161593 283812 161829
rect 284048 161593 284090 161829
rect 283770 161509 284090 161593
rect 283770 161273 283812 161509
rect 284048 161273 284090 161509
rect 283770 161241 284090 161273
rect 299909 161829 300229 161861
rect 299909 161593 299951 161829
rect 300187 161593 300229 161829
rect 299909 161509 300229 161593
rect 299909 161273 299951 161509
rect 300187 161273 300229 161509
rect 299909 161241 300229 161273
rect 305840 161829 306160 161861
rect 305840 161593 305882 161829
rect 306118 161593 306160 161829
rect 305840 161509 306160 161593
rect 305840 161273 305882 161509
rect 306118 161273 306160 161509
rect 305840 161241 306160 161273
rect 311770 161829 312090 161861
rect 311770 161593 311812 161829
rect 312048 161593 312090 161829
rect 311770 161509 312090 161593
rect 311770 161273 311812 161509
rect 312048 161273 312090 161509
rect 311770 161241 312090 161273
rect 327909 161829 328229 161861
rect 327909 161593 327951 161829
rect 328187 161593 328229 161829
rect 327909 161509 328229 161593
rect 327909 161273 327951 161509
rect 328187 161273 328229 161509
rect 327909 161241 328229 161273
rect 333840 161829 334160 161861
rect 333840 161593 333882 161829
rect 334118 161593 334160 161829
rect 333840 161509 334160 161593
rect 333840 161273 333882 161509
rect 334118 161273 334160 161509
rect 333840 161241 334160 161273
rect 339770 161829 340090 161861
rect 339770 161593 339812 161829
rect 340048 161593 340090 161829
rect 339770 161509 340090 161593
rect 339770 161273 339812 161509
rect 340048 161273 340090 161509
rect 339770 161241 340090 161273
rect 355909 161829 356229 161861
rect 355909 161593 355951 161829
rect 356187 161593 356229 161829
rect 355909 161509 356229 161593
rect 355909 161273 355951 161509
rect 356187 161273 356229 161509
rect 355909 161241 356229 161273
rect 361840 161829 362160 161861
rect 361840 161593 361882 161829
rect 362118 161593 362160 161829
rect 361840 161509 362160 161593
rect 361840 161273 361882 161509
rect 362118 161273 362160 161509
rect 361840 161241 362160 161273
rect 367770 161829 368090 161861
rect 367770 161593 367812 161829
rect 368048 161593 368090 161829
rect 367770 161509 368090 161593
rect 367770 161273 367812 161509
rect 368048 161273 368090 161509
rect 367770 161241 368090 161273
rect 383909 161829 384229 161861
rect 383909 161593 383951 161829
rect 384187 161593 384229 161829
rect 383909 161509 384229 161593
rect 383909 161273 383951 161509
rect 384187 161273 384229 161509
rect 383909 161241 384229 161273
rect 389840 161829 390160 161861
rect 389840 161593 389882 161829
rect 390118 161593 390160 161829
rect 389840 161509 390160 161593
rect 389840 161273 389882 161509
rect 390118 161273 390160 161509
rect 389840 161241 390160 161273
rect 395770 161829 396090 161861
rect 395770 161593 395812 161829
rect 396048 161593 396090 161829
rect 395770 161509 396090 161593
rect 395770 161273 395812 161509
rect 396048 161273 396090 161509
rect 395770 161241 396090 161273
rect 411909 161829 412229 161861
rect 411909 161593 411951 161829
rect 412187 161593 412229 161829
rect 411909 161509 412229 161593
rect 411909 161273 411951 161509
rect 412187 161273 412229 161509
rect 411909 161241 412229 161273
rect 417840 161829 418160 161861
rect 417840 161593 417882 161829
rect 418118 161593 418160 161829
rect 417840 161509 418160 161593
rect 417840 161273 417882 161509
rect 418118 161273 418160 161509
rect 417840 161241 418160 161273
rect 423770 161829 424090 161861
rect 423770 161593 423812 161829
rect 424048 161593 424090 161829
rect 423770 161509 424090 161593
rect 423770 161273 423812 161509
rect 424048 161273 424090 161509
rect 423770 161241 424090 161273
rect 439909 161829 440229 161861
rect 439909 161593 439951 161829
rect 440187 161593 440229 161829
rect 439909 161509 440229 161593
rect 439909 161273 439951 161509
rect 440187 161273 440229 161509
rect 439909 161241 440229 161273
rect 445840 161829 446160 161861
rect 445840 161593 445882 161829
rect 446118 161593 446160 161829
rect 445840 161509 446160 161593
rect 445840 161273 445882 161509
rect 446118 161273 446160 161509
rect 445840 161241 446160 161273
rect 451770 161829 452090 161861
rect 451770 161593 451812 161829
rect 452048 161593 452090 161829
rect 451770 161509 452090 161593
rect 451770 161273 451812 161509
rect 452048 161273 452090 161509
rect 451770 161241 452090 161273
rect 467909 161829 468229 161861
rect 467909 161593 467951 161829
rect 468187 161593 468229 161829
rect 467909 161509 468229 161593
rect 467909 161273 467951 161509
rect 468187 161273 468229 161509
rect 467909 161241 468229 161273
rect 473840 161829 474160 161861
rect 473840 161593 473882 161829
rect 474118 161593 474160 161829
rect 473840 161509 474160 161593
rect 473840 161273 473882 161509
rect 474118 161273 474160 161509
rect 473840 161241 474160 161273
rect 479770 161829 480090 161861
rect 479770 161593 479812 161829
rect 480048 161593 480090 161829
rect 479770 161509 480090 161593
rect 479770 161273 479812 161509
rect 480048 161273 480090 161509
rect 479770 161241 480090 161273
rect 495909 161829 496229 161861
rect 495909 161593 495951 161829
rect 496187 161593 496229 161829
rect 495909 161509 496229 161593
rect 495909 161273 495951 161509
rect 496187 161273 496229 161509
rect 495909 161241 496229 161273
rect 501840 161829 502160 161861
rect 501840 161593 501882 161829
rect 502118 161593 502160 161829
rect 501840 161509 502160 161593
rect 501840 161273 501882 161509
rect 502118 161273 502160 161509
rect 501840 161241 502160 161273
rect 507770 161829 508090 161861
rect 507770 161593 507812 161829
rect 508048 161593 508090 161829
rect 507770 161509 508090 161593
rect 507770 161273 507812 161509
rect 508048 161273 508090 161509
rect 507770 161241 508090 161273
rect 523909 161829 524229 161861
rect 523909 161593 523951 161829
rect 524187 161593 524229 161829
rect 523909 161509 524229 161593
rect 523909 161273 523951 161509
rect 524187 161273 524229 161509
rect 523909 161241 524229 161273
rect 529840 161829 530160 161861
rect 529840 161593 529882 161829
rect 530118 161593 530160 161829
rect 529840 161509 530160 161593
rect 529840 161273 529882 161509
rect 530118 161273 530160 161509
rect 529840 161241 530160 161273
rect 535770 161829 536090 161861
rect 535770 161593 535812 161829
rect 536048 161593 536090 161829
rect 535770 161509 536090 161593
rect 535770 161273 535812 161509
rect 536048 161273 536090 161509
rect 535770 161241 536090 161273
rect 551909 161829 552229 161861
rect 551909 161593 551951 161829
rect 552187 161593 552229 161829
rect 551909 161509 552229 161593
rect 551909 161273 551951 161509
rect 552187 161273 552229 161509
rect 551909 161241 552229 161273
rect 557840 161829 558160 161861
rect 557840 161593 557882 161829
rect 558118 161593 558160 161829
rect 557840 161509 558160 161593
rect 557840 161273 557882 161509
rect 558118 161273 558160 161509
rect 557840 161241 558160 161273
rect 563770 161829 564090 161861
rect 563770 161593 563812 161829
rect 564048 161593 564090 161829
rect 563770 161509 564090 161593
rect 563770 161273 563812 161509
rect 564048 161273 564090 161509
rect 563770 161241 564090 161273
rect 573494 161829 574114 188273
rect 573494 161593 573526 161829
rect 573762 161593 573846 161829
rect 574082 161593 574114 161829
rect 573494 161509 574114 161593
rect 573494 161273 573526 161509
rect 573762 161273 573846 161509
rect 574082 161273 574114 161509
rect 22875 158454 23195 158486
rect 22875 158218 22917 158454
rect 23153 158218 23195 158454
rect 22875 158134 23195 158218
rect 22875 157898 22917 158134
rect 23153 157898 23195 158134
rect 22875 157866 23195 157898
rect 28806 158454 29126 158486
rect 28806 158218 28848 158454
rect 29084 158218 29126 158454
rect 28806 158134 29126 158218
rect 28806 157898 28848 158134
rect 29084 157898 29126 158134
rect 28806 157866 29126 157898
rect 50875 158454 51195 158486
rect 50875 158218 50917 158454
rect 51153 158218 51195 158454
rect 50875 158134 51195 158218
rect 50875 157898 50917 158134
rect 51153 157898 51195 158134
rect 50875 157866 51195 157898
rect 56806 158454 57126 158486
rect 56806 158218 56848 158454
rect 57084 158218 57126 158454
rect 56806 158134 57126 158218
rect 56806 157898 56848 158134
rect 57084 157898 57126 158134
rect 56806 157866 57126 157898
rect 78875 158454 79195 158486
rect 78875 158218 78917 158454
rect 79153 158218 79195 158454
rect 78875 158134 79195 158218
rect 78875 157898 78917 158134
rect 79153 157898 79195 158134
rect 78875 157866 79195 157898
rect 84806 158454 85126 158486
rect 84806 158218 84848 158454
rect 85084 158218 85126 158454
rect 84806 158134 85126 158218
rect 84806 157898 84848 158134
rect 85084 157898 85126 158134
rect 84806 157866 85126 157898
rect 106875 158454 107195 158486
rect 106875 158218 106917 158454
rect 107153 158218 107195 158454
rect 106875 158134 107195 158218
rect 106875 157898 106917 158134
rect 107153 157898 107195 158134
rect 106875 157866 107195 157898
rect 112806 158454 113126 158486
rect 112806 158218 112848 158454
rect 113084 158218 113126 158454
rect 112806 158134 113126 158218
rect 112806 157898 112848 158134
rect 113084 157898 113126 158134
rect 112806 157866 113126 157898
rect 134875 158454 135195 158486
rect 134875 158218 134917 158454
rect 135153 158218 135195 158454
rect 134875 158134 135195 158218
rect 134875 157898 134917 158134
rect 135153 157898 135195 158134
rect 134875 157866 135195 157898
rect 140806 158454 141126 158486
rect 140806 158218 140848 158454
rect 141084 158218 141126 158454
rect 140806 158134 141126 158218
rect 140806 157898 140848 158134
rect 141084 157898 141126 158134
rect 140806 157866 141126 157898
rect 162875 158454 163195 158486
rect 162875 158218 162917 158454
rect 163153 158218 163195 158454
rect 162875 158134 163195 158218
rect 162875 157898 162917 158134
rect 163153 157898 163195 158134
rect 162875 157866 163195 157898
rect 168806 158454 169126 158486
rect 168806 158218 168848 158454
rect 169084 158218 169126 158454
rect 168806 158134 169126 158218
rect 168806 157898 168848 158134
rect 169084 157898 169126 158134
rect 168806 157866 169126 157898
rect 190875 158454 191195 158486
rect 190875 158218 190917 158454
rect 191153 158218 191195 158454
rect 190875 158134 191195 158218
rect 190875 157898 190917 158134
rect 191153 157898 191195 158134
rect 190875 157866 191195 157898
rect 196806 158454 197126 158486
rect 196806 158218 196848 158454
rect 197084 158218 197126 158454
rect 196806 158134 197126 158218
rect 196806 157898 196848 158134
rect 197084 157898 197126 158134
rect 196806 157866 197126 157898
rect 218875 158454 219195 158486
rect 218875 158218 218917 158454
rect 219153 158218 219195 158454
rect 218875 158134 219195 158218
rect 218875 157898 218917 158134
rect 219153 157898 219195 158134
rect 218875 157866 219195 157898
rect 224806 158454 225126 158486
rect 224806 158218 224848 158454
rect 225084 158218 225126 158454
rect 224806 158134 225126 158218
rect 224806 157898 224848 158134
rect 225084 157898 225126 158134
rect 224806 157866 225126 157898
rect 246875 158454 247195 158486
rect 246875 158218 246917 158454
rect 247153 158218 247195 158454
rect 246875 158134 247195 158218
rect 246875 157898 246917 158134
rect 247153 157898 247195 158134
rect 246875 157866 247195 157898
rect 252806 158454 253126 158486
rect 252806 158218 252848 158454
rect 253084 158218 253126 158454
rect 252806 158134 253126 158218
rect 252806 157898 252848 158134
rect 253084 157898 253126 158134
rect 252806 157866 253126 157898
rect 274875 158454 275195 158486
rect 274875 158218 274917 158454
rect 275153 158218 275195 158454
rect 274875 158134 275195 158218
rect 274875 157898 274917 158134
rect 275153 157898 275195 158134
rect 274875 157866 275195 157898
rect 280806 158454 281126 158486
rect 280806 158218 280848 158454
rect 281084 158218 281126 158454
rect 280806 158134 281126 158218
rect 280806 157898 280848 158134
rect 281084 157898 281126 158134
rect 280806 157866 281126 157898
rect 302875 158454 303195 158486
rect 302875 158218 302917 158454
rect 303153 158218 303195 158454
rect 302875 158134 303195 158218
rect 302875 157898 302917 158134
rect 303153 157898 303195 158134
rect 302875 157866 303195 157898
rect 308806 158454 309126 158486
rect 308806 158218 308848 158454
rect 309084 158218 309126 158454
rect 308806 158134 309126 158218
rect 308806 157898 308848 158134
rect 309084 157898 309126 158134
rect 308806 157866 309126 157898
rect 330875 158454 331195 158486
rect 330875 158218 330917 158454
rect 331153 158218 331195 158454
rect 330875 158134 331195 158218
rect 330875 157898 330917 158134
rect 331153 157898 331195 158134
rect 330875 157866 331195 157898
rect 336806 158454 337126 158486
rect 336806 158218 336848 158454
rect 337084 158218 337126 158454
rect 336806 158134 337126 158218
rect 336806 157898 336848 158134
rect 337084 157898 337126 158134
rect 336806 157866 337126 157898
rect 358875 158454 359195 158486
rect 358875 158218 358917 158454
rect 359153 158218 359195 158454
rect 358875 158134 359195 158218
rect 358875 157898 358917 158134
rect 359153 157898 359195 158134
rect 358875 157866 359195 157898
rect 364806 158454 365126 158486
rect 364806 158218 364848 158454
rect 365084 158218 365126 158454
rect 364806 158134 365126 158218
rect 364806 157898 364848 158134
rect 365084 157898 365126 158134
rect 364806 157866 365126 157898
rect 386875 158454 387195 158486
rect 386875 158218 386917 158454
rect 387153 158218 387195 158454
rect 386875 158134 387195 158218
rect 386875 157898 386917 158134
rect 387153 157898 387195 158134
rect 386875 157866 387195 157898
rect 392806 158454 393126 158486
rect 392806 158218 392848 158454
rect 393084 158218 393126 158454
rect 392806 158134 393126 158218
rect 392806 157898 392848 158134
rect 393084 157898 393126 158134
rect 392806 157866 393126 157898
rect 414875 158454 415195 158486
rect 414875 158218 414917 158454
rect 415153 158218 415195 158454
rect 414875 158134 415195 158218
rect 414875 157898 414917 158134
rect 415153 157898 415195 158134
rect 414875 157866 415195 157898
rect 420806 158454 421126 158486
rect 420806 158218 420848 158454
rect 421084 158218 421126 158454
rect 420806 158134 421126 158218
rect 420806 157898 420848 158134
rect 421084 157898 421126 158134
rect 420806 157866 421126 157898
rect 442875 158454 443195 158486
rect 442875 158218 442917 158454
rect 443153 158218 443195 158454
rect 442875 158134 443195 158218
rect 442875 157898 442917 158134
rect 443153 157898 443195 158134
rect 442875 157866 443195 157898
rect 448806 158454 449126 158486
rect 448806 158218 448848 158454
rect 449084 158218 449126 158454
rect 448806 158134 449126 158218
rect 448806 157898 448848 158134
rect 449084 157898 449126 158134
rect 448806 157866 449126 157898
rect 470875 158454 471195 158486
rect 470875 158218 470917 158454
rect 471153 158218 471195 158454
rect 470875 158134 471195 158218
rect 470875 157898 470917 158134
rect 471153 157898 471195 158134
rect 470875 157866 471195 157898
rect 476806 158454 477126 158486
rect 476806 158218 476848 158454
rect 477084 158218 477126 158454
rect 476806 158134 477126 158218
rect 476806 157898 476848 158134
rect 477084 157898 477126 158134
rect 476806 157866 477126 157898
rect 498875 158454 499195 158486
rect 498875 158218 498917 158454
rect 499153 158218 499195 158454
rect 498875 158134 499195 158218
rect 498875 157898 498917 158134
rect 499153 157898 499195 158134
rect 498875 157866 499195 157898
rect 504806 158454 505126 158486
rect 504806 158218 504848 158454
rect 505084 158218 505126 158454
rect 504806 158134 505126 158218
rect 504806 157898 504848 158134
rect 505084 157898 505126 158134
rect 504806 157866 505126 157898
rect 526875 158454 527195 158486
rect 526875 158218 526917 158454
rect 527153 158218 527195 158454
rect 526875 158134 527195 158218
rect 526875 157898 526917 158134
rect 527153 157898 527195 158134
rect 526875 157866 527195 157898
rect 532806 158454 533126 158486
rect 532806 158218 532848 158454
rect 533084 158218 533126 158454
rect 532806 158134 533126 158218
rect 532806 157898 532848 158134
rect 533084 157898 533126 158134
rect 532806 157866 533126 157898
rect 554875 158454 555195 158486
rect 554875 158218 554917 158454
rect 555153 158218 555195 158454
rect 554875 158134 555195 158218
rect 554875 157898 554917 158134
rect 555153 157898 555195 158134
rect 554875 157866 555195 157898
rect 560806 158454 561126 158486
rect 560806 158218 560848 158454
rect 561084 158218 561126 158454
rect 560806 158134 561126 158218
rect 560806 157898 560848 158134
rect 561084 157898 561126 158134
rect 560806 157866 561126 157898
rect -2006 134593 -1974 134829
rect -1738 134593 -1654 134829
rect -1418 134593 -1386 134829
rect -2006 134509 -1386 134593
rect -2006 134273 -1974 134509
rect -1738 134273 -1654 134509
rect -1418 134273 -1386 134509
rect -2006 107829 -1386 134273
rect 19910 134829 20230 134861
rect 19910 134593 19952 134829
rect 20188 134593 20230 134829
rect 19910 134509 20230 134593
rect 19910 134273 19952 134509
rect 20188 134273 20230 134509
rect 19910 134241 20230 134273
rect 25840 134829 26160 134861
rect 25840 134593 25882 134829
rect 26118 134593 26160 134829
rect 25840 134509 26160 134593
rect 25840 134273 25882 134509
rect 26118 134273 26160 134509
rect 25840 134241 26160 134273
rect 31771 134829 32091 134861
rect 31771 134593 31813 134829
rect 32049 134593 32091 134829
rect 31771 134509 32091 134593
rect 31771 134273 31813 134509
rect 32049 134273 32091 134509
rect 31771 134241 32091 134273
rect 47910 134829 48230 134861
rect 47910 134593 47952 134829
rect 48188 134593 48230 134829
rect 47910 134509 48230 134593
rect 47910 134273 47952 134509
rect 48188 134273 48230 134509
rect 47910 134241 48230 134273
rect 53840 134829 54160 134861
rect 53840 134593 53882 134829
rect 54118 134593 54160 134829
rect 53840 134509 54160 134593
rect 53840 134273 53882 134509
rect 54118 134273 54160 134509
rect 53840 134241 54160 134273
rect 59771 134829 60091 134861
rect 59771 134593 59813 134829
rect 60049 134593 60091 134829
rect 59771 134509 60091 134593
rect 59771 134273 59813 134509
rect 60049 134273 60091 134509
rect 59771 134241 60091 134273
rect 75910 134829 76230 134861
rect 75910 134593 75952 134829
rect 76188 134593 76230 134829
rect 75910 134509 76230 134593
rect 75910 134273 75952 134509
rect 76188 134273 76230 134509
rect 75910 134241 76230 134273
rect 81840 134829 82160 134861
rect 81840 134593 81882 134829
rect 82118 134593 82160 134829
rect 81840 134509 82160 134593
rect 81840 134273 81882 134509
rect 82118 134273 82160 134509
rect 81840 134241 82160 134273
rect 87771 134829 88091 134861
rect 87771 134593 87813 134829
rect 88049 134593 88091 134829
rect 87771 134509 88091 134593
rect 87771 134273 87813 134509
rect 88049 134273 88091 134509
rect 87771 134241 88091 134273
rect 103910 134829 104230 134861
rect 103910 134593 103952 134829
rect 104188 134593 104230 134829
rect 103910 134509 104230 134593
rect 103910 134273 103952 134509
rect 104188 134273 104230 134509
rect 103910 134241 104230 134273
rect 109840 134829 110160 134861
rect 109840 134593 109882 134829
rect 110118 134593 110160 134829
rect 109840 134509 110160 134593
rect 109840 134273 109882 134509
rect 110118 134273 110160 134509
rect 109840 134241 110160 134273
rect 115771 134829 116091 134861
rect 115771 134593 115813 134829
rect 116049 134593 116091 134829
rect 115771 134509 116091 134593
rect 115771 134273 115813 134509
rect 116049 134273 116091 134509
rect 115771 134241 116091 134273
rect 131910 134829 132230 134861
rect 131910 134593 131952 134829
rect 132188 134593 132230 134829
rect 131910 134509 132230 134593
rect 131910 134273 131952 134509
rect 132188 134273 132230 134509
rect 131910 134241 132230 134273
rect 137840 134829 138160 134861
rect 137840 134593 137882 134829
rect 138118 134593 138160 134829
rect 137840 134509 138160 134593
rect 137840 134273 137882 134509
rect 138118 134273 138160 134509
rect 137840 134241 138160 134273
rect 143771 134829 144091 134861
rect 143771 134593 143813 134829
rect 144049 134593 144091 134829
rect 143771 134509 144091 134593
rect 143771 134273 143813 134509
rect 144049 134273 144091 134509
rect 143771 134241 144091 134273
rect 159910 134829 160230 134861
rect 159910 134593 159952 134829
rect 160188 134593 160230 134829
rect 159910 134509 160230 134593
rect 159910 134273 159952 134509
rect 160188 134273 160230 134509
rect 159910 134241 160230 134273
rect 165840 134829 166160 134861
rect 165840 134593 165882 134829
rect 166118 134593 166160 134829
rect 165840 134509 166160 134593
rect 165840 134273 165882 134509
rect 166118 134273 166160 134509
rect 165840 134241 166160 134273
rect 171771 134829 172091 134861
rect 171771 134593 171813 134829
rect 172049 134593 172091 134829
rect 171771 134509 172091 134593
rect 171771 134273 171813 134509
rect 172049 134273 172091 134509
rect 171771 134241 172091 134273
rect 187910 134829 188230 134861
rect 187910 134593 187952 134829
rect 188188 134593 188230 134829
rect 187910 134509 188230 134593
rect 187910 134273 187952 134509
rect 188188 134273 188230 134509
rect 187910 134241 188230 134273
rect 193840 134829 194160 134861
rect 193840 134593 193882 134829
rect 194118 134593 194160 134829
rect 193840 134509 194160 134593
rect 193840 134273 193882 134509
rect 194118 134273 194160 134509
rect 193840 134241 194160 134273
rect 199771 134829 200091 134861
rect 199771 134593 199813 134829
rect 200049 134593 200091 134829
rect 199771 134509 200091 134593
rect 199771 134273 199813 134509
rect 200049 134273 200091 134509
rect 199771 134241 200091 134273
rect 215910 134829 216230 134861
rect 215910 134593 215952 134829
rect 216188 134593 216230 134829
rect 215910 134509 216230 134593
rect 215910 134273 215952 134509
rect 216188 134273 216230 134509
rect 215910 134241 216230 134273
rect 221840 134829 222160 134861
rect 221840 134593 221882 134829
rect 222118 134593 222160 134829
rect 221840 134509 222160 134593
rect 221840 134273 221882 134509
rect 222118 134273 222160 134509
rect 221840 134241 222160 134273
rect 227771 134829 228091 134861
rect 227771 134593 227813 134829
rect 228049 134593 228091 134829
rect 227771 134509 228091 134593
rect 227771 134273 227813 134509
rect 228049 134273 228091 134509
rect 227771 134241 228091 134273
rect 243910 134829 244230 134861
rect 243910 134593 243952 134829
rect 244188 134593 244230 134829
rect 243910 134509 244230 134593
rect 243910 134273 243952 134509
rect 244188 134273 244230 134509
rect 243910 134241 244230 134273
rect 249840 134829 250160 134861
rect 249840 134593 249882 134829
rect 250118 134593 250160 134829
rect 249840 134509 250160 134593
rect 249840 134273 249882 134509
rect 250118 134273 250160 134509
rect 249840 134241 250160 134273
rect 255771 134829 256091 134861
rect 255771 134593 255813 134829
rect 256049 134593 256091 134829
rect 255771 134509 256091 134593
rect 255771 134273 255813 134509
rect 256049 134273 256091 134509
rect 255771 134241 256091 134273
rect 271910 134829 272230 134861
rect 271910 134593 271952 134829
rect 272188 134593 272230 134829
rect 271910 134509 272230 134593
rect 271910 134273 271952 134509
rect 272188 134273 272230 134509
rect 271910 134241 272230 134273
rect 277840 134829 278160 134861
rect 277840 134593 277882 134829
rect 278118 134593 278160 134829
rect 277840 134509 278160 134593
rect 277840 134273 277882 134509
rect 278118 134273 278160 134509
rect 277840 134241 278160 134273
rect 283771 134829 284091 134861
rect 283771 134593 283813 134829
rect 284049 134593 284091 134829
rect 283771 134509 284091 134593
rect 283771 134273 283813 134509
rect 284049 134273 284091 134509
rect 283771 134241 284091 134273
rect 299910 134829 300230 134861
rect 299910 134593 299952 134829
rect 300188 134593 300230 134829
rect 299910 134509 300230 134593
rect 299910 134273 299952 134509
rect 300188 134273 300230 134509
rect 299910 134241 300230 134273
rect 305840 134829 306160 134861
rect 305840 134593 305882 134829
rect 306118 134593 306160 134829
rect 305840 134509 306160 134593
rect 305840 134273 305882 134509
rect 306118 134273 306160 134509
rect 305840 134241 306160 134273
rect 311771 134829 312091 134861
rect 311771 134593 311813 134829
rect 312049 134593 312091 134829
rect 311771 134509 312091 134593
rect 311771 134273 311813 134509
rect 312049 134273 312091 134509
rect 311771 134241 312091 134273
rect 327910 134829 328230 134861
rect 327910 134593 327952 134829
rect 328188 134593 328230 134829
rect 327910 134509 328230 134593
rect 327910 134273 327952 134509
rect 328188 134273 328230 134509
rect 327910 134241 328230 134273
rect 333840 134829 334160 134861
rect 333840 134593 333882 134829
rect 334118 134593 334160 134829
rect 333840 134509 334160 134593
rect 333840 134273 333882 134509
rect 334118 134273 334160 134509
rect 333840 134241 334160 134273
rect 339771 134829 340091 134861
rect 339771 134593 339813 134829
rect 340049 134593 340091 134829
rect 339771 134509 340091 134593
rect 339771 134273 339813 134509
rect 340049 134273 340091 134509
rect 339771 134241 340091 134273
rect 355910 134829 356230 134861
rect 355910 134593 355952 134829
rect 356188 134593 356230 134829
rect 355910 134509 356230 134593
rect 355910 134273 355952 134509
rect 356188 134273 356230 134509
rect 355910 134241 356230 134273
rect 361840 134829 362160 134861
rect 361840 134593 361882 134829
rect 362118 134593 362160 134829
rect 361840 134509 362160 134593
rect 361840 134273 361882 134509
rect 362118 134273 362160 134509
rect 361840 134241 362160 134273
rect 367771 134829 368091 134861
rect 367771 134593 367813 134829
rect 368049 134593 368091 134829
rect 367771 134509 368091 134593
rect 367771 134273 367813 134509
rect 368049 134273 368091 134509
rect 367771 134241 368091 134273
rect 383910 134829 384230 134861
rect 383910 134593 383952 134829
rect 384188 134593 384230 134829
rect 383910 134509 384230 134593
rect 383910 134273 383952 134509
rect 384188 134273 384230 134509
rect 383910 134241 384230 134273
rect 389840 134829 390160 134861
rect 389840 134593 389882 134829
rect 390118 134593 390160 134829
rect 389840 134509 390160 134593
rect 389840 134273 389882 134509
rect 390118 134273 390160 134509
rect 389840 134241 390160 134273
rect 395771 134829 396091 134861
rect 395771 134593 395813 134829
rect 396049 134593 396091 134829
rect 395771 134509 396091 134593
rect 395771 134273 395813 134509
rect 396049 134273 396091 134509
rect 395771 134241 396091 134273
rect 411910 134829 412230 134861
rect 411910 134593 411952 134829
rect 412188 134593 412230 134829
rect 411910 134509 412230 134593
rect 411910 134273 411952 134509
rect 412188 134273 412230 134509
rect 411910 134241 412230 134273
rect 417840 134829 418160 134861
rect 417840 134593 417882 134829
rect 418118 134593 418160 134829
rect 417840 134509 418160 134593
rect 417840 134273 417882 134509
rect 418118 134273 418160 134509
rect 417840 134241 418160 134273
rect 423771 134829 424091 134861
rect 423771 134593 423813 134829
rect 424049 134593 424091 134829
rect 423771 134509 424091 134593
rect 423771 134273 423813 134509
rect 424049 134273 424091 134509
rect 423771 134241 424091 134273
rect 439910 134829 440230 134861
rect 439910 134593 439952 134829
rect 440188 134593 440230 134829
rect 439910 134509 440230 134593
rect 439910 134273 439952 134509
rect 440188 134273 440230 134509
rect 439910 134241 440230 134273
rect 445840 134829 446160 134861
rect 445840 134593 445882 134829
rect 446118 134593 446160 134829
rect 445840 134509 446160 134593
rect 445840 134273 445882 134509
rect 446118 134273 446160 134509
rect 445840 134241 446160 134273
rect 451771 134829 452091 134861
rect 451771 134593 451813 134829
rect 452049 134593 452091 134829
rect 451771 134509 452091 134593
rect 451771 134273 451813 134509
rect 452049 134273 452091 134509
rect 451771 134241 452091 134273
rect 467910 134829 468230 134861
rect 467910 134593 467952 134829
rect 468188 134593 468230 134829
rect 467910 134509 468230 134593
rect 467910 134273 467952 134509
rect 468188 134273 468230 134509
rect 467910 134241 468230 134273
rect 473840 134829 474160 134861
rect 473840 134593 473882 134829
rect 474118 134593 474160 134829
rect 473840 134509 474160 134593
rect 473840 134273 473882 134509
rect 474118 134273 474160 134509
rect 473840 134241 474160 134273
rect 479771 134829 480091 134861
rect 479771 134593 479813 134829
rect 480049 134593 480091 134829
rect 479771 134509 480091 134593
rect 479771 134273 479813 134509
rect 480049 134273 480091 134509
rect 479771 134241 480091 134273
rect 495910 134829 496230 134861
rect 495910 134593 495952 134829
rect 496188 134593 496230 134829
rect 495910 134509 496230 134593
rect 495910 134273 495952 134509
rect 496188 134273 496230 134509
rect 495910 134241 496230 134273
rect 501840 134829 502160 134861
rect 501840 134593 501882 134829
rect 502118 134593 502160 134829
rect 501840 134509 502160 134593
rect 501840 134273 501882 134509
rect 502118 134273 502160 134509
rect 501840 134241 502160 134273
rect 507771 134829 508091 134861
rect 507771 134593 507813 134829
rect 508049 134593 508091 134829
rect 507771 134509 508091 134593
rect 507771 134273 507813 134509
rect 508049 134273 508091 134509
rect 507771 134241 508091 134273
rect 523910 134829 524230 134861
rect 523910 134593 523952 134829
rect 524188 134593 524230 134829
rect 523910 134509 524230 134593
rect 523910 134273 523952 134509
rect 524188 134273 524230 134509
rect 523910 134241 524230 134273
rect 529840 134829 530160 134861
rect 529840 134593 529882 134829
rect 530118 134593 530160 134829
rect 529840 134509 530160 134593
rect 529840 134273 529882 134509
rect 530118 134273 530160 134509
rect 529840 134241 530160 134273
rect 535771 134829 536091 134861
rect 535771 134593 535813 134829
rect 536049 134593 536091 134829
rect 535771 134509 536091 134593
rect 535771 134273 535813 134509
rect 536049 134273 536091 134509
rect 535771 134241 536091 134273
rect 551910 134829 552230 134861
rect 551910 134593 551952 134829
rect 552188 134593 552230 134829
rect 551910 134509 552230 134593
rect 551910 134273 551952 134509
rect 552188 134273 552230 134509
rect 551910 134241 552230 134273
rect 557840 134829 558160 134861
rect 557840 134593 557882 134829
rect 558118 134593 558160 134829
rect 557840 134509 558160 134593
rect 557840 134273 557882 134509
rect 558118 134273 558160 134509
rect 557840 134241 558160 134273
rect 563771 134829 564091 134861
rect 563771 134593 563813 134829
rect 564049 134593 564091 134829
rect 563771 134509 564091 134593
rect 563771 134273 563813 134509
rect 564049 134273 564091 134509
rect 563771 134241 564091 134273
rect 573494 134829 574114 161273
rect 573494 134593 573526 134829
rect 573762 134593 573846 134829
rect 574082 134593 574114 134829
rect 573494 134509 574114 134593
rect 573494 134273 573526 134509
rect 573762 134273 573846 134509
rect 574082 134273 574114 134509
rect 22874 131454 23194 131486
rect 22874 131218 22916 131454
rect 23152 131218 23194 131454
rect 22874 131134 23194 131218
rect 22874 130898 22916 131134
rect 23152 130898 23194 131134
rect 22874 130866 23194 130898
rect 28805 131454 29125 131486
rect 28805 131218 28847 131454
rect 29083 131218 29125 131454
rect 28805 131134 29125 131218
rect 28805 130898 28847 131134
rect 29083 130898 29125 131134
rect 28805 130866 29125 130898
rect 50874 131454 51194 131486
rect 50874 131218 50916 131454
rect 51152 131218 51194 131454
rect 50874 131134 51194 131218
rect 50874 130898 50916 131134
rect 51152 130898 51194 131134
rect 50874 130866 51194 130898
rect 56805 131454 57125 131486
rect 56805 131218 56847 131454
rect 57083 131218 57125 131454
rect 56805 131134 57125 131218
rect 56805 130898 56847 131134
rect 57083 130898 57125 131134
rect 56805 130866 57125 130898
rect 78874 131454 79194 131486
rect 78874 131218 78916 131454
rect 79152 131218 79194 131454
rect 78874 131134 79194 131218
rect 78874 130898 78916 131134
rect 79152 130898 79194 131134
rect 78874 130866 79194 130898
rect 84805 131454 85125 131486
rect 84805 131218 84847 131454
rect 85083 131218 85125 131454
rect 84805 131134 85125 131218
rect 84805 130898 84847 131134
rect 85083 130898 85125 131134
rect 84805 130866 85125 130898
rect 106874 131454 107194 131486
rect 106874 131218 106916 131454
rect 107152 131218 107194 131454
rect 106874 131134 107194 131218
rect 106874 130898 106916 131134
rect 107152 130898 107194 131134
rect 106874 130866 107194 130898
rect 112805 131454 113125 131486
rect 112805 131218 112847 131454
rect 113083 131218 113125 131454
rect 112805 131134 113125 131218
rect 112805 130898 112847 131134
rect 113083 130898 113125 131134
rect 112805 130866 113125 130898
rect 134874 131454 135194 131486
rect 134874 131218 134916 131454
rect 135152 131218 135194 131454
rect 134874 131134 135194 131218
rect 134874 130898 134916 131134
rect 135152 130898 135194 131134
rect 134874 130866 135194 130898
rect 140805 131454 141125 131486
rect 140805 131218 140847 131454
rect 141083 131218 141125 131454
rect 140805 131134 141125 131218
rect 140805 130898 140847 131134
rect 141083 130898 141125 131134
rect 140805 130866 141125 130898
rect 162874 131454 163194 131486
rect 162874 131218 162916 131454
rect 163152 131218 163194 131454
rect 162874 131134 163194 131218
rect 162874 130898 162916 131134
rect 163152 130898 163194 131134
rect 162874 130866 163194 130898
rect 168805 131454 169125 131486
rect 168805 131218 168847 131454
rect 169083 131218 169125 131454
rect 168805 131134 169125 131218
rect 168805 130898 168847 131134
rect 169083 130898 169125 131134
rect 168805 130866 169125 130898
rect 190874 131454 191194 131486
rect 190874 131218 190916 131454
rect 191152 131218 191194 131454
rect 190874 131134 191194 131218
rect 190874 130898 190916 131134
rect 191152 130898 191194 131134
rect 190874 130866 191194 130898
rect 196805 131454 197125 131486
rect 196805 131218 196847 131454
rect 197083 131218 197125 131454
rect 196805 131134 197125 131218
rect 196805 130898 196847 131134
rect 197083 130898 197125 131134
rect 196805 130866 197125 130898
rect 218874 131454 219194 131486
rect 218874 131218 218916 131454
rect 219152 131218 219194 131454
rect 218874 131134 219194 131218
rect 218874 130898 218916 131134
rect 219152 130898 219194 131134
rect 218874 130866 219194 130898
rect 224805 131454 225125 131486
rect 224805 131218 224847 131454
rect 225083 131218 225125 131454
rect 224805 131134 225125 131218
rect 224805 130898 224847 131134
rect 225083 130898 225125 131134
rect 224805 130866 225125 130898
rect 246874 131454 247194 131486
rect 246874 131218 246916 131454
rect 247152 131218 247194 131454
rect 246874 131134 247194 131218
rect 246874 130898 246916 131134
rect 247152 130898 247194 131134
rect 246874 130866 247194 130898
rect 252805 131454 253125 131486
rect 252805 131218 252847 131454
rect 253083 131218 253125 131454
rect 252805 131134 253125 131218
rect 252805 130898 252847 131134
rect 253083 130898 253125 131134
rect 252805 130866 253125 130898
rect 274874 131454 275194 131486
rect 274874 131218 274916 131454
rect 275152 131218 275194 131454
rect 274874 131134 275194 131218
rect 274874 130898 274916 131134
rect 275152 130898 275194 131134
rect 274874 130866 275194 130898
rect 280805 131454 281125 131486
rect 280805 131218 280847 131454
rect 281083 131218 281125 131454
rect 280805 131134 281125 131218
rect 280805 130898 280847 131134
rect 281083 130898 281125 131134
rect 280805 130866 281125 130898
rect 302874 131454 303194 131486
rect 302874 131218 302916 131454
rect 303152 131218 303194 131454
rect 302874 131134 303194 131218
rect 302874 130898 302916 131134
rect 303152 130898 303194 131134
rect 302874 130866 303194 130898
rect 308805 131454 309125 131486
rect 308805 131218 308847 131454
rect 309083 131218 309125 131454
rect 308805 131134 309125 131218
rect 308805 130898 308847 131134
rect 309083 130898 309125 131134
rect 308805 130866 309125 130898
rect 330874 131454 331194 131486
rect 330874 131218 330916 131454
rect 331152 131218 331194 131454
rect 330874 131134 331194 131218
rect 330874 130898 330916 131134
rect 331152 130898 331194 131134
rect 330874 130866 331194 130898
rect 336805 131454 337125 131486
rect 336805 131218 336847 131454
rect 337083 131218 337125 131454
rect 336805 131134 337125 131218
rect 336805 130898 336847 131134
rect 337083 130898 337125 131134
rect 336805 130866 337125 130898
rect 358874 131454 359194 131486
rect 358874 131218 358916 131454
rect 359152 131218 359194 131454
rect 358874 131134 359194 131218
rect 358874 130898 358916 131134
rect 359152 130898 359194 131134
rect 358874 130866 359194 130898
rect 364805 131454 365125 131486
rect 364805 131218 364847 131454
rect 365083 131218 365125 131454
rect 364805 131134 365125 131218
rect 364805 130898 364847 131134
rect 365083 130898 365125 131134
rect 364805 130866 365125 130898
rect 386874 131454 387194 131486
rect 386874 131218 386916 131454
rect 387152 131218 387194 131454
rect 386874 131134 387194 131218
rect 386874 130898 386916 131134
rect 387152 130898 387194 131134
rect 386874 130866 387194 130898
rect 392805 131454 393125 131486
rect 392805 131218 392847 131454
rect 393083 131218 393125 131454
rect 392805 131134 393125 131218
rect 392805 130898 392847 131134
rect 393083 130898 393125 131134
rect 392805 130866 393125 130898
rect 414874 131454 415194 131486
rect 414874 131218 414916 131454
rect 415152 131218 415194 131454
rect 414874 131134 415194 131218
rect 414874 130898 414916 131134
rect 415152 130898 415194 131134
rect 414874 130866 415194 130898
rect 420805 131454 421125 131486
rect 420805 131218 420847 131454
rect 421083 131218 421125 131454
rect 420805 131134 421125 131218
rect 420805 130898 420847 131134
rect 421083 130898 421125 131134
rect 420805 130866 421125 130898
rect 442874 131454 443194 131486
rect 442874 131218 442916 131454
rect 443152 131218 443194 131454
rect 442874 131134 443194 131218
rect 442874 130898 442916 131134
rect 443152 130898 443194 131134
rect 442874 130866 443194 130898
rect 448805 131454 449125 131486
rect 448805 131218 448847 131454
rect 449083 131218 449125 131454
rect 448805 131134 449125 131218
rect 448805 130898 448847 131134
rect 449083 130898 449125 131134
rect 448805 130866 449125 130898
rect 470874 131454 471194 131486
rect 470874 131218 470916 131454
rect 471152 131218 471194 131454
rect 470874 131134 471194 131218
rect 470874 130898 470916 131134
rect 471152 130898 471194 131134
rect 470874 130866 471194 130898
rect 476805 131454 477125 131486
rect 476805 131218 476847 131454
rect 477083 131218 477125 131454
rect 476805 131134 477125 131218
rect 476805 130898 476847 131134
rect 477083 130898 477125 131134
rect 476805 130866 477125 130898
rect 498874 131454 499194 131486
rect 498874 131218 498916 131454
rect 499152 131218 499194 131454
rect 498874 131134 499194 131218
rect 498874 130898 498916 131134
rect 499152 130898 499194 131134
rect 498874 130866 499194 130898
rect 504805 131454 505125 131486
rect 504805 131218 504847 131454
rect 505083 131218 505125 131454
rect 504805 131134 505125 131218
rect 504805 130898 504847 131134
rect 505083 130898 505125 131134
rect 504805 130866 505125 130898
rect 526874 131454 527194 131486
rect 526874 131218 526916 131454
rect 527152 131218 527194 131454
rect 526874 131134 527194 131218
rect 526874 130898 526916 131134
rect 527152 130898 527194 131134
rect 526874 130866 527194 130898
rect 532805 131454 533125 131486
rect 532805 131218 532847 131454
rect 533083 131218 533125 131454
rect 532805 131134 533125 131218
rect 532805 130898 532847 131134
rect 533083 130898 533125 131134
rect 532805 130866 533125 130898
rect 554874 131454 555194 131486
rect 554874 131218 554916 131454
rect 555152 131218 555194 131454
rect 554874 131134 555194 131218
rect 554874 130898 554916 131134
rect 555152 130898 555194 131134
rect 554874 130866 555194 130898
rect 560805 131454 561125 131486
rect 560805 131218 560847 131454
rect 561083 131218 561125 131454
rect 560805 131134 561125 131218
rect 560805 130898 560847 131134
rect 561083 130898 561125 131134
rect 560805 130866 561125 130898
rect -2006 107593 -1974 107829
rect -1738 107593 -1654 107829
rect -1418 107593 -1386 107829
rect -2006 107509 -1386 107593
rect -2006 107273 -1974 107509
rect -1738 107273 -1654 107509
rect -1418 107273 -1386 107509
rect -2006 80829 -1386 107273
rect 19909 107829 20229 107861
rect 19909 107593 19951 107829
rect 20187 107593 20229 107829
rect 19909 107509 20229 107593
rect 19909 107273 19951 107509
rect 20187 107273 20229 107509
rect 19909 107241 20229 107273
rect 25840 107829 26160 107861
rect 25840 107593 25882 107829
rect 26118 107593 26160 107829
rect 25840 107509 26160 107593
rect 25840 107273 25882 107509
rect 26118 107273 26160 107509
rect 25840 107241 26160 107273
rect 31770 107829 32090 107861
rect 31770 107593 31812 107829
rect 32048 107593 32090 107829
rect 31770 107509 32090 107593
rect 31770 107273 31812 107509
rect 32048 107273 32090 107509
rect 31770 107241 32090 107273
rect 47909 107829 48229 107861
rect 47909 107593 47951 107829
rect 48187 107593 48229 107829
rect 47909 107509 48229 107593
rect 47909 107273 47951 107509
rect 48187 107273 48229 107509
rect 47909 107241 48229 107273
rect 53840 107829 54160 107861
rect 53840 107593 53882 107829
rect 54118 107593 54160 107829
rect 53840 107509 54160 107593
rect 53840 107273 53882 107509
rect 54118 107273 54160 107509
rect 53840 107241 54160 107273
rect 59770 107829 60090 107861
rect 59770 107593 59812 107829
rect 60048 107593 60090 107829
rect 59770 107509 60090 107593
rect 59770 107273 59812 107509
rect 60048 107273 60090 107509
rect 59770 107241 60090 107273
rect 75909 107829 76229 107861
rect 75909 107593 75951 107829
rect 76187 107593 76229 107829
rect 75909 107509 76229 107593
rect 75909 107273 75951 107509
rect 76187 107273 76229 107509
rect 75909 107241 76229 107273
rect 81840 107829 82160 107861
rect 81840 107593 81882 107829
rect 82118 107593 82160 107829
rect 81840 107509 82160 107593
rect 81840 107273 81882 107509
rect 82118 107273 82160 107509
rect 81840 107241 82160 107273
rect 87770 107829 88090 107861
rect 87770 107593 87812 107829
rect 88048 107593 88090 107829
rect 87770 107509 88090 107593
rect 87770 107273 87812 107509
rect 88048 107273 88090 107509
rect 87770 107241 88090 107273
rect 103909 107829 104229 107861
rect 103909 107593 103951 107829
rect 104187 107593 104229 107829
rect 103909 107509 104229 107593
rect 103909 107273 103951 107509
rect 104187 107273 104229 107509
rect 103909 107241 104229 107273
rect 109840 107829 110160 107861
rect 109840 107593 109882 107829
rect 110118 107593 110160 107829
rect 109840 107509 110160 107593
rect 109840 107273 109882 107509
rect 110118 107273 110160 107509
rect 109840 107241 110160 107273
rect 115770 107829 116090 107861
rect 115770 107593 115812 107829
rect 116048 107593 116090 107829
rect 115770 107509 116090 107593
rect 115770 107273 115812 107509
rect 116048 107273 116090 107509
rect 115770 107241 116090 107273
rect 131168 107829 131488 107861
rect 131168 107593 131210 107829
rect 131446 107593 131488 107829
rect 131168 107509 131488 107593
rect 131168 107273 131210 107509
rect 131446 107273 131488 107509
rect 131168 107241 131488 107273
rect 135616 107829 135936 107861
rect 135616 107593 135658 107829
rect 135894 107593 135936 107829
rect 135616 107509 135936 107593
rect 135616 107273 135658 107509
rect 135894 107273 135936 107509
rect 135616 107241 135936 107273
rect 140064 107829 140384 107861
rect 140064 107593 140106 107829
rect 140342 107593 140384 107829
rect 140064 107509 140384 107593
rect 140064 107273 140106 107509
rect 140342 107273 140384 107509
rect 140064 107241 140384 107273
rect 144512 107829 144832 107861
rect 144512 107593 144554 107829
rect 144790 107593 144832 107829
rect 144512 107509 144832 107593
rect 144512 107273 144554 107509
rect 144790 107273 144832 107509
rect 144512 107241 144832 107273
rect 159909 107829 160229 107861
rect 159909 107593 159951 107829
rect 160187 107593 160229 107829
rect 159909 107509 160229 107593
rect 159909 107273 159951 107509
rect 160187 107273 160229 107509
rect 159909 107241 160229 107273
rect 165840 107829 166160 107861
rect 165840 107593 165882 107829
rect 166118 107593 166160 107829
rect 165840 107509 166160 107593
rect 165840 107273 165882 107509
rect 166118 107273 166160 107509
rect 165840 107241 166160 107273
rect 171770 107829 172090 107861
rect 171770 107593 171812 107829
rect 172048 107593 172090 107829
rect 171770 107509 172090 107593
rect 171770 107273 171812 107509
rect 172048 107273 172090 107509
rect 171770 107241 172090 107273
rect 187909 107829 188229 107861
rect 187909 107593 187951 107829
rect 188187 107593 188229 107829
rect 187909 107509 188229 107593
rect 187909 107273 187951 107509
rect 188187 107273 188229 107509
rect 187909 107241 188229 107273
rect 193840 107829 194160 107861
rect 193840 107593 193882 107829
rect 194118 107593 194160 107829
rect 193840 107509 194160 107593
rect 193840 107273 193882 107509
rect 194118 107273 194160 107509
rect 193840 107241 194160 107273
rect 199770 107829 200090 107861
rect 199770 107593 199812 107829
rect 200048 107593 200090 107829
rect 199770 107509 200090 107593
rect 199770 107273 199812 107509
rect 200048 107273 200090 107509
rect 199770 107241 200090 107273
rect 215168 107829 215488 107861
rect 215168 107593 215210 107829
rect 215446 107593 215488 107829
rect 215168 107509 215488 107593
rect 215168 107273 215210 107509
rect 215446 107273 215488 107509
rect 215168 107241 215488 107273
rect 219616 107829 219936 107861
rect 219616 107593 219658 107829
rect 219894 107593 219936 107829
rect 219616 107509 219936 107593
rect 219616 107273 219658 107509
rect 219894 107273 219936 107509
rect 219616 107241 219936 107273
rect 224064 107829 224384 107861
rect 224064 107593 224106 107829
rect 224342 107593 224384 107829
rect 224064 107509 224384 107593
rect 224064 107273 224106 107509
rect 224342 107273 224384 107509
rect 224064 107241 224384 107273
rect 228512 107829 228832 107861
rect 228512 107593 228554 107829
rect 228790 107593 228832 107829
rect 228512 107509 228832 107593
rect 228512 107273 228554 107509
rect 228790 107273 228832 107509
rect 228512 107241 228832 107273
rect 243909 107829 244229 107861
rect 243909 107593 243951 107829
rect 244187 107593 244229 107829
rect 243909 107509 244229 107593
rect 243909 107273 243951 107509
rect 244187 107273 244229 107509
rect 243909 107241 244229 107273
rect 249840 107829 250160 107861
rect 249840 107593 249882 107829
rect 250118 107593 250160 107829
rect 249840 107509 250160 107593
rect 249840 107273 249882 107509
rect 250118 107273 250160 107509
rect 249840 107241 250160 107273
rect 255770 107829 256090 107861
rect 255770 107593 255812 107829
rect 256048 107593 256090 107829
rect 255770 107509 256090 107593
rect 255770 107273 255812 107509
rect 256048 107273 256090 107509
rect 255770 107241 256090 107273
rect 271909 107829 272229 107861
rect 271909 107593 271951 107829
rect 272187 107593 272229 107829
rect 271909 107509 272229 107593
rect 271909 107273 271951 107509
rect 272187 107273 272229 107509
rect 271909 107241 272229 107273
rect 277840 107829 278160 107861
rect 277840 107593 277882 107829
rect 278118 107593 278160 107829
rect 277840 107509 278160 107593
rect 277840 107273 277882 107509
rect 278118 107273 278160 107509
rect 277840 107241 278160 107273
rect 283770 107829 284090 107861
rect 283770 107593 283812 107829
rect 284048 107593 284090 107829
rect 283770 107509 284090 107593
rect 283770 107273 283812 107509
rect 284048 107273 284090 107509
rect 283770 107241 284090 107273
rect 299909 107829 300229 107861
rect 299909 107593 299951 107829
rect 300187 107593 300229 107829
rect 299909 107509 300229 107593
rect 299909 107273 299951 107509
rect 300187 107273 300229 107509
rect 299909 107241 300229 107273
rect 305840 107829 306160 107861
rect 305840 107593 305882 107829
rect 306118 107593 306160 107829
rect 305840 107509 306160 107593
rect 305840 107273 305882 107509
rect 306118 107273 306160 107509
rect 305840 107241 306160 107273
rect 311770 107829 312090 107861
rect 311770 107593 311812 107829
rect 312048 107593 312090 107829
rect 311770 107509 312090 107593
rect 311770 107273 311812 107509
rect 312048 107273 312090 107509
rect 311770 107241 312090 107273
rect 327909 107829 328229 107861
rect 327909 107593 327951 107829
rect 328187 107593 328229 107829
rect 327909 107509 328229 107593
rect 327909 107273 327951 107509
rect 328187 107273 328229 107509
rect 327909 107241 328229 107273
rect 333840 107829 334160 107861
rect 333840 107593 333882 107829
rect 334118 107593 334160 107829
rect 333840 107509 334160 107593
rect 333840 107273 333882 107509
rect 334118 107273 334160 107509
rect 333840 107241 334160 107273
rect 339770 107829 340090 107861
rect 339770 107593 339812 107829
rect 340048 107593 340090 107829
rect 339770 107509 340090 107593
rect 339770 107273 339812 107509
rect 340048 107273 340090 107509
rect 339770 107241 340090 107273
rect 355909 107829 356229 107861
rect 355909 107593 355951 107829
rect 356187 107593 356229 107829
rect 355909 107509 356229 107593
rect 355909 107273 355951 107509
rect 356187 107273 356229 107509
rect 355909 107241 356229 107273
rect 361840 107829 362160 107861
rect 361840 107593 361882 107829
rect 362118 107593 362160 107829
rect 361840 107509 362160 107593
rect 361840 107273 361882 107509
rect 362118 107273 362160 107509
rect 361840 107241 362160 107273
rect 367770 107829 368090 107861
rect 367770 107593 367812 107829
rect 368048 107593 368090 107829
rect 367770 107509 368090 107593
rect 367770 107273 367812 107509
rect 368048 107273 368090 107509
rect 367770 107241 368090 107273
rect 383909 107829 384229 107861
rect 383909 107593 383951 107829
rect 384187 107593 384229 107829
rect 383909 107509 384229 107593
rect 383909 107273 383951 107509
rect 384187 107273 384229 107509
rect 383909 107241 384229 107273
rect 389840 107829 390160 107861
rect 389840 107593 389882 107829
rect 390118 107593 390160 107829
rect 389840 107509 390160 107593
rect 389840 107273 389882 107509
rect 390118 107273 390160 107509
rect 389840 107241 390160 107273
rect 395770 107829 396090 107861
rect 395770 107593 395812 107829
rect 396048 107593 396090 107829
rect 395770 107509 396090 107593
rect 395770 107273 395812 107509
rect 396048 107273 396090 107509
rect 395770 107241 396090 107273
rect 411909 107829 412229 107861
rect 411909 107593 411951 107829
rect 412187 107593 412229 107829
rect 411909 107509 412229 107593
rect 411909 107273 411951 107509
rect 412187 107273 412229 107509
rect 411909 107241 412229 107273
rect 417840 107829 418160 107861
rect 417840 107593 417882 107829
rect 418118 107593 418160 107829
rect 417840 107509 418160 107593
rect 417840 107273 417882 107509
rect 418118 107273 418160 107509
rect 417840 107241 418160 107273
rect 423770 107829 424090 107861
rect 423770 107593 423812 107829
rect 424048 107593 424090 107829
rect 423770 107509 424090 107593
rect 423770 107273 423812 107509
rect 424048 107273 424090 107509
rect 423770 107241 424090 107273
rect 439909 107829 440229 107861
rect 439909 107593 439951 107829
rect 440187 107593 440229 107829
rect 439909 107509 440229 107593
rect 439909 107273 439951 107509
rect 440187 107273 440229 107509
rect 439909 107241 440229 107273
rect 445840 107829 446160 107861
rect 445840 107593 445882 107829
rect 446118 107593 446160 107829
rect 445840 107509 446160 107593
rect 445840 107273 445882 107509
rect 446118 107273 446160 107509
rect 445840 107241 446160 107273
rect 451770 107829 452090 107861
rect 451770 107593 451812 107829
rect 452048 107593 452090 107829
rect 451770 107509 452090 107593
rect 451770 107273 451812 107509
rect 452048 107273 452090 107509
rect 451770 107241 452090 107273
rect 467909 107829 468229 107861
rect 467909 107593 467951 107829
rect 468187 107593 468229 107829
rect 467909 107509 468229 107593
rect 467909 107273 467951 107509
rect 468187 107273 468229 107509
rect 467909 107241 468229 107273
rect 473840 107829 474160 107861
rect 473840 107593 473882 107829
rect 474118 107593 474160 107829
rect 473840 107509 474160 107593
rect 473840 107273 473882 107509
rect 474118 107273 474160 107509
rect 473840 107241 474160 107273
rect 479770 107829 480090 107861
rect 479770 107593 479812 107829
rect 480048 107593 480090 107829
rect 479770 107509 480090 107593
rect 479770 107273 479812 107509
rect 480048 107273 480090 107509
rect 479770 107241 480090 107273
rect 495909 107829 496229 107861
rect 495909 107593 495951 107829
rect 496187 107593 496229 107829
rect 495909 107509 496229 107593
rect 495909 107273 495951 107509
rect 496187 107273 496229 107509
rect 495909 107241 496229 107273
rect 501840 107829 502160 107861
rect 501840 107593 501882 107829
rect 502118 107593 502160 107829
rect 501840 107509 502160 107593
rect 501840 107273 501882 107509
rect 502118 107273 502160 107509
rect 501840 107241 502160 107273
rect 507770 107829 508090 107861
rect 507770 107593 507812 107829
rect 508048 107593 508090 107829
rect 507770 107509 508090 107593
rect 507770 107273 507812 107509
rect 508048 107273 508090 107509
rect 507770 107241 508090 107273
rect 523909 107829 524229 107861
rect 523909 107593 523951 107829
rect 524187 107593 524229 107829
rect 523909 107509 524229 107593
rect 523909 107273 523951 107509
rect 524187 107273 524229 107509
rect 523909 107241 524229 107273
rect 529840 107829 530160 107861
rect 529840 107593 529882 107829
rect 530118 107593 530160 107829
rect 529840 107509 530160 107593
rect 529840 107273 529882 107509
rect 530118 107273 530160 107509
rect 529840 107241 530160 107273
rect 535770 107829 536090 107861
rect 535770 107593 535812 107829
rect 536048 107593 536090 107829
rect 535770 107509 536090 107593
rect 535770 107273 535812 107509
rect 536048 107273 536090 107509
rect 535770 107241 536090 107273
rect 551909 107829 552229 107861
rect 551909 107593 551951 107829
rect 552187 107593 552229 107829
rect 551909 107509 552229 107593
rect 551909 107273 551951 107509
rect 552187 107273 552229 107509
rect 551909 107241 552229 107273
rect 557840 107829 558160 107861
rect 557840 107593 557882 107829
rect 558118 107593 558160 107829
rect 557840 107509 558160 107593
rect 557840 107273 557882 107509
rect 558118 107273 558160 107509
rect 557840 107241 558160 107273
rect 563770 107829 564090 107861
rect 563770 107593 563812 107829
rect 564048 107593 564090 107829
rect 563770 107509 564090 107593
rect 563770 107273 563812 107509
rect 564048 107273 564090 107509
rect 563770 107241 564090 107273
rect 573494 107829 574114 134273
rect 573494 107593 573526 107829
rect 573762 107593 573846 107829
rect 574082 107593 574114 107829
rect 573494 107509 574114 107593
rect 573494 107273 573526 107509
rect 573762 107273 573846 107509
rect 574082 107273 574114 107509
rect 22875 104454 23195 104486
rect 22875 104218 22917 104454
rect 23153 104218 23195 104454
rect 22875 104134 23195 104218
rect 22875 103898 22917 104134
rect 23153 103898 23195 104134
rect 22875 103866 23195 103898
rect 28806 104454 29126 104486
rect 28806 104218 28848 104454
rect 29084 104218 29126 104454
rect 28806 104134 29126 104218
rect 28806 103898 28848 104134
rect 29084 103898 29126 104134
rect 28806 103866 29126 103898
rect 50875 104454 51195 104486
rect 50875 104218 50917 104454
rect 51153 104218 51195 104454
rect 50875 104134 51195 104218
rect 50875 103898 50917 104134
rect 51153 103898 51195 104134
rect 50875 103866 51195 103898
rect 56806 104454 57126 104486
rect 56806 104218 56848 104454
rect 57084 104218 57126 104454
rect 56806 104134 57126 104218
rect 56806 103898 56848 104134
rect 57084 103898 57126 104134
rect 56806 103866 57126 103898
rect 78875 104454 79195 104486
rect 78875 104218 78917 104454
rect 79153 104218 79195 104454
rect 78875 104134 79195 104218
rect 78875 103898 78917 104134
rect 79153 103898 79195 104134
rect 78875 103866 79195 103898
rect 84806 104454 85126 104486
rect 84806 104218 84848 104454
rect 85084 104218 85126 104454
rect 84806 104134 85126 104218
rect 84806 103898 84848 104134
rect 85084 103898 85126 104134
rect 84806 103866 85126 103898
rect 106875 104454 107195 104486
rect 106875 104218 106917 104454
rect 107153 104218 107195 104454
rect 106875 104134 107195 104218
rect 106875 103898 106917 104134
rect 107153 103898 107195 104134
rect 106875 103866 107195 103898
rect 112806 104454 113126 104486
rect 112806 104218 112848 104454
rect 113084 104218 113126 104454
rect 112806 104134 113126 104218
rect 112806 103898 112848 104134
rect 113084 103898 113126 104134
rect 112806 103866 113126 103898
rect 133392 104454 133712 104486
rect 133392 104218 133434 104454
rect 133670 104218 133712 104454
rect 133392 104134 133712 104218
rect 133392 103898 133434 104134
rect 133670 103898 133712 104134
rect 133392 103866 133712 103898
rect 137840 104454 138160 104486
rect 137840 104218 137882 104454
rect 138118 104218 138160 104454
rect 137840 104134 138160 104218
rect 137840 103898 137882 104134
rect 138118 103898 138160 104134
rect 137840 103866 138160 103898
rect 142288 104454 142608 104486
rect 142288 104218 142330 104454
rect 142566 104218 142608 104454
rect 142288 104134 142608 104218
rect 142288 103898 142330 104134
rect 142566 103898 142608 104134
rect 142288 103866 142608 103898
rect 162875 104454 163195 104486
rect 162875 104218 162917 104454
rect 163153 104218 163195 104454
rect 162875 104134 163195 104218
rect 162875 103898 162917 104134
rect 163153 103898 163195 104134
rect 162875 103866 163195 103898
rect 168806 104454 169126 104486
rect 168806 104218 168848 104454
rect 169084 104218 169126 104454
rect 168806 104134 169126 104218
rect 168806 103898 168848 104134
rect 169084 103898 169126 104134
rect 168806 103866 169126 103898
rect 190875 104454 191195 104486
rect 190875 104218 190917 104454
rect 191153 104218 191195 104454
rect 190875 104134 191195 104218
rect 190875 103898 190917 104134
rect 191153 103898 191195 104134
rect 190875 103866 191195 103898
rect 196806 104454 197126 104486
rect 196806 104218 196848 104454
rect 197084 104218 197126 104454
rect 196806 104134 197126 104218
rect 196806 103898 196848 104134
rect 197084 103898 197126 104134
rect 196806 103866 197126 103898
rect 217392 104454 217712 104486
rect 217392 104218 217434 104454
rect 217670 104218 217712 104454
rect 217392 104134 217712 104218
rect 217392 103898 217434 104134
rect 217670 103898 217712 104134
rect 217392 103866 217712 103898
rect 221840 104454 222160 104486
rect 221840 104218 221882 104454
rect 222118 104218 222160 104454
rect 221840 104134 222160 104218
rect 221840 103898 221882 104134
rect 222118 103898 222160 104134
rect 221840 103866 222160 103898
rect 226288 104454 226608 104486
rect 226288 104218 226330 104454
rect 226566 104218 226608 104454
rect 226288 104134 226608 104218
rect 226288 103898 226330 104134
rect 226566 103898 226608 104134
rect 226288 103866 226608 103898
rect 246875 104454 247195 104486
rect 246875 104218 246917 104454
rect 247153 104218 247195 104454
rect 246875 104134 247195 104218
rect 246875 103898 246917 104134
rect 247153 103898 247195 104134
rect 246875 103866 247195 103898
rect 252806 104454 253126 104486
rect 252806 104218 252848 104454
rect 253084 104218 253126 104454
rect 252806 104134 253126 104218
rect 252806 103898 252848 104134
rect 253084 103898 253126 104134
rect 252806 103866 253126 103898
rect 274875 104454 275195 104486
rect 274875 104218 274917 104454
rect 275153 104218 275195 104454
rect 274875 104134 275195 104218
rect 274875 103898 274917 104134
rect 275153 103898 275195 104134
rect 274875 103866 275195 103898
rect 280806 104454 281126 104486
rect 280806 104218 280848 104454
rect 281084 104218 281126 104454
rect 280806 104134 281126 104218
rect 280806 103898 280848 104134
rect 281084 103898 281126 104134
rect 280806 103866 281126 103898
rect 302875 104454 303195 104486
rect 302875 104218 302917 104454
rect 303153 104218 303195 104454
rect 302875 104134 303195 104218
rect 302875 103898 302917 104134
rect 303153 103898 303195 104134
rect 302875 103866 303195 103898
rect 308806 104454 309126 104486
rect 308806 104218 308848 104454
rect 309084 104218 309126 104454
rect 308806 104134 309126 104218
rect 308806 103898 308848 104134
rect 309084 103898 309126 104134
rect 308806 103866 309126 103898
rect 330875 104454 331195 104486
rect 330875 104218 330917 104454
rect 331153 104218 331195 104454
rect 330875 104134 331195 104218
rect 330875 103898 330917 104134
rect 331153 103898 331195 104134
rect 330875 103866 331195 103898
rect 336806 104454 337126 104486
rect 336806 104218 336848 104454
rect 337084 104218 337126 104454
rect 336806 104134 337126 104218
rect 336806 103898 336848 104134
rect 337084 103898 337126 104134
rect 336806 103866 337126 103898
rect 358875 104454 359195 104486
rect 358875 104218 358917 104454
rect 359153 104218 359195 104454
rect 358875 104134 359195 104218
rect 358875 103898 358917 104134
rect 359153 103898 359195 104134
rect 358875 103866 359195 103898
rect 364806 104454 365126 104486
rect 364806 104218 364848 104454
rect 365084 104218 365126 104454
rect 364806 104134 365126 104218
rect 364806 103898 364848 104134
rect 365084 103898 365126 104134
rect 364806 103866 365126 103898
rect 386875 104454 387195 104486
rect 386875 104218 386917 104454
rect 387153 104218 387195 104454
rect 386875 104134 387195 104218
rect 386875 103898 386917 104134
rect 387153 103898 387195 104134
rect 386875 103866 387195 103898
rect 392806 104454 393126 104486
rect 392806 104218 392848 104454
rect 393084 104218 393126 104454
rect 392806 104134 393126 104218
rect 392806 103898 392848 104134
rect 393084 103898 393126 104134
rect 392806 103866 393126 103898
rect 414875 104454 415195 104486
rect 414875 104218 414917 104454
rect 415153 104218 415195 104454
rect 414875 104134 415195 104218
rect 414875 103898 414917 104134
rect 415153 103898 415195 104134
rect 414875 103866 415195 103898
rect 420806 104454 421126 104486
rect 420806 104218 420848 104454
rect 421084 104218 421126 104454
rect 420806 104134 421126 104218
rect 420806 103898 420848 104134
rect 421084 103898 421126 104134
rect 420806 103866 421126 103898
rect 442875 104454 443195 104486
rect 442875 104218 442917 104454
rect 443153 104218 443195 104454
rect 442875 104134 443195 104218
rect 442875 103898 442917 104134
rect 443153 103898 443195 104134
rect 442875 103866 443195 103898
rect 448806 104454 449126 104486
rect 448806 104218 448848 104454
rect 449084 104218 449126 104454
rect 448806 104134 449126 104218
rect 448806 103898 448848 104134
rect 449084 103898 449126 104134
rect 448806 103866 449126 103898
rect 470875 104454 471195 104486
rect 470875 104218 470917 104454
rect 471153 104218 471195 104454
rect 470875 104134 471195 104218
rect 470875 103898 470917 104134
rect 471153 103898 471195 104134
rect 470875 103866 471195 103898
rect 476806 104454 477126 104486
rect 476806 104218 476848 104454
rect 477084 104218 477126 104454
rect 476806 104134 477126 104218
rect 476806 103898 476848 104134
rect 477084 103898 477126 104134
rect 476806 103866 477126 103898
rect 498875 104454 499195 104486
rect 498875 104218 498917 104454
rect 499153 104218 499195 104454
rect 498875 104134 499195 104218
rect 498875 103898 498917 104134
rect 499153 103898 499195 104134
rect 498875 103866 499195 103898
rect 504806 104454 505126 104486
rect 504806 104218 504848 104454
rect 505084 104218 505126 104454
rect 504806 104134 505126 104218
rect 504806 103898 504848 104134
rect 505084 103898 505126 104134
rect 504806 103866 505126 103898
rect 526875 104454 527195 104486
rect 526875 104218 526917 104454
rect 527153 104218 527195 104454
rect 526875 104134 527195 104218
rect 526875 103898 526917 104134
rect 527153 103898 527195 104134
rect 526875 103866 527195 103898
rect 532806 104454 533126 104486
rect 532806 104218 532848 104454
rect 533084 104218 533126 104454
rect 532806 104134 533126 104218
rect 532806 103898 532848 104134
rect 533084 103898 533126 104134
rect 532806 103866 533126 103898
rect 554875 104454 555195 104486
rect 554875 104218 554917 104454
rect 555153 104218 555195 104454
rect 554875 104134 555195 104218
rect 554875 103898 554917 104134
rect 555153 103898 555195 104134
rect 554875 103866 555195 103898
rect 560806 104454 561126 104486
rect 560806 104218 560848 104454
rect 561084 104218 561126 104454
rect 560806 104134 561126 104218
rect 560806 103898 560848 104134
rect 561084 103898 561126 104134
rect 560806 103866 561126 103898
rect -2006 80593 -1974 80829
rect -1738 80593 -1654 80829
rect -1418 80593 -1386 80829
rect -2006 80509 -1386 80593
rect -2006 80273 -1974 80509
rect -1738 80273 -1654 80509
rect -1418 80273 -1386 80509
rect -2006 53829 -1386 80273
rect 19910 80829 20230 80861
rect 19910 80593 19952 80829
rect 20188 80593 20230 80829
rect 19910 80509 20230 80593
rect 19910 80273 19952 80509
rect 20188 80273 20230 80509
rect 19910 80241 20230 80273
rect 25840 80829 26160 80861
rect 25840 80593 25882 80829
rect 26118 80593 26160 80829
rect 25840 80509 26160 80593
rect 25840 80273 25882 80509
rect 26118 80273 26160 80509
rect 25840 80241 26160 80273
rect 31771 80829 32091 80861
rect 31771 80593 31813 80829
rect 32049 80593 32091 80829
rect 31771 80509 32091 80593
rect 31771 80273 31813 80509
rect 32049 80273 32091 80509
rect 31771 80241 32091 80273
rect 47910 80829 48230 80861
rect 47910 80593 47952 80829
rect 48188 80593 48230 80829
rect 47910 80509 48230 80593
rect 47910 80273 47952 80509
rect 48188 80273 48230 80509
rect 47910 80241 48230 80273
rect 53840 80829 54160 80861
rect 53840 80593 53882 80829
rect 54118 80593 54160 80829
rect 53840 80509 54160 80593
rect 53840 80273 53882 80509
rect 54118 80273 54160 80509
rect 53840 80241 54160 80273
rect 59771 80829 60091 80861
rect 59771 80593 59813 80829
rect 60049 80593 60091 80829
rect 59771 80509 60091 80593
rect 59771 80273 59813 80509
rect 60049 80273 60091 80509
rect 59771 80241 60091 80273
rect 75910 80829 76230 80861
rect 75910 80593 75952 80829
rect 76188 80593 76230 80829
rect 75910 80509 76230 80593
rect 75910 80273 75952 80509
rect 76188 80273 76230 80509
rect 75910 80241 76230 80273
rect 81840 80829 82160 80861
rect 81840 80593 81882 80829
rect 82118 80593 82160 80829
rect 81840 80509 82160 80593
rect 81840 80273 81882 80509
rect 82118 80273 82160 80509
rect 81840 80241 82160 80273
rect 87771 80829 88091 80861
rect 87771 80593 87813 80829
rect 88049 80593 88091 80829
rect 87771 80509 88091 80593
rect 87771 80273 87813 80509
rect 88049 80273 88091 80509
rect 87771 80241 88091 80273
rect 103910 80829 104230 80861
rect 103910 80593 103952 80829
rect 104188 80593 104230 80829
rect 103910 80509 104230 80593
rect 103910 80273 103952 80509
rect 104188 80273 104230 80509
rect 103910 80241 104230 80273
rect 109840 80829 110160 80861
rect 109840 80593 109882 80829
rect 110118 80593 110160 80829
rect 109840 80509 110160 80593
rect 109840 80273 109882 80509
rect 110118 80273 110160 80509
rect 109840 80241 110160 80273
rect 115771 80829 116091 80861
rect 115771 80593 115813 80829
rect 116049 80593 116091 80829
rect 115771 80509 116091 80593
rect 115771 80273 115813 80509
rect 116049 80273 116091 80509
rect 115771 80241 116091 80273
rect 131910 80829 132230 80861
rect 131910 80593 131952 80829
rect 132188 80593 132230 80829
rect 131910 80509 132230 80593
rect 131910 80273 131952 80509
rect 132188 80273 132230 80509
rect 131910 80241 132230 80273
rect 137840 80829 138160 80861
rect 137840 80593 137882 80829
rect 138118 80593 138160 80829
rect 137840 80509 138160 80593
rect 137840 80273 137882 80509
rect 138118 80273 138160 80509
rect 137840 80241 138160 80273
rect 143771 80829 144091 80861
rect 143771 80593 143813 80829
rect 144049 80593 144091 80829
rect 143771 80509 144091 80593
rect 143771 80273 143813 80509
rect 144049 80273 144091 80509
rect 143771 80241 144091 80273
rect 159910 80829 160230 80861
rect 159910 80593 159952 80829
rect 160188 80593 160230 80829
rect 159910 80509 160230 80593
rect 159910 80273 159952 80509
rect 160188 80273 160230 80509
rect 159910 80241 160230 80273
rect 165840 80829 166160 80861
rect 165840 80593 165882 80829
rect 166118 80593 166160 80829
rect 165840 80509 166160 80593
rect 165840 80273 165882 80509
rect 166118 80273 166160 80509
rect 165840 80241 166160 80273
rect 171771 80829 172091 80861
rect 171771 80593 171813 80829
rect 172049 80593 172091 80829
rect 171771 80509 172091 80593
rect 171771 80273 171813 80509
rect 172049 80273 172091 80509
rect 171771 80241 172091 80273
rect 187910 80829 188230 80861
rect 187910 80593 187952 80829
rect 188188 80593 188230 80829
rect 187910 80509 188230 80593
rect 187910 80273 187952 80509
rect 188188 80273 188230 80509
rect 187910 80241 188230 80273
rect 193840 80829 194160 80861
rect 193840 80593 193882 80829
rect 194118 80593 194160 80829
rect 193840 80509 194160 80593
rect 193840 80273 193882 80509
rect 194118 80273 194160 80509
rect 193840 80241 194160 80273
rect 199771 80829 200091 80861
rect 199771 80593 199813 80829
rect 200049 80593 200091 80829
rect 199771 80509 200091 80593
rect 199771 80273 199813 80509
rect 200049 80273 200091 80509
rect 199771 80241 200091 80273
rect 215910 80829 216230 80861
rect 215910 80593 215952 80829
rect 216188 80593 216230 80829
rect 215910 80509 216230 80593
rect 215910 80273 215952 80509
rect 216188 80273 216230 80509
rect 215910 80241 216230 80273
rect 221840 80829 222160 80861
rect 221840 80593 221882 80829
rect 222118 80593 222160 80829
rect 221840 80509 222160 80593
rect 221840 80273 221882 80509
rect 222118 80273 222160 80509
rect 221840 80241 222160 80273
rect 227771 80829 228091 80861
rect 227771 80593 227813 80829
rect 228049 80593 228091 80829
rect 227771 80509 228091 80593
rect 227771 80273 227813 80509
rect 228049 80273 228091 80509
rect 227771 80241 228091 80273
rect 243910 80829 244230 80861
rect 243910 80593 243952 80829
rect 244188 80593 244230 80829
rect 243910 80509 244230 80593
rect 243910 80273 243952 80509
rect 244188 80273 244230 80509
rect 243910 80241 244230 80273
rect 249840 80829 250160 80861
rect 249840 80593 249882 80829
rect 250118 80593 250160 80829
rect 249840 80509 250160 80593
rect 249840 80273 249882 80509
rect 250118 80273 250160 80509
rect 249840 80241 250160 80273
rect 255771 80829 256091 80861
rect 255771 80593 255813 80829
rect 256049 80593 256091 80829
rect 255771 80509 256091 80593
rect 255771 80273 255813 80509
rect 256049 80273 256091 80509
rect 255771 80241 256091 80273
rect 271910 80829 272230 80861
rect 271910 80593 271952 80829
rect 272188 80593 272230 80829
rect 271910 80509 272230 80593
rect 271910 80273 271952 80509
rect 272188 80273 272230 80509
rect 271910 80241 272230 80273
rect 277840 80829 278160 80861
rect 277840 80593 277882 80829
rect 278118 80593 278160 80829
rect 277840 80509 278160 80593
rect 277840 80273 277882 80509
rect 278118 80273 278160 80509
rect 277840 80241 278160 80273
rect 283771 80829 284091 80861
rect 283771 80593 283813 80829
rect 284049 80593 284091 80829
rect 283771 80509 284091 80593
rect 283771 80273 283813 80509
rect 284049 80273 284091 80509
rect 283771 80241 284091 80273
rect 299910 80829 300230 80861
rect 299910 80593 299952 80829
rect 300188 80593 300230 80829
rect 299910 80509 300230 80593
rect 299910 80273 299952 80509
rect 300188 80273 300230 80509
rect 299910 80241 300230 80273
rect 305840 80829 306160 80861
rect 305840 80593 305882 80829
rect 306118 80593 306160 80829
rect 305840 80509 306160 80593
rect 305840 80273 305882 80509
rect 306118 80273 306160 80509
rect 305840 80241 306160 80273
rect 311771 80829 312091 80861
rect 311771 80593 311813 80829
rect 312049 80593 312091 80829
rect 311771 80509 312091 80593
rect 311771 80273 311813 80509
rect 312049 80273 312091 80509
rect 311771 80241 312091 80273
rect 327910 80829 328230 80861
rect 327910 80593 327952 80829
rect 328188 80593 328230 80829
rect 327910 80509 328230 80593
rect 327910 80273 327952 80509
rect 328188 80273 328230 80509
rect 327910 80241 328230 80273
rect 333840 80829 334160 80861
rect 333840 80593 333882 80829
rect 334118 80593 334160 80829
rect 333840 80509 334160 80593
rect 333840 80273 333882 80509
rect 334118 80273 334160 80509
rect 333840 80241 334160 80273
rect 339771 80829 340091 80861
rect 339771 80593 339813 80829
rect 340049 80593 340091 80829
rect 339771 80509 340091 80593
rect 339771 80273 339813 80509
rect 340049 80273 340091 80509
rect 339771 80241 340091 80273
rect 355910 80829 356230 80861
rect 355910 80593 355952 80829
rect 356188 80593 356230 80829
rect 355910 80509 356230 80593
rect 355910 80273 355952 80509
rect 356188 80273 356230 80509
rect 355910 80241 356230 80273
rect 361840 80829 362160 80861
rect 361840 80593 361882 80829
rect 362118 80593 362160 80829
rect 361840 80509 362160 80593
rect 361840 80273 361882 80509
rect 362118 80273 362160 80509
rect 361840 80241 362160 80273
rect 367771 80829 368091 80861
rect 367771 80593 367813 80829
rect 368049 80593 368091 80829
rect 367771 80509 368091 80593
rect 367771 80273 367813 80509
rect 368049 80273 368091 80509
rect 367771 80241 368091 80273
rect 383910 80829 384230 80861
rect 383910 80593 383952 80829
rect 384188 80593 384230 80829
rect 383910 80509 384230 80593
rect 383910 80273 383952 80509
rect 384188 80273 384230 80509
rect 383910 80241 384230 80273
rect 389840 80829 390160 80861
rect 389840 80593 389882 80829
rect 390118 80593 390160 80829
rect 389840 80509 390160 80593
rect 389840 80273 389882 80509
rect 390118 80273 390160 80509
rect 389840 80241 390160 80273
rect 395771 80829 396091 80861
rect 395771 80593 395813 80829
rect 396049 80593 396091 80829
rect 395771 80509 396091 80593
rect 395771 80273 395813 80509
rect 396049 80273 396091 80509
rect 395771 80241 396091 80273
rect 411910 80829 412230 80861
rect 411910 80593 411952 80829
rect 412188 80593 412230 80829
rect 411910 80509 412230 80593
rect 411910 80273 411952 80509
rect 412188 80273 412230 80509
rect 411910 80241 412230 80273
rect 417840 80829 418160 80861
rect 417840 80593 417882 80829
rect 418118 80593 418160 80829
rect 417840 80509 418160 80593
rect 417840 80273 417882 80509
rect 418118 80273 418160 80509
rect 417840 80241 418160 80273
rect 423771 80829 424091 80861
rect 423771 80593 423813 80829
rect 424049 80593 424091 80829
rect 423771 80509 424091 80593
rect 423771 80273 423813 80509
rect 424049 80273 424091 80509
rect 423771 80241 424091 80273
rect 439910 80829 440230 80861
rect 439910 80593 439952 80829
rect 440188 80593 440230 80829
rect 439910 80509 440230 80593
rect 439910 80273 439952 80509
rect 440188 80273 440230 80509
rect 439910 80241 440230 80273
rect 445840 80829 446160 80861
rect 445840 80593 445882 80829
rect 446118 80593 446160 80829
rect 445840 80509 446160 80593
rect 445840 80273 445882 80509
rect 446118 80273 446160 80509
rect 445840 80241 446160 80273
rect 451771 80829 452091 80861
rect 451771 80593 451813 80829
rect 452049 80593 452091 80829
rect 451771 80509 452091 80593
rect 451771 80273 451813 80509
rect 452049 80273 452091 80509
rect 451771 80241 452091 80273
rect 467910 80829 468230 80861
rect 467910 80593 467952 80829
rect 468188 80593 468230 80829
rect 467910 80509 468230 80593
rect 467910 80273 467952 80509
rect 468188 80273 468230 80509
rect 467910 80241 468230 80273
rect 473840 80829 474160 80861
rect 473840 80593 473882 80829
rect 474118 80593 474160 80829
rect 473840 80509 474160 80593
rect 473840 80273 473882 80509
rect 474118 80273 474160 80509
rect 473840 80241 474160 80273
rect 479771 80829 480091 80861
rect 479771 80593 479813 80829
rect 480049 80593 480091 80829
rect 479771 80509 480091 80593
rect 479771 80273 479813 80509
rect 480049 80273 480091 80509
rect 479771 80241 480091 80273
rect 495910 80829 496230 80861
rect 495910 80593 495952 80829
rect 496188 80593 496230 80829
rect 495910 80509 496230 80593
rect 495910 80273 495952 80509
rect 496188 80273 496230 80509
rect 495910 80241 496230 80273
rect 501840 80829 502160 80861
rect 501840 80593 501882 80829
rect 502118 80593 502160 80829
rect 501840 80509 502160 80593
rect 501840 80273 501882 80509
rect 502118 80273 502160 80509
rect 501840 80241 502160 80273
rect 507771 80829 508091 80861
rect 507771 80593 507813 80829
rect 508049 80593 508091 80829
rect 507771 80509 508091 80593
rect 507771 80273 507813 80509
rect 508049 80273 508091 80509
rect 507771 80241 508091 80273
rect 523910 80829 524230 80861
rect 523910 80593 523952 80829
rect 524188 80593 524230 80829
rect 523910 80509 524230 80593
rect 523910 80273 523952 80509
rect 524188 80273 524230 80509
rect 523910 80241 524230 80273
rect 529840 80829 530160 80861
rect 529840 80593 529882 80829
rect 530118 80593 530160 80829
rect 529840 80509 530160 80593
rect 529840 80273 529882 80509
rect 530118 80273 530160 80509
rect 529840 80241 530160 80273
rect 535771 80829 536091 80861
rect 535771 80593 535813 80829
rect 536049 80593 536091 80829
rect 535771 80509 536091 80593
rect 535771 80273 535813 80509
rect 536049 80273 536091 80509
rect 535771 80241 536091 80273
rect 551910 80829 552230 80861
rect 551910 80593 551952 80829
rect 552188 80593 552230 80829
rect 551910 80509 552230 80593
rect 551910 80273 551952 80509
rect 552188 80273 552230 80509
rect 551910 80241 552230 80273
rect 557840 80829 558160 80861
rect 557840 80593 557882 80829
rect 558118 80593 558160 80829
rect 557840 80509 558160 80593
rect 557840 80273 557882 80509
rect 558118 80273 558160 80509
rect 557840 80241 558160 80273
rect 563771 80829 564091 80861
rect 563771 80593 563813 80829
rect 564049 80593 564091 80829
rect 563771 80509 564091 80593
rect 563771 80273 563813 80509
rect 564049 80273 564091 80509
rect 563771 80241 564091 80273
rect 573494 80829 574114 107273
rect 573494 80593 573526 80829
rect 573762 80593 573846 80829
rect 574082 80593 574114 80829
rect 573494 80509 574114 80593
rect 573494 80273 573526 80509
rect 573762 80273 573846 80509
rect 574082 80273 574114 80509
rect 22874 77454 23194 77486
rect 22874 77218 22916 77454
rect 23152 77218 23194 77454
rect 22874 77134 23194 77218
rect 22874 76898 22916 77134
rect 23152 76898 23194 77134
rect 22874 76866 23194 76898
rect 28805 77454 29125 77486
rect 28805 77218 28847 77454
rect 29083 77218 29125 77454
rect 28805 77134 29125 77218
rect 28805 76898 28847 77134
rect 29083 76898 29125 77134
rect 28805 76866 29125 76898
rect 50874 77454 51194 77486
rect 50874 77218 50916 77454
rect 51152 77218 51194 77454
rect 50874 77134 51194 77218
rect 50874 76898 50916 77134
rect 51152 76898 51194 77134
rect 50874 76866 51194 76898
rect 56805 77454 57125 77486
rect 56805 77218 56847 77454
rect 57083 77218 57125 77454
rect 56805 77134 57125 77218
rect 56805 76898 56847 77134
rect 57083 76898 57125 77134
rect 56805 76866 57125 76898
rect 78874 77454 79194 77486
rect 78874 77218 78916 77454
rect 79152 77218 79194 77454
rect 78874 77134 79194 77218
rect 78874 76898 78916 77134
rect 79152 76898 79194 77134
rect 78874 76866 79194 76898
rect 84805 77454 85125 77486
rect 84805 77218 84847 77454
rect 85083 77218 85125 77454
rect 84805 77134 85125 77218
rect 84805 76898 84847 77134
rect 85083 76898 85125 77134
rect 84805 76866 85125 76898
rect 106874 77454 107194 77486
rect 106874 77218 106916 77454
rect 107152 77218 107194 77454
rect 106874 77134 107194 77218
rect 106874 76898 106916 77134
rect 107152 76898 107194 77134
rect 106874 76866 107194 76898
rect 112805 77454 113125 77486
rect 112805 77218 112847 77454
rect 113083 77218 113125 77454
rect 112805 77134 113125 77218
rect 112805 76898 112847 77134
rect 113083 76898 113125 77134
rect 112805 76866 113125 76898
rect 134874 77454 135194 77486
rect 134874 77218 134916 77454
rect 135152 77218 135194 77454
rect 134874 77134 135194 77218
rect 134874 76898 134916 77134
rect 135152 76898 135194 77134
rect 134874 76866 135194 76898
rect 140805 77454 141125 77486
rect 140805 77218 140847 77454
rect 141083 77218 141125 77454
rect 140805 77134 141125 77218
rect 140805 76898 140847 77134
rect 141083 76898 141125 77134
rect 140805 76866 141125 76898
rect 162874 77454 163194 77486
rect 162874 77218 162916 77454
rect 163152 77218 163194 77454
rect 162874 77134 163194 77218
rect 162874 76898 162916 77134
rect 163152 76898 163194 77134
rect 162874 76866 163194 76898
rect 168805 77454 169125 77486
rect 168805 77218 168847 77454
rect 169083 77218 169125 77454
rect 168805 77134 169125 77218
rect 168805 76898 168847 77134
rect 169083 76898 169125 77134
rect 168805 76866 169125 76898
rect 190874 77454 191194 77486
rect 190874 77218 190916 77454
rect 191152 77218 191194 77454
rect 190874 77134 191194 77218
rect 190874 76898 190916 77134
rect 191152 76898 191194 77134
rect 190874 76866 191194 76898
rect 196805 77454 197125 77486
rect 196805 77218 196847 77454
rect 197083 77218 197125 77454
rect 196805 77134 197125 77218
rect 196805 76898 196847 77134
rect 197083 76898 197125 77134
rect 196805 76866 197125 76898
rect 218874 77454 219194 77486
rect 218874 77218 218916 77454
rect 219152 77218 219194 77454
rect 218874 77134 219194 77218
rect 218874 76898 218916 77134
rect 219152 76898 219194 77134
rect 218874 76866 219194 76898
rect 224805 77454 225125 77486
rect 224805 77218 224847 77454
rect 225083 77218 225125 77454
rect 224805 77134 225125 77218
rect 224805 76898 224847 77134
rect 225083 76898 225125 77134
rect 224805 76866 225125 76898
rect 246874 77454 247194 77486
rect 246874 77218 246916 77454
rect 247152 77218 247194 77454
rect 246874 77134 247194 77218
rect 246874 76898 246916 77134
rect 247152 76898 247194 77134
rect 246874 76866 247194 76898
rect 252805 77454 253125 77486
rect 252805 77218 252847 77454
rect 253083 77218 253125 77454
rect 252805 77134 253125 77218
rect 252805 76898 252847 77134
rect 253083 76898 253125 77134
rect 252805 76866 253125 76898
rect 274874 77454 275194 77486
rect 274874 77218 274916 77454
rect 275152 77218 275194 77454
rect 274874 77134 275194 77218
rect 274874 76898 274916 77134
rect 275152 76898 275194 77134
rect 274874 76866 275194 76898
rect 280805 77454 281125 77486
rect 280805 77218 280847 77454
rect 281083 77218 281125 77454
rect 280805 77134 281125 77218
rect 280805 76898 280847 77134
rect 281083 76898 281125 77134
rect 280805 76866 281125 76898
rect 302874 77454 303194 77486
rect 302874 77218 302916 77454
rect 303152 77218 303194 77454
rect 302874 77134 303194 77218
rect 302874 76898 302916 77134
rect 303152 76898 303194 77134
rect 302874 76866 303194 76898
rect 308805 77454 309125 77486
rect 308805 77218 308847 77454
rect 309083 77218 309125 77454
rect 308805 77134 309125 77218
rect 308805 76898 308847 77134
rect 309083 76898 309125 77134
rect 308805 76866 309125 76898
rect 330874 77454 331194 77486
rect 330874 77218 330916 77454
rect 331152 77218 331194 77454
rect 330874 77134 331194 77218
rect 330874 76898 330916 77134
rect 331152 76898 331194 77134
rect 330874 76866 331194 76898
rect 336805 77454 337125 77486
rect 336805 77218 336847 77454
rect 337083 77218 337125 77454
rect 336805 77134 337125 77218
rect 336805 76898 336847 77134
rect 337083 76898 337125 77134
rect 336805 76866 337125 76898
rect 358874 77454 359194 77486
rect 358874 77218 358916 77454
rect 359152 77218 359194 77454
rect 358874 77134 359194 77218
rect 358874 76898 358916 77134
rect 359152 76898 359194 77134
rect 358874 76866 359194 76898
rect 364805 77454 365125 77486
rect 364805 77218 364847 77454
rect 365083 77218 365125 77454
rect 364805 77134 365125 77218
rect 364805 76898 364847 77134
rect 365083 76898 365125 77134
rect 364805 76866 365125 76898
rect 386874 77454 387194 77486
rect 386874 77218 386916 77454
rect 387152 77218 387194 77454
rect 386874 77134 387194 77218
rect 386874 76898 386916 77134
rect 387152 76898 387194 77134
rect 386874 76866 387194 76898
rect 392805 77454 393125 77486
rect 392805 77218 392847 77454
rect 393083 77218 393125 77454
rect 392805 77134 393125 77218
rect 392805 76898 392847 77134
rect 393083 76898 393125 77134
rect 392805 76866 393125 76898
rect 414874 77454 415194 77486
rect 414874 77218 414916 77454
rect 415152 77218 415194 77454
rect 414874 77134 415194 77218
rect 414874 76898 414916 77134
rect 415152 76898 415194 77134
rect 414874 76866 415194 76898
rect 420805 77454 421125 77486
rect 420805 77218 420847 77454
rect 421083 77218 421125 77454
rect 420805 77134 421125 77218
rect 420805 76898 420847 77134
rect 421083 76898 421125 77134
rect 420805 76866 421125 76898
rect 442874 77454 443194 77486
rect 442874 77218 442916 77454
rect 443152 77218 443194 77454
rect 442874 77134 443194 77218
rect 442874 76898 442916 77134
rect 443152 76898 443194 77134
rect 442874 76866 443194 76898
rect 448805 77454 449125 77486
rect 448805 77218 448847 77454
rect 449083 77218 449125 77454
rect 448805 77134 449125 77218
rect 448805 76898 448847 77134
rect 449083 76898 449125 77134
rect 448805 76866 449125 76898
rect 470874 77454 471194 77486
rect 470874 77218 470916 77454
rect 471152 77218 471194 77454
rect 470874 77134 471194 77218
rect 470874 76898 470916 77134
rect 471152 76898 471194 77134
rect 470874 76866 471194 76898
rect 476805 77454 477125 77486
rect 476805 77218 476847 77454
rect 477083 77218 477125 77454
rect 476805 77134 477125 77218
rect 476805 76898 476847 77134
rect 477083 76898 477125 77134
rect 476805 76866 477125 76898
rect 498874 77454 499194 77486
rect 498874 77218 498916 77454
rect 499152 77218 499194 77454
rect 498874 77134 499194 77218
rect 498874 76898 498916 77134
rect 499152 76898 499194 77134
rect 498874 76866 499194 76898
rect 504805 77454 505125 77486
rect 504805 77218 504847 77454
rect 505083 77218 505125 77454
rect 504805 77134 505125 77218
rect 504805 76898 504847 77134
rect 505083 76898 505125 77134
rect 504805 76866 505125 76898
rect 526874 77454 527194 77486
rect 526874 77218 526916 77454
rect 527152 77218 527194 77454
rect 526874 77134 527194 77218
rect 526874 76898 526916 77134
rect 527152 76898 527194 77134
rect 526874 76866 527194 76898
rect 532805 77454 533125 77486
rect 532805 77218 532847 77454
rect 533083 77218 533125 77454
rect 532805 77134 533125 77218
rect 532805 76898 532847 77134
rect 533083 76898 533125 77134
rect 532805 76866 533125 76898
rect 554874 77454 555194 77486
rect 554874 77218 554916 77454
rect 555152 77218 555194 77454
rect 554874 77134 555194 77218
rect 554874 76898 554916 77134
rect 555152 76898 555194 77134
rect 554874 76866 555194 76898
rect 560805 77454 561125 77486
rect 560805 77218 560847 77454
rect 561083 77218 561125 77454
rect 560805 77134 561125 77218
rect 560805 76898 560847 77134
rect 561083 76898 561125 77134
rect 560805 76866 561125 76898
rect -2006 53593 -1974 53829
rect -1738 53593 -1654 53829
rect -1418 53593 -1386 53829
rect -2006 53509 -1386 53593
rect -2006 53273 -1974 53509
rect -1738 53273 -1654 53509
rect -1418 53273 -1386 53509
rect -2006 26829 -1386 53273
rect 19909 53829 20229 53861
rect 19909 53593 19951 53829
rect 20187 53593 20229 53829
rect 19909 53509 20229 53593
rect 19909 53273 19951 53509
rect 20187 53273 20229 53509
rect 19909 53241 20229 53273
rect 25840 53829 26160 53861
rect 25840 53593 25882 53829
rect 26118 53593 26160 53829
rect 25840 53509 26160 53593
rect 25840 53273 25882 53509
rect 26118 53273 26160 53509
rect 25840 53241 26160 53273
rect 31770 53829 32090 53861
rect 31770 53593 31812 53829
rect 32048 53593 32090 53829
rect 31770 53509 32090 53593
rect 31770 53273 31812 53509
rect 32048 53273 32090 53509
rect 31770 53241 32090 53273
rect 47909 53829 48229 53861
rect 47909 53593 47951 53829
rect 48187 53593 48229 53829
rect 47909 53509 48229 53593
rect 47909 53273 47951 53509
rect 48187 53273 48229 53509
rect 47909 53241 48229 53273
rect 53840 53829 54160 53861
rect 53840 53593 53882 53829
rect 54118 53593 54160 53829
rect 53840 53509 54160 53593
rect 53840 53273 53882 53509
rect 54118 53273 54160 53509
rect 53840 53241 54160 53273
rect 59770 53829 60090 53861
rect 59770 53593 59812 53829
rect 60048 53593 60090 53829
rect 59770 53509 60090 53593
rect 59770 53273 59812 53509
rect 60048 53273 60090 53509
rect 59770 53241 60090 53273
rect 75909 53829 76229 53861
rect 75909 53593 75951 53829
rect 76187 53593 76229 53829
rect 75909 53509 76229 53593
rect 75909 53273 75951 53509
rect 76187 53273 76229 53509
rect 75909 53241 76229 53273
rect 81840 53829 82160 53861
rect 81840 53593 81882 53829
rect 82118 53593 82160 53829
rect 81840 53509 82160 53593
rect 81840 53273 81882 53509
rect 82118 53273 82160 53509
rect 81840 53241 82160 53273
rect 87770 53829 88090 53861
rect 87770 53593 87812 53829
rect 88048 53593 88090 53829
rect 87770 53509 88090 53593
rect 87770 53273 87812 53509
rect 88048 53273 88090 53509
rect 87770 53241 88090 53273
rect 103909 53829 104229 53861
rect 103909 53593 103951 53829
rect 104187 53593 104229 53829
rect 103909 53509 104229 53593
rect 103909 53273 103951 53509
rect 104187 53273 104229 53509
rect 103909 53241 104229 53273
rect 109840 53829 110160 53861
rect 109840 53593 109882 53829
rect 110118 53593 110160 53829
rect 109840 53509 110160 53593
rect 109840 53273 109882 53509
rect 110118 53273 110160 53509
rect 109840 53241 110160 53273
rect 115770 53829 116090 53861
rect 115770 53593 115812 53829
rect 116048 53593 116090 53829
rect 115770 53509 116090 53593
rect 115770 53273 115812 53509
rect 116048 53273 116090 53509
rect 115770 53241 116090 53273
rect 131909 53829 132229 53861
rect 131909 53593 131951 53829
rect 132187 53593 132229 53829
rect 131909 53509 132229 53593
rect 131909 53273 131951 53509
rect 132187 53273 132229 53509
rect 131909 53241 132229 53273
rect 137840 53829 138160 53861
rect 137840 53593 137882 53829
rect 138118 53593 138160 53829
rect 137840 53509 138160 53593
rect 137840 53273 137882 53509
rect 138118 53273 138160 53509
rect 137840 53241 138160 53273
rect 143770 53829 144090 53861
rect 143770 53593 143812 53829
rect 144048 53593 144090 53829
rect 143770 53509 144090 53593
rect 143770 53273 143812 53509
rect 144048 53273 144090 53509
rect 143770 53241 144090 53273
rect 159909 53829 160229 53861
rect 159909 53593 159951 53829
rect 160187 53593 160229 53829
rect 159909 53509 160229 53593
rect 159909 53273 159951 53509
rect 160187 53273 160229 53509
rect 159909 53241 160229 53273
rect 165840 53829 166160 53861
rect 165840 53593 165882 53829
rect 166118 53593 166160 53829
rect 165840 53509 166160 53593
rect 165840 53273 165882 53509
rect 166118 53273 166160 53509
rect 165840 53241 166160 53273
rect 171770 53829 172090 53861
rect 171770 53593 171812 53829
rect 172048 53593 172090 53829
rect 171770 53509 172090 53593
rect 171770 53273 171812 53509
rect 172048 53273 172090 53509
rect 171770 53241 172090 53273
rect 187909 53829 188229 53861
rect 187909 53593 187951 53829
rect 188187 53593 188229 53829
rect 187909 53509 188229 53593
rect 187909 53273 187951 53509
rect 188187 53273 188229 53509
rect 187909 53241 188229 53273
rect 193840 53829 194160 53861
rect 193840 53593 193882 53829
rect 194118 53593 194160 53829
rect 193840 53509 194160 53593
rect 193840 53273 193882 53509
rect 194118 53273 194160 53509
rect 193840 53241 194160 53273
rect 199770 53829 200090 53861
rect 199770 53593 199812 53829
rect 200048 53593 200090 53829
rect 199770 53509 200090 53593
rect 199770 53273 199812 53509
rect 200048 53273 200090 53509
rect 199770 53241 200090 53273
rect 215909 53829 216229 53861
rect 215909 53593 215951 53829
rect 216187 53593 216229 53829
rect 215909 53509 216229 53593
rect 215909 53273 215951 53509
rect 216187 53273 216229 53509
rect 215909 53241 216229 53273
rect 221840 53829 222160 53861
rect 221840 53593 221882 53829
rect 222118 53593 222160 53829
rect 221840 53509 222160 53593
rect 221840 53273 221882 53509
rect 222118 53273 222160 53509
rect 221840 53241 222160 53273
rect 227770 53829 228090 53861
rect 227770 53593 227812 53829
rect 228048 53593 228090 53829
rect 227770 53509 228090 53593
rect 227770 53273 227812 53509
rect 228048 53273 228090 53509
rect 227770 53241 228090 53273
rect 243909 53829 244229 53861
rect 243909 53593 243951 53829
rect 244187 53593 244229 53829
rect 243909 53509 244229 53593
rect 243909 53273 243951 53509
rect 244187 53273 244229 53509
rect 243909 53241 244229 53273
rect 249840 53829 250160 53861
rect 249840 53593 249882 53829
rect 250118 53593 250160 53829
rect 249840 53509 250160 53593
rect 249840 53273 249882 53509
rect 250118 53273 250160 53509
rect 249840 53241 250160 53273
rect 255770 53829 256090 53861
rect 255770 53593 255812 53829
rect 256048 53593 256090 53829
rect 255770 53509 256090 53593
rect 255770 53273 255812 53509
rect 256048 53273 256090 53509
rect 255770 53241 256090 53273
rect 271909 53829 272229 53861
rect 271909 53593 271951 53829
rect 272187 53593 272229 53829
rect 271909 53509 272229 53593
rect 271909 53273 271951 53509
rect 272187 53273 272229 53509
rect 271909 53241 272229 53273
rect 277840 53829 278160 53861
rect 277840 53593 277882 53829
rect 278118 53593 278160 53829
rect 277840 53509 278160 53593
rect 277840 53273 277882 53509
rect 278118 53273 278160 53509
rect 277840 53241 278160 53273
rect 283770 53829 284090 53861
rect 283770 53593 283812 53829
rect 284048 53593 284090 53829
rect 283770 53509 284090 53593
rect 283770 53273 283812 53509
rect 284048 53273 284090 53509
rect 283770 53241 284090 53273
rect 299909 53829 300229 53861
rect 299909 53593 299951 53829
rect 300187 53593 300229 53829
rect 299909 53509 300229 53593
rect 299909 53273 299951 53509
rect 300187 53273 300229 53509
rect 299909 53241 300229 53273
rect 305840 53829 306160 53861
rect 305840 53593 305882 53829
rect 306118 53593 306160 53829
rect 305840 53509 306160 53593
rect 305840 53273 305882 53509
rect 306118 53273 306160 53509
rect 305840 53241 306160 53273
rect 311770 53829 312090 53861
rect 311770 53593 311812 53829
rect 312048 53593 312090 53829
rect 311770 53509 312090 53593
rect 311770 53273 311812 53509
rect 312048 53273 312090 53509
rect 311770 53241 312090 53273
rect 327909 53829 328229 53861
rect 327909 53593 327951 53829
rect 328187 53593 328229 53829
rect 327909 53509 328229 53593
rect 327909 53273 327951 53509
rect 328187 53273 328229 53509
rect 327909 53241 328229 53273
rect 333840 53829 334160 53861
rect 333840 53593 333882 53829
rect 334118 53593 334160 53829
rect 333840 53509 334160 53593
rect 333840 53273 333882 53509
rect 334118 53273 334160 53509
rect 333840 53241 334160 53273
rect 339770 53829 340090 53861
rect 339770 53593 339812 53829
rect 340048 53593 340090 53829
rect 339770 53509 340090 53593
rect 339770 53273 339812 53509
rect 340048 53273 340090 53509
rect 339770 53241 340090 53273
rect 355909 53829 356229 53861
rect 355909 53593 355951 53829
rect 356187 53593 356229 53829
rect 355909 53509 356229 53593
rect 355909 53273 355951 53509
rect 356187 53273 356229 53509
rect 355909 53241 356229 53273
rect 361840 53829 362160 53861
rect 361840 53593 361882 53829
rect 362118 53593 362160 53829
rect 361840 53509 362160 53593
rect 361840 53273 361882 53509
rect 362118 53273 362160 53509
rect 361840 53241 362160 53273
rect 367770 53829 368090 53861
rect 367770 53593 367812 53829
rect 368048 53593 368090 53829
rect 367770 53509 368090 53593
rect 367770 53273 367812 53509
rect 368048 53273 368090 53509
rect 367770 53241 368090 53273
rect 383909 53829 384229 53861
rect 383909 53593 383951 53829
rect 384187 53593 384229 53829
rect 383909 53509 384229 53593
rect 383909 53273 383951 53509
rect 384187 53273 384229 53509
rect 383909 53241 384229 53273
rect 389840 53829 390160 53861
rect 389840 53593 389882 53829
rect 390118 53593 390160 53829
rect 389840 53509 390160 53593
rect 389840 53273 389882 53509
rect 390118 53273 390160 53509
rect 389840 53241 390160 53273
rect 395770 53829 396090 53861
rect 395770 53593 395812 53829
rect 396048 53593 396090 53829
rect 395770 53509 396090 53593
rect 395770 53273 395812 53509
rect 396048 53273 396090 53509
rect 395770 53241 396090 53273
rect 411909 53829 412229 53861
rect 411909 53593 411951 53829
rect 412187 53593 412229 53829
rect 411909 53509 412229 53593
rect 411909 53273 411951 53509
rect 412187 53273 412229 53509
rect 411909 53241 412229 53273
rect 417840 53829 418160 53861
rect 417840 53593 417882 53829
rect 418118 53593 418160 53829
rect 417840 53509 418160 53593
rect 417840 53273 417882 53509
rect 418118 53273 418160 53509
rect 417840 53241 418160 53273
rect 423770 53829 424090 53861
rect 423770 53593 423812 53829
rect 424048 53593 424090 53829
rect 423770 53509 424090 53593
rect 423770 53273 423812 53509
rect 424048 53273 424090 53509
rect 423770 53241 424090 53273
rect 439909 53829 440229 53861
rect 439909 53593 439951 53829
rect 440187 53593 440229 53829
rect 439909 53509 440229 53593
rect 439909 53273 439951 53509
rect 440187 53273 440229 53509
rect 439909 53241 440229 53273
rect 445840 53829 446160 53861
rect 445840 53593 445882 53829
rect 446118 53593 446160 53829
rect 445840 53509 446160 53593
rect 445840 53273 445882 53509
rect 446118 53273 446160 53509
rect 445840 53241 446160 53273
rect 451770 53829 452090 53861
rect 451770 53593 451812 53829
rect 452048 53593 452090 53829
rect 451770 53509 452090 53593
rect 451770 53273 451812 53509
rect 452048 53273 452090 53509
rect 451770 53241 452090 53273
rect 467909 53829 468229 53861
rect 467909 53593 467951 53829
rect 468187 53593 468229 53829
rect 467909 53509 468229 53593
rect 467909 53273 467951 53509
rect 468187 53273 468229 53509
rect 467909 53241 468229 53273
rect 473840 53829 474160 53861
rect 473840 53593 473882 53829
rect 474118 53593 474160 53829
rect 473840 53509 474160 53593
rect 473840 53273 473882 53509
rect 474118 53273 474160 53509
rect 473840 53241 474160 53273
rect 479770 53829 480090 53861
rect 479770 53593 479812 53829
rect 480048 53593 480090 53829
rect 479770 53509 480090 53593
rect 479770 53273 479812 53509
rect 480048 53273 480090 53509
rect 479770 53241 480090 53273
rect 495909 53829 496229 53861
rect 495909 53593 495951 53829
rect 496187 53593 496229 53829
rect 495909 53509 496229 53593
rect 495909 53273 495951 53509
rect 496187 53273 496229 53509
rect 495909 53241 496229 53273
rect 501840 53829 502160 53861
rect 501840 53593 501882 53829
rect 502118 53593 502160 53829
rect 501840 53509 502160 53593
rect 501840 53273 501882 53509
rect 502118 53273 502160 53509
rect 501840 53241 502160 53273
rect 507770 53829 508090 53861
rect 507770 53593 507812 53829
rect 508048 53593 508090 53829
rect 507770 53509 508090 53593
rect 507770 53273 507812 53509
rect 508048 53273 508090 53509
rect 507770 53241 508090 53273
rect 523909 53829 524229 53861
rect 523909 53593 523951 53829
rect 524187 53593 524229 53829
rect 523909 53509 524229 53593
rect 523909 53273 523951 53509
rect 524187 53273 524229 53509
rect 523909 53241 524229 53273
rect 529840 53829 530160 53861
rect 529840 53593 529882 53829
rect 530118 53593 530160 53829
rect 529840 53509 530160 53593
rect 529840 53273 529882 53509
rect 530118 53273 530160 53509
rect 529840 53241 530160 53273
rect 535770 53829 536090 53861
rect 535770 53593 535812 53829
rect 536048 53593 536090 53829
rect 535770 53509 536090 53593
rect 535770 53273 535812 53509
rect 536048 53273 536090 53509
rect 535770 53241 536090 53273
rect 551909 53829 552229 53861
rect 551909 53593 551951 53829
rect 552187 53593 552229 53829
rect 551909 53509 552229 53593
rect 551909 53273 551951 53509
rect 552187 53273 552229 53509
rect 551909 53241 552229 53273
rect 557840 53829 558160 53861
rect 557840 53593 557882 53829
rect 558118 53593 558160 53829
rect 557840 53509 558160 53593
rect 557840 53273 557882 53509
rect 558118 53273 558160 53509
rect 557840 53241 558160 53273
rect 563770 53829 564090 53861
rect 563770 53593 563812 53829
rect 564048 53593 564090 53829
rect 563770 53509 564090 53593
rect 563770 53273 563812 53509
rect 564048 53273 564090 53509
rect 563770 53241 564090 53273
rect 573494 53829 574114 80273
rect 573494 53593 573526 53829
rect 573762 53593 573846 53829
rect 574082 53593 574114 53829
rect 573494 53509 574114 53593
rect 573494 53273 573526 53509
rect 573762 53273 573846 53509
rect 574082 53273 574114 53509
rect 22875 50454 23195 50486
rect 22875 50218 22917 50454
rect 23153 50218 23195 50454
rect 22875 50134 23195 50218
rect 22875 49898 22917 50134
rect 23153 49898 23195 50134
rect 22875 49866 23195 49898
rect 28806 50454 29126 50486
rect 28806 50218 28848 50454
rect 29084 50218 29126 50454
rect 28806 50134 29126 50218
rect 28806 49898 28848 50134
rect 29084 49898 29126 50134
rect 28806 49866 29126 49898
rect 50875 50454 51195 50486
rect 50875 50218 50917 50454
rect 51153 50218 51195 50454
rect 50875 50134 51195 50218
rect 50875 49898 50917 50134
rect 51153 49898 51195 50134
rect 50875 49866 51195 49898
rect 56806 50454 57126 50486
rect 56806 50218 56848 50454
rect 57084 50218 57126 50454
rect 56806 50134 57126 50218
rect 56806 49898 56848 50134
rect 57084 49898 57126 50134
rect 56806 49866 57126 49898
rect 78875 50454 79195 50486
rect 78875 50218 78917 50454
rect 79153 50218 79195 50454
rect 78875 50134 79195 50218
rect 78875 49898 78917 50134
rect 79153 49898 79195 50134
rect 78875 49866 79195 49898
rect 84806 50454 85126 50486
rect 84806 50218 84848 50454
rect 85084 50218 85126 50454
rect 84806 50134 85126 50218
rect 84806 49898 84848 50134
rect 85084 49898 85126 50134
rect 84806 49866 85126 49898
rect 106875 50454 107195 50486
rect 106875 50218 106917 50454
rect 107153 50218 107195 50454
rect 106875 50134 107195 50218
rect 106875 49898 106917 50134
rect 107153 49898 107195 50134
rect 106875 49866 107195 49898
rect 112806 50454 113126 50486
rect 112806 50218 112848 50454
rect 113084 50218 113126 50454
rect 112806 50134 113126 50218
rect 112806 49898 112848 50134
rect 113084 49898 113126 50134
rect 112806 49866 113126 49898
rect 134875 50454 135195 50486
rect 134875 50218 134917 50454
rect 135153 50218 135195 50454
rect 134875 50134 135195 50218
rect 134875 49898 134917 50134
rect 135153 49898 135195 50134
rect 134875 49866 135195 49898
rect 140806 50454 141126 50486
rect 140806 50218 140848 50454
rect 141084 50218 141126 50454
rect 140806 50134 141126 50218
rect 140806 49898 140848 50134
rect 141084 49898 141126 50134
rect 140806 49866 141126 49898
rect 162875 50454 163195 50486
rect 162875 50218 162917 50454
rect 163153 50218 163195 50454
rect 162875 50134 163195 50218
rect 162875 49898 162917 50134
rect 163153 49898 163195 50134
rect 162875 49866 163195 49898
rect 168806 50454 169126 50486
rect 168806 50218 168848 50454
rect 169084 50218 169126 50454
rect 168806 50134 169126 50218
rect 168806 49898 168848 50134
rect 169084 49898 169126 50134
rect 168806 49866 169126 49898
rect 190875 50454 191195 50486
rect 190875 50218 190917 50454
rect 191153 50218 191195 50454
rect 190875 50134 191195 50218
rect 190875 49898 190917 50134
rect 191153 49898 191195 50134
rect 190875 49866 191195 49898
rect 196806 50454 197126 50486
rect 196806 50218 196848 50454
rect 197084 50218 197126 50454
rect 196806 50134 197126 50218
rect 196806 49898 196848 50134
rect 197084 49898 197126 50134
rect 196806 49866 197126 49898
rect 218875 50454 219195 50486
rect 218875 50218 218917 50454
rect 219153 50218 219195 50454
rect 218875 50134 219195 50218
rect 218875 49898 218917 50134
rect 219153 49898 219195 50134
rect 218875 49866 219195 49898
rect 224806 50454 225126 50486
rect 224806 50218 224848 50454
rect 225084 50218 225126 50454
rect 224806 50134 225126 50218
rect 224806 49898 224848 50134
rect 225084 49898 225126 50134
rect 224806 49866 225126 49898
rect 246875 50454 247195 50486
rect 246875 50218 246917 50454
rect 247153 50218 247195 50454
rect 246875 50134 247195 50218
rect 246875 49898 246917 50134
rect 247153 49898 247195 50134
rect 246875 49866 247195 49898
rect 252806 50454 253126 50486
rect 252806 50218 252848 50454
rect 253084 50218 253126 50454
rect 252806 50134 253126 50218
rect 252806 49898 252848 50134
rect 253084 49898 253126 50134
rect 252806 49866 253126 49898
rect 274875 50454 275195 50486
rect 274875 50218 274917 50454
rect 275153 50218 275195 50454
rect 274875 50134 275195 50218
rect 274875 49898 274917 50134
rect 275153 49898 275195 50134
rect 274875 49866 275195 49898
rect 280806 50454 281126 50486
rect 280806 50218 280848 50454
rect 281084 50218 281126 50454
rect 280806 50134 281126 50218
rect 280806 49898 280848 50134
rect 281084 49898 281126 50134
rect 280806 49866 281126 49898
rect 302875 50454 303195 50486
rect 302875 50218 302917 50454
rect 303153 50218 303195 50454
rect 302875 50134 303195 50218
rect 302875 49898 302917 50134
rect 303153 49898 303195 50134
rect 302875 49866 303195 49898
rect 308806 50454 309126 50486
rect 308806 50218 308848 50454
rect 309084 50218 309126 50454
rect 308806 50134 309126 50218
rect 308806 49898 308848 50134
rect 309084 49898 309126 50134
rect 308806 49866 309126 49898
rect 330875 50454 331195 50486
rect 330875 50218 330917 50454
rect 331153 50218 331195 50454
rect 330875 50134 331195 50218
rect 330875 49898 330917 50134
rect 331153 49898 331195 50134
rect 330875 49866 331195 49898
rect 336806 50454 337126 50486
rect 336806 50218 336848 50454
rect 337084 50218 337126 50454
rect 336806 50134 337126 50218
rect 336806 49898 336848 50134
rect 337084 49898 337126 50134
rect 336806 49866 337126 49898
rect 358875 50454 359195 50486
rect 358875 50218 358917 50454
rect 359153 50218 359195 50454
rect 358875 50134 359195 50218
rect 358875 49898 358917 50134
rect 359153 49898 359195 50134
rect 358875 49866 359195 49898
rect 364806 50454 365126 50486
rect 364806 50218 364848 50454
rect 365084 50218 365126 50454
rect 364806 50134 365126 50218
rect 364806 49898 364848 50134
rect 365084 49898 365126 50134
rect 364806 49866 365126 49898
rect 386875 50454 387195 50486
rect 386875 50218 386917 50454
rect 387153 50218 387195 50454
rect 386875 50134 387195 50218
rect 386875 49898 386917 50134
rect 387153 49898 387195 50134
rect 386875 49866 387195 49898
rect 392806 50454 393126 50486
rect 392806 50218 392848 50454
rect 393084 50218 393126 50454
rect 392806 50134 393126 50218
rect 392806 49898 392848 50134
rect 393084 49898 393126 50134
rect 392806 49866 393126 49898
rect 414875 50454 415195 50486
rect 414875 50218 414917 50454
rect 415153 50218 415195 50454
rect 414875 50134 415195 50218
rect 414875 49898 414917 50134
rect 415153 49898 415195 50134
rect 414875 49866 415195 49898
rect 420806 50454 421126 50486
rect 420806 50218 420848 50454
rect 421084 50218 421126 50454
rect 420806 50134 421126 50218
rect 420806 49898 420848 50134
rect 421084 49898 421126 50134
rect 420806 49866 421126 49898
rect 442875 50454 443195 50486
rect 442875 50218 442917 50454
rect 443153 50218 443195 50454
rect 442875 50134 443195 50218
rect 442875 49898 442917 50134
rect 443153 49898 443195 50134
rect 442875 49866 443195 49898
rect 448806 50454 449126 50486
rect 448806 50218 448848 50454
rect 449084 50218 449126 50454
rect 448806 50134 449126 50218
rect 448806 49898 448848 50134
rect 449084 49898 449126 50134
rect 448806 49866 449126 49898
rect 470875 50454 471195 50486
rect 470875 50218 470917 50454
rect 471153 50218 471195 50454
rect 470875 50134 471195 50218
rect 470875 49898 470917 50134
rect 471153 49898 471195 50134
rect 470875 49866 471195 49898
rect 476806 50454 477126 50486
rect 476806 50218 476848 50454
rect 477084 50218 477126 50454
rect 476806 50134 477126 50218
rect 476806 49898 476848 50134
rect 477084 49898 477126 50134
rect 476806 49866 477126 49898
rect 498875 50454 499195 50486
rect 498875 50218 498917 50454
rect 499153 50218 499195 50454
rect 498875 50134 499195 50218
rect 498875 49898 498917 50134
rect 499153 49898 499195 50134
rect 498875 49866 499195 49898
rect 504806 50454 505126 50486
rect 504806 50218 504848 50454
rect 505084 50218 505126 50454
rect 504806 50134 505126 50218
rect 504806 49898 504848 50134
rect 505084 49898 505126 50134
rect 504806 49866 505126 49898
rect 526875 50454 527195 50486
rect 526875 50218 526917 50454
rect 527153 50218 527195 50454
rect 526875 50134 527195 50218
rect 526875 49898 526917 50134
rect 527153 49898 527195 50134
rect 526875 49866 527195 49898
rect 532806 50454 533126 50486
rect 532806 50218 532848 50454
rect 533084 50218 533126 50454
rect 532806 50134 533126 50218
rect 532806 49898 532848 50134
rect 533084 49898 533126 50134
rect 532806 49866 533126 49898
rect 554875 50454 555195 50486
rect 554875 50218 554917 50454
rect 555153 50218 555195 50454
rect 554875 50134 555195 50218
rect 554875 49898 554917 50134
rect 555153 49898 555195 50134
rect 554875 49866 555195 49898
rect 560806 50454 561126 50486
rect 560806 50218 560848 50454
rect 561084 50218 561126 50454
rect 560806 50134 561126 50218
rect 560806 49898 560848 50134
rect 561084 49898 561126 50134
rect 560806 49866 561126 49898
rect 48083 42124 48149 42125
rect 48083 42060 48084 42124
rect 48148 42060 48149 42124
rect 48083 42059 48149 42060
rect 42747 35324 42813 35325
rect 42747 35260 42748 35324
rect 42812 35260 42813 35324
rect 42747 35259 42813 35260
rect -2006 26593 -1974 26829
rect -1738 26593 -1654 26829
rect -1418 26593 -1386 26829
rect -2006 26509 -1386 26593
rect -2006 26273 -1974 26509
rect -1738 26273 -1654 26509
rect -1418 26273 -1386 26509
rect -2006 -346 -1386 26273
rect 22418 26829 22738 26861
rect 22418 26593 22460 26829
rect 22696 26593 22738 26829
rect 22418 26509 22738 26593
rect 22418 26273 22460 26509
rect 22696 26273 22738 26509
rect 22418 26241 22738 26273
rect 33366 26829 33686 26861
rect 33366 26593 33408 26829
rect 33644 26593 33686 26829
rect 33366 26509 33686 26593
rect 33366 26273 33408 26509
rect 33644 26273 33686 26509
rect 33366 26241 33686 26273
rect 27892 23454 28212 23486
rect 27892 23218 27934 23454
rect 28170 23218 28212 23454
rect 27892 23134 28212 23218
rect 27892 22898 27934 23134
rect 28170 22898 28212 23134
rect 27892 22866 28212 22898
rect 38840 23454 39160 23486
rect 38840 23218 38882 23454
rect 39118 23218 39160 23454
rect 38840 23134 39160 23218
rect 38840 22898 38882 23134
rect 39118 22898 39160 23134
rect 38840 22866 39160 22898
rect 42750 5677 42810 35259
rect 44314 26829 44634 26861
rect 44314 26593 44356 26829
rect 44592 26593 44634 26829
rect 44314 26509 44634 26593
rect 44314 26273 44356 26509
rect 44592 26273 44634 26509
rect 44314 26241 44634 26273
rect 48086 16557 48146 42059
rect 55262 26829 55582 26861
rect 55262 26593 55304 26829
rect 55540 26593 55582 26829
rect 55262 26509 55582 26593
rect 55262 26273 55304 26509
rect 55540 26273 55582 26509
rect 55262 26241 55582 26273
rect 49788 23454 50108 23486
rect 49788 23218 49830 23454
rect 50066 23218 50108 23454
rect 49788 23134 50108 23218
rect 49788 22898 49830 23134
rect 50066 22898 50108 23134
rect 49788 22866 50108 22898
rect 60736 23454 61056 23486
rect 60736 23218 60778 23454
rect 61014 23218 61056 23454
rect 60736 23134 61056 23218
rect 60736 22898 60778 23134
rect 61014 22898 61056 23134
rect 60736 22866 61056 22898
rect 65994 23454 66614 41000
rect 75910 26829 76230 26861
rect 75910 26593 75952 26829
rect 76188 26593 76230 26829
rect 75910 26509 76230 26593
rect 75910 26273 75952 26509
rect 76188 26273 76230 26509
rect 75910 26241 76230 26273
rect 81840 26829 82160 26861
rect 81840 26593 81882 26829
rect 82118 26593 82160 26829
rect 81840 26509 82160 26593
rect 81840 26273 81882 26509
rect 82118 26273 82160 26509
rect 81840 26241 82160 26273
rect 87771 26829 88091 26861
rect 87771 26593 87813 26829
rect 88049 26593 88091 26829
rect 87771 26509 88091 26593
rect 87771 26273 87813 26509
rect 88049 26273 88091 26509
rect 87771 26241 88091 26273
rect 103910 26829 104230 26861
rect 103910 26593 103952 26829
rect 104188 26593 104230 26829
rect 103910 26509 104230 26593
rect 103910 26273 103952 26509
rect 104188 26273 104230 26509
rect 103910 26241 104230 26273
rect 109840 26829 110160 26861
rect 109840 26593 109882 26829
rect 110118 26593 110160 26829
rect 109840 26509 110160 26593
rect 109840 26273 109882 26509
rect 110118 26273 110160 26509
rect 109840 26241 110160 26273
rect 115771 26829 116091 26861
rect 115771 26593 115813 26829
rect 116049 26593 116091 26829
rect 115771 26509 116091 26593
rect 115771 26273 115813 26509
rect 116049 26273 116091 26509
rect 115771 26241 116091 26273
rect 131910 26829 132230 26861
rect 131910 26593 131952 26829
rect 132188 26593 132230 26829
rect 131910 26509 132230 26593
rect 131910 26273 131952 26509
rect 132188 26273 132230 26509
rect 131910 26241 132230 26273
rect 137840 26829 138160 26861
rect 137840 26593 137882 26829
rect 138118 26593 138160 26829
rect 137840 26509 138160 26593
rect 137840 26273 137882 26509
rect 138118 26273 138160 26509
rect 137840 26241 138160 26273
rect 143771 26829 144091 26861
rect 143771 26593 143813 26829
rect 144049 26593 144091 26829
rect 143771 26509 144091 26593
rect 143771 26273 143813 26509
rect 144049 26273 144091 26509
rect 143771 26241 144091 26273
rect 159910 26829 160230 26861
rect 159910 26593 159952 26829
rect 160188 26593 160230 26829
rect 159910 26509 160230 26593
rect 159910 26273 159952 26509
rect 160188 26273 160230 26509
rect 159910 26241 160230 26273
rect 165840 26829 166160 26861
rect 165840 26593 165882 26829
rect 166118 26593 166160 26829
rect 165840 26509 166160 26593
rect 165840 26273 165882 26509
rect 166118 26273 166160 26509
rect 165840 26241 166160 26273
rect 171771 26829 172091 26861
rect 171771 26593 171813 26829
rect 172049 26593 172091 26829
rect 171771 26509 172091 26593
rect 171771 26273 171813 26509
rect 172049 26273 172091 26509
rect 171771 26241 172091 26273
rect 187910 26829 188230 26861
rect 187910 26593 187952 26829
rect 188188 26593 188230 26829
rect 187910 26509 188230 26593
rect 187910 26273 187952 26509
rect 188188 26273 188230 26509
rect 187910 26241 188230 26273
rect 193840 26829 194160 26861
rect 193840 26593 193882 26829
rect 194118 26593 194160 26829
rect 193840 26509 194160 26593
rect 193840 26273 193882 26509
rect 194118 26273 194160 26509
rect 193840 26241 194160 26273
rect 199771 26829 200091 26861
rect 199771 26593 199813 26829
rect 200049 26593 200091 26829
rect 199771 26509 200091 26593
rect 199771 26273 199813 26509
rect 200049 26273 200091 26509
rect 199771 26241 200091 26273
rect 215910 26829 216230 26861
rect 215910 26593 215952 26829
rect 216188 26593 216230 26829
rect 215910 26509 216230 26593
rect 215910 26273 215952 26509
rect 216188 26273 216230 26509
rect 215910 26241 216230 26273
rect 221840 26829 222160 26861
rect 221840 26593 221882 26829
rect 222118 26593 222160 26829
rect 221840 26509 222160 26593
rect 221840 26273 221882 26509
rect 222118 26273 222160 26509
rect 221840 26241 222160 26273
rect 227771 26829 228091 26861
rect 227771 26593 227813 26829
rect 228049 26593 228091 26829
rect 227771 26509 228091 26593
rect 227771 26273 227813 26509
rect 228049 26273 228091 26509
rect 227771 26241 228091 26273
rect 243910 26829 244230 26861
rect 243910 26593 243952 26829
rect 244188 26593 244230 26829
rect 243910 26509 244230 26593
rect 243910 26273 243952 26509
rect 244188 26273 244230 26509
rect 243910 26241 244230 26273
rect 249840 26829 250160 26861
rect 249840 26593 249882 26829
rect 250118 26593 250160 26829
rect 249840 26509 250160 26593
rect 249840 26273 249882 26509
rect 250118 26273 250160 26509
rect 249840 26241 250160 26273
rect 255771 26829 256091 26861
rect 255771 26593 255813 26829
rect 256049 26593 256091 26829
rect 255771 26509 256091 26593
rect 255771 26273 255813 26509
rect 256049 26273 256091 26509
rect 255771 26241 256091 26273
rect 271910 26829 272230 26861
rect 271910 26593 271952 26829
rect 272188 26593 272230 26829
rect 271910 26509 272230 26593
rect 271910 26273 271952 26509
rect 272188 26273 272230 26509
rect 271910 26241 272230 26273
rect 277840 26829 278160 26861
rect 277840 26593 277882 26829
rect 278118 26593 278160 26829
rect 277840 26509 278160 26593
rect 277840 26273 277882 26509
rect 278118 26273 278160 26509
rect 277840 26241 278160 26273
rect 283771 26829 284091 26861
rect 283771 26593 283813 26829
rect 284049 26593 284091 26829
rect 283771 26509 284091 26593
rect 283771 26273 283813 26509
rect 284049 26273 284091 26509
rect 283771 26241 284091 26273
rect 299910 26829 300230 26861
rect 299910 26593 299952 26829
rect 300188 26593 300230 26829
rect 299910 26509 300230 26593
rect 299910 26273 299952 26509
rect 300188 26273 300230 26509
rect 299910 26241 300230 26273
rect 305840 26829 306160 26861
rect 305840 26593 305882 26829
rect 306118 26593 306160 26829
rect 305840 26509 306160 26593
rect 305840 26273 305882 26509
rect 306118 26273 306160 26509
rect 305840 26241 306160 26273
rect 311771 26829 312091 26861
rect 311771 26593 311813 26829
rect 312049 26593 312091 26829
rect 311771 26509 312091 26593
rect 311771 26273 311813 26509
rect 312049 26273 312091 26509
rect 311771 26241 312091 26273
rect 327910 26829 328230 26861
rect 327910 26593 327952 26829
rect 328188 26593 328230 26829
rect 327910 26509 328230 26593
rect 327910 26273 327952 26509
rect 328188 26273 328230 26509
rect 327910 26241 328230 26273
rect 333840 26829 334160 26861
rect 333840 26593 333882 26829
rect 334118 26593 334160 26829
rect 333840 26509 334160 26593
rect 333840 26273 333882 26509
rect 334118 26273 334160 26509
rect 333840 26241 334160 26273
rect 339771 26829 340091 26861
rect 339771 26593 339813 26829
rect 340049 26593 340091 26829
rect 339771 26509 340091 26593
rect 339771 26273 339813 26509
rect 340049 26273 340091 26509
rect 339771 26241 340091 26273
rect 355910 26829 356230 26861
rect 355910 26593 355952 26829
rect 356188 26593 356230 26829
rect 355910 26509 356230 26593
rect 355910 26273 355952 26509
rect 356188 26273 356230 26509
rect 355910 26241 356230 26273
rect 361840 26829 362160 26861
rect 361840 26593 361882 26829
rect 362118 26593 362160 26829
rect 361840 26509 362160 26593
rect 361840 26273 361882 26509
rect 362118 26273 362160 26509
rect 361840 26241 362160 26273
rect 367771 26829 368091 26861
rect 367771 26593 367813 26829
rect 368049 26593 368091 26829
rect 367771 26509 368091 26593
rect 367771 26273 367813 26509
rect 368049 26273 368091 26509
rect 367771 26241 368091 26273
rect 383910 26829 384230 26861
rect 383910 26593 383952 26829
rect 384188 26593 384230 26829
rect 383910 26509 384230 26593
rect 383910 26273 383952 26509
rect 384188 26273 384230 26509
rect 383910 26241 384230 26273
rect 389840 26829 390160 26861
rect 389840 26593 389882 26829
rect 390118 26593 390160 26829
rect 389840 26509 390160 26593
rect 389840 26273 389882 26509
rect 390118 26273 390160 26509
rect 389840 26241 390160 26273
rect 395771 26829 396091 26861
rect 395771 26593 395813 26829
rect 396049 26593 396091 26829
rect 395771 26509 396091 26593
rect 395771 26273 395813 26509
rect 396049 26273 396091 26509
rect 395771 26241 396091 26273
rect 411910 26829 412230 26861
rect 411910 26593 411952 26829
rect 412188 26593 412230 26829
rect 411910 26509 412230 26593
rect 411910 26273 411952 26509
rect 412188 26273 412230 26509
rect 411910 26241 412230 26273
rect 417840 26829 418160 26861
rect 417840 26593 417882 26829
rect 418118 26593 418160 26829
rect 417840 26509 418160 26593
rect 417840 26273 417882 26509
rect 418118 26273 418160 26509
rect 417840 26241 418160 26273
rect 423771 26829 424091 26861
rect 423771 26593 423813 26829
rect 424049 26593 424091 26829
rect 423771 26509 424091 26593
rect 423771 26273 423813 26509
rect 424049 26273 424091 26509
rect 423771 26241 424091 26273
rect 439910 26829 440230 26861
rect 439910 26593 439952 26829
rect 440188 26593 440230 26829
rect 439910 26509 440230 26593
rect 439910 26273 439952 26509
rect 440188 26273 440230 26509
rect 439910 26241 440230 26273
rect 445840 26829 446160 26861
rect 445840 26593 445882 26829
rect 446118 26593 446160 26829
rect 445840 26509 446160 26593
rect 445840 26273 445882 26509
rect 446118 26273 446160 26509
rect 445840 26241 446160 26273
rect 451771 26829 452091 26861
rect 451771 26593 451813 26829
rect 452049 26593 452091 26829
rect 451771 26509 452091 26593
rect 451771 26273 451813 26509
rect 452049 26273 452091 26509
rect 451771 26241 452091 26273
rect 467910 26829 468230 26861
rect 467910 26593 467952 26829
rect 468188 26593 468230 26829
rect 467910 26509 468230 26593
rect 467910 26273 467952 26509
rect 468188 26273 468230 26509
rect 467910 26241 468230 26273
rect 473840 26829 474160 26861
rect 473840 26593 473882 26829
rect 474118 26593 474160 26829
rect 473840 26509 474160 26593
rect 473840 26273 473882 26509
rect 474118 26273 474160 26509
rect 473840 26241 474160 26273
rect 479771 26829 480091 26861
rect 479771 26593 479813 26829
rect 480049 26593 480091 26829
rect 479771 26509 480091 26593
rect 479771 26273 479813 26509
rect 480049 26273 480091 26509
rect 479771 26241 480091 26273
rect 495910 26829 496230 26861
rect 495910 26593 495952 26829
rect 496188 26593 496230 26829
rect 495910 26509 496230 26593
rect 495910 26273 495952 26509
rect 496188 26273 496230 26509
rect 495910 26241 496230 26273
rect 501840 26829 502160 26861
rect 501840 26593 501882 26829
rect 502118 26593 502160 26829
rect 501840 26509 502160 26593
rect 501840 26273 501882 26509
rect 502118 26273 502160 26509
rect 501840 26241 502160 26273
rect 507771 26829 508091 26861
rect 507771 26593 507813 26829
rect 508049 26593 508091 26829
rect 507771 26509 508091 26593
rect 507771 26273 507813 26509
rect 508049 26273 508091 26509
rect 507771 26241 508091 26273
rect 523910 26829 524230 26861
rect 523910 26593 523952 26829
rect 524188 26593 524230 26829
rect 523910 26509 524230 26593
rect 523910 26273 523952 26509
rect 524188 26273 524230 26509
rect 523910 26241 524230 26273
rect 529840 26829 530160 26861
rect 529840 26593 529882 26829
rect 530118 26593 530160 26829
rect 529840 26509 530160 26593
rect 529840 26273 529882 26509
rect 530118 26273 530160 26509
rect 529840 26241 530160 26273
rect 535771 26829 536091 26861
rect 535771 26593 535813 26829
rect 536049 26593 536091 26829
rect 535771 26509 536091 26593
rect 535771 26273 535813 26509
rect 536049 26273 536091 26509
rect 535771 26241 536091 26273
rect 551910 26829 552230 26861
rect 551910 26593 551952 26829
rect 552188 26593 552230 26829
rect 551910 26509 552230 26593
rect 551910 26273 551952 26509
rect 552188 26273 552230 26509
rect 551910 26241 552230 26273
rect 557840 26829 558160 26861
rect 557840 26593 557882 26829
rect 558118 26593 558160 26829
rect 557840 26509 558160 26593
rect 557840 26273 557882 26509
rect 558118 26273 558160 26509
rect 557840 26241 558160 26273
rect 563771 26829 564091 26861
rect 563771 26593 563813 26829
rect 564049 26593 564091 26829
rect 563771 26509 564091 26593
rect 563771 26273 563813 26509
rect 564049 26273 564091 26509
rect 563771 26241 564091 26273
rect 573494 26829 574114 53273
rect 573494 26593 573526 26829
rect 573762 26593 573846 26829
rect 574082 26593 574114 26829
rect 573494 26509 574114 26593
rect 573494 26273 573526 26509
rect 573762 26273 573846 26509
rect 574082 26273 574114 26509
rect 65994 23218 66026 23454
rect 66262 23218 66346 23454
rect 66582 23218 66614 23454
rect 65994 23134 66614 23218
rect 65994 22898 66026 23134
rect 66262 22898 66346 23134
rect 66582 22898 66614 23134
rect 48083 16556 48149 16557
rect 48083 16492 48084 16556
rect 48148 16492 48149 16556
rect 48083 16491 48149 16492
rect 42747 5676 42813 5677
rect 42747 5612 42748 5676
rect 42812 5612 42813 5676
rect 42747 5611 42813 5612
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 65994 -1306 66614 22898
rect 78874 23454 79194 23486
rect 78874 23218 78916 23454
rect 79152 23218 79194 23454
rect 78874 23134 79194 23218
rect 78874 22898 78916 23134
rect 79152 22898 79194 23134
rect 78874 22866 79194 22898
rect 84805 23454 85125 23486
rect 84805 23218 84847 23454
rect 85083 23218 85125 23454
rect 84805 23134 85125 23218
rect 84805 22898 84847 23134
rect 85083 22898 85125 23134
rect 84805 22866 85125 22898
rect 106874 23454 107194 23486
rect 106874 23218 106916 23454
rect 107152 23218 107194 23454
rect 106874 23134 107194 23218
rect 106874 22898 106916 23134
rect 107152 22898 107194 23134
rect 106874 22866 107194 22898
rect 112805 23454 113125 23486
rect 112805 23218 112847 23454
rect 113083 23218 113125 23454
rect 112805 23134 113125 23218
rect 112805 22898 112847 23134
rect 113083 22898 113125 23134
rect 112805 22866 113125 22898
rect 134874 23454 135194 23486
rect 134874 23218 134916 23454
rect 135152 23218 135194 23454
rect 134874 23134 135194 23218
rect 134874 22898 134916 23134
rect 135152 22898 135194 23134
rect 134874 22866 135194 22898
rect 140805 23454 141125 23486
rect 140805 23218 140847 23454
rect 141083 23218 141125 23454
rect 140805 23134 141125 23218
rect 140805 22898 140847 23134
rect 141083 22898 141125 23134
rect 140805 22866 141125 22898
rect 162874 23454 163194 23486
rect 162874 23218 162916 23454
rect 163152 23218 163194 23454
rect 162874 23134 163194 23218
rect 162874 22898 162916 23134
rect 163152 22898 163194 23134
rect 162874 22866 163194 22898
rect 168805 23454 169125 23486
rect 168805 23218 168847 23454
rect 169083 23218 169125 23454
rect 168805 23134 169125 23218
rect 168805 22898 168847 23134
rect 169083 22898 169125 23134
rect 168805 22866 169125 22898
rect 190874 23454 191194 23486
rect 190874 23218 190916 23454
rect 191152 23218 191194 23454
rect 190874 23134 191194 23218
rect 190874 22898 190916 23134
rect 191152 22898 191194 23134
rect 190874 22866 191194 22898
rect 196805 23454 197125 23486
rect 196805 23218 196847 23454
rect 197083 23218 197125 23454
rect 196805 23134 197125 23218
rect 196805 22898 196847 23134
rect 197083 22898 197125 23134
rect 196805 22866 197125 22898
rect 218874 23454 219194 23486
rect 218874 23218 218916 23454
rect 219152 23218 219194 23454
rect 218874 23134 219194 23218
rect 218874 22898 218916 23134
rect 219152 22898 219194 23134
rect 218874 22866 219194 22898
rect 224805 23454 225125 23486
rect 224805 23218 224847 23454
rect 225083 23218 225125 23454
rect 224805 23134 225125 23218
rect 224805 22898 224847 23134
rect 225083 22898 225125 23134
rect 224805 22866 225125 22898
rect 246874 23454 247194 23486
rect 246874 23218 246916 23454
rect 247152 23218 247194 23454
rect 246874 23134 247194 23218
rect 246874 22898 246916 23134
rect 247152 22898 247194 23134
rect 246874 22866 247194 22898
rect 252805 23454 253125 23486
rect 252805 23218 252847 23454
rect 253083 23218 253125 23454
rect 252805 23134 253125 23218
rect 252805 22898 252847 23134
rect 253083 22898 253125 23134
rect 252805 22866 253125 22898
rect 274874 23454 275194 23486
rect 274874 23218 274916 23454
rect 275152 23218 275194 23454
rect 274874 23134 275194 23218
rect 274874 22898 274916 23134
rect 275152 22898 275194 23134
rect 274874 22866 275194 22898
rect 280805 23454 281125 23486
rect 280805 23218 280847 23454
rect 281083 23218 281125 23454
rect 280805 23134 281125 23218
rect 280805 22898 280847 23134
rect 281083 22898 281125 23134
rect 280805 22866 281125 22898
rect 302874 23454 303194 23486
rect 302874 23218 302916 23454
rect 303152 23218 303194 23454
rect 302874 23134 303194 23218
rect 302874 22898 302916 23134
rect 303152 22898 303194 23134
rect 302874 22866 303194 22898
rect 308805 23454 309125 23486
rect 308805 23218 308847 23454
rect 309083 23218 309125 23454
rect 308805 23134 309125 23218
rect 308805 22898 308847 23134
rect 309083 22898 309125 23134
rect 308805 22866 309125 22898
rect 330874 23454 331194 23486
rect 330874 23218 330916 23454
rect 331152 23218 331194 23454
rect 330874 23134 331194 23218
rect 330874 22898 330916 23134
rect 331152 22898 331194 23134
rect 330874 22866 331194 22898
rect 336805 23454 337125 23486
rect 336805 23218 336847 23454
rect 337083 23218 337125 23454
rect 336805 23134 337125 23218
rect 336805 22898 336847 23134
rect 337083 22898 337125 23134
rect 336805 22866 337125 22898
rect 358874 23454 359194 23486
rect 358874 23218 358916 23454
rect 359152 23218 359194 23454
rect 358874 23134 359194 23218
rect 358874 22898 358916 23134
rect 359152 22898 359194 23134
rect 358874 22866 359194 22898
rect 364805 23454 365125 23486
rect 364805 23218 364847 23454
rect 365083 23218 365125 23454
rect 364805 23134 365125 23218
rect 364805 22898 364847 23134
rect 365083 22898 365125 23134
rect 364805 22866 365125 22898
rect 386874 23454 387194 23486
rect 386874 23218 386916 23454
rect 387152 23218 387194 23454
rect 386874 23134 387194 23218
rect 386874 22898 386916 23134
rect 387152 22898 387194 23134
rect 386874 22866 387194 22898
rect 392805 23454 393125 23486
rect 392805 23218 392847 23454
rect 393083 23218 393125 23454
rect 392805 23134 393125 23218
rect 392805 22898 392847 23134
rect 393083 22898 393125 23134
rect 392805 22866 393125 22898
rect 414874 23454 415194 23486
rect 414874 23218 414916 23454
rect 415152 23218 415194 23454
rect 414874 23134 415194 23218
rect 414874 22898 414916 23134
rect 415152 22898 415194 23134
rect 414874 22866 415194 22898
rect 420805 23454 421125 23486
rect 420805 23218 420847 23454
rect 421083 23218 421125 23454
rect 420805 23134 421125 23218
rect 420805 22898 420847 23134
rect 421083 22898 421125 23134
rect 420805 22866 421125 22898
rect 442874 23454 443194 23486
rect 442874 23218 442916 23454
rect 443152 23218 443194 23454
rect 442874 23134 443194 23218
rect 442874 22898 442916 23134
rect 443152 22898 443194 23134
rect 442874 22866 443194 22898
rect 448805 23454 449125 23486
rect 448805 23218 448847 23454
rect 449083 23218 449125 23454
rect 448805 23134 449125 23218
rect 448805 22898 448847 23134
rect 449083 22898 449125 23134
rect 448805 22866 449125 22898
rect 470874 23454 471194 23486
rect 470874 23218 470916 23454
rect 471152 23218 471194 23454
rect 470874 23134 471194 23218
rect 470874 22898 470916 23134
rect 471152 22898 471194 23134
rect 470874 22866 471194 22898
rect 476805 23454 477125 23486
rect 476805 23218 476847 23454
rect 477083 23218 477125 23454
rect 476805 23134 477125 23218
rect 476805 22898 476847 23134
rect 477083 22898 477125 23134
rect 476805 22866 477125 22898
rect 498874 23454 499194 23486
rect 498874 23218 498916 23454
rect 499152 23218 499194 23454
rect 498874 23134 499194 23218
rect 498874 22898 498916 23134
rect 499152 22898 499194 23134
rect 498874 22866 499194 22898
rect 504805 23454 505125 23486
rect 504805 23218 504847 23454
rect 505083 23218 505125 23454
rect 504805 23134 505125 23218
rect 504805 22898 504847 23134
rect 505083 22898 505125 23134
rect 504805 22866 505125 22898
rect 526874 23454 527194 23486
rect 526874 23218 526916 23454
rect 527152 23218 527194 23454
rect 526874 23134 527194 23218
rect 526874 22898 526916 23134
rect 527152 22898 527194 23134
rect 526874 22866 527194 22898
rect 532805 23454 533125 23486
rect 532805 23218 532847 23454
rect 533083 23218 533125 23454
rect 532805 23134 533125 23218
rect 532805 22898 532847 23134
rect 533083 22898 533125 23134
rect 532805 22866 533125 22898
rect 554874 23454 555194 23486
rect 554874 23218 554916 23454
rect 555152 23218 555194 23454
rect 554874 23134 555194 23218
rect 554874 22898 554916 23134
rect 555152 22898 555194 23134
rect 554874 22866 555194 22898
rect 560805 23454 561125 23486
rect 560805 23218 560847 23454
rect 561083 23218 561125 23454
rect 560805 23134 561125 23218
rect 560805 22898 560847 23134
rect 561083 22898 561125 23134
rect 560805 22866 561125 22898
rect 65994 -1542 66026 -1306
rect 66262 -1542 66346 -1306
rect 66582 -1542 66614 -1306
rect 65994 -1626 66614 -1542
rect 65994 -1862 66026 -1626
rect 66262 -1862 66346 -1626
rect 66582 -1862 66614 -1626
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 65994 -7654 66614 -1862
rect 573494 -346 574114 26273
rect 580214 13429 580274 670651
rect 585310 647829 585930 674273
rect 585310 647593 585342 647829
rect 585578 647593 585662 647829
rect 585898 647593 585930 647829
rect 585310 647509 585930 647593
rect 585310 647273 585342 647509
rect 585578 647273 585662 647509
rect 585898 647273 585930 647509
rect 580395 644060 580461 644061
rect 580395 643996 580396 644060
rect 580460 643996 580461 644060
rect 580395 643995 580461 643996
rect 580211 13428 580277 13429
rect 580211 13364 580212 13428
rect 580276 13364 580277 13428
rect 580211 13363 580277 13364
rect 580398 13157 580458 643995
rect 585310 620829 585930 647273
rect 585310 620593 585342 620829
rect 585578 620593 585662 620829
rect 585898 620593 585930 620829
rect 585310 620509 585930 620593
rect 585310 620273 585342 620509
rect 585578 620273 585662 620509
rect 585898 620273 585930 620509
rect 580579 617540 580645 617541
rect 580579 617476 580580 617540
rect 580644 617476 580645 617540
rect 580579 617475 580645 617476
rect 580582 13565 580642 617475
rect 585310 593829 585930 620273
rect 585310 593593 585342 593829
rect 585578 593593 585662 593829
rect 585898 593593 585930 593829
rect 585310 593509 585930 593593
rect 585310 593273 585342 593509
rect 585578 593273 585662 593509
rect 585898 593273 585930 593509
rect 585310 566829 585930 593273
rect 585310 566593 585342 566829
rect 585578 566593 585662 566829
rect 585898 566593 585930 566829
rect 585310 566509 585930 566593
rect 585310 566273 585342 566509
rect 585578 566273 585662 566509
rect 585898 566273 585930 566509
rect 580763 564364 580829 564365
rect 580763 564300 580764 564364
rect 580828 564300 580829 564364
rect 580763 564299 580829 564300
rect 580766 37909 580826 564299
rect 585310 539829 585930 566273
rect 585310 539593 585342 539829
rect 585578 539593 585662 539829
rect 585898 539593 585930 539829
rect 585310 539509 585930 539593
rect 585310 539273 585342 539509
rect 585578 539273 585662 539509
rect 585898 539273 585930 539509
rect 585310 512829 585930 539273
rect 585310 512593 585342 512829
rect 585578 512593 585662 512829
rect 585898 512593 585930 512829
rect 585310 512509 585930 512593
rect 585310 512273 585342 512509
rect 585578 512273 585662 512509
rect 585898 512273 585930 512509
rect 585310 485829 585930 512273
rect 585310 485593 585342 485829
rect 585578 485593 585662 485829
rect 585898 485593 585930 485829
rect 585310 485509 585930 485593
rect 585310 485273 585342 485509
rect 585578 485273 585662 485509
rect 585898 485273 585930 485509
rect 585310 458829 585930 485273
rect 585310 458593 585342 458829
rect 585578 458593 585662 458829
rect 585898 458593 585930 458829
rect 585310 458509 585930 458593
rect 585310 458273 585342 458509
rect 585578 458273 585662 458509
rect 585898 458273 585930 458509
rect 585310 431829 585930 458273
rect 585310 431593 585342 431829
rect 585578 431593 585662 431829
rect 585898 431593 585930 431829
rect 585310 431509 585930 431593
rect 585310 431273 585342 431509
rect 585578 431273 585662 431509
rect 585898 431273 585930 431509
rect 585310 404829 585930 431273
rect 585310 404593 585342 404829
rect 585578 404593 585662 404829
rect 585898 404593 585930 404829
rect 585310 404509 585930 404593
rect 585310 404273 585342 404509
rect 585578 404273 585662 404509
rect 585898 404273 585930 404509
rect 585310 377829 585930 404273
rect 585310 377593 585342 377829
rect 585578 377593 585662 377829
rect 585898 377593 585930 377829
rect 585310 377509 585930 377593
rect 585310 377273 585342 377509
rect 585578 377273 585662 377509
rect 585898 377273 585930 377509
rect 585310 350829 585930 377273
rect 585310 350593 585342 350829
rect 585578 350593 585662 350829
rect 585898 350593 585930 350829
rect 585310 350509 585930 350593
rect 585310 350273 585342 350509
rect 585578 350273 585662 350509
rect 585898 350273 585930 350509
rect 585310 323829 585930 350273
rect 585310 323593 585342 323829
rect 585578 323593 585662 323829
rect 585898 323593 585930 323829
rect 585310 323509 585930 323593
rect 585310 323273 585342 323509
rect 585578 323273 585662 323509
rect 585898 323273 585930 323509
rect 585310 296829 585930 323273
rect 585310 296593 585342 296829
rect 585578 296593 585662 296829
rect 585898 296593 585930 296829
rect 585310 296509 585930 296593
rect 585310 296273 585342 296509
rect 585578 296273 585662 296509
rect 585898 296273 585930 296509
rect 585310 269829 585930 296273
rect 585310 269593 585342 269829
rect 585578 269593 585662 269829
rect 585898 269593 585930 269829
rect 585310 269509 585930 269593
rect 585310 269273 585342 269509
rect 585578 269273 585662 269509
rect 585898 269273 585930 269509
rect 585310 242829 585930 269273
rect 585310 242593 585342 242829
rect 585578 242593 585662 242829
rect 585898 242593 585930 242829
rect 585310 242509 585930 242593
rect 585310 242273 585342 242509
rect 585578 242273 585662 242509
rect 585898 242273 585930 242509
rect 585310 215829 585930 242273
rect 585310 215593 585342 215829
rect 585578 215593 585662 215829
rect 585898 215593 585930 215829
rect 585310 215509 585930 215593
rect 585310 215273 585342 215509
rect 585578 215273 585662 215509
rect 585898 215273 585930 215509
rect 585310 188829 585930 215273
rect 585310 188593 585342 188829
rect 585578 188593 585662 188829
rect 585898 188593 585930 188829
rect 585310 188509 585930 188593
rect 585310 188273 585342 188509
rect 585578 188273 585662 188509
rect 585898 188273 585930 188509
rect 585310 161829 585930 188273
rect 585310 161593 585342 161829
rect 585578 161593 585662 161829
rect 585898 161593 585930 161829
rect 585310 161509 585930 161593
rect 585310 161273 585342 161509
rect 585578 161273 585662 161509
rect 585898 161273 585930 161509
rect 585310 134829 585930 161273
rect 585310 134593 585342 134829
rect 585578 134593 585662 134829
rect 585898 134593 585930 134829
rect 585310 134509 585930 134593
rect 585310 134273 585342 134509
rect 585578 134273 585662 134509
rect 585898 134273 585930 134509
rect 585310 107829 585930 134273
rect 585310 107593 585342 107829
rect 585578 107593 585662 107829
rect 585898 107593 585930 107829
rect 585310 107509 585930 107593
rect 585310 107273 585342 107509
rect 585578 107273 585662 107509
rect 585898 107273 585930 107509
rect 585310 80829 585930 107273
rect 585310 80593 585342 80829
rect 585578 80593 585662 80829
rect 585898 80593 585930 80829
rect 585310 80509 585930 80593
rect 585310 80273 585342 80509
rect 585578 80273 585662 80509
rect 585898 80273 585930 80509
rect 585310 53829 585930 80273
rect 585310 53593 585342 53829
rect 585578 53593 585662 53829
rect 585898 53593 585930 53829
rect 585310 53509 585930 53593
rect 585310 53273 585342 53509
rect 585578 53273 585662 53509
rect 585898 53273 585930 53509
rect 580763 37908 580829 37909
rect 580763 37844 580764 37908
rect 580828 37844 580829 37908
rect 580763 37843 580829 37844
rect 585310 26829 585930 53273
rect 585310 26593 585342 26829
rect 585578 26593 585662 26829
rect 585898 26593 585930 26829
rect 585310 26509 585930 26593
rect 585310 26273 585342 26509
rect 585578 26273 585662 26509
rect 585898 26273 585930 26509
rect 580579 13564 580645 13565
rect 580579 13500 580580 13564
rect 580644 13500 580645 13564
rect 580579 13499 580645 13500
rect 580395 13156 580461 13157
rect 580395 13092 580396 13156
rect 580460 13092 580461 13156
rect 580395 13091 580461 13092
rect 573494 -582 573526 -346
rect 573762 -582 573846 -346
rect 574082 -582 574114 -346
rect 573494 -666 574114 -582
rect 573494 -902 573526 -666
rect 573762 -902 573846 -666
rect 574082 -902 574114 -666
rect 573494 -7654 574114 -902
rect 585310 -346 585930 26273
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 698454 586890 705242
rect 586270 698218 586302 698454
rect 586538 698218 586622 698454
rect 586858 698218 586890 698454
rect 586270 698134 586890 698218
rect 586270 697898 586302 698134
rect 586538 697898 586622 698134
rect 586858 697898 586890 698134
rect 586270 671454 586890 697898
rect 586270 671218 586302 671454
rect 586538 671218 586622 671454
rect 586858 671218 586890 671454
rect 586270 671134 586890 671218
rect 586270 670898 586302 671134
rect 586538 670898 586622 671134
rect 586858 670898 586890 671134
rect 586270 644454 586890 670898
rect 586270 644218 586302 644454
rect 586538 644218 586622 644454
rect 586858 644218 586890 644454
rect 586270 644134 586890 644218
rect 586270 643898 586302 644134
rect 586538 643898 586622 644134
rect 586858 643898 586890 644134
rect 586270 617454 586890 643898
rect 586270 617218 586302 617454
rect 586538 617218 586622 617454
rect 586858 617218 586890 617454
rect 586270 617134 586890 617218
rect 586270 616898 586302 617134
rect 586538 616898 586622 617134
rect 586858 616898 586890 617134
rect 586270 590454 586890 616898
rect 586270 590218 586302 590454
rect 586538 590218 586622 590454
rect 586858 590218 586890 590454
rect 586270 590134 586890 590218
rect 586270 589898 586302 590134
rect 586538 589898 586622 590134
rect 586858 589898 586890 590134
rect 586270 563454 586890 589898
rect 586270 563218 586302 563454
rect 586538 563218 586622 563454
rect 586858 563218 586890 563454
rect 586270 563134 586890 563218
rect 586270 562898 586302 563134
rect 586538 562898 586622 563134
rect 586858 562898 586890 563134
rect 586270 536454 586890 562898
rect 586270 536218 586302 536454
rect 586538 536218 586622 536454
rect 586858 536218 586890 536454
rect 586270 536134 586890 536218
rect 586270 535898 586302 536134
rect 586538 535898 586622 536134
rect 586858 535898 586890 536134
rect 586270 509454 586890 535898
rect 586270 509218 586302 509454
rect 586538 509218 586622 509454
rect 586858 509218 586890 509454
rect 586270 509134 586890 509218
rect 586270 508898 586302 509134
rect 586538 508898 586622 509134
rect 586858 508898 586890 509134
rect 586270 482454 586890 508898
rect 586270 482218 586302 482454
rect 586538 482218 586622 482454
rect 586858 482218 586890 482454
rect 586270 482134 586890 482218
rect 586270 481898 586302 482134
rect 586538 481898 586622 482134
rect 586858 481898 586890 482134
rect 586270 455454 586890 481898
rect 586270 455218 586302 455454
rect 586538 455218 586622 455454
rect 586858 455218 586890 455454
rect 586270 455134 586890 455218
rect 586270 454898 586302 455134
rect 586538 454898 586622 455134
rect 586858 454898 586890 455134
rect 586270 428454 586890 454898
rect 586270 428218 586302 428454
rect 586538 428218 586622 428454
rect 586858 428218 586890 428454
rect 586270 428134 586890 428218
rect 586270 427898 586302 428134
rect 586538 427898 586622 428134
rect 586858 427898 586890 428134
rect 586270 401454 586890 427898
rect 586270 401218 586302 401454
rect 586538 401218 586622 401454
rect 586858 401218 586890 401454
rect 586270 401134 586890 401218
rect 586270 400898 586302 401134
rect 586538 400898 586622 401134
rect 586858 400898 586890 401134
rect 586270 374454 586890 400898
rect 586270 374218 586302 374454
rect 586538 374218 586622 374454
rect 586858 374218 586890 374454
rect 586270 374134 586890 374218
rect 586270 373898 586302 374134
rect 586538 373898 586622 374134
rect 586858 373898 586890 374134
rect 586270 347454 586890 373898
rect 586270 347218 586302 347454
rect 586538 347218 586622 347454
rect 586858 347218 586890 347454
rect 586270 347134 586890 347218
rect 586270 346898 586302 347134
rect 586538 346898 586622 347134
rect 586858 346898 586890 347134
rect 586270 320454 586890 346898
rect 586270 320218 586302 320454
rect 586538 320218 586622 320454
rect 586858 320218 586890 320454
rect 586270 320134 586890 320218
rect 586270 319898 586302 320134
rect 586538 319898 586622 320134
rect 586858 319898 586890 320134
rect 586270 293454 586890 319898
rect 586270 293218 586302 293454
rect 586538 293218 586622 293454
rect 586858 293218 586890 293454
rect 586270 293134 586890 293218
rect 586270 292898 586302 293134
rect 586538 292898 586622 293134
rect 586858 292898 586890 293134
rect 586270 266454 586890 292898
rect 586270 266218 586302 266454
rect 586538 266218 586622 266454
rect 586858 266218 586890 266454
rect 586270 266134 586890 266218
rect 586270 265898 586302 266134
rect 586538 265898 586622 266134
rect 586858 265898 586890 266134
rect 586270 239454 586890 265898
rect 586270 239218 586302 239454
rect 586538 239218 586622 239454
rect 586858 239218 586890 239454
rect 586270 239134 586890 239218
rect 586270 238898 586302 239134
rect 586538 238898 586622 239134
rect 586858 238898 586890 239134
rect 586270 212454 586890 238898
rect 586270 212218 586302 212454
rect 586538 212218 586622 212454
rect 586858 212218 586890 212454
rect 586270 212134 586890 212218
rect 586270 211898 586302 212134
rect 586538 211898 586622 212134
rect 586858 211898 586890 212134
rect 586270 185454 586890 211898
rect 586270 185218 586302 185454
rect 586538 185218 586622 185454
rect 586858 185218 586890 185454
rect 586270 185134 586890 185218
rect 586270 184898 586302 185134
rect 586538 184898 586622 185134
rect 586858 184898 586890 185134
rect 586270 158454 586890 184898
rect 586270 158218 586302 158454
rect 586538 158218 586622 158454
rect 586858 158218 586890 158454
rect 586270 158134 586890 158218
rect 586270 157898 586302 158134
rect 586538 157898 586622 158134
rect 586858 157898 586890 158134
rect 586270 131454 586890 157898
rect 586270 131218 586302 131454
rect 586538 131218 586622 131454
rect 586858 131218 586890 131454
rect 586270 131134 586890 131218
rect 586270 130898 586302 131134
rect 586538 130898 586622 131134
rect 586858 130898 586890 131134
rect 586270 104454 586890 130898
rect 586270 104218 586302 104454
rect 586538 104218 586622 104454
rect 586858 104218 586890 104454
rect 586270 104134 586890 104218
rect 586270 103898 586302 104134
rect 586538 103898 586622 104134
rect 586858 103898 586890 104134
rect 586270 77454 586890 103898
rect 586270 77218 586302 77454
rect 586538 77218 586622 77454
rect 586858 77218 586890 77454
rect 586270 77134 586890 77218
rect 586270 76898 586302 77134
rect 586538 76898 586622 77134
rect 586858 76898 586890 77134
rect 586270 50454 586890 76898
rect 586270 50218 586302 50454
rect 586538 50218 586622 50454
rect 586858 50218 586890 50454
rect 586270 50134 586890 50218
rect 586270 49898 586302 50134
rect 586538 49898 586622 50134
rect 586858 49898 586890 50134
rect 586270 23454 586890 49898
rect 586270 23218 586302 23454
rect 586538 23218 586622 23454
rect 586858 23218 586890 23454
rect 586270 23134 586890 23218
rect 586270 22898 586302 23134
rect 586538 22898 586622 23134
rect 586858 22898 586890 23134
rect 586270 -1306 586890 22898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 -2266 587850 706202
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 -3226 588810 707162
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 -4186 589770 708122
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 -5146 590730 709082
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 -6106 591690 710042
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 -7066 592650 711002
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect 38026 705562 38262 705798
rect 38346 705562 38582 705798
rect 38026 705242 38262 705478
rect 38346 705242 38582 705478
rect -2934 698218 -2698 698454
rect -2614 698218 -2378 698454
rect -2934 697898 -2698 698134
rect -2614 697898 -2378 698134
rect -2934 671218 -2698 671454
rect -2614 671218 -2378 671454
rect -2934 670898 -2698 671134
rect -2614 670898 -2378 671134
rect -2934 644218 -2698 644454
rect -2614 644218 -2378 644454
rect -2934 643898 -2698 644134
rect -2614 643898 -2378 644134
rect -2934 617218 -2698 617454
rect -2614 617218 -2378 617454
rect -2934 616898 -2698 617134
rect -2614 616898 -2378 617134
rect -2934 590218 -2698 590454
rect -2614 590218 -2378 590454
rect -2934 589898 -2698 590134
rect -2614 589898 -2378 590134
rect -2934 563218 -2698 563454
rect -2614 563218 -2378 563454
rect -2934 562898 -2698 563134
rect -2614 562898 -2378 563134
rect -2934 536218 -2698 536454
rect -2614 536218 -2378 536454
rect -2934 535898 -2698 536134
rect -2614 535898 -2378 536134
rect -2934 509218 -2698 509454
rect -2614 509218 -2378 509454
rect -2934 508898 -2698 509134
rect -2614 508898 -2378 509134
rect -2934 482218 -2698 482454
rect -2614 482218 -2378 482454
rect -2934 481898 -2698 482134
rect -2614 481898 -2378 482134
rect -2934 455218 -2698 455454
rect -2614 455218 -2378 455454
rect -2934 454898 -2698 455134
rect -2614 454898 -2378 455134
rect -2934 428218 -2698 428454
rect -2614 428218 -2378 428454
rect -2934 427898 -2698 428134
rect -2614 427898 -2378 428134
rect -2934 401218 -2698 401454
rect -2614 401218 -2378 401454
rect -2934 400898 -2698 401134
rect -2614 400898 -2378 401134
rect -2934 374218 -2698 374454
rect -2614 374218 -2378 374454
rect -2934 373898 -2698 374134
rect -2614 373898 -2378 374134
rect -2934 347218 -2698 347454
rect -2614 347218 -2378 347454
rect -2934 346898 -2698 347134
rect -2614 346898 -2378 347134
rect -2934 320218 -2698 320454
rect -2614 320218 -2378 320454
rect -2934 319898 -2698 320134
rect -2614 319898 -2378 320134
rect -2934 293218 -2698 293454
rect -2614 293218 -2378 293454
rect -2934 292898 -2698 293134
rect -2614 292898 -2378 293134
rect -2934 266218 -2698 266454
rect -2614 266218 -2378 266454
rect -2934 265898 -2698 266134
rect -2614 265898 -2378 266134
rect -2934 239218 -2698 239454
rect -2614 239218 -2378 239454
rect -2934 238898 -2698 239134
rect -2614 238898 -2378 239134
rect -2934 212218 -2698 212454
rect -2614 212218 -2378 212454
rect -2934 211898 -2698 212134
rect -2614 211898 -2378 212134
rect -2934 185218 -2698 185454
rect -2614 185218 -2378 185454
rect -2934 184898 -2698 185134
rect -2614 184898 -2378 185134
rect -2934 158218 -2698 158454
rect -2614 158218 -2378 158454
rect -2934 157898 -2698 158134
rect -2614 157898 -2378 158134
rect -2934 131218 -2698 131454
rect -2614 131218 -2378 131454
rect -2934 130898 -2698 131134
rect -2614 130898 -2378 131134
rect -2934 104218 -2698 104454
rect -2614 104218 -2378 104454
rect -2934 103898 -2698 104134
rect -2614 103898 -2378 104134
rect -2934 77218 -2698 77454
rect -2614 77218 -2378 77454
rect -2934 76898 -2698 77134
rect -2614 76898 -2378 77134
rect -2934 50218 -2698 50454
rect -2614 50218 -2378 50454
rect -2934 49898 -2698 50134
rect -2614 49898 -2378 50134
rect -2934 23218 -2698 23454
rect -2614 23218 -2378 23454
rect -2934 22898 -2698 23134
rect -2614 22898 -2378 23134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 701593 -1738 701829
rect -1654 701593 -1418 701829
rect -1974 701273 -1738 701509
rect -1654 701273 -1418 701509
rect 38026 698218 38262 698454
rect 38346 698218 38582 698454
rect 38026 697898 38262 698134
rect 38346 697898 38582 698134
rect 41526 704602 41762 704838
rect 41846 704602 42082 704838
rect 41526 704282 41762 704518
rect 41846 704282 42082 704518
rect 41526 701593 41762 701829
rect 41846 701593 42082 701829
rect 41526 701273 41762 701509
rect 41846 701273 42082 701509
rect 66026 705562 66262 705798
rect 66346 705562 66582 705798
rect 66026 705242 66262 705478
rect 66346 705242 66582 705478
rect 66026 698218 66262 698454
rect 66346 698218 66582 698454
rect 66026 697898 66262 698134
rect 66346 697898 66582 698134
rect 69526 704602 69762 704838
rect 69846 704602 70082 704838
rect 69526 704282 69762 704518
rect 69846 704282 70082 704518
rect 69526 701593 69762 701829
rect 69846 701593 70082 701829
rect 69526 701273 69762 701509
rect 69846 701273 70082 701509
rect 94026 705562 94262 705798
rect 94346 705562 94582 705798
rect 94026 705242 94262 705478
rect 94346 705242 94582 705478
rect 94026 698218 94262 698454
rect 94346 698218 94582 698454
rect 94026 697898 94262 698134
rect 94346 697898 94582 698134
rect 97526 704602 97762 704838
rect 97846 704602 98082 704838
rect 97526 704282 97762 704518
rect 97846 704282 98082 704518
rect 97526 701593 97762 701829
rect 97846 701593 98082 701829
rect 97526 701273 97762 701509
rect 97846 701273 98082 701509
rect 122026 705562 122262 705798
rect 122346 705562 122582 705798
rect 122026 705242 122262 705478
rect 122346 705242 122582 705478
rect 122026 698218 122262 698454
rect 122346 698218 122582 698454
rect 122026 697898 122262 698134
rect 122346 697898 122582 698134
rect 125526 704602 125762 704838
rect 125846 704602 126082 704838
rect 125526 704282 125762 704518
rect 125846 704282 126082 704518
rect 125526 701593 125762 701829
rect 125846 701593 126082 701829
rect 125526 701273 125762 701509
rect 125846 701273 126082 701509
rect 150026 705562 150262 705798
rect 150346 705562 150582 705798
rect 150026 705242 150262 705478
rect 150346 705242 150582 705478
rect 150026 698218 150262 698454
rect 150346 698218 150582 698454
rect 150026 697898 150262 698134
rect 150346 697898 150582 698134
rect 153526 704602 153762 704838
rect 153846 704602 154082 704838
rect 153526 704282 153762 704518
rect 153846 704282 154082 704518
rect 153526 701593 153762 701829
rect 153846 701593 154082 701829
rect 153526 701273 153762 701509
rect 153846 701273 154082 701509
rect 178026 705562 178262 705798
rect 178346 705562 178582 705798
rect 178026 705242 178262 705478
rect 178346 705242 178582 705478
rect 178026 698218 178262 698454
rect 178346 698218 178582 698454
rect 178026 697898 178262 698134
rect 178346 697898 178582 698134
rect 181526 704602 181762 704838
rect 181846 704602 182082 704838
rect 181526 704282 181762 704518
rect 181846 704282 182082 704518
rect 181526 701593 181762 701829
rect 181846 701593 182082 701829
rect 181526 701273 181762 701509
rect 181846 701273 182082 701509
rect 206026 705562 206262 705798
rect 206346 705562 206582 705798
rect 206026 705242 206262 705478
rect 206346 705242 206582 705478
rect 206026 698218 206262 698454
rect 206346 698218 206582 698454
rect 206026 697898 206262 698134
rect 206346 697898 206582 698134
rect 209526 704602 209762 704838
rect 209846 704602 210082 704838
rect 209526 704282 209762 704518
rect 209846 704282 210082 704518
rect 209526 701593 209762 701829
rect 209846 701593 210082 701829
rect 209526 701273 209762 701509
rect 209846 701273 210082 701509
rect 234026 705562 234262 705798
rect 234346 705562 234582 705798
rect 234026 705242 234262 705478
rect 234346 705242 234582 705478
rect 234026 698218 234262 698454
rect 234346 698218 234582 698454
rect 234026 697898 234262 698134
rect 234346 697898 234582 698134
rect 237526 704602 237762 704838
rect 237846 704602 238082 704838
rect 237526 704282 237762 704518
rect 237846 704282 238082 704518
rect 237526 701593 237762 701829
rect 237846 701593 238082 701829
rect 237526 701273 237762 701509
rect 237846 701273 238082 701509
rect 262026 705562 262262 705798
rect 262346 705562 262582 705798
rect 262026 705242 262262 705478
rect 262346 705242 262582 705478
rect 262026 698218 262262 698454
rect 262346 698218 262582 698454
rect 262026 697898 262262 698134
rect 262346 697898 262582 698134
rect 265526 704602 265762 704838
rect 265846 704602 266082 704838
rect 265526 704282 265762 704518
rect 265846 704282 266082 704518
rect 265526 701593 265762 701829
rect 265846 701593 266082 701829
rect 265526 701273 265762 701509
rect 265846 701273 266082 701509
rect 290026 705562 290262 705798
rect 290346 705562 290582 705798
rect 290026 705242 290262 705478
rect 290346 705242 290582 705478
rect 290026 698218 290262 698454
rect 290346 698218 290582 698454
rect 290026 697898 290262 698134
rect 290346 697898 290582 698134
rect 293526 704602 293762 704838
rect 293846 704602 294082 704838
rect 293526 704282 293762 704518
rect 293846 704282 294082 704518
rect 293526 701593 293762 701829
rect 293846 701593 294082 701829
rect 293526 701273 293762 701509
rect 293846 701273 294082 701509
rect 318026 705562 318262 705798
rect 318346 705562 318582 705798
rect 318026 705242 318262 705478
rect 318346 705242 318582 705478
rect 318026 698218 318262 698454
rect 318346 698218 318582 698454
rect 318026 697898 318262 698134
rect 318346 697898 318582 698134
rect 321526 704602 321762 704838
rect 321846 704602 322082 704838
rect 321526 704282 321762 704518
rect 321846 704282 322082 704518
rect 321526 701593 321762 701829
rect 321846 701593 322082 701829
rect 321526 701273 321762 701509
rect 321846 701273 322082 701509
rect 346026 705562 346262 705798
rect 346346 705562 346582 705798
rect 346026 705242 346262 705478
rect 346346 705242 346582 705478
rect 346026 698218 346262 698454
rect 346346 698218 346582 698454
rect 346026 697898 346262 698134
rect 346346 697898 346582 698134
rect 349526 704602 349762 704838
rect 349846 704602 350082 704838
rect 349526 704282 349762 704518
rect 349846 704282 350082 704518
rect 349526 701593 349762 701829
rect 349846 701593 350082 701829
rect 349526 701273 349762 701509
rect 349846 701273 350082 701509
rect 374026 705562 374262 705798
rect 374346 705562 374582 705798
rect 374026 705242 374262 705478
rect 374346 705242 374582 705478
rect 374026 698218 374262 698454
rect 374346 698218 374582 698454
rect 374026 697898 374262 698134
rect 374346 697898 374582 698134
rect 377526 704602 377762 704838
rect 377846 704602 378082 704838
rect 377526 704282 377762 704518
rect 377846 704282 378082 704518
rect 377526 701593 377762 701829
rect 377846 701593 378082 701829
rect 377526 701273 377762 701509
rect 377846 701273 378082 701509
rect 402026 705562 402262 705798
rect 402346 705562 402582 705798
rect 402026 705242 402262 705478
rect 402346 705242 402582 705478
rect 402026 698218 402262 698454
rect 402346 698218 402582 698454
rect 402026 697898 402262 698134
rect 402346 697898 402582 698134
rect 405526 704602 405762 704838
rect 405846 704602 406082 704838
rect 405526 704282 405762 704518
rect 405846 704282 406082 704518
rect 405526 701593 405762 701829
rect 405846 701593 406082 701829
rect 405526 701273 405762 701509
rect 405846 701273 406082 701509
rect 430026 705562 430262 705798
rect 430346 705562 430582 705798
rect 430026 705242 430262 705478
rect 430346 705242 430582 705478
rect 430026 698218 430262 698454
rect 430346 698218 430582 698454
rect 430026 697898 430262 698134
rect 430346 697898 430582 698134
rect 433526 704602 433762 704838
rect 433846 704602 434082 704838
rect 433526 704282 433762 704518
rect 433846 704282 434082 704518
rect 433526 701593 433762 701829
rect 433846 701593 434082 701829
rect 433526 701273 433762 701509
rect 433846 701273 434082 701509
rect 458026 705562 458262 705798
rect 458346 705562 458582 705798
rect 458026 705242 458262 705478
rect 458346 705242 458582 705478
rect 458026 698218 458262 698454
rect 458346 698218 458582 698454
rect 458026 697898 458262 698134
rect 458346 697898 458582 698134
rect 461526 704602 461762 704838
rect 461846 704602 462082 704838
rect 461526 704282 461762 704518
rect 461846 704282 462082 704518
rect 461526 701593 461762 701829
rect 461846 701593 462082 701829
rect 461526 701273 461762 701509
rect 461846 701273 462082 701509
rect 486026 705562 486262 705798
rect 486346 705562 486582 705798
rect 486026 705242 486262 705478
rect 486346 705242 486582 705478
rect 486026 698218 486262 698454
rect 486346 698218 486582 698454
rect 486026 697898 486262 698134
rect 486346 697898 486582 698134
rect 489526 704602 489762 704838
rect 489846 704602 490082 704838
rect 489526 704282 489762 704518
rect 489846 704282 490082 704518
rect 489526 701593 489762 701829
rect 489846 701593 490082 701829
rect 489526 701273 489762 701509
rect 489846 701273 490082 701509
rect 514026 705562 514262 705798
rect 514346 705562 514582 705798
rect 514026 705242 514262 705478
rect 514346 705242 514582 705478
rect 514026 698218 514262 698454
rect 514346 698218 514582 698454
rect 514026 697898 514262 698134
rect 514346 697898 514582 698134
rect 517526 704602 517762 704838
rect 517846 704602 518082 704838
rect 517526 704282 517762 704518
rect 517846 704282 518082 704518
rect 517526 701593 517762 701829
rect 517846 701593 518082 701829
rect 517526 701273 517762 701509
rect 517846 701273 518082 701509
rect 542026 705562 542262 705798
rect 542346 705562 542582 705798
rect 542026 705242 542262 705478
rect 542346 705242 542582 705478
rect 542026 698218 542262 698454
rect 542346 698218 542582 698454
rect 542026 697898 542262 698134
rect 542346 697898 542582 698134
rect 545526 704602 545762 704838
rect 545846 704602 546082 704838
rect 545526 704282 545762 704518
rect 545846 704282 546082 704518
rect 545526 701593 545762 701829
rect 545846 701593 546082 701829
rect 545526 701273 545762 701509
rect 545846 701273 546082 701509
rect 570026 705562 570262 705798
rect 570346 705562 570582 705798
rect 570026 705242 570262 705478
rect 570346 705242 570582 705478
rect 570026 698218 570262 698454
rect 570346 698218 570582 698454
rect 570026 697898 570262 698134
rect 570346 697898 570582 698134
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 573526 704602 573762 704838
rect 573846 704602 574082 704838
rect 573526 704282 573762 704518
rect 573846 704282 574082 704518
rect 573526 701593 573762 701829
rect 573846 701593 574082 701829
rect 573526 701273 573762 701509
rect 573846 701273 574082 701509
rect -1974 674593 -1738 674829
rect -1654 674593 -1418 674829
rect -1974 674273 -1738 674509
rect -1654 674273 -1418 674509
rect 19952 674593 20188 674829
rect 19952 674273 20188 674509
rect 25882 674593 26118 674829
rect 25882 674273 26118 674509
rect 31813 674593 32049 674829
rect 31813 674273 32049 674509
rect 47952 674593 48188 674829
rect 47952 674273 48188 674509
rect 53882 674593 54118 674829
rect 53882 674273 54118 674509
rect 59813 674593 60049 674829
rect 59813 674273 60049 674509
rect 75952 674593 76188 674829
rect 75952 674273 76188 674509
rect 81882 674593 82118 674829
rect 81882 674273 82118 674509
rect 87813 674593 88049 674829
rect 87813 674273 88049 674509
rect 103952 674593 104188 674829
rect 103952 674273 104188 674509
rect 109882 674593 110118 674829
rect 109882 674273 110118 674509
rect 115813 674593 116049 674829
rect 115813 674273 116049 674509
rect 131952 674593 132188 674829
rect 131952 674273 132188 674509
rect 137882 674593 138118 674829
rect 137882 674273 138118 674509
rect 143813 674593 144049 674829
rect 143813 674273 144049 674509
rect 159952 674593 160188 674829
rect 159952 674273 160188 674509
rect 165882 674593 166118 674829
rect 165882 674273 166118 674509
rect 171813 674593 172049 674829
rect 171813 674273 172049 674509
rect 187952 674593 188188 674829
rect 187952 674273 188188 674509
rect 193882 674593 194118 674829
rect 193882 674273 194118 674509
rect 199813 674593 200049 674829
rect 199813 674273 200049 674509
rect 215952 674593 216188 674829
rect 215952 674273 216188 674509
rect 221882 674593 222118 674829
rect 221882 674273 222118 674509
rect 227813 674593 228049 674829
rect 227813 674273 228049 674509
rect 243952 674593 244188 674829
rect 243952 674273 244188 674509
rect 249882 674593 250118 674829
rect 249882 674273 250118 674509
rect 255813 674593 256049 674829
rect 255813 674273 256049 674509
rect 271952 674593 272188 674829
rect 271952 674273 272188 674509
rect 277882 674593 278118 674829
rect 277882 674273 278118 674509
rect 283813 674593 284049 674829
rect 283813 674273 284049 674509
rect 299952 674593 300188 674829
rect 299952 674273 300188 674509
rect 305882 674593 306118 674829
rect 305882 674273 306118 674509
rect 311813 674593 312049 674829
rect 311813 674273 312049 674509
rect 327952 674593 328188 674829
rect 327952 674273 328188 674509
rect 333882 674593 334118 674829
rect 333882 674273 334118 674509
rect 339813 674593 340049 674829
rect 339813 674273 340049 674509
rect 355952 674593 356188 674829
rect 355952 674273 356188 674509
rect 361882 674593 362118 674829
rect 361882 674273 362118 674509
rect 367813 674593 368049 674829
rect 367813 674273 368049 674509
rect 383952 674593 384188 674829
rect 383952 674273 384188 674509
rect 389882 674593 390118 674829
rect 389882 674273 390118 674509
rect 395813 674593 396049 674829
rect 395813 674273 396049 674509
rect 411952 674593 412188 674829
rect 411952 674273 412188 674509
rect 417882 674593 418118 674829
rect 417882 674273 418118 674509
rect 423813 674593 424049 674829
rect 423813 674273 424049 674509
rect 439952 674593 440188 674829
rect 439952 674273 440188 674509
rect 445882 674593 446118 674829
rect 445882 674273 446118 674509
rect 451813 674593 452049 674829
rect 451813 674273 452049 674509
rect 467952 674593 468188 674829
rect 467952 674273 468188 674509
rect 473882 674593 474118 674829
rect 473882 674273 474118 674509
rect 479813 674593 480049 674829
rect 479813 674273 480049 674509
rect 495952 674593 496188 674829
rect 495952 674273 496188 674509
rect 501882 674593 502118 674829
rect 501882 674273 502118 674509
rect 507813 674593 508049 674829
rect 507813 674273 508049 674509
rect 523952 674593 524188 674829
rect 523952 674273 524188 674509
rect 529882 674593 530118 674829
rect 529882 674273 530118 674509
rect 535813 674593 536049 674829
rect 535813 674273 536049 674509
rect 551952 674593 552188 674829
rect 551952 674273 552188 674509
rect 557882 674593 558118 674829
rect 557882 674273 558118 674509
rect 563813 674593 564049 674829
rect 563813 674273 564049 674509
rect 573526 674593 573762 674829
rect 573846 674593 574082 674829
rect 573526 674273 573762 674509
rect 573846 674273 574082 674509
rect 22916 671218 23152 671454
rect 22916 670898 23152 671134
rect 28847 671218 29083 671454
rect 28847 670898 29083 671134
rect 50916 671218 51152 671454
rect 50916 670898 51152 671134
rect 56847 671218 57083 671454
rect 56847 670898 57083 671134
rect 78916 671218 79152 671454
rect 78916 670898 79152 671134
rect 84847 671218 85083 671454
rect 84847 670898 85083 671134
rect 106916 671218 107152 671454
rect 106916 670898 107152 671134
rect 112847 671218 113083 671454
rect 112847 670898 113083 671134
rect 134916 671218 135152 671454
rect 134916 670898 135152 671134
rect 140847 671218 141083 671454
rect 140847 670898 141083 671134
rect 162916 671218 163152 671454
rect 162916 670898 163152 671134
rect 168847 671218 169083 671454
rect 168847 670898 169083 671134
rect 190916 671218 191152 671454
rect 190916 670898 191152 671134
rect 196847 671218 197083 671454
rect 196847 670898 197083 671134
rect 218916 671218 219152 671454
rect 218916 670898 219152 671134
rect 224847 671218 225083 671454
rect 224847 670898 225083 671134
rect 246916 671218 247152 671454
rect 246916 670898 247152 671134
rect 252847 671218 253083 671454
rect 252847 670898 253083 671134
rect 274916 671218 275152 671454
rect 274916 670898 275152 671134
rect 280847 671218 281083 671454
rect 280847 670898 281083 671134
rect 302916 671218 303152 671454
rect 302916 670898 303152 671134
rect 308847 671218 309083 671454
rect 308847 670898 309083 671134
rect 330916 671218 331152 671454
rect 330916 670898 331152 671134
rect 336847 671218 337083 671454
rect 336847 670898 337083 671134
rect 358916 671218 359152 671454
rect 358916 670898 359152 671134
rect 364847 671218 365083 671454
rect 364847 670898 365083 671134
rect 386916 671218 387152 671454
rect 386916 670898 387152 671134
rect 392847 671218 393083 671454
rect 392847 670898 393083 671134
rect 414916 671218 415152 671454
rect 414916 670898 415152 671134
rect 420847 671218 421083 671454
rect 420847 670898 421083 671134
rect 442916 671218 443152 671454
rect 442916 670898 443152 671134
rect 448847 671218 449083 671454
rect 448847 670898 449083 671134
rect 470916 671218 471152 671454
rect 470916 670898 471152 671134
rect 476847 671218 477083 671454
rect 476847 670898 477083 671134
rect 498916 671218 499152 671454
rect 498916 670898 499152 671134
rect 504847 671218 505083 671454
rect 504847 670898 505083 671134
rect 526916 671218 527152 671454
rect 526916 670898 527152 671134
rect 532847 671218 533083 671454
rect 532847 670898 533083 671134
rect 554916 671218 555152 671454
rect 554916 670898 555152 671134
rect 560847 671218 561083 671454
rect 560847 670898 561083 671134
rect -1974 647593 -1738 647829
rect -1654 647593 -1418 647829
rect -1974 647273 -1738 647509
rect -1654 647273 -1418 647509
rect 19951 647593 20187 647829
rect 19951 647273 20187 647509
rect 25882 647593 26118 647829
rect 25882 647273 26118 647509
rect 31812 647593 32048 647829
rect 31812 647273 32048 647509
rect 47951 647593 48187 647829
rect 47951 647273 48187 647509
rect 53882 647593 54118 647829
rect 53882 647273 54118 647509
rect 59812 647593 60048 647829
rect 59812 647273 60048 647509
rect 75951 647593 76187 647829
rect 75951 647273 76187 647509
rect 81882 647593 82118 647829
rect 81882 647273 82118 647509
rect 87812 647593 88048 647829
rect 87812 647273 88048 647509
rect 103951 647593 104187 647829
rect 103951 647273 104187 647509
rect 109882 647593 110118 647829
rect 109882 647273 110118 647509
rect 115812 647593 116048 647829
rect 115812 647273 116048 647509
rect 131951 647593 132187 647829
rect 131951 647273 132187 647509
rect 137882 647593 138118 647829
rect 137882 647273 138118 647509
rect 143812 647593 144048 647829
rect 143812 647273 144048 647509
rect 159951 647593 160187 647829
rect 159951 647273 160187 647509
rect 165882 647593 166118 647829
rect 165882 647273 166118 647509
rect 171812 647593 172048 647829
rect 171812 647273 172048 647509
rect 187951 647593 188187 647829
rect 187951 647273 188187 647509
rect 193882 647593 194118 647829
rect 193882 647273 194118 647509
rect 199812 647593 200048 647829
rect 199812 647273 200048 647509
rect 215951 647593 216187 647829
rect 215951 647273 216187 647509
rect 221882 647593 222118 647829
rect 221882 647273 222118 647509
rect 227812 647593 228048 647829
rect 227812 647273 228048 647509
rect 243951 647593 244187 647829
rect 243951 647273 244187 647509
rect 249882 647593 250118 647829
rect 249882 647273 250118 647509
rect 255812 647593 256048 647829
rect 255812 647273 256048 647509
rect 271951 647593 272187 647829
rect 271951 647273 272187 647509
rect 277882 647593 278118 647829
rect 277882 647273 278118 647509
rect 283812 647593 284048 647829
rect 283812 647273 284048 647509
rect 299951 647593 300187 647829
rect 299951 647273 300187 647509
rect 305882 647593 306118 647829
rect 305882 647273 306118 647509
rect 311812 647593 312048 647829
rect 311812 647273 312048 647509
rect 327951 647593 328187 647829
rect 327951 647273 328187 647509
rect 333882 647593 334118 647829
rect 333882 647273 334118 647509
rect 339812 647593 340048 647829
rect 339812 647273 340048 647509
rect 355951 647593 356187 647829
rect 355951 647273 356187 647509
rect 361882 647593 362118 647829
rect 361882 647273 362118 647509
rect 367812 647593 368048 647829
rect 367812 647273 368048 647509
rect 383951 647593 384187 647829
rect 383951 647273 384187 647509
rect 389882 647593 390118 647829
rect 389882 647273 390118 647509
rect 395812 647593 396048 647829
rect 395812 647273 396048 647509
rect 411951 647593 412187 647829
rect 411951 647273 412187 647509
rect 417882 647593 418118 647829
rect 417882 647273 418118 647509
rect 423812 647593 424048 647829
rect 423812 647273 424048 647509
rect 439951 647593 440187 647829
rect 439951 647273 440187 647509
rect 445882 647593 446118 647829
rect 445882 647273 446118 647509
rect 451812 647593 452048 647829
rect 451812 647273 452048 647509
rect 467951 647593 468187 647829
rect 467951 647273 468187 647509
rect 473882 647593 474118 647829
rect 473882 647273 474118 647509
rect 479812 647593 480048 647829
rect 479812 647273 480048 647509
rect 495951 647593 496187 647829
rect 495951 647273 496187 647509
rect 501882 647593 502118 647829
rect 501882 647273 502118 647509
rect 507812 647593 508048 647829
rect 507812 647273 508048 647509
rect 523951 647593 524187 647829
rect 523951 647273 524187 647509
rect 529882 647593 530118 647829
rect 529882 647273 530118 647509
rect 535812 647593 536048 647829
rect 535812 647273 536048 647509
rect 551951 647593 552187 647829
rect 551951 647273 552187 647509
rect 557882 647593 558118 647829
rect 557882 647273 558118 647509
rect 563812 647593 564048 647829
rect 563812 647273 564048 647509
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 701593 585578 701829
rect 585662 701593 585898 701829
rect 585342 701273 585578 701509
rect 585662 701273 585898 701509
rect 585342 674593 585578 674829
rect 585662 674593 585898 674829
rect 585342 674273 585578 674509
rect 585662 674273 585898 674509
rect 573526 647593 573762 647829
rect 573846 647593 574082 647829
rect 573526 647273 573762 647509
rect 573846 647273 574082 647509
rect 22917 644218 23153 644454
rect 22917 643898 23153 644134
rect 28848 644218 29084 644454
rect 28848 643898 29084 644134
rect 50917 644218 51153 644454
rect 50917 643898 51153 644134
rect 56848 644218 57084 644454
rect 56848 643898 57084 644134
rect 78917 644218 79153 644454
rect 78917 643898 79153 644134
rect 84848 644218 85084 644454
rect 84848 643898 85084 644134
rect 106917 644218 107153 644454
rect 106917 643898 107153 644134
rect 112848 644218 113084 644454
rect 112848 643898 113084 644134
rect 134917 644218 135153 644454
rect 134917 643898 135153 644134
rect 140848 644218 141084 644454
rect 140848 643898 141084 644134
rect 162917 644218 163153 644454
rect 162917 643898 163153 644134
rect 168848 644218 169084 644454
rect 168848 643898 169084 644134
rect 190917 644218 191153 644454
rect 190917 643898 191153 644134
rect 196848 644218 197084 644454
rect 196848 643898 197084 644134
rect 218917 644218 219153 644454
rect 218917 643898 219153 644134
rect 224848 644218 225084 644454
rect 224848 643898 225084 644134
rect 246917 644218 247153 644454
rect 246917 643898 247153 644134
rect 252848 644218 253084 644454
rect 252848 643898 253084 644134
rect 274917 644218 275153 644454
rect 274917 643898 275153 644134
rect 280848 644218 281084 644454
rect 280848 643898 281084 644134
rect 302917 644218 303153 644454
rect 302917 643898 303153 644134
rect 308848 644218 309084 644454
rect 308848 643898 309084 644134
rect 330917 644218 331153 644454
rect 330917 643898 331153 644134
rect 336848 644218 337084 644454
rect 336848 643898 337084 644134
rect 358917 644218 359153 644454
rect 358917 643898 359153 644134
rect 364848 644218 365084 644454
rect 364848 643898 365084 644134
rect 386917 644218 387153 644454
rect 386917 643898 387153 644134
rect 392848 644218 393084 644454
rect 392848 643898 393084 644134
rect 414917 644218 415153 644454
rect 414917 643898 415153 644134
rect 420848 644218 421084 644454
rect 420848 643898 421084 644134
rect 442917 644218 443153 644454
rect 442917 643898 443153 644134
rect 448848 644218 449084 644454
rect 448848 643898 449084 644134
rect 470917 644218 471153 644454
rect 470917 643898 471153 644134
rect 476848 644218 477084 644454
rect 476848 643898 477084 644134
rect 498917 644218 499153 644454
rect 498917 643898 499153 644134
rect 504848 644218 505084 644454
rect 504848 643898 505084 644134
rect 526917 644218 527153 644454
rect 526917 643898 527153 644134
rect 532848 644218 533084 644454
rect 532848 643898 533084 644134
rect 554917 644218 555153 644454
rect 554917 643898 555153 644134
rect 560848 644218 561084 644454
rect 560848 643898 561084 644134
rect -1974 620593 -1738 620829
rect -1654 620593 -1418 620829
rect -1974 620273 -1738 620509
rect -1654 620273 -1418 620509
rect 19952 620593 20188 620829
rect 19952 620273 20188 620509
rect 25882 620593 26118 620829
rect 25882 620273 26118 620509
rect 31813 620593 32049 620829
rect 31813 620273 32049 620509
rect 47952 620593 48188 620829
rect 47952 620273 48188 620509
rect 53882 620593 54118 620829
rect 53882 620273 54118 620509
rect 59813 620593 60049 620829
rect 59813 620273 60049 620509
rect 75952 620593 76188 620829
rect 75952 620273 76188 620509
rect 81882 620593 82118 620829
rect 81882 620273 82118 620509
rect 87813 620593 88049 620829
rect 87813 620273 88049 620509
rect 103952 620593 104188 620829
rect 103952 620273 104188 620509
rect 109882 620593 110118 620829
rect 109882 620273 110118 620509
rect 115813 620593 116049 620829
rect 115813 620273 116049 620509
rect 131952 620593 132188 620829
rect 131952 620273 132188 620509
rect 137882 620593 138118 620829
rect 137882 620273 138118 620509
rect 143813 620593 144049 620829
rect 143813 620273 144049 620509
rect 159952 620593 160188 620829
rect 159952 620273 160188 620509
rect 165882 620593 166118 620829
rect 165882 620273 166118 620509
rect 171813 620593 172049 620829
rect 171813 620273 172049 620509
rect 187952 620593 188188 620829
rect 187952 620273 188188 620509
rect 193882 620593 194118 620829
rect 193882 620273 194118 620509
rect 199813 620593 200049 620829
rect 199813 620273 200049 620509
rect 215952 620593 216188 620829
rect 215952 620273 216188 620509
rect 221882 620593 222118 620829
rect 221882 620273 222118 620509
rect 227813 620593 228049 620829
rect 227813 620273 228049 620509
rect 243952 620593 244188 620829
rect 243952 620273 244188 620509
rect 249882 620593 250118 620829
rect 249882 620273 250118 620509
rect 255813 620593 256049 620829
rect 255813 620273 256049 620509
rect 271952 620593 272188 620829
rect 271952 620273 272188 620509
rect 277882 620593 278118 620829
rect 277882 620273 278118 620509
rect 283813 620593 284049 620829
rect 283813 620273 284049 620509
rect 299952 620593 300188 620829
rect 299952 620273 300188 620509
rect 305882 620593 306118 620829
rect 305882 620273 306118 620509
rect 311813 620593 312049 620829
rect 311813 620273 312049 620509
rect 327952 620593 328188 620829
rect 327952 620273 328188 620509
rect 333882 620593 334118 620829
rect 333882 620273 334118 620509
rect 339813 620593 340049 620829
rect 339813 620273 340049 620509
rect 355952 620593 356188 620829
rect 355952 620273 356188 620509
rect 361882 620593 362118 620829
rect 361882 620273 362118 620509
rect 367813 620593 368049 620829
rect 367813 620273 368049 620509
rect 383952 620593 384188 620829
rect 383952 620273 384188 620509
rect 389882 620593 390118 620829
rect 389882 620273 390118 620509
rect 395813 620593 396049 620829
rect 395813 620273 396049 620509
rect 411952 620593 412188 620829
rect 411952 620273 412188 620509
rect 417882 620593 418118 620829
rect 417882 620273 418118 620509
rect 423813 620593 424049 620829
rect 423813 620273 424049 620509
rect 439952 620593 440188 620829
rect 439952 620273 440188 620509
rect 445882 620593 446118 620829
rect 445882 620273 446118 620509
rect 451813 620593 452049 620829
rect 451813 620273 452049 620509
rect 467952 620593 468188 620829
rect 467952 620273 468188 620509
rect 473882 620593 474118 620829
rect 473882 620273 474118 620509
rect 479813 620593 480049 620829
rect 479813 620273 480049 620509
rect 495952 620593 496188 620829
rect 495952 620273 496188 620509
rect 501882 620593 502118 620829
rect 501882 620273 502118 620509
rect 507813 620593 508049 620829
rect 507813 620273 508049 620509
rect 523952 620593 524188 620829
rect 523952 620273 524188 620509
rect 529882 620593 530118 620829
rect 529882 620273 530118 620509
rect 535813 620593 536049 620829
rect 535813 620273 536049 620509
rect 551952 620593 552188 620829
rect 551952 620273 552188 620509
rect 557882 620593 558118 620829
rect 557882 620273 558118 620509
rect 563813 620593 564049 620829
rect 563813 620273 564049 620509
rect 573526 620593 573762 620829
rect 573846 620593 574082 620829
rect 573526 620273 573762 620509
rect 573846 620273 574082 620509
rect 22916 617218 23152 617454
rect 22916 616898 23152 617134
rect 28847 617218 29083 617454
rect 28847 616898 29083 617134
rect 50916 617218 51152 617454
rect 50916 616898 51152 617134
rect 56847 617218 57083 617454
rect 56847 616898 57083 617134
rect 78916 617218 79152 617454
rect 78916 616898 79152 617134
rect 84847 617218 85083 617454
rect 84847 616898 85083 617134
rect 106916 617218 107152 617454
rect 106916 616898 107152 617134
rect 112847 617218 113083 617454
rect 112847 616898 113083 617134
rect 134916 617218 135152 617454
rect 134916 616898 135152 617134
rect 140847 617218 141083 617454
rect 140847 616898 141083 617134
rect 162916 617218 163152 617454
rect 162916 616898 163152 617134
rect 168847 617218 169083 617454
rect 168847 616898 169083 617134
rect 190916 617218 191152 617454
rect 190916 616898 191152 617134
rect 196847 617218 197083 617454
rect 196847 616898 197083 617134
rect 218916 617218 219152 617454
rect 218916 616898 219152 617134
rect 224847 617218 225083 617454
rect 224847 616898 225083 617134
rect 246916 617218 247152 617454
rect 246916 616898 247152 617134
rect 252847 617218 253083 617454
rect 252847 616898 253083 617134
rect 274916 617218 275152 617454
rect 274916 616898 275152 617134
rect 280847 617218 281083 617454
rect 280847 616898 281083 617134
rect 302916 617218 303152 617454
rect 302916 616898 303152 617134
rect 308847 617218 309083 617454
rect 308847 616898 309083 617134
rect 330916 617218 331152 617454
rect 330916 616898 331152 617134
rect 336847 617218 337083 617454
rect 336847 616898 337083 617134
rect 358916 617218 359152 617454
rect 358916 616898 359152 617134
rect 364847 617218 365083 617454
rect 364847 616898 365083 617134
rect 386916 617218 387152 617454
rect 386916 616898 387152 617134
rect 392847 617218 393083 617454
rect 392847 616898 393083 617134
rect 414916 617218 415152 617454
rect 414916 616898 415152 617134
rect 420847 617218 421083 617454
rect 420847 616898 421083 617134
rect 442916 617218 443152 617454
rect 442916 616898 443152 617134
rect 448847 617218 449083 617454
rect 448847 616898 449083 617134
rect 470916 617218 471152 617454
rect 470916 616898 471152 617134
rect 476847 617218 477083 617454
rect 476847 616898 477083 617134
rect 498916 617218 499152 617454
rect 498916 616898 499152 617134
rect 504847 617218 505083 617454
rect 504847 616898 505083 617134
rect 526916 617218 527152 617454
rect 526916 616898 527152 617134
rect 532847 617218 533083 617454
rect 532847 616898 533083 617134
rect 554916 617218 555152 617454
rect 554916 616898 555152 617134
rect 560847 617218 561083 617454
rect 560847 616898 561083 617134
rect -1974 593593 -1738 593829
rect -1654 593593 -1418 593829
rect -1974 593273 -1738 593509
rect -1654 593273 -1418 593509
rect 19951 593593 20187 593829
rect 19951 593273 20187 593509
rect 25882 593593 26118 593829
rect 25882 593273 26118 593509
rect 31812 593593 32048 593829
rect 31812 593273 32048 593509
rect 47951 593593 48187 593829
rect 47951 593273 48187 593509
rect 53882 593593 54118 593829
rect 53882 593273 54118 593509
rect 59812 593593 60048 593829
rect 59812 593273 60048 593509
rect 75951 593593 76187 593829
rect 75951 593273 76187 593509
rect 81882 593593 82118 593829
rect 81882 593273 82118 593509
rect 87812 593593 88048 593829
rect 87812 593273 88048 593509
rect 103951 593593 104187 593829
rect 103951 593273 104187 593509
rect 109882 593593 110118 593829
rect 109882 593273 110118 593509
rect 115812 593593 116048 593829
rect 115812 593273 116048 593509
rect 131951 593593 132187 593829
rect 131951 593273 132187 593509
rect 137882 593593 138118 593829
rect 137882 593273 138118 593509
rect 143812 593593 144048 593829
rect 143812 593273 144048 593509
rect 159951 593593 160187 593829
rect 159951 593273 160187 593509
rect 165882 593593 166118 593829
rect 165882 593273 166118 593509
rect 171812 593593 172048 593829
rect 171812 593273 172048 593509
rect 187951 593593 188187 593829
rect 187951 593273 188187 593509
rect 193882 593593 194118 593829
rect 193882 593273 194118 593509
rect 199812 593593 200048 593829
rect 199812 593273 200048 593509
rect 215951 593593 216187 593829
rect 215951 593273 216187 593509
rect 221882 593593 222118 593829
rect 221882 593273 222118 593509
rect 227812 593593 228048 593829
rect 227812 593273 228048 593509
rect 243951 593593 244187 593829
rect 243951 593273 244187 593509
rect 249882 593593 250118 593829
rect 249882 593273 250118 593509
rect 255812 593593 256048 593829
rect 255812 593273 256048 593509
rect 271951 593593 272187 593829
rect 271951 593273 272187 593509
rect 277882 593593 278118 593829
rect 277882 593273 278118 593509
rect 283812 593593 284048 593829
rect 283812 593273 284048 593509
rect 299951 593593 300187 593829
rect 299951 593273 300187 593509
rect 305882 593593 306118 593829
rect 305882 593273 306118 593509
rect 311812 593593 312048 593829
rect 311812 593273 312048 593509
rect 327951 593593 328187 593829
rect 327951 593273 328187 593509
rect 333882 593593 334118 593829
rect 333882 593273 334118 593509
rect 339812 593593 340048 593829
rect 339812 593273 340048 593509
rect 355951 593593 356187 593829
rect 355951 593273 356187 593509
rect 361882 593593 362118 593829
rect 361882 593273 362118 593509
rect 367812 593593 368048 593829
rect 367812 593273 368048 593509
rect 383951 593593 384187 593829
rect 383951 593273 384187 593509
rect 389882 593593 390118 593829
rect 389882 593273 390118 593509
rect 395812 593593 396048 593829
rect 395812 593273 396048 593509
rect 411951 593593 412187 593829
rect 411951 593273 412187 593509
rect 417882 593593 418118 593829
rect 417882 593273 418118 593509
rect 423812 593593 424048 593829
rect 423812 593273 424048 593509
rect 439951 593593 440187 593829
rect 439951 593273 440187 593509
rect 445882 593593 446118 593829
rect 445882 593273 446118 593509
rect 451812 593593 452048 593829
rect 451812 593273 452048 593509
rect 467951 593593 468187 593829
rect 467951 593273 468187 593509
rect 473882 593593 474118 593829
rect 473882 593273 474118 593509
rect 479812 593593 480048 593829
rect 479812 593273 480048 593509
rect 495951 593593 496187 593829
rect 495951 593273 496187 593509
rect 501882 593593 502118 593829
rect 501882 593273 502118 593509
rect 507812 593593 508048 593829
rect 507812 593273 508048 593509
rect 523951 593593 524187 593829
rect 523951 593273 524187 593509
rect 529882 593593 530118 593829
rect 529882 593273 530118 593509
rect 535812 593593 536048 593829
rect 535812 593273 536048 593509
rect 551951 593593 552187 593829
rect 551951 593273 552187 593509
rect 557882 593593 558118 593829
rect 557882 593273 558118 593509
rect 563812 593593 564048 593829
rect 563812 593273 564048 593509
rect 573526 593593 573762 593829
rect 573846 593593 574082 593829
rect 573526 593273 573762 593509
rect 573846 593273 574082 593509
rect 22917 590218 23153 590454
rect 22917 589898 23153 590134
rect 28848 590218 29084 590454
rect 28848 589898 29084 590134
rect 50917 590218 51153 590454
rect 50917 589898 51153 590134
rect 56848 590218 57084 590454
rect 56848 589898 57084 590134
rect 78917 590218 79153 590454
rect 78917 589898 79153 590134
rect 84848 590218 85084 590454
rect 84848 589898 85084 590134
rect 106917 590218 107153 590454
rect 106917 589898 107153 590134
rect 112848 590218 113084 590454
rect 112848 589898 113084 590134
rect 134917 590218 135153 590454
rect 134917 589898 135153 590134
rect 140848 590218 141084 590454
rect 140848 589898 141084 590134
rect 162917 590218 163153 590454
rect 162917 589898 163153 590134
rect 168848 590218 169084 590454
rect 168848 589898 169084 590134
rect 190917 590218 191153 590454
rect 190917 589898 191153 590134
rect 196848 590218 197084 590454
rect 196848 589898 197084 590134
rect 218917 590218 219153 590454
rect 218917 589898 219153 590134
rect 224848 590218 225084 590454
rect 224848 589898 225084 590134
rect 246917 590218 247153 590454
rect 246917 589898 247153 590134
rect 252848 590218 253084 590454
rect 252848 589898 253084 590134
rect 274917 590218 275153 590454
rect 274917 589898 275153 590134
rect 280848 590218 281084 590454
rect 280848 589898 281084 590134
rect 302917 590218 303153 590454
rect 302917 589898 303153 590134
rect 308848 590218 309084 590454
rect 308848 589898 309084 590134
rect 330917 590218 331153 590454
rect 330917 589898 331153 590134
rect 336848 590218 337084 590454
rect 336848 589898 337084 590134
rect 358917 590218 359153 590454
rect 358917 589898 359153 590134
rect 364848 590218 365084 590454
rect 364848 589898 365084 590134
rect 386917 590218 387153 590454
rect 386917 589898 387153 590134
rect 392848 590218 393084 590454
rect 392848 589898 393084 590134
rect 414917 590218 415153 590454
rect 414917 589898 415153 590134
rect 420848 590218 421084 590454
rect 420848 589898 421084 590134
rect 442917 590218 443153 590454
rect 442917 589898 443153 590134
rect 448848 590218 449084 590454
rect 448848 589898 449084 590134
rect 470917 590218 471153 590454
rect 470917 589898 471153 590134
rect 476848 590218 477084 590454
rect 476848 589898 477084 590134
rect 498917 590218 499153 590454
rect 498917 589898 499153 590134
rect 504848 590218 505084 590454
rect 504848 589898 505084 590134
rect 526917 590218 527153 590454
rect 526917 589898 527153 590134
rect 532848 590218 533084 590454
rect 532848 589898 533084 590134
rect 554917 590218 555153 590454
rect 554917 589898 555153 590134
rect 560848 590218 561084 590454
rect 560848 589898 561084 590134
rect -1974 566593 -1738 566829
rect -1654 566593 -1418 566829
rect -1974 566273 -1738 566509
rect -1654 566273 -1418 566509
rect 19952 566593 20188 566829
rect 19952 566273 20188 566509
rect 25882 566593 26118 566829
rect 25882 566273 26118 566509
rect 31813 566593 32049 566829
rect 31813 566273 32049 566509
rect 47952 566593 48188 566829
rect 47952 566273 48188 566509
rect 53882 566593 54118 566829
rect 53882 566273 54118 566509
rect 59813 566593 60049 566829
rect 59813 566273 60049 566509
rect 75952 566593 76188 566829
rect 75952 566273 76188 566509
rect 81882 566593 82118 566829
rect 81882 566273 82118 566509
rect 87813 566593 88049 566829
rect 87813 566273 88049 566509
rect 103952 566593 104188 566829
rect 103952 566273 104188 566509
rect 109882 566593 110118 566829
rect 109882 566273 110118 566509
rect 115813 566593 116049 566829
rect 115813 566273 116049 566509
rect 131952 566593 132188 566829
rect 131952 566273 132188 566509
rect 137882 566593 138118 566829
rect 137882 566273 138118 566509
rect 143813 566593 144049 566829
rect 143813 566273 144049 566509
rect 159952 566593 160188 566829
rect 159952 566273 160188 566509
rect 165882 566593 166118 566829
rect 165882 566273 166118 566509
rect 171813 566593 172049 566829
rect 171813 566273 172049 566509
rect 187952 566593 188188 566829
rect 187952 566273 188188 566509
rect 193882 566593 194118 566829
rect 193882 566273 194118 566509
rect 199813 566593 200049 566829
rect 199813 566273 200049 566509
rect 215952 566593 216188 566829
rect 215952 566273 216188 566509
rect 221882 566593 222118 566829
rect 221882 566273 222118 566509
rect 227813 566593 228049 566829
rect 227813 566273 228049 566509
rect 243952 566593 244188 566829
rect 243952 566273 244188 566509
rect 249882 566593 250118 566829
rect 249882 566273 250118 566509
rect 255813 566593 256049 566829
rect 255813 566273 256049 566509
rect 271952 566593 272188 566829
rect 271952 566273 272188 566509
rect 277882 566593 278118 566829
rect 277882 566273 278118 566509
rect 283813 566593 284049 566829
rect 283813 566273 284049 566509
rect 299952 566593 300188 566829
rect 299952 566273 300188 566509
rect 305882 566593 306118 566829
rect 305882 566273 306118 566509
rect 311813 566593 312049 566829
rect 311813 566273 312049 566509
rect 327952 566593 328188 566829
rect 327952 566273 328188 566509
rect 333882 566593 334118 566829
rect 333882 566273 334118 566509
rect 339813 566593 340049 566829
rect 339813 566273 340049 566509
rect 355952 566593 356188 566829
rect 355952 566273 356188 566509
rect 361882 566593 362118 566829
rect 361882 566273 362118 566509
rect 367813 566593 368049 566829
rect 367813 566273 368049 566509
rect 383952 566593 384188 566829
rect 383952 566273 384188 566509
rect 389882 566593 390118 566829
rect 389882 566273 390118 566509
rect 395813 566593 396049 566829
rect 395813 566273 396049 566509
rect 411952 566593 412188 566829
rect 411952 566273 412188 566509
rect 417882 566593 418118 566829
rect 417882 566273 418118 566509
rect 423813 566593 424049 566829
rect 423813 566273 424049 566509
rect 439952 566593 440188 566829
rect 439952 566273 440188 566509
rect 445882 566593 446118 566829
rect 445882 566273 446118 566509
rect 451813 566593 452049 566829
rect 451813 566273 452049 566509
rect 467952 566593 468188 566829
rect 467952 566273 468188 566509
rect 473882 566593 474118 566829
rect 473882 566273 474118 566509
rect 479813 566593 480049 566829
rect 479813 566273 480049 566509
rect 495952 566593 496188 566829
rect 495952 566273 496188 566509
rect 501882 566593 502118 566829
rect 501882 566273 502118 566509
rect 507813 566593 508049 566829
rect 507813 566273 508049 566509
rect 523952 566593 524188 566829
rect 523952 566273 524188 566509
rect 529882 566593 530118 566829
rect 529882 566273 530118 566509
rect 535813 566593 536049 566829
rect 535813 566273 536049 566509
rect 551952 566593 552188 566829
rect 551952 566273 552188 566509
rect 557882 566593 558118 566829
rect 557882 566273 558118 566509
rect 563813 566593 564049 566829
rect 563813 566273 564049 566509
rect 573526 566593 573762 566829
rect 573846 566593 574082 566829
rect 573526 566273 573762 566509
rect 573846 566273 574082 566509
rect 22916 563218 23152 563454
rect 22916 562898 23152 563134
rect 28847 563218 29083 563454
rect 28847 562898 29083 563134
rect 50916 563218 51152 563454
rect 50916 562898 51152 563134
rect 56847 563218 57083 563454
rect 56847 562898 57083 563134
rect 78916 563218 79152 563454
rect 78916 562898 79152 563134
rect 84847 563218 85083 563454
rect 84847 562898 85083 563134
rect 106916 563218 107152 563454
rect 106916 562898 107152 563134
rect 112847 563218 113083 563454
rect 112847 562898 113083 563134
rect 134916 563218 135152 563454
rect 134916 562898 135152 563134
rect 140847 563218 141083 563454
rect 140847 562898 141083 563134
rect 162916 563218 163152 563454
rect 162916 562898 163152 563134
rect 168847 563218 169083 563454
rect 168847 562898 169083 563134
rect 190916 563218 191152 563454
rect 190916 562898 191152 563134
rect 196847 563218 197083 563454
rect 196847 562898 197083 563134
rect 218916 563218 219152 563454
rect 218916 562898 219152 563134
rect 224847 563218 225083 563454
rect 224847 562898 225083 563134
rect 246916 563218 247152 563454
rect 246916 562898 247152 563134
rect 252847 563218 253083 563454
rect 252847 562898 253083 563134
rect 274916 563218 275152 563454
rect 274916 562898 275152 563134
rect 280847 563218 281083 563454
rect 280847 562898 281083 563134
rect 302916 563218 303152 563454
rect 302916 562898 303152 563134
rect 308847 563218 309083 563454
rect 308847 562898 309083 563134
rect 330916 563218 331152 563454
rect 330916 562898 331152 563134
rect 336847 563218 337083 563454
rect 336847 562898 337083 563134
rect 358916 563218 359152 563454
rect 358916 562898 359152 563134
rect 364847 563218 365083 563454
rect 364847 562898 365083 563134
rect 386916 563218 387152 563454
rect 386916 562898 387152 563134
rect 392847 563218 393083 563454
rect 392847 562898 393083 563134
rect 414916 563218 415152 563454
rect 414916 562898 415152 563134
rect 420847 563218 421083 563454
rect 420847 562898 421083 563134
rect 442916 563218 443152 563454
rect 442916 562898 443152 563134
rect 448847 563218 449083 563454
rect 448847 562898 449083 563134
rect 470916 563218 471152 563454
rect 470916 562898 471152 563134
rect 476847 563218 477083 563454
rect 476847 562898 477083 563134
rect 498916 563218 499152 563454
rect 498916 562898 499152 563134
rect 504847 563218 505083 563454
rect 504847 562898 505083 563134
rect 526916 563218 527152 563454
rect 526916 562898 527152 563134
rect 532847 563218 533083 563454
rect 532847 562898 533083 563134
rect 554916 563218 555152 563454
rect 554916 562898 555152 563134
rect 560847 563218 561083 563454
rect 560847 562898 561083 563134
rect -1974 539593 -1738 539829
rect -1654 539593 -1418 539829
rect -1974 539273 -1738 539509
rect -1654 539273 -1418 539509
rect 19951 539593 20187 539829
rect 19951 539273 20187 539509
rect 25882 539593 26118 539829
rect 25882 539273 26118 539509
rect 31812 539593 32048 539829
rect 31812 539273 32048 539509
rect 47951 539593 48187 539829
rect 47951 539273 48187 539509
rect 53882 539593 54118 539829
rect 53882 539273 54118 539509
rect 59812 539593 60048 539829
rect 59812 539273 60048 539509
rect 75951 539593 76187 539829
rect 75951 539273 76187 539509
rect 81882 539593 82118 539829
rect 81882 539273 82118 539509
rect 87812 539593 88048 539829
rect 87812 539273 88048 539509
rect 103951 539593 104187 539829
rect 103951 539273 104187 539509
rect 109882 539593 110118 539829
rect 109882 539273 110118 539509
rect 115812 539593 116048 539829
rect 115812 539273 116048 539509
rect 131951 539593 132187 539829
rect 131951 539273 132187 539509
rect 137882 539593 138118 539829
rect 137882 539273 138118 539509
rect 143812 539593 144048 539829
rect 143812 539273 144048 539509
rect 159951 539593 160187 539829
rect 159951 539273 160187 539509
rect 165882 539593 166118 539829
rect 165882 539273 166118 539509
rect 171812 539593 172048 539829
rect 171812 539273 172048 539509
rect 187951 539593 188187 539829
rect 187951 539273 188187 539509
rect 193882 539593 194118 539829
rect 193882 539273 194118 539509
rect 199812 539593 200048 539829
rect 199812 539273 200048 539509
rect 215951 539593 216187 539829
rect 215951 539273 216187 539509
rect 221882 539593 222118 539829
rect 221882 539273 222118 539509
rect 227812 539593 228048 539829
rect 227812 539273 228048 539509
rect 243951 539593 244187 539829
rect 243951 539273 244187 539509
rect 249882 539593 250118 539829
rect 249882 539273 250118 539509
rect 255812 539593 256048 539829
rect 255812 539273 256048 539509
rect 271951 539593 272187 539829
rect 271951 539273 272187 539509
rect 277882 539593 278118 539829
rect 277882 539273 278118 539509
rect 283812 539593 284048 539829
rect 283812 539273 284048 539509
rect 299951 539593 300187 539829
rect 299951 539273 300187 539509
rect 305882 539593 306118 539829
rect 305882 539273 306118 539509
rect 311812 539593 312048 539829
rect 311812 539273 312048 539509
rect 327951 539593 328187 539829
rect 327951 539273 328187 539509
rect 333882 539593 334118 539829
rect 333882 539273 334118 539509
rect 339812 539593 340048 539829
rect 339812 539273 340048 539509
rect 355951 539593 356187 539829
rect 355951 539273 356187 539509
rect 361882 539593 362118 539829
rect 361882 539273 362118 539509
rect 367812 539593 368048 539829
rect 367812 539273 368048 539509
rect 383951 539593 384187 539829
rect 383951 539273 384187 539509
rect 389882 539593 390118 539829
rect 389882 539273 390118 539509
rect 395812 539593 396048 539829
rect 395812 539273 396048 539509
rect 411951 539593 412187 539829
rect 411951 539273 412187 539509
rect 417882 539593 418118 539829
rect 417882 539273 418118 539509
rect 423812 539593 424048 539829
rect 423812 539273 424048 539509
rect 439951 539593 440187 539829
rect 439951 539273 440187 539509
rect 445882 539593 446118 539829
rect 445882 539273 446118 539509
rect 451812 539593 452048 539829
rect 451812 539273 452048 539509
rect 467951 539593 468187 539829
rect 467951 539273 468187 539509
rect 473882 539593 474118 539829
rect 473882 539273 474118 539509
rect 479812 539593 480048 539829
rect 479812 539273 480048 539509
rect 495951 539593 496187 539829
rect 495951 539273 496187 539509
rect 501882 539593 502118 539829
rect 501882 539273 502118 539509
rect 507812 539593 508048 539829
rect 507812 539273 508048 539509
rect 523951 539593 524187 539829
rect 523951 539273 524187 539509
rect 529882 539593 530118 539829
rect 529882 539273 530118 539509
rect 535812 539593 536048 539829
rect 535812 539273 536048 539509
rect 551951 539593 552187 539829
rect 551951 539273 552187 539509
rect 557882 539593 558118 539829
rect 557882 539273 558118 539509
rect 563812 539593 564048 539829
rect 563812 539273 564048 539509
rect 573526 539593 573762 539829
rect 573846 539593 574082 539829
rect 573526 539273 573762 539509
rect 573846 539273 574082 539509
rect 22917 536218 23153 536454
rect 22917 535898 23153 536134
rect 28848 536218 29084 536454
rect 28848 535898 29084 536134
rect 50917 536218 51153 536454
rect 50917 535898 51153 536134
rect 56848 536218 57084 536454
rect 56848 535898 57084 536134
rect 78917 536218 79153 536454
rect 78917 535898 79153 536134
rect 84848 536218 85084 536454
rect 84848 535898 85084 536134
rect 106917 536218 107153 536454
rect 106917 535898 107153 536134
rect 112848 536218 113084 536454
rect 112848 535898 113084 536134
rect 134917 536218 135153 536454
rect 134917 535898 135153 536134
rect 140848 536218 141084 536454
rect 140848 535898 141084 536134
rect 162917 536218 163153 536454
rect 162917 535898 163153 536134
rect 168848 536218 169084 536454
rect 168848 535898 169084 536134
rect 190917 536218 191153 536454
rect 190917 535898 191153 536134
rect 196848 536218 197084 536454
rect 196848 535898 197084 536134
rect 218917 536218 219153 536454
rect 218917 535898 219153 536134
rect 224848 536218 225084 536454
rect 224848 535898 225084 536134
rect 246917 536218 247153 536454
rect 246917 535898 247153 536134
rect 252848 536218 253084 536454
rect 252848 535898 253084 536134
rect 274917 536218 275153 536454
rect 274917 535898 275153 536134
rect 280848 536218 281084 536454
rect 280848 535898 281084 536134
rect 302917 536218 303153 536454
rect 302917 535898 303153 536134
rect 308848 536218 309084 536454
rect 308848 535898 309084 536134
rect 330917 536218 331153 536454
rect 330917 535898 331153 536134
rect 336848 536218 337084 536454
rect 336848 535898 337084 536134
rect 358917 536218 359153 536454
rect 358917 535898 359153 536134
rect 364848 536218 365084 536454
rect 364848 535898 365084 536134
rect 386917 536218 387153 536454
rect 386917 535898 387153 536134
rect 392848 536218 393084 536454
rect 392848 535898 393084 536134
rect 414917 536218 415153 536454
rect 414917 535898 415153 536134
rect 420848 536218 421084 536454
rect 420848 535898 421084 536134
rect 442917 536218 443153 536454
rect 442917 535898 443153 536134
rect 448848 536218 449084 536454
rect 448848 535898 449084 536134
rect 470917 536218 471153 536454
rect 470917 535898 471153 536134
rect 476848 536218 477084 536454
rect 476848 535898 477084 536134
rect 498917 536218 499153 536454
rect 498917 535898 499153 536134
rect 504848 536218 505084 536454
rect 504848 535898 505084 536134
rect 526917 536218 527153 536454
rect 526917 535898 527153 536134
rect 532848 536218 533084 536454
rect 532848 535898 533084 536134
rect 554917 536218 555153 536454
rect 554917 535898 555153 536134
rect 560848 536218 561084 536454
rect 560848 535898 561084 536134
rect -1974 512593 -1738 512829
rect -1654 512593 -1418 512829
rect -1974 512273 -1738 512509
rect -1654 512273 -1418 512509
rect 19952 512593 20188 512829
rect 19952 512273 20188 512509
rect 25882 512593 26118 512829
rect 25882 512273 26118 512509
rect 31813 512593 32049 512829
rect 31813 512273 32049 512509
rect 47952 512593 48188 512829
rect 47952 512273 48188 512509
rect 53882 512593 54118 512829
rect 53882 512273 54118 512509
rect 59813 512593 60049 512829
rect 59813 512273 60049 512509
rect 75952 512593 76188 512829
rect 75952 512273 76188 512509
rect 81882 512593 82118 512829
rect 81882 512273 82118 512509
rect 87813 512593 88049 512829
rect 87813 512273 88049 512509
rect 103952 512593 104188 512829
rect 103952 512273 104188 512509
rect 109882 512593 110118 512829
rect 109882 512273 110118 512509
rect 115813 512593 116049 512829
rect 115813 512273 116049 512509
rect 131952 512593 132188 512829
rect 131952 512273 132188 512509
rect 137882 512593 138118 512829
rect 137882 512273 138118 512509
rect 143813 512593 144049 512829
rect 143813 512273 144049 512509
rect 159952 512593 160188 512829
rect 159952 512273 160188 512509
rect 165882 512593 166118 512829
rect 165882 512273 166118 512509
rect 171813 512593 172049 512829
rect 171813 512273 172049 512509
rect 187952 512593 188188 512829
rect 187952 512273 188188 512509
rect 193882 512593 194118 512829
rect 193882 512273 194118 512509
rect 199813 512593 200049 512829
rect 199813 512273 200049 512509
rect 215952 512593 216188 512829
rect 215952 512273 216188 512509
rect 221882 512593 222118 512829
rect 221882 512273 222118 512509
rect 227813 512593 228049 512829
rect 227813 512273 228049 512509
rect 243952 512593 244188 512829
rect 243952 512273 244188 512509
rect 249882 512593 250118 512829
rect 249882 512273 250118 512509
rect 255813 512593 256049 512829
rect 255813 512273 256049 512509
rect 271952 512593 272188 512829
rect 271952 512273 272188 512509
rect 277882 512593 278118 512829
rect 277882 512273 278118 512509
rect 283813 512593 284049 512829
rect 283813 512273 284049 512509
rect 299952 512593 300188 512829
rect 299952 512273 300188 512509
rect 305882 512593 306118 512829
rect 305882 512273 306118 512509
rect 311813 512593 312049 512829
rect 311813 512273 312049 512509
rect 327952 512593 328188 512829
rect 327952 512273 328188 512509
rect 333882 512593 334118 512829
rect 333882 512273 334118 512509
rect 339813 512593 340049 512829
rect 339813 512273 340049 512509
rect 355952 512593 356188 512829
rect 355952 512273 356188 512509
rect 361882 512593 362118 512829
rect 361882 512273 362118 512509
rect 367813 512593 368049 512829
rect 367813 512273 368049 512509
rect 383952 512593 384188 512829
rect 383952 512273 384188 512509
rect 389882 512593 390118 512829
rect 389882 512273 390118 512509
rect 395813 512593 396049 512829
rect 395813 512273 396049 512509
rect 411952 512593 412188 512829
rect 411952 512273 412188 512509
rect 417882 512593 418118 512829
rect 417882 512273 418118 512509
rect 423813 512593 424049 512829
rect 423813 512273 424049 512509
rect 439952 512593 440188 512829
rect 439952 512273 440188 512509
rect 445882 512593 446118 512829
rect 445882 512273 446118 512509
rect 451813 512593 452049 512829
rect 451813 512273 452049 512509
rect 467952 512593 468188 512829
rect 467952 512273 468188 512509
rect 473882 512593 474118 512829
rect 473882 512273 474118 512509
rect 479813 512593 480049 512829
rect 479813 512273 480049 512509
rect 495952 512593 496188 512829
rect 495952 512273 496188 512509
rect 501882 512593 502118 512829
rect 501882 512273 502118 512509
rect 507813 512593 508049 512829
rect 507813 512273 508049 512509
rect 523952 512593 524188 512829
rect 523952 512273 524188 512509
rect 529882 512593 530118 512829
rect 529882 512273 530118 512509
rect 535813 512593 536049 512829
rect 535813 512273 536049 512509
rect 551952 512593 552188 512829
rect 551952 512273 552188 512509
rect 557882 512593 558118 512829
rect 557882 512273 558118 512509
rect 563813 512593 564049 512829
rect 563813 512273 564049 512509
rect 573526 512593 573762 512829
rect 573846 512593 574082 512829
rect 573526 512273 573762 512509
rect 573846 512273 574082 512509
rect 22916 509218 23152 509454
rect 22916 508898 23152 509134
rect 28847 509218 29083 509454
rect 28847 508898 29083 509134
rect 50916 509218 51152 509454
rect 50916 508898 51152 509134
rect 56847 509218 57083 509454
rect 56847 508898 57083 509134
rect 78916 509218 79152 509454
rect 78916 508898 79152 509134
rect 84847 509218 85083 509454
rect 84847 508898 85083 509134
rect 106916 509218 107152 509454
rect 106916 508898 107152 509134
rect 112847 509218 113083 509454
rect 112847 508898 113083 509134
rect 134916 509218 135152 509454
rect 134916 508898 135152 509134
rect 140847 509218 141083 509454
rect 140847 508898 141083 509134
rect 162916 509218 163152 509454
rect 162916 508898 163152 509134
rect 168847 509218 169083 509454
rect 168847 508898 169083 509134
rect 190916 509218 191152 509454
rect 190916 508898 191152 509134
rect 196847 509218 197083 509454
rect 196847 508898 197083 509134
rect 218916 509218 219152 509454
rect 218916 508898 219152 509134
rect 224847 509218 225083 509454
rect 224847 508898 225083 509134
rect 246916 509218 247152 509454
rect 246916 508898 247152 509134
rect 252847 509218 253083 509454
rect 252847 508898 253083 509134
rect 274916 509218 275152 509454
rect 274916 508898 275152 509134
rect 280847 509218 281083 509454
rect 280847 508898 281083 509134
rect 302916 509218 303152 509454
rect 302916 508898 303152 509134
rect 308847 509218 309083 509454
rect 308847 508898 309083 509134
rect 330916 509218 331152 509454
rect 330916 508898 331152 509134
rect 336847 509218 337083 509454
rect 336847 508898 337083 509134
rect 358916 509218 359152 509454
rect 358916 508898 359152 509134
rect 364847 509218 365083 509454
rect 364847 508898 365083 509134
rect 386916 509218 387152 509454
rect 386916 508898 387152 509134
rect 392847 509218 393083 509454
rect 392847 508898 393083 509134
rect 414916 509218 415152 509454
rect 414916 508898 415152 509134
rect 420847 509218 421083 509454
rect 420847 508898 421083 509134
rect 442916 509218 443152 509454
rect 442916 508898 443152 509134
rect 448847 509218 449083 509454
rect 448847 508898 449083 509134
rect 470916 509218 471152 509454
rect 470916 508898 471152 509134
rect 476847 509218 477083 509454
rect 476847 508898 477083 509134
rect 498916 509218 499152 509454
rect 498916 508898 499152 509134
rect 504847 509218 505083 509454
rect 504847 508898 505083 509134
rect 526916 509218 527152 509454
rect 526916 508898 527152 509134
rect 532847 509218 533083 509454
rect 532847 508898 533083 509134
rect 554916 509218 555152 509454
rect 554916 508898 555152 509134
rect 560847 509218 561083 509454
rect 560847 508898 561083 509134
rect -1974 485593 -1738 485829
rect -1654 485593 -1418 485829
rect -1974 485273 -1738 485509
rect -1654 485273 -1418 485509
rect 19951 485593 20187 485829
rect 19951 485273 20187 485509
rect 25882 485593 26118 485829
rect 25882 485273 26118 485509
rect 31812 485593 32048 485829
rect 31812 485273 32048 485509
rect 47951 485593 48187 485829
rect 47951 485273 48187 485509
rect 53882 485593 54118 485829
rect 53882 485273 54118 485509
rect 59812 485593 60048 485829
rect 59812 485273 60048 485509
rect 75951 485593 76187 485829
rect 75951 485273 76187 485509
rect 81882 485593 82118 485829
rect 81882 485273 82118 485509
rect 87812 485593 88048 485829
rect 87812 485273 88048 485509
rect 103951 485593 104187 485829
rect 103951 485273 104187 485509
rect 109882 485593 110118 485829
rect 109882 485273 110118 485509
rect 115812 485593 116048 485829
rect 115812 485273 116048 485509
rect 131951 485593 132187 485829
rect 131951 485273 132187 485509
rect 137882 485593 138118 485829
rect 137882 485273 138118 485509
rect 143812 485593 144048 485829
rect 143812 485273 144048 485509
rect 159951 485593 160187 485829
rect 159951 485273 160187 485509
rect 165882 485593 166118 485829
rect 165882 485273 166118 485509
rect 171812 485593 172048 485829
rect 171812 485273 172048 485509
rect 187951 485593 188187 485829
rect 187951 485273 188187 485509
rect 193882 485593 194118 485829
rect 193882 485273 194118 485509
rect 199812 485593 200048 485829
rect 199812 485273 200048 485509
rect 215951 485593 216187 485829
rect 215951 485273 216187 485509
rect 221882 485593 222118 485829
rect 221882 485273 222118 485509
rect 227812 485593 228048 485829
rect 227812 485273 228048 485509
rect 243951 485593 244187 485829
rect 243951 485273 244187 485509
rect 249882 485593 250118 485829
rect 249882 485273 250118 485509
rect 255812 485593 256048 485829
rect 255812 485273 256048 485509
rect 271951 485593 272187 485829
rect 271951 485273 272187 485509
rect 277882 485593 278118 485829
rect 277882 485273 278118 485509
rect 283812 485593 284048 485829
rect 283812 485273 284048 485509
rect 299951 485593 300187 485829
rect 299951 485273 300187 485509
rect 305882 485593 306118 485829
rect 305882 485273 306118 485509
rect 311812 485593 312048 485829
rect 311812 485273 312048 485509
rect 327951 485593 328187 485829
rect 327951 485273 328187 485509
rect 333882 485593 334118 485829
rect 333882 485273 334118 485509
rect 339812 485593 340048 485829
rect 339812 485273 340048 485509
rect 355951 485593 356187 485829
rect 355951 485273 356187 485509
rect 361882 485593 362118 485829
rect 361882 485273 362118 485509
rect 367812 485593 368048 485829
rect 367812 485273 368048 485509
rect 383951 485593 384187 485829
rect 383951 485273 384187 485509
rect 389882 485593 390118 485829
rect 389882 485273 390118 485509
rect 395812 485593 396048 485829
rect 395812 485273 396048 485509
rect 411951 485593 412187 485829
rect 411951 485273 412187 485509
rect 417882 485593 418118 485829
rect 417882 485273 418118 485509
rect 423812 485593 424048 485829
rect 423812 485273 424048 485509
rect 439951 485593 440187 485829
rect 439951 485273 440187 485509
rect 445882 485593 446118 485829
rect 445882 485273 446118 485509
rect 451812 485593 452048 485829
rect 451812 485273 452048 485509
rect 467951 485593 468187 485829
rect 467951 485273 468187 485509
rect 473882 485593 474118 485829
rect 473882 485273 474118 485509
rect 479812 485593 480048 485829
rect 479812 485273 480048 485509
rect 495951 485593 496187 485829
rect 495951 485273 496187 485509
rect 501882 485593 502118 485829
rect 501882 485273 502118 485509
rect 507812 485593 508048 485829
rect 507812 485273 508048 485509
rect 523951 485593 524187 485829
rect 523951 485273 524187 485509
rect 529882 485593 530118 485829
rect 529882 485273 530118 485509
rect 535812 485593 536048 485829
rect 535812 485273 536048 485509
rect 551951 485593 552187 485829
rect 551951 485273 552187 485509
rect 557882 485593 558118 485829
rect 557882 485273 558118 485509
rect 563812 485593 564048 485829
rect 563812 485273 564048 485509
rect 573526 485593 573762 485829
rect 573846 485593 574082 485829
rect 573526 485273 573762 485509
rect 573846 485273 574082 485509
rect 22917 482218 23153 482454
rect 22917 481898 23153 482134
rect 28848 482218 29084 482454
rect 28848 481898 29084 482134
rect 50917 482218 51153 482454
rect 50917 481898 51153 482134
rect 56848 482218 57084 482454
rect 56848 481898 57084 482134
rect 78917 482218 79153 482454
rect 78917 481898 79153 482134
rect 84848 482218 85084 482454
rect 84848 481898 85084 482134
rect 106917 482218 107153 482454
rect 106917 481898 107153 482134
rect 112848 482218 113084 482454
rect 112848 481898 113084 482134
rect 134917 482218 135153 482454
rect 134917 481898 135153 482134
rect 140848 482218 141084 482454
rect 140848 481898 141084 482134
rect 162917 482218 163153 482454
rect 162917 481898 163153 482134
rect 168848 482218 169084 482454
rect 168848 481898 169084 482134
rect 190917 482218 191153 482454
rect 190917 481898 191153 482134
rect 196848 482218 197084 482454
rect 196848 481898 197084 482134
rect 218917 482218 219153 482454
rect 218917 481898 219153 482134
rect 224848 482218 225084 482454
rect 224848 481898 225084 482134
rect 246917 482218 247153 482454
rect 246917 481898 247153 482134
rect 252848 482218 253084 482454
rect 252848 481898 253084 482134
rect 274917 482218 275153 482454
rect 274917 481898 275153 482134
rect 280848 482218 281084 482454
rect 280848 481898 281084 482134
rect 302917 482218 303153 482454
rect 302917 481898 303153 482134
rect 308848 482218 309084 482454
rect 308848 481898 309084 482134
rect 330917 482218 331153 482454
rect 330917 481898 331153 482134
rect 336848 482218 337084 482454
rect 336848 481898 337084 482134
rect 358917 482218 359153 482454
rect 358917 481898 359153 482134
rect 364848 482218 365084 482454
rect 364848 481898 365084 482134
rect 386917 482218 387153 482454
rect 386917 481898 387153 482134
rect 392848 482218 393084 482454
rect 392848 481898 393084 482134
rect 414917 482218 415153 482454
rect 414917 481898 415153 482134
rect 420848 482218 421084 482454
rect 420848 481898 421084 482134
rect 442917 482218 443153 482454
rect 442917 481898 443153 482134
rect 448848 482218 449084 482454
rect 448848 481898 449084 482134
rect 470917 482218 471153 482454
rect 470917 481898 471153 482134
rect 476848 482218 477084 482454
rect 476848 481898 477084 482134
rect 498917 482218 499153 482454
rect 498917 481898 499153 482134
rect 504848 482218 505084 482454
rect 504848 481898 505084 482134
rect 526917 482218 527153 482454
rect 526917 481898 527153 482134
rect 532848 482218 533084 482454
rect 532848 481898 533084 482134
rect 554917 482218 555153 482454
rect 554917 481898 555153 482134
rect 560848 482218 561084 482454
rect 560848 481898 561084 482134
rect -1974 458593 -1738 458829
rect -1654 458593 -1418 458829
rect -1974 458273 -1738 458509
rect -1654 458273 -1418 458509
rect 19952 458593 20188 458829
rect 19952 458273 20188 458509
rect 25882 458593 26118 458829
rect 25882 458273 26118 458509
rect 31813 458593 32049 458829
rect 31813 458273 32049 458509
rect 47952 458593 48188 458829
rect 47952 458273 48188 458509
rect 53882 458593 54118 458829
rect 53882 458273 54118 458509
rect 59813 458593 60049 458829
rect 59813 458273 60049 458509
rect 75952 458593 76188 458829
rect 75952 458273 76188 458509
rect 81882 458593 82118 458829
rect 81882 458273 82118 458509
rect 87813 458593 88049 458829
rect 87813 458273 88049 458509
rect 103952 458593 104188 458829
rect 103952 458273 104188 458509
rect 109882 458593 110118 458829
rect 109882 458273 110118 458509
rect 115813 458593 116049 458829
rect 115813 458273 116049 458509
rect 131952 458593 132188 458829
rect 131952 458273 132188 458509
rect 137882 458593 138118 458829
rect 137882 458273 138118 458509
rect 143813 458593 144049 458829
rect 143813 458273 144049 458509
rect 159952 458593 160188 458829
rect 159952 458273 160188 458509
rect 165882 458593 166118 458829
rect 165882 458273 166118 458509
rect 171813 458593 172049 458829
rect 171813 458273 172049 458509
rect 187952 458593 188188 458829
rect 187952 458273 188188 458509
rect 193882 458593 194118 458829
rect 193882 458273 194118 458509
rect 199813 458593 200049 458829
rect 199813 458273 200049 458509
rect 215952 458593 216188 458829
rect 215952 458273 216188 458509
rect 221882 458593 222118 458829
rect 221882 458273 222118 458509
rect 227813 458593 228049 458829
rect 227813 458273 228049 458509
rect 243952 458593 244188 458829
rect 243952 458273 244188 458509
rect 249882 458593 250118 458829
rect 249882 458273 250118 458509
rect 255813 458593 256049 458829
rect 255813 458273 256049 458509
rect 271952 458593 272188 458829
rect 271952 458273 272188 458509
rect 277882 458593 278118 458829
rect 277882 458273 278118 458509
rect 283813 458593 284049 458829
rect 283813 458273 284049 458509
rect 299952 458593 300188 458829
rect 299952 458273 300188 458509
rect 305882 458593 306118 458829
rect 305882 458273 306118 458509
rect 311813 458593 312049 458829
rect 311813 458273 312049 458509
rect 327952 458593 328188 458829
rect 327952 458273 328188 458509
rect 333882 458593 334118 458829
rect 333882 458273 334118 458509
rect 339813 458593 340049 458829
rect 339813 458273 340049 458509
rect 355952 458593 356188 458829
rect 355952 458273 356188 458509
rect 361882 458593 362118 458829
rect 361882 458273 362118 458509
rect 367813 458593 368049 458829
rect 367813 458273 368049 458509
rect 383952 458593 384188 458829
rect 383952 458273 384188 458509
rect 389882 458593 390118 458829
rect 389882 458273 390118 458509
rect 395813 458593 396049 458829
rect 395813 458273 396049 458509
rect 411952 458593 412188 458829
rect 411952 458273 412188 458509
rect 417882 458593 418118 458829
rect 417882 458273 418118 458509
rect 423813 458593 424049 458829
rect 423813 458273 424049 458509
rect 439952 458593 440188 458829
rect 439952 458273 440188 458509
rect 445882 458593 446118 458829
rect 445882 458273 446118 458509
rect 451813 458593 452049 458829
rect 451813 458273 452049 458509
rect 467952 458593 468188 458829
rect 467952 458273 468188 458509
rect 473882 458593 474118 458829
rect 473882 458273 474118 458509
rect 479813 458593 480049 458829
rect 479813 458273 480049 458509
rect 495952 458593 496188 458829
rect 495952 458273 496188 458509
rect 501882 458593 502118 458829
rect 501882 458273 502118 458509
rect 507813 458593 508049 458829
rect 507813 458273 508049 458509
rect 523952 458593 524188 458829
rect 523952 458273 524188 458509
rect 529882 458593 530118 458829
rect 529882 458273 530118 458509
rect 535813 458593 536049 458829
rect 535813 458273 536049 458509
rect 551952 458593 552188 458829
rect 551952 458273 552188 458509
rect 557882 458593 558118 458829
rect 557882 458273 558118 458509
rect 563813 458593 564049 458829
rect 563813 458273 564049 458509
rect 573526 458593 573762 458829
rect 573846 458593 574082 458829
rect 573526 458273 573762 458509
rect 573846 458273 574082 458509
rect 22916 455218 23152 455454
rect 22916 454898 23152 455134
rect 28847 455218 29083 455454
rect 28847 454898 29083 455134
rect 50916 455218 51152 455454
rect 50916 454898 51152 455134
rect 56847 455218 57083 455454
rect 56847 454898 57083 455134
rect 78916 455218 79152 455454
rect 78916 454898 79152 455134
rect 84847 455218 85083 455454
rect 84847 454898 85083 455134
rect 106916 455218 107152 455454
rect 106916 454898 107152 455134
rect 112847 455218 113083 455454
rect 112847 454898 113083 455134
rect 134916 455218 135152 455454
rect 134916 454898 135152 455134
rect 140847 455218 141083 455454
rect 140847 454898 141083 455134
rect 162916 455218 163152 455454
rect 162916 454898 163152 455134
rect 168847 455218 169083 455454
rect 168847 454898 169083 455134
rect 190916 455218 191152 455454
rect 190916 454898 191152 455134
rect 196847 455218 197083 455454
rect 196847 454898 197083 455134
rect 218916 455218 219152 455454
rect 218916 454898 219152 455134
rect 224847 455218 225083 455454
rect 224847 454898 225083 455134
rect 246916 455218 247152 455454
rect 246916 454898 247152 455134
rect 252847 455218 253083 455454
rect 252847 454898 253083 455134
rect 274916 455218 275152 455454
rect 274916 454898 275152 455134
rect 280847 455218 281083 455454
rect 280847 454898 281083 455134
rect 302916 455218 303152 455454
rect 302916 454898 303152 455134
rect 308847 455218 309083 455454
rect 308847 454898 309083 455134
rect 330916 455218 331152 455454
rect 330916 454898 331152 455134
rect 336847 455218 337083 455454
rect 336847 454898 337083 455134
rect 358916 455218 359152 455454
rect 358916 454898 359152 455134
rect 364847 455218 365083 455454
rect 364847 454898 365083 455134
rect 386916 455218 387152 455454
rect 386916 454898 387152 455134
rect 392847 455218 393083 455454
rect 392847 454898 393083 455134
rect 414916 455218 415152 455454
rect 414916 454898 415152 455134
rect 420847 455218 421083 455454
rect 420847 454898 421083 455134
rect 442916 455218 443152 455454
rect 442916 454898 443152 455134
rect 448847 455218 449083 455454
rect 448847 454898 449083 455134
rect 470916 455218 471152 455454
rect 470916 454898 471152 455134
rect 476847 455218 477083 455454
rect 476847 454898 477083 455134
rect 498916 455218 499152 455454
rect 498916 454898 499152 455134
rect 504847 455218 505083 455454
rect 504847 454898 505083 455134
rect 526916 455218 527152 455454
rect 526916 454898 527152 455134
rect 532847 455218 533083 455454
rect 532847 454898 533083 455134
rect 554916 455218 555152 455454
rect 554916 454898 555152 455134
rect 560847 455218 561083 455454
rect 560847 454898 561083 455134
rect -1974 431593 -1738 431829
rect -1654 431593 -1418 431829
rect -1974 431273 -1738 431509
rect -1654 431273 -1418 431509
rect 19951 431593 20187 431829
rect 19951 431273 20187 431509
rect 25882 431593 26118 431829
rect 25882 431273 26118 431509
rect 31812 431593 32048 431829
rect 31812 431273 32048 431509
rect 47951 431593 48187 431829
rect 47951 431273 48187 431509
rect 53882 431593 54118 431829
rect 53882 431273 54118 431509
rect 59812 431593 60048 431829
rect 59812 431273 60048 431509
rect 75951 431593 76187 431829
rect 75951 431273 76187 431509
rect 81882 431593 82118 431829
rect 81882 431273 82118 431509
rect 87812 431593 88048 431829
rect 87812 431273 88048 431509
rect 103951 431593 104187 431829
rect 103951 431273 104187 431509
rect 109882 431593 110118 431829
rect 109882 431273 110118 431509
rect 115812 431593 116048 431829
rect 115812 431273 116048 431509
rect 131951 431593 132187 431829
rect 131951 431273 132187 431509
rect 137882 431593 138118 431829
rect 137882 431273 138118 431509
rect 143812 431593 144048 431829
rect 143812 431273 144048 431509
rect 159951 431593 160187 431829
rect 159951 431273 160187 431509
rect 165882 431593 166118 431829
rect 165882 431273 166118 431509
rect 171812 431593 172048 431829
rect 171812 431273 172048 431509
rect 187951 431593 188187 431829
rect 187951 431273 188187 431509
rect 193882 431593 194118 431829
rect 193882 431273 194118 431509
rect 199812 431593 200048 431829
rect 199812 431273 200048 431509
rect 215951 431593 216187 431829
rect 215951 431273 216187 431509
rect 221882 431593 222118 431829
rect 221882 431273 222118 431509
rect 227812 431593 228048 431829
rect 227812 431273 228048 431509
rect 243951 431593 244187 431829
rect 243951 431273 244187 431509
rect 249882 431593 250118 431829
rect 249882 431273 250118 431509
rect 255812 431593 256048 431829
rect 255812 431273 256048 431509
rect 271951 431593 272187 431829
rect 271951 431273 272187 431509
rect 277882 431593 278118 431829
rect 277882 431273 278118 431509
rect 283812 431593 284048 431829
rect 283812 431273 284048 431509
rect 299951 431593 300187 431829
rect 299951 431273 300187 431509
rect 305882 431593 306118 431829
rect 305882 431273 306118 431509
rect 311812 431593 312048 431829
rect 311812 431273 312048 431509
rect 327951 431593 328187 431829
rect 327951 431273 328187 431509
rect 333882 431593 334118 431829
rect 333882 431273 334118 431509
rect 339812 431593 340048 431829
rect 339812 431273 340048 431509
rect 355951 431593 356187 431829
rect 355951 431273 356187 431509
rect 361882 431593 362118 431829
rect 361882 431273 362118 431509
rect 367812 431593 368048 431829
rect 367812 431273 368048 431509
rect 383951 431593 384187 431829
rect 383951 431273 384187 431509
rect 389882 431593 390118 431829
rect 389882 431273 390118 431509
rect 395812 431593 396048 431829
rect 395812 431273 396048 431509
rect 411951 431593 412187 431829
rect 411951 431273 412187 431509
rect 417882 431593 418118 431829
rect 417882 431273 418118 431509
rect 423812 431593 424048 431829
rect 423812 431273 424048 431509
rect 439951 431593 440187 431829
rect 439951 431273 440187 431509
rect 445882 431593 446118 431829
rect 445882 431273 446118 431509
rect 451812 431593 452048 431829
rect 451812 431273 452048 431509
rect 467951 431593 468187 431829
rect 467951 431273 468187 431509
rect 473882 431593 474118 431829
rect 473882 431273 474118 431509
rect 479812 431593 480048 431829
rect 479812 431273 480048 431509
rect 495951 431593 496187 431829
rect 495951 431273 496187 431509
rect 501882 431593 502118 431829
rect 501882 431273 502118 431509
rect 507812 431593 508048 431829
rect 507812 431273 508048 431509
rect 523951 431593 524187 431829
rect 523951 431273 524187 431509
rect 529882 431593 530118 431829
rect 529882 431273 530118 431509
rect 535812 431593 536048 431829
rect 535812 431273 536048 431509
rect 551951 431593 552187 431829
rect 551951 431273 552187 431509
rect 557882 431593 558118 431829
rect 557882 431273 558118 431509
rect 563812 431593 564048 431829
rect 563812 431273 564048 431509
rect 573526 431593 573762 431829
rect 573846 431593 574082 431829
rect 573526 431273 573762 431509
rect 573846 431273 574082 431509
rect 22917 428218 23153 428454
rect 22917 427898 23153 428134
rect 28848 428218 29084 428454
rect 28848 427898 29084 428134
rect 50917 428218 51153 428454
rect 50917 427898 51153 428134
rect 56848 428218 57084 428454
rect 56848 427898 57084 428134
rect 78917 428218 79153 428454
rect 78917 427898 79153 428134
rect 84848 428218 85084 428454
rect 84848 427898 85084 428134
rect 106917 428218 107153 428454
rect 106917 427898 107153 428134
rect 112848 428218 113084 428454
rect 112848 427898 113084 428134
rect 134917 428218 135153 428454
rect 134917 427898 135153 428134
rect 140848 428218 141084 428454
rect 140848 427898 141084 428134
rect 162917 428218 163153 428454
rect 162917 427898 163153 428134
rect 168848 428218 169084 428454
rect 168848 427898 169084 428134
rect 190917 428218 191153 428454
rect 190917 427898 191153 428134
rect 196848 428218 197084 428454
rect 196848 427898 197084 428134
rect 218917 428218 219153 428454
rect 218917 427898 219153 428134
rect 224848 428218 225084 428454
rect 224848 427898 225084 428134
rect 246917 428218 247153 428454
rect 246917 427898 247153 428134
rect 252848 428218 253084 428454
rect 252848 427898 253084 428134
rect 274917 428218 275153 428454
rect 274917 427898 275153 428134
rect 280848 428218 281084 428454
rect 280848 427898 281084 428134
rect 302917 428218 303153 428454
rect 302917 427898 303153 428134
rect 308848 428218 309084 428454
rect 308848 427898 309084 428134
rect 330917 428218 331153 428454
rect 330917 427898 331153 428134
rect 336848 428218 337084 428454
rect 336848 427898 337084 428134
rect 358917 428218 359153 428454
rect 358917 427898 359153 428134
rect 364848 428218 365084 428454
rect 364848 427898 365084 428134
rect 386917 428218 387153 428454
rect 386917 427898 387153 428134
rect 392848 428218 393084 428454
rect 392848 427898 393084 428134
rect 414917 428218 415153 428454
rect 414917 427898 415153 428134
rect 420848 428218 421084 428454
rect 420848 427898 421084 428134
rect 442917 428218 443153 428454
rect 442917 427898 443153 428134
rect 448848 428218 449084 428454
rect 448848 427898 449084 428134
rect 470917 428218 471153 428454
rect 470917 427898 471153 428134
rect 476848 428218 477084 428454
rect 476848 427898 477084 428134
rect 498917 428218 499153 428454
rect 498917 427898 499153 428134
rect 504848 428218 505084 428454
rect 504848 427898 505084 428134
rect 526917 428218 527153 428454
rect 526917 427898 527153 428134
rect 532848 428218 533084 428454
rect 532848 427898 533084 428134
rect 554917 428218 555153 428454
rect 554917 427898 555153 428134
rect 560848 428218 561084 428454
rect 560848 427898 561084 428134
rect -1974 404593 -1738 404829
rect -1654 404593 -1418 404829
rect -1974 404273 -1738 404509
rect -1654 404273 -1418 404509
rect 19952 404593 20188 404829
rect 19952 404273 20188 404509
rect 25882 404593 26118 404829
rect 25882 404273 26118 404509
rect 31813 404593 32049 404829
rect 31813 404273 32049 404509
rect 47952 404593 48188 404829
rect 47952 404273 48188 404509
rect 53882 404593 54118 404829
rect 53882 404273 54118 404509
rect 59813 404593 60049 404829
rect 59813 404273 60049 404509
rect 75952 404593 76188 404829
rect 75952 404273 76188 404509
rect 81882 404593 82118 404829
rect 81882 404273 82118 404509
rect 87813 404593 88049 404829
rect 87813 404273 88049 404509
rect 103952 404593 104188 404829
rect 103952 404273 104188 404509
rect 109882 404593 110118 404829
rect 109882 404273 110118 404509
rect 115813 404593 116049 404829
rect 115813 404273 116049 404509
rect 131952 404593 132188 404829
rect 131952 404273 132188 404509
rect 137882 404593 138118 404829
rect 137882 404273 138118 404509
rect 143813 404593 144049 404829
rect 143813 404273 144049 404509
rect 159952 404593 160188 404829
rect 159952 404273 160188 404509
rect 165882 404593 166118 404829
rect 165882 404273 166118 404509
rect 171813 404593 172049 404829
rect 171813 404273 172049 404509
rect 187952 404593 188188 404829
rect 187952 404273 188188 404509
rect 193882 404593 194118 404829
rect 193882 404273 194118 404509
rect 199813 404593 200049 404829
rect 199813 404273 200049 404509
rect 215952 404593 216188 404829
rect 215952 404273 216188 404509
rect 221882 404593 222118 404829
rect 221882 404273 222118 404509
rect 227813 404593 228049 404829
rect 227813 404273 228049 404509
rect 243952 404593 244188 404829
rect 243952 404273 244188 404509
rect 249882 404593 250118 404829
rect 249882 404273 250118 404509
rect 255813 404593 256049 404829
rect 255813 404273 256049 404509
rect 271952 404593 272188 404829
rect 271952 404273 272188 404509
rect 277882 404593 278118 404829
rect 277882 404273 278118 404509
rect 283813 404593 284049 404829
rect 283813 404273 284049 404509
rect 299952 404593 300188 404829
rect 299952 404273 300188 404509
rect 305882 404593 306118 404829
rect 305882 404273 306118 404509
rect 311813 404593 312049 404829
rect 311813 404273 312049 404509
rect 327952 404593 328188 404829
rect 327952 404273 328188 404509
rect 333882 404593 334118 404829
rect 333882 404273 334118 404509
rect 339813 404593 340049 404829
rect 339813 404273 340049 404509
rect 355952 404593 356188 404829
rect 355952 404273 356188 404509
rect 361882 404593 362118 404829
rect 361882 404273 362118 404509
rect 367813 404593 368049 404829
rect 367813 404273 368049 404509
rect 383952 404593 384188 404829
rect 383952 404273 384188 404509
rect 389882 404593 390118 404829
rect 389882 404273 390118 404509
rect 395813 404593 396049 404829
rect 395813 404273 396049 404509
rect 411952 404593 412188 404829
rect 411952 404273 412188 404509
rect 417882 404593 418118 404829
rect 417882 404273 418118 404509
rect 423813 404593 424049 404829
rect 423813 404273 424049 404509
rect 439952 404593 440188 404829
rect 439952 404273 440188 404509
rect 445882 404593 446118 404829
rect 445882 404273 446118 404509
rect 451813 404593 452049 404829
rect 451813 404273 452049 404509
rect 467952 404593 468188 404829
rect 467952 404273 468188 404509
rect 473882 404593 474118 404829
rect 473882 404273 474118 404509
rect 479813 404593 480049 404829
rect 479813 404273 480049 404509
rect 495952 404593 496188 404829
rect 495952 404273 496188 404509
rect 501882 404593 502118 404829
rect 501882 404273 502118 404509
rect 507813 404593 508049 404829
rect 507813 404273 508049 404509
rect 523952 404593 524188 404829
rect 523952 404273 524188 404509
rect 529882 404593 530118 404829
rect 529882 404273 530118 404509
rect 535813 404593 536049 404829
rect 535813 404273 536049 404509
rect 551952 404593 552188 404829
rect 551952 404273 552188 404509
rect 557882 404593 558118 404829
rect 557882 404273 558118 404509
rect 563813 404593 564049 404829
rect 563813 404273 564049 404509
rect 573526 404593 573762 404829
rect 573846 404593 574082 404829
rect 573526 404273 573762 404509
rect 573846 404273 574082 404509
rect 22916 401218 23152 401454
rect 22916 400898 23152 401134
rect 28847 401218 29083 401454
rect 28847 400898 29083 401134
rect 50916 401218 51152 401454
rect 50916 400898 51152 401134
rect 56847 401218 57083 401454
rect 56847 400898 57083 401134
rect 78916 401218 79152 401454
rect 78916 400898 79152 401134
rect 84847 401218 85083 401454
rect 84847 400898 85083 401134
rect 106916 401218 107152 401454
rect 106916 400898 107152 401134
rect 112847 401218 113083 401454
rect 112847 400898 113083 401134
rect 134916 401218 135152 401454
rect 134916 400898 135152 401134
rect 140847 401218 141083 401454
rect 140847 400898 141083 401134
rect 162916 401218 163152 401454
rect 162916 400898 163152 401134
rect 168847 401218 169083 401454
rect 168847 400898 169083 401134
rect 190916 401218 191152 401454
rect 190916 400898 191152 401134
rect 196847 401218 197083 401454
rect 196847 400898 197083 401134
rect 218916 401218 219152 401454
rect 218916 400898 219152 401134
rect 224847 401218 225083 401454
rect 224847 400898 225083 401134
rect 246916 401218 247152 401454
rect 246916 400898 247152 401134
rect 252847 401218 253083 401454
rect 252847 400898 253083 401134
rect 274916 401218 275152 401454
rect 274916 400898 275152 401134
rect 280847 401218 281083 401454
rect 280847 400898 281083 401134
rect 302916 401218 303152 401454
rect 302916 400898 303152 401134
rect 308847 401218 309083 401454
rect 308847 400898 309083 401134
rect 330916 401218 331152 401454
rect 330916 400898 331152 401134
rect 336847 401218 337083 401454
rect 336847 400898 337083 401134
rect 358916 401218 359152 401454
rect 358916 400898 359152 401134
rect 364847 401218 365083 401454
rect 364847 400898 365083 401134
rect 386916 401218 387152 401454
rect 386916 400898 387152 401134
rect 392847 401218 393083 401454
rect 392847 400898 393083 401134
rect 414916 401218 415152 401454
rect 414916 400898 415152 401134
rect 420847 401218 421083 401454
rect 420847 400898 421083 401134
rect 442916 401218 443152 401454
rect 442916 400898 443152 401134
rect 448847 401218 449083 401454
rect 448847 400898 449083 401134
rect 470916 401218 471152 401454
rect 470916 400898 471152 401134
rect 476847 401218 477083 401454
rect 476847 400898 477083 401134
rect 498916 401218 499152 401454
rect 498916 400898 499152 401134
rect 504847 401218 505083 401454
rect 504847 400898 505083 401134
rect 526916 401218 527152 401454
rect 526916 400898 527152 401134
rect 532847 401218 533083 401454
rect 532847 400898 533083 401134
rect 554916 401218 555152 401454
rect 554916 400898 555152 401134
rect 560847 401218 561083 401454
rect 560847 400898 561083 401134
rect -1974 377593 -1738 377829
rect -1654 377593 -1418 377829
rect -1974 377273 -1738 377509
rect -1654 377273 -1418 377509
rect 19951 377593 20187 377829
rect 19951 377273 20187 377509
rect 25882 377593 26118 377829
rect 25882 377273 26118 377509
rect 31812 377593 32048 377829
rect 31812 377273 32048 377509
rect 47951 377593 48187 377829
rect 47951 377273 48187 377509
rect 53882 377593 54118 377829
rect 53882 377273 54118 377509
rect 59812 377593 60048 377829
rect 59812 377273 60048 377509
rect 75951 377593 76187 377829
rect 75951 377273 76187 377509
rect 81882 377593 82118 377829
rect 81882 377273 82118 377509
rect 87812 377593 88048 377829
rect 87812 377273 88048 377509
rect 103951 377593 104187 377829
rect 103951 377273 104187 377509
rect 109882 377593 110118 377829
rect 109882 377273 110118 377509
rect 115812 377593 116048 377829
rect 115812 377273 116048 377509
rect 131951 377593 132187 377829
rect 131951 377273 132187 377509
rect 137882 377593 138118 377829
rect 137882 377273 138118 377509
rect 143812 377593 144048 377829
rect 143812 377273 144048 377509
rect 159951 377593 160187 377829
rect 159951 377273 160187 377509
rect 165882 377593 166118 377829
rect 165882 377273 166118 377509
rect 171812 377593 172048 377829
rect 171812 377273 172048 377509
rect 187951 377593 188187 377829
rect 187951 377273 188187 377509
rect 193882 377593 194118 377829
rect 193882 377273 194118 377509
rect 199812 377593 200048 377829
rect 199812 377273 200048 377509
rect 215951 377593 216187 377829
rect 215951 377273 216187 377509
rect 221882 377593 222118 377829
rect 221882 377273 222118 377509
rect 227812 377593 228048 377829
rect 227812 377273 228048 377509
rect 243951 377593 244187 377829
rect 243951 377273 244187 377509
rect 249882 377593 250118 377829
rect 249882 377273 250118 377509
rect 255812 377593 256048 377829
rect 255812 377273 256048 377509
rect 271951 377593 272187 377829
rect 271951 377273 272187 377509
rect 277882 377593 278118 377829
rect 277882 377273 278118 377509
rect 283812 377593 284048 377829
rect 283812 377273 284048 377509
rect 299951 377593 300187 377829
rect 299951 377273 300187 377509
rect 305882 377593 306118 377829
rect 305882 377273 306118 377509
rect 311812 377593 312048 377829
rect 311812 377273 312048 377509
rect 327951 377593 328187 377829
rect 327951 377273 328187 377509
rect 333882 377593 334118 377829
rect 333882 377273 334118 377509
rect 339812 377593 340048 377829
rect 339812 377273 340048 377509
rect 355951 377593 356187 377829
rect 355951 377273 356187 377509
rect 361882 377593 362118 377829
rect 361882 377273 362118 377509
rect 367812 377593 368048 377829
rect 367812 377273 368048 377509
rect 383951 377593 384187 377829
rect 383951 377273 384187 377509
rect 389882 377593 390118 377829
rect 389882 377273 390118 377509
rect 395812 377593 396048 377829
rect 395812 377273 396048 377509
rect 411951 377593 412187 377829
rect 411951 377273 412187 377509
rect 417882 377593 418118 377829
rect 417882 377273 418118 377509
rect 423812 377593 424048 377829
rect 423812 377273 424048 377509
rect 439951 377593 440187 377829
rect 439951 377273 440187 377509
rect 445882 377593 446118 377829
rect 445882 377273 446118 377509
rect 451812 377593 452048 377829
rect 451812 377273 452048 377509
rect 467951 377593 468187 377829
rect 467951 377273 468187 377509
rect 473882 377593 474118 377829
rect 473882 377273 474118 377509
rect 479812 377593 480048 377829
rect 479812 377273 480048 377509
rect 495951 377593 496187 377829
rect 495951 377273 496187 377509
rect 501882 377593 502118 377829
rect 501882 377273 502118 377509
rect 507812 377593 508048 377829
rect 507812 377273 508048 377509
rect 523951 377593 524187 377829
rect 523951 377273 524187 377509
rect 529882 377593 530118 377829
rect 529882 377273 530118 377509
rect 535812 377593 536048 377829
rect 535812 377273 536048 377509
rect 551951 377593 552187 377829
rect 551951 377273 552187 377509
rect 557882 377593 558118 377829
rect 557882 377273 558118 377509
rect 563812 377593 564048 377829
rect 563812 377273 564048 377509
rect 573526 377593 573762 377829
rect 573846 377593 574082 377829
rect 573526 377273 573762 377509
rect 573846 377273 574082 377509
rect 22917 374218 23153 374454
rect 22917 373898 23153 374134
rect 28848 374218 29084 374454
rect 28848 373898 29084 374134
rect 50917 374218 51153 374454
rect 50917 373898 51153 374134
rect 56848 374218 57084 374454
rect 56848 373898 57084 374134
rect 78917 374218 79153 374454
rect 78917 373898 79153 374134
rect 84848 374218 85084 374454
rect 84848 373898 85084 374134
rect 106917 374218 107153 374454
rect 106917 373898 107153 374134
rect 112848 374218 113084 374454
rect 112848 373898 113084 374134
rect 134917 374218 135153 374454
rect 134917 373898 135153 374134
rect 140848 374218 141084 374454
rect 140848 373898 141084 374134
rect 162917 374218 163153 374454
rect 162917 373898 163153 374134
rect 168848 374218 169084 374454
rect 168848 373898 169084 374134
rect 190917 374218 191153 374454
rect 190917 373898 191153 374134
rect 196848 374218 197084 374454
rect 196848 373898 197084 374134
rect 218917 374218 219153 374454
rect 218917 373898 219153 374134
rect 224848 374218 225084 374454
rect 224848 373898 225084 374134
rect 246917 374218 247153 374454
rect 246917 373898 247153 374134
rect 252848 374218 253084 374454
rect 252848 373898 253084 374134
rect 274917 374218 275153 374454
rect 274917 373898 275153 374134
rect 280848 374218 281084 374454
rect 280848 373898 281084 374134
rect 302917 374218 303153 374454
rect 302917 373898 303153 374134
rect 308848 374218 309084 374454
rect 308848 373898 309084 374134
rect 330917 374218 331153 374454
rect 330917 373898 331153 374134
rect 336848 374218 337084 374454
rect 336848 373898 337084 374134
rect 358917 374218 359153 374454
rect 358917 373898 359153 374134
rect 364848 374218 365084 374454
rect 364848 373898 365084 374134
rect 386917 374218 387153 374454
rect 386917 373898 387153 374134
rect 392848 374218 393084 374454
rect 392848 373898 393084 374134
rect 414917 374218 415153 374454
rect 414917 373898 415153 374134
rect 420848 374218 421084 374454
rect 420848 373898 421084 374134
rect 442917 374218 443153 374454
rect 442917 373898 443153 374134
rect 448848 374218 449084 374454
rect 448848 373898 449084 374134
rect 470917 374218 471153 374454
rect 470917 373898 471153 374134
rect 476848 374218 477084 374454
rect 476848 373898 477084 374134
rect 498917 374218 499153 374454
rect 498917 373898 499153 374134
rect 504848 374218 505084 374454
rect 504848 373898 505084 374134
rect 526917 374218 527153 374454
rect 526917 373898 527153 374134
rect 532848 374218 533084 374454
rect 532848 373898 533084 374134
rect 554917 374218 555153 374454
rect 554917 373898 555153 374134
rect 560848 374218 561084 374454
rect 560848 373898 561084 374134
rect -1974 350593 -1738 350829
rect -1654 350593 -1418 350829
rect -1974 350273 -1738 350509
rect -1654 350273 -1418 350509
rect 19952 350593 20188 350829
rect 19952 350273 20188 350509
rect 25882 350593 26118 350829
rect 25882 350273 26118 350509
rect 31813 350593 32049 350829
rect 31813 350273 32049 350509
rect 47952 350593 48188 350829
rect 47952 350273 48188 350509
rect 53882 350593 54118 350829
rect 53882 350273 54118 350509
rect 59813 350593 60049 350829
rect 59813 350273 60049 350509
rect 75952 350593 76188 350829
rect 75952 350273 76188 350509
rect 81882 350593 82118 350829
rect 81882 350273 82118 350509
rect 87813 350593 88049 350829
rect 87813 350273 88049 350509
rect 103952 350593 104188 350829
rect 103952 350273 104188 350509
rect 109882 350593 110118 350829
rect 109882 350273 110118 350509
rect 115813 350593 116049 350829
rect 115813 350273 116049 350509
rect 131952 350593 132188 350829
rect 131952 350273 132188 350509
rect 137882 350593 138118 350829
rect 137882 350273 138118 350509
rect 143813 350593 144049 350829
rect 143813 350273 144049 350509
rect 159952 350593 160188 350829
rect 159952 350273 160188 350509
rect 165882 350593 166118 350829
rect 165882 350273 166118 350509
rect 171813 350593 172049 350829
rect 171813 350273 172049 350509
rect 187952 350593 188188 350829
rect 187952 350273 188188 350509
rect 193882 350593 194118 350829
rect 193882 350273 194118 350509
rect 199813 350593 200049 350829
rect 199813 350273 200049 350509
rect 215952 350593 216188 350829
rect 215952 350273 216188 350509
rect 221882 350593 222118 350829
rect 221882 350273 222118 350509
rect 227813 350593 228049 350829
rect 227813 350273 228049 350509
rect 243952 350593 244188 350829
rect 243952 350273 244188 350509
rect 249882 350593 250118 350829
rect 249882 350273 250118 350509
rect 255813 350593 256049 350829
rect 255813 350273 256049 350509
rect 271952 350593 272188 350829
rect 271952 350273 272188 350509
rect 277882 350593 278118 350829
rect 277882 350273 278118 350509
rect 283813 350593 284049 350829
rect 283813 350273 284049 350509
rect 299952 350593 300188 350829
rect 299952 350273 300188 350509
rect 305882 350593 306118 350829
rect 305882 350273 306118 350509
rect 311813 350593 312049 350829
rect 311813 350273 312049 350509
rect 327952 350593 328188 350829
rect 327952 350273 328188 350509
rect 333882 350593 334118 350829
rect 333882 350273 334118 350509
rect 339813 350593 340049 350829
rect 339813 350273 340049 350509
rect 355952 350593 356188 350829
rect 355952 350273 356188 350509
rect 361882 350593 362118 350829
rect 361882 350273 362118 350509
rect 367813 350593 368049 350829
rect 367813 350273 368049 350509
rect 383952 350593 384188 350829
rect 383952 350273 384188 350509
rect 389882 350593 390118 350829
rect 389882 350273 390118 350509
rect 395813 350593 396049 350829
rect 395813 350273 396049 350509
rect 411952 350593 412188 350829
rect 411952 350273 412188 350509
rect 417882 350593 418118 350829
rect 417882 350273 418118 350509
rect 423813 350593 424049 350829
rect 423813 350273 424049 350509
rect 439952 350593 440188 350829
rect 439952 350273 440188 350509
rect 445882 350593 446118 350829
rect 445882 350273 446118 350509
rect 451813 350593 452049 350829
rect 451813 350273 452049 350509
rect 467952 350593 468188 350829
rect 467952 350273 468188 350509
rect 473882 350593 474118 350829
rect 473882 350273 474118 350509
rect 479813 350593 480049 350829
rect 479813 350273 480049 350509
rect 495952 350593 496188 350829
rect 495952 350273 496188 350509
rect 501882 350593 502118 350829
rect 501882 350273 502118 350509
rect 507813 350593 508049 350829
rect 507813 350273 508049 350509
rect 523952 350593 524188 350829
rect 523952 350273 524188 350509
rect 529882 350593 530118 350829
rect 529882 350273 530118 350509
rect 535813 350593 536049 350829
rect 535813 350273 536049 350509
rect 551952 350593 552188 350829
rect 551952 350273 552188 350509
rect 557882 350593 558118 350829
rect 557882 350273 558118 350509
rect 563813 350593 564049 350829
rect 563813 350273 564049 350509
rect 573526 350593 573762 350829
rect 573846 350593 574082 350829
rect 573526 350273 573762 350509
rect 573846 350273 574082 350509
rect 22916 347218 23152 347454
rect 22916 346898 23152 347134
rect 28847 347218 29083 347454
rect 28847 346898 29083 347134
rect 50916 347218 51152 347454
rect 50916 346898 51152 347134
rect 56847 347218 57083 347454
rect 56847 346898 57083 347134
rect 78916 347218 79152 347454
rect 78916 346898 79152 347134
rect 84847 347218 85083 347454
rect 84847 346898 85083 347134
rect 106916 347218 107152 347454
rect 106916 346898 107152 347134
rect 112847 347218 113083 347454
rect 112847 346898 113083 347134
rect 134916 347218 135152 347454
rect 134916 346898 135152 347134
rect 140847 347218 141083 347454
rect 140847 346898 141083 347134
rect 162916 347218 163152 347454
rect 162916 346898 163152 347134
rect 168847 347218 169083 347454
rect 168847 346898 169083 347134
rect 190916 347218 191152 347454
rect 190916 346898 191152 347134
rect 196847 347218 197083 347454
rect 196847 346898 197083 347134
rect 218916 347218 219152 347454
rect 218916 346898 219152 347134
rect 224847 347218 225083 347454
rect 224847 346898 225083 347134
rect 246916 347218 247152 347454
rect 246916 346898 247152 347134
rect 252847 347218 253083 347454
rect 252847 346898 253083 347134
rect 274916 347218 275152 347454
rect 274916 346898 275152 347134
rect 280847 347218 281083 347454
rect 280847 346898 281083 347134
rect 302916 347218 303152 347454
rect 302916 346898 303152 347134
rect 308847 347218 309083 347454
rect 308847 346898 309083 347134
rect 330916 347218 331152 347454
rect 330916 346898 331152 347134
rect 336847 347218 337083 347454
rect 336847 346898 337083 347134
rect 358916 347218 359152 347454
rect 358916 346898 359152 347134
rect 364847 347218 365083 347454
rect 364847 346898 365083 347134
rect 386916 347218 387152 347454
rect 386916 346898 387152 347134
rect 392847 347218 393083 347454
rect 392847 346898 393083 347134
rect 414916 347218 415152 347454
rect 414916 346898 415152 347134
rect 420847 347218 421083 347454
rect 420847 346898 421083 347134
rect 442916 347218 443152 347454
rect 442916 346898 443152 347134
rect 448847 347218 449083 347454
rect 448847 346898 449083 347134
rect 470916 347218 471152 347454
rect 470916 346898 471152 347134
rect 476847 347218 477083 347454
rect 476847 346898 477083 347134
rect 498916 347218 499152 347454
rect 498916 346898 499152 347134
rect 504847 347218 505083 347454
rect 504847 346898 505083 347134
rect 526916 347218 527152 347454
rect 526916 346898 527152 347134
rect 532847 347218 533083 347454
rect 532847 346898 533083 347134
rect 554916 347218 555152 347454
rect 554916 346898 555152 347134
rect 560847 347218 561083 347454
rect 560847 346898 561083 347134
rect -1974 323593 -1738 323829
rect -1654 323593 -1418 323829
rect -1974 323273 -1738 323509
rect -1654 323273 -1418 323509
rect 19951 323593 20187 323829
rect 19951 323273 20187 323509
rect 25882 323593 26118 323829
rect 25882 323273 26118 323509
rect 31812 323593 32048 323829
rect 31812 323273 32048 323509
rect 47951 323593 48187 323829
rect 47951 323273 48187 323509
rect 53882 323593 54118 323829
rect 53882 323273 54118 323509
rect 59812 323593 60048 323829
rect 59812 323273 60048 323509
rect 75951 323593 76187 323829
rect 75951 323273 76187 323509
rect 81882 323593 82118 323829
rect 81882 323273 82118 323509
rect 87812 323593 88048 323829
rect 87812 323273 88048 323509
rect 103951 323593 104187 323829
rect 103951 323273 104187 323509
rect 109882 323593 110118 323829
rect 109882 323273 110118 323509
rect 115812 323593 116048 323829
rect 115812 323273 116048 323509
rect 131951 323593 132187 323829
rect 131951 323273 132187 323509
rect 137882 323593 138118 323829
rect 137882 323273 138118 323509
rect 143812 323593 144048 323829
rect 143812 323273 144048 323509
rect 159951 323593 160187 323829
rect 159951 323273 160187 323509
rect 165882 323593 166118 323829
rect 165882 323273 166118 323509
rect 171812 323593 172048 323829
rect 171812 323273 172048 323509
rect 187951 323593 188187 323829
rect 187951 323273 188187 323509
rect 193882 323593 194118 323829
rect 193882 323273 194118 323509
rect 199812 323593 200048 323829
rect 199812 323273 200048 323509
rect 215951 323593 216187 323829
rect 215951 323273 216187 323509
rect 221882 323593 222118 323829
rect 221882 323273 222118 323509
rect 227812 323593 228048 323829
rect 227812 323273 228048 323509
rect 243951 323593 244187 323829
rect 243951 323273 244187 323509
rect 249882 323593 250118 323829
rect 249882 323273 250118 323509
rect 255812 323593 256048 323829
rect 255812 323273 256048 323509
rect 271951 323593 272187 323829
rect 271951 323273 272187 323509
rect 277882 323593 278118 323829
rect 277882 323273 278118 323509
rect 283812 323593 284048 323829
rect 283812 323273 284048 323509
rect 299951 323593 300187 323829
rect 299951 323273 300187 323509
rect 305882 323593 306118 323829
rect 305882 323273 306118 323509
rect 311812 323593 312048 323829
rect 311812 323273 312048 323509
rect 327951 323593 328187 323829
rect 327951 323273 328187 323509
rect 333882 323593 334118 323829
rect 333882 323273 334118 323509
rect 339812 323593 340048 323829
rect 339812 323273 340048 323509
rect 355951 323593 356187 323829
rect 355951 323273 356187 323509
rect 361882 323593 362118 323829
rect 361882 323273 362118 323509
rect 367812 323593 368048 323829
rect 367812 323273 368048 323509
rect 383951 323593 384187 323829
rect 383951 323273 384187 323509
rect 389882 323593 390118 323829
rect 389882 323273 390118 323509
rect 395812 323593 396048 323829
rect 395812 323273 396048 323509
rect 411951 323593 412187 323829
rect 411951 323273 412187 323509
rect 417882 323593 418118 323829
rect 417882 323273 418118 323509
rect 423812 323593 424048 323829
rect 423812 323273 424048 323509
rect 439951 323593 440187 323829
rect 439951 323273 440187 323509
rect 445882 323593 446118 323829
rect 445882 323273 446118 323509
rect 451812 323593 452048 323829
rect 451812 323273 452048 323509
rect 467951 323593 468187 323829
rect 467951 323273 468187 323509
rect 473882 323593 474118 323829
rect 473882 323273 474118 323509
rect 479812 323593 480048 323829
rect 479812 323273 480048 323509
rect 495951 323593 496187 323829
rect 495951 323273 496187 323509
rect 501882 323593 502118 323829
rect 501882 323273 502118 323509
rect 507812 323593 508048 323829
rect 507812 323273 508048 323509
rect 523951 323593 524187 323829
rect 523951 323273 524187 323509
rect 529882 323593 530118 323829
rect 529882 323273 530118 323509
rect 535812 323593 536048 323829
rect 535812 323273 536048 323509
rect 551951 323593 552187 323829
rect 551951 323273 552187 323509
rect 557882 323593 558118 323829
rect 557882 323273 558118 323509
rect 563812 323593 564048 323829
rect 563812 323273 564048 323509
rect 573526 323593 573762 323829
rect 573846 323593 574082 323829
rect 573526 323273 573762 323509
rect 573846 323273 574082 323509
rect 22917 320218 23153 320454
rect 22917 319898 23153 320134
rect 28848 320218 29084 320454
rect 28848 319898 29084 320134
rect 50917 320218 51153 320454
rect 50917 319898 51153 320134
rect 56848 320218 57084 320454
rect 56848 319898 57084 320134
rect 78917 320218 79153 320454
rect 78917 319898 79153 320134
rect 84848 320218 85084 320454
rect 84848 319898 85084 320134
rect 106917 320218 107153 320454
rect 106917 319898 107153 320134
rect 112848 320218 113084 320454
rect 112848 319898 113084 320134
rect 134917 320218 135153 320454
rect 134917 319898 135153 320134
rect 140848 320218 141084 320454
rect 140848 319898 141084 320134
rect 162917 320218 163153 320454
rect 162917 319898 163153 320134
rect 168848 320218 169084 320454
rect 168848 319898 169084 320134
rect 190917 320218 191153 320454
rect 190917 319898 191153 320134
rect 196848 320218 197084 320454
rect 196848 319898 197084 320134
rect 218917 320218 219153 320454
rect 218917 319898 219153 320134
rect 224848 320218 225084 320454
rect 224848 319898 225084 320134
rect 246917 320218 247153 320454
rect 246917 319898 247153 320134
rect 252848 320218 253084 320454
rect 252848 319898 253084 320134
rect 274917 320218 275153 320454
rect 274917 319898 275153 320134
rect 280848 320218 281084 320454
rect 280848 319898 281084 320134
rect 302917 320218 303153 320454
rect 302917 319898 303153 320134
rect 308848 320218 309084 320454
rect 308848 319898 309084 320134
rect 330917 320218 331153 320454
rect 330917 319898 331153 320134
rect 336848 320218 337084 320454
rect 336848 319898 337084 320134
rect 358917 320218 359153 320454
rect 358917 319898 359153 320134
rect 364848 320218 365084 320454
rect 364848 319898 365084 320134
rect 386917 320218 387153 320454
rect 386917 319898 387153 320134
rect 392848 320218 393084 320454
rect 392848 319898 393084 320134
rect 414917 320218 415153 320454
rect 414917 319898 415153 320134
rect 420848 320218 421084 320454
rect 420848 319898 421084 320134
rect 442917 320218 443153 320454
rect 442917 319898 443153 320134
rect 448848 320218 449084 320454
rect 448848 319898 449084 320134
rect 470917 320218 471153 320454
rect 470917 319898 471153 320134
rect 476848 320218 477084 320454
rect 476848 319898 477084 320134
rect 498917 320218 499153 320454
rect 498917 319898 499153 320134
rect 504848 320218 505084 320454
rect 504848 319898 505084 320134
rect 526917 320218 527153 320454
rect 526917 319898 527153 320134
rect 532848 320218 533084 320454
rect 532848 319898 533084 320134
rect 554917 320218 555153 320454
rect 554917 319898 555153 320134
rect 560848 320218 561084 320454
rect 560848 319898 561084 320134
rect -1974 296593 -1738 296829
rect -1654 296593 -1418 296829
rect -1974 296273 -1738 296509
rect -1654 296273 -1418 296509
rect 19952 296593 20188 296829
rect 19952 296273 20188 296509
rect 25882 296593 26118 296829
rect 25882 296273 26118 296509
rect 31813 296593 32049 296829
rect 31813 296273 32049 296509
rect 47952 296593 48188 296829
rect 47952 296273 48188 296509
rect 53882 296593 54118 296829
rect 53882 296273 54118 296509
rect 59813 296593 60049 296829
rect 59813 296273 60049 296509
rect 75952 296593 76188 296829
rect 75952 296273 76188 296509
rect 81882 296593 82118 296829
rect 81882 296273 82118 296509
rect 87813 296593 88049 296829
rect 87813 296273 88049 296509
rect 103952 296593 104188 296829
rect 103952 296273 104188 296509
rect 109882 296593 110118 296829
rect 109882 296273 110118 296509
rect 115813 296593 116049 296829
rect 115813 296273 116049 296509
rect 131952 296593 132188 296829
rect 131952 296273 132188 296509
rect 137882 296593 138118 296829
rect 137882 296273 138118 296509
rect 143813 296593 144049 296829
rect 143813 296273 144049 296509
rect 159952 296593 160188 296829
rect 159952 296273 160188 296509
rect 165882 296593 166118 296829
rect 165882 296273 166118 296509
rect 171813 296593 172049 296829
rect 171813 296273 172049 296509
rect 187952 296593 188188 296829
rect 187952 296273 188188 296509
rect 193882 296593 194118 296829
rect 193882 296273 194118 296509
rect 199813 296593 200049 296829
rect 199813 296273 200049 296509
rect 215952 296593 216188 296829
rect 215952 296273 216188 296509
rect 221882 296593 222118 296829
rect 221882 296273 222118 296509
rect 227813 296593 228049 296829
rect 227813 296273 228049 296509
rect 243952 296593 244188 296829
rect 243952 296273 244188 296509
rect 249882 296593 250118 296829
rect 249882 296273 250118 296509
rect 255813 296593 256049 296829
rect 255813 296273 256049 296509
rect 271952 296593 272188 296829
rect 271952 296273 272188 296509
rect 277882 296593 278118 296829
rect 277882 296273 278118 296509
rect 283813 296593 284049 296829
rect 283813 296273 284049 296509
rect 299952 296593 300188 296829
rect 299952 296273 300188 296509
rect 305882 296593 306118 296829
rect 305882 296273 306118 296509
rect 311813 296593 312049 296829
rect 311813 296273 312049 296509
rect 327952 296593 328188 296829
rect 327952 296273 328188 296509
rect 333882 296593 334118 296829
rect 333882 296273 334118 296509
rect 339813 296593 340049 296829
rect 339813 296273 340049 296509
rect 355952 296593 356188 296829
rect 355952 296273 356188 296509
rect 361882 296593 362118 296829
rect 361882 296273 362118 296509
rect 367813 296593 368049 296829
rect 367813 296273 368049 296509
rect 383952 296593 384188 296829
rect 383952 296273 384188 296509
rect 389882 296593 390118 296829
rect 389882 296273 390118 296509
rect 395813 296593 396049 296829
rect 395813 296273 396049 296509
rect 411952 296593 412188 296829
rect 411952 296273 412188 296509
rect 417882 296593 418118 296829
rect 417882 296273 418118 296509
rect 423813 296593 424049 296829
rect 423813 296273 424049 296509
rect 439952 296593 440188 296829
rect 439952 296273 440188 296509
rect 445882 296593 446118 296829
rect 445882 296273 446118 296509
rect 451813 296593 452049 296829
rect 451813 296273 452049 296509
rect 467952 296593 468188 296829
rect 467952 296273 468188 296509
rect 473882 296593 474118 296829
rect 473882 296273 474118 296509
rect 479813 296593 480049 296829
rect 479813 296273 480049 296509
rect 495952 296593 496188 296829
rect 495952 296273 496188 296509
rect 501882 296593 502118 296829
rect 501882 296273 502118 296509
rect 507813 296593 508049 296829
rect 507813 296273 508049 296509
rect 523952 296593 524188 296829
rect 523952 296273 524188 296509
rect 529882 296593 530118 296829
rect 529882 296273 530118 296509
rect 535813 296593 536049 296829
rect 535813 296273 536049 296509
rect 551952 296593 552188 296829
rect 551952 296273 552188 296509
rect 557882 296593 558118 296829
rect 557882 296273 558118 296509
rect 563813 296593 564049 296829
rect 563813 296273 564049 296509
rect 573526 296593 573762 296829
rect 573846 296593 574082 296829
rect 573526 296273 573762 296509
rect 573846 296273 574082 296509
rect 22916 293218 23152 293454
rect 22916 292898 23152 293134
rect 28847 293218 29083 293454
rect 28847 292898 29083 293134
rect 50916 293218 51152 293454
rect 50916 292898 51152 293134
rect 56847 293218 57083 293454
rect 56847 292898 57083 293134
rect 78916 293218 79152 293454
rect 78916 292898 79152 293134
rect 84847 293218 85083 293454
rect 84847 292898 85083 293134
rect 106916 293218 107152 293454
rect 106916 292898 107152 293134
rect 112847 293218 113083 293454
rect 112847 292898 113083 293134
rect 134916 293218 135152 293454
rect 134916 292898 135152 293134
rect 140847 293218 141083 293454
rect 140847 292898 141083 293134
rect 162916 293218 163152 293454
rect 162916 292898 163152 293134
rect 168847 293218 169083 293454
rect 168847 292898 169083 293134
rect 190916 293218 191152 293454
rect 190916 292898 191152 293134
rect 196847 293218 197083 293454
rect 196847 292898 197083 293134
rect 218916 293218 219152 293454
rect 218916 292898 219152 293134
rect 224847 293218 225083 293454
rect 224847 292898 225083 293134
rect 246916 293218 247152 293454
rect 246916 292898 247152 293134
rect 252847 293218 253083 293454
rect 252847 292898 253083 293134
rect 274916 293218 275152 293454
rect 274916 292898 275152 293134
rect 280847 293218 281083 293454
rect 280847 292898 281083 293134
rect 302916 293218 303152 293454
rect 302916 292898 303152 293134
rect 308847 293218 309083 293454
rect 308847 292898 309083 293134
rect 330916 293218 331152 293454
rect 330916 292898 331152 293134
rect 336847 293218 337083 293454
rect 336847 292898 337083 293134
rect 358916 293218 359152 293454
rect 358916 292898 359152 293134
rect 364847 293218 365083 293454
rect 364847 292898 365083 293134
rect 386916 293218 387152 293454
rect 386916 292898 387152 293134
rect 392847 293218 393083 293454
rect 392847 292898 393083 293134
rect 414916 293218 415152 293454
rect 414916 292898 415152 293134
rect 420847 293218 421083 293454
rect 420847 292898 421083 293134
rect 442916 293218 443152 293454
rect 442916 292898 443152 293134
rect 448847 293218 449083 293454
rect 448847 292898 449083 293134
rect 470916 293218 471152 293454
rect 470916 292898 471152 293134
rect 476847 293218 477083 293454
rect 476847 292898 477083 293134
rect 498916 293218 499152 293454
rect 498916 292898 499152 293134
rect 504847 293218 505083 293454
rect 504847 292898 505083 293134
rect 526916 293218 527152 293454
rect 526916 292898 527152 293134
rect 532847 293218 533083 293454
rect 532847 292898 533083 293134
rect 554916 293218 555152 293454
rect 554916 292898 555152 293134
rect 560847 293218 561083 293454
rect 560847 292898 561083 293134
rect -1974 269593 -1738 269829
rect -1654 269593 -1418 269829
rect -1974 269273 -1738 269509
rect -1654 269273 -1418 269509
rect 19951 269593 20187 269829
rect 19951 269273 20187 269509
rect 25882 269593 26118 269829
rect 25882 269273 26118 269509
rect 31812 269593 32048 269829
rect 31812 269273 32048 269509
rect 47951 269593 48187 269829
rect 47951 269273 48187 269509
rect 53882 269593 54118 269829
rect 53882 269273 54118 269509
rect 59812 269593 60048 269829
rect 59812 269273 60048 269509
rect 75951 269593 76187 269829
rect 75951 269273 76187 269509
rect 81882 269593 82118 269829
rect 81882 269273 82118 269509
rect 87812 269593 88048 269829
rect 87812 269273 88048 269509
rect 103951 269593 104187 269829
rect 103951 269273 104187 269509
rect 109882 269593 110118 269829
rect 109882 269273 110118 269509
rect 115812 269593 116048 269829
rect 115812 269273 116048 269509
rect 131951 269593 132187 269829
rect 131951 269273 132187 269509
rect 137882 269593 138118 269829
rect 137882 269273 138118 269509
rect 143812 269593 144048 269829
rect 143812 269273 144048 269509
rect 159951 269593 160187 269829
rect 159951 269273 160187 269509
rect 165882 269593 166118 269829
rect 165882 269273 166118 269509
rect 171812 269593 172048 269829
rect 171812 269273 172048 269509
rect 187951 269593 188187 269829
rect 187951 269273 188187 269509
rect 193882 269593 194118 269829
rect 193882 269273 194118 269509
rect 199812 269593 200048 269829
rect 199812 269273 200048 269509
rect 215951 269593 216187 269829
rect 215951 269273 216187 269509
rect 221882 269593 222118 269829
rect 221882 269273 222118 269509
rect 227812 269593 228048 269829
rect 227812 269273 228048 269509
rect 243951 269593 244187 269829
rect 243951 269273 244187 269509
rect 249882 269593 250118 269829
rect 249882 269273 250118 269509
rect 255812 269593 256048 269829
rect 255812 269273 256048 269509
rect 271951 269593 272187 269829
rect 271951 269273 272187 269509
rect 277882 269593 278118 269829
rect 277882 269273 278118 269509
rect 283812 269593 284048 269829
rect 283812 269273 284048 269509
rect 299951 269593 300187 269829
rect 299951 269273 300187 269509
rect 305882 269593 306118 269829
rect 305882 269273 306118 269509
rect 311812 269593 312048 269829
rect 311812 269273 312048 269509
rect 327951 269593 328187 269829
rect 327951 269273 328187 269509
rect 333882 269593 334118 269829
rect 333882 269273 334118 269509
rect 339812 269593 340048 269829
rect 339812 269273 340048 269509
rect 355951 269593 356187 269829
rect 355951 269273 356187 269509
rect 361882 269593 362118 269829
rect 361882 269273 362118 269509
rect 367812 269593 368048 269829
rect 367812 269273 368048 269509
rect 383951 269593 384187 269829
rect 383951 269273 384187 269509
rect 389882 269593 390118 269829
rect 389882 269273 390118 269509
rect 395812 269593 396048 269829
rect 395812 269273 396048 269509
rect 411951 269593 412187 269829
rect 411951 269273 412187 269509
rect 417882 269593 418118 269829
rect 417882 269273 418118 269509
rect 423812 269593 424048 269829
rect 423812 269273 424048 269509
rect 439951 269593 440187 269829
rect 439951 269273 440187 269509
rect 445882 269593 446118 269829
rect 445882 269273 446118 269509
rect 451812 269593 452048 269829
rect 451812 269273 452048 269509
rect 467951 269593 468187 269829
rect 467951 269273 468187 269509
rect 473882 269593 474118 269829
rect 473882 269273 474118 269509
rect 479812 269593 480048 269829
rect 479812 269273 480048 269509
rect 495951 269593 496187 269829
rect 495951 269273 496187 269509
rect 501882 269593 502118 269829
rect 501882 269273 502118 269509
rect 507812 269593 508048 269829
rect 507812 269273 508048 269509
rect 523951 269593 524187 269829
rect 523951 269273 524187 269509
rect 529882 269593 530118 269829
rect 529882 269273 530118 269509
rect 535812 269593 536048 269829
rect 535812 269273 536048 269509
rect 551951 269593 552187 269829
rect 551951 269273 552187 269509
rect 557882 269593 558118 269829
rect 557882 269273 558118 269509
rect 563812 269593 564048 269829
rect 563812 269273 564048 269509
rect 573526 269593 573762 269829
rect 573846 269593 574082 269829
rect 573526 269273 573762 269509
rect 573846 269273 574082 269509
rect 22917 266218 23153 266454
rect 22917 265898 23153 266134
rect 28848 266218 29084 266454
rect 28848 265898 29084 266134
rect 50917 266218 51153 266454
rect 50917 265898 51153 266134
rect 56848 266218 57084 266454
rect 56848 265898 57084 266134
rect 78917 266218 79153 266454
rect 78917 265898 79153 266134
rect 84848 266218 85084 266454
rect 84848 265898 85084 266134
rect 106917 266218 107153 266454
rect 106917 265898 107153 266134
rect 112848 266218 113084 266454
rect 112848 265898 113084 266134
rect 134917 266218 135153 266454
rect 134917 265898 135153 266134
rect 140848 266218 141084 266454
rect 140848 265898 141084 266134
rect 162917 266218 163153 266454
rect 162917 265898 163153 266134
rect 168848 266218 169084 266454
rect 168848 265898 169084 266134
rect 190917 266218 191153 266454
rect 190917 265898 191153 266134
rect 196848 266218 197084 266454
rect 196848 265898 197084 266134
rect 218917 266218 219153 266454
rect 218917 265898 219153 266134
rect 224848 266218 225084 266454
rect 224848 265898 225084 266134
rect 246917 266218 247153 266454
rect 246917 265898 247153 266134
rect 252848 266218 253084 266454
rect 252848 265898 253084 266134
rect 274917 266218 275153 266454
rect 274917 265898 275153 266134
rect 280848 266218 281084 266454
rect 280848 265898 281084 266134
rect 302917 266218 303153 266454
rect 302917 265898 303153 266134
rect 308848 266218 309084 266454
rect 308848 265898 309084 266134
rect 330917 266218 331153 266454
rect 330917 265898 331153 266134
rect 336848 266218 337084 266454
rect 336848 265898 337084 266134
rect 358917 266218 359153 266454
rect 358917 265898 359153 266134
rect 364848 266218 365084 266454
rect 364848 265898 365084 266134
rect 386917 266218 387153 266454
rect 386917 265898 387153 266134
rect 392848 266218 393084 266454
rect 392848 265898 393084 266134
rect 414917 266218 415153 266454
rect 414917 265898 415153 266134
rect 420848 266218 421084 266454
rect 420848 265898 421084 266134
rect 442917 266218 443153 266454
rect 442917 265898 443153 266134
rect 448848 266218 449084 266454
rect 448848 265898 449084 266134
rect 470917 266218 471153 266454
rect 470917 265898 471153 266134
rect 476848 266218 477084 266454
rect 476848 265898 477084 266134
rect 498917 266218 499153 266454
rect 498917 265898 499153 266134
rect 504848 266218 505084 266454
rect 504848 265898 505084 266134
rect 526917 266218 527153 266454
rect 526917 265898 527153 266134
rect 532848 266218 533084 266454
rect 532848 265898 533084 266134
rect 554917 266218 555153 266454
rect 554917 265898 555153 266134
rect 560848 266218 561084 266454
rect 560848 265898 561084 266134
rect -1974 242593 -1738 242829
rect -1654 242593 -1418 242829
rect -1974 242273 -1738 242509
rect -1654 242273 -1418 242509
rect 19952 242593 20188 242829
rect 19952 242273 20188 242509
rect 25882 242593 26118 242829
rect 25882 242273 26118 242509
rect 31813 242593 32049 242829
rect 31813 242273 32049 242509
rect 47952 242593 48188 242829
rect 47952 242273 48188 242509
rect 53882 242593 54118 242829
rect 53882 242273 54118 242509
rect 59813 242593 60049 242829
rect 59813 242273 60049 242509
rect 75952 242593 76188 242829
rect 75952 242273 76188 242509
rect 81882 242593 82118 242829
rect 81882 242273 82118 242509
rect 87813 242593 88049 242829
rect 87813 242273 88049 242509
rect 103952 242593 104188 242829
rect 103952 242273 104188 242509
rect 109882 242593 110118 242829
rect 109882 242273 110118 242509
rect 115813 242593 116049 242829
rect 115813 242273 116049 242509
rect 131952 242593 132188 242829
rect 131952 242273 132188 242509
rect 137882 242593 138118 242829
rect 137882 242273 138118 242509
rect 143813 242593 144049 242829
rect 143813 242273 144049 242509
rect 159952 242593 160188 242829
rect 159952 242273 160188 242509
rect 165882 242593 166118 242829
rect 165882 242273 166118 242509
rect 171813 242593 172049 242829
rect 171813 242273 172049 242509
rect 187952 242593 188188 242829
rect 187952 242273 188188 242509
rect 193882 242593 194118 242829
rect 193882 242273 194118 242509
rect 199813 242593 200049 242829
rect 199813 242273 200049 242509
rect 215952 242593 216188 242829
rect 215952 242273 216188 242509
rect 221882 242593 222118 242829
rect 221882 242273 222118 242509
rect 227813 242593 228049 242829
rect 227813 242273 228049 242509
rect 243952 242593 244188 242829
rect 243952 242273 244188 242509
rect 249882 242593 250118 242829
rect 249882 242273 250118 242509
rect 255813 242593 256049 242829
rect 255813 242273 256049 242509
rect 271952 242593 272188 242829
rect 271952 242273 272188 242509
rect 277882 242593 278118 242829
rect 277882 242273 278118 242509
rect 283813 242593 284049 242829
rect 283813 242273 284049 242509
rect 299952 242593 300188 242829
rect 299952 242273 300188 242509
rect 305882 242593 306118 242829
rect 305882 242273 306118 242509
rect 311813 242593 312049 242829
rect 311813 242273 312049 242509
rect 327952 242593 328188 242829
rect 327952 242273 328188 242509
rect 333882 242593 334118 242829
rect 333882 242273 334118 242509
rect 339813 242593 340049 242829
rect 339813 242273 340049 242509
rect 355952 242593 356188 242829
rect 355952 242273 356188 242509
rect 361882 242593 362118 242829
rect 361882 242273 362118 242509
rect 367813 242593 368049 242829
rect 367813 242273 368049 242509
rect 383952 242593 384188 242829
rect 383952 242273 384188 242509
rect 389882 242593 390118 242829
rect 389882 242273 390118 242509
rect 395813 242593 396049 242829
rect 395813 242273 396049 242509
rect 411952 242593 412188 242829
rect 411952 242273 412188 242509
rect 417882 242593 418118 242829
rect 417882 242273 418118 242509
rect 423813 242593 424049 242829
rect 423813 242273 424049 242509
rect 439952 242593 440188 242829
rect 439952 242273 440188 242509
rect 445882 242593 446118 242829
rect 445882 242273 446118 242509
rect 451813 242593 452049 242829
rect 451813 242273 452049 242509
rect 467952 242593 468188 242829
rect 467952 242273 468188 242509
rect 473882 242593 474118 242829
rect 473882 242273 474118 242509
rect 479813 242593 480049 242829
rect 479813 242273 480049 242509
rect 495952 242593 496188 242829
rect 495952 242273 496188 242509
rect 501882 242593 502118 242829
rect 501882 242273 502118 242509
rect 507813 242593 508049 242829
rect 507813 242273 508049 242509
rect 523952 242593 524188 242829
rect 523952 242273 524188 242509
rect 529882 242593 530118 242829
rect 529882 242273 530118 242509
rect 535813 242593 536049 242829
rect 535813 242273 536049 242509
rect 551952 242593 552188 242829
rect 551952 242273 552188 242509
rect 557882 242593 558118 242829
rect 557882 242273 558118 242509
rect 563813 242593 564049 242829
rect 563813 242273 564049 242509
rect 573526 242593 573762 242829
rect 573846 242593 574082 242829
rect 573526 242273 573762 242509
rect 573846 242273 574082 242509
rect 22916 239218 23152 239454
rect 22916 238898 23152 239134
rect 28847 239218 29083 239454
rect 28847 238898 29083 239134
rect 50916 239218 51152 239454
rect 50916 238898 51152 239134
rect 56847 239218 57083 239454
rect 56847 238898 57083 239134
rect 78916 239218 79152 239454
rect 78916 238898 79152 239134
rect 84847 239218 85083 239454
rect 84847 238898 85083 239134
rect 106916 239218 107152 239454
rect 106916 238898 107152 239134
rect 112847 239218 113083 239454
rect 112847 238898 113083 239134
rect 134916 239218 135152 239454
rect 134916 238898 135152 239134
rect 140847 239218 141083 239454
rect 140847 238898 141083 239134
rect 162916 239218 163152 239454
rect 162916 238898 163152 239134
rect 168847 239218 169083 239454
rect 168847 238898 169083 239134
rect 190916 239218 191152 239454
rect 190916 238898 191152 239134
rect 196847 239218 197083 239454
rect 196847 238898 197083 239134
rect 218916 239218 219152 239454
rect 218916 238898 219152 239134
rect 224847 239218 225083 239454
rect 224847 238898 225083 239134
rect 246916 239218 247152 239454
rect 246916 238898 247152 239134
rect 252847 239218 253083 239454
rect 252847 238898 253083 239134
rect 274916 239218 275152 239454
rect 274916 238898 275152 239134
rect 280847 239218 281083 239454
rect 280847 238898 281083 239134
rect 302916 239218 303152 239454
rect 302916 238898 303152 239134
rect 308847 239218 309083 239454
rect 308847 238898 309083 239134
rect 330916 239218 331152 239454
rect 330916 238898 331152 239134
rect 336847 239218 337083 239454
rect 336847 238898 337083 239134
rect 358916 239218 359152 239454
rect 358916 238898 359152 239134
rect 364847 239218 365083 239454
rect 364847 238898 365083 239134
rect 386916 239218 387152 239454
rect 386916 238898 387152 239134
rect 392847 239218 393083 239454
rect 392847 238898 393083 239134
rect 414916 239218 415152 239454
rect 414916 238898 415152 239134
rect 420847 239218 421083 239454
rect 420847 238898 421083 239134
rect 442916 239218 443152 239454
rect 442916 238898 443152 239134
rect 448847 239218 449083 239454
rect 448847 238898 449083 239134
rect 470916 239218 471152 239454
rect 470916 238898 471152 239134
rect 476847 239218 477083 239454
rect 476847 238898 477083 239134
rect 498916 239218 499152 239454
rect 498916 238898 499152 239134
rect 504847 239218 505083 239454
rect 504847 238898 505083 239134
rect 526916 239218 527152 239454
rect 526916 238898 527152 239134
rect 532847 239218 533083 239454
rect 532847 238898 533083 239134
rect 554916 239218 555152 239454
rect 554916 238898 555152 239134
rect 560847 239218 561083 239454
rect 560847 238898 561083 239134
rect -1974 215593 -1738 215829
rect -1654 215593 -1418 215829
rect -1974 215273 -1738 215509
rect -1654 215273 -1418 215509
rect 19951 215593 20187 215829
rect 19951 215273 20187 215509
rect 25882 215593 26118 215829
rect 25882 215273 26118 215509
rect 31812 215593 32048 215829
rect 31812 215273 32048 215509
rect 47951 215593 48187 215829
rect 47951 215273 48187 215509
rect 53882 215593 54118 215829
rect 53882 215273 54118 215509
rect 59812 215593 60048 215829
rect 59812 215273 60048 215509
rect 75951 215593 76187 215829
rect 75951 215273 76187 215509
rect 81882 215593 82118 215829
rect 81882 215273 82118 215509
rect 87812 215593 88048 215829
rect 87812 215273 88048 215509
rect 103951 215593 104187 215829
rect 103951 215273 104187 215509
rect 109882 215593 110118 215829
rect 109882 215273 110118 215509
rect 115812 215593 116048 215829
rect 115812 215273 116048 215509
rect 131951 215593 132187 215829
rect 131951 215273 132187 215509
rect 137882 215593 138118 215829
rect 137882 215273 138118 215509
rect 143812 215593 144048 215829
rect 143812 215273 144048 215509
rect 159951 215593 160187 215829
rect 159951 215273 160187 215509
rect 165882 215593 166118 215829
rect 165882 215273 166118 215509
rect 171812 215593 172048 215829
rect 171812 215273 172048 215509
rect 187951 215593 188187 215829
rect 187951 215273 188187 215509
rect 193882 215593 194118 215829
rect 193882 215273 194118 215509
rect 199812 215593 200048 215829
rect 199812 215273 200048 215509
rect 215951 215593 216187 215829
rect 215951 215273 216187 215509
rect 221882 215593 222118 215829
rect 221882 215273 222118 215509
rect 227812 215593 228048 215829
rect 227812 215273 228048 215509
rect 243951 215593 244187 215829
rect 243951 215273 244187 215509
rect 249882 215593 250118 215829
rect 249882 215273 250118 215509
rect 255812 215593 256048 215829
rect 255812 215273 256048 215509
rect 271951 215593 272187 215829
rect 271951 215273 272187 215509
rect 277882 215593 278118 215829
rect 277882 215273 278118 215509
rect 283812 215593 284048 215829
rect 283812 215273 284048 215509
rect 299951 215593 300187 215829
rect 299951 215273 300187 215509
rect 305882 215593 306118 215829
rect 305882 215273 306118 215509
rect 311812 215593 312048 215829
rect 311812 215273 312048 215509
rect 327951 215593 328187 215829
rect 327951 215273 328187 215509
rect 333882 215593 334118 215829
rect 333882 215273 334118 215509
rect 339812 215593 340048 215829
rect 339812 215273 340048 215509
rect 355951 215593 356187 215829
rect 355951 215273 356187 215509
rect 361882 215593 362118 215829
rect 361882 215273 362118 215509
rect 367812 215593 368048 215829
rect 367812 215273 368048 215509
rect 383951 215593 384187 215829
rect 383951 215273 384187 215509
rect 389882 215593 390118 215829
rect 389882 215273 390118 215509
rect 395812 215593 396048 215829
rect 395812 215273 396048 215509
rect 411951 215593 412187 215829
rect 411951 215273 412187 215509
rect 417882 215593 418118 215829
rect 417882 215273 418118 215509
rect 423812 215593 424048 215829
rect 423812 215273 424048 215509
rect 439951 215593 440187 215829
rect 439951 215273 440187 215509
rect 445882 215593 446118 215829
rect 445882 215273 446118 215509
rect 451812 215593 452048 215829
rect 451812 215273 452048 215509
rect 467951 215593 468187 215829
rect 467951 215273 468187 215509
rect 473882 215593 474118 215829
rect 473882 215273 474118 215509
rect 479812 215593 480048 215829
rect 479812 215273 480048 215509
rect 495951 215593 496187 215829
rect 495951 215273 496187 215509
rect 501882 215593 502118 215829
rect 501882 215273 502118 215509
rect 507812 215593 508048 215829
rect 507812 215273 508048 215509
rect 523951 215593 524187 215829
rect 523951 215273 524187 215509
rect 529882 215593 530118 215829
rect 529882 215273 530118 215509
rect 535812 215593 536048 215829
rect 535812 215273 536048 215509
rect 551951 215593 552187 215829
rect 551951 215273 552187 215509
rect 557882 215593 558118 215829
rect 557882 215273 558118 215509
rect 563812 215593 564048 215829
rect 563812 215273 564048 215509
rect 573526 215593 573762 215829
rect 573846 215593 574082 215829
rect 573526 215273 573762 215509
rect 573846 215273 574082 215509
rect 22917 212218 23153 212454
rect 22917 211898 23153 212134
rect 28848 212218 29084 212454
rect 28848 211898 29084 212134
rect 50917 212218 51153 212454
rect 50917 211898 51153 212134
rect 56848 212218 57084 212454
rect 56848 211898 57084 212134
rect 78917 212218 79153 212454
rect 78917 211898 79153 212134
rect 84848 212218 85084 212454
rect 84848 211898 85084 212134
rect 106917 212218 107153 212454
rect 106917 211898 107153 212134
rect 112848 212218 113084 212454
rect 112848 211898 113084 212134
rect 134917 212218 135153 212454
rect 134917 211898 135153 212134
rect 140848 212218 141084 212454
rect 140848 211898 141084 212134
rect 162917 212218 163153 212454
rect 162917 211898 163153 212134
rect 168848 212218 169084 212454
rect 168848 211898 169084 212134
rect 190917 212218 191153 212454
rect 190917 211898 191153 212134
rect 196848 212218 197084 212454
rect 196848 211898 197084 212134
rect 218917 212218 219153 212454
rect 218917 211898 219153 212134
rect 224848 212218 225084 212454
rect 224848 211898 225084 212134
rect 246917 212218 247153 212454
rect 246917 211898 247153 212134
rect 252848 212218 253084 212454
rect 252848 211898 253084 212134
rect 274917 212218 275153 212454
rect 274917 211898 275153 212134
rect 280848 212218 281084 212454
rect 280848 211898 281084 212134
rect 302917 212218 303153 212454
rect 302917 211898 303153 212134
rect 308848 212218 309084 212454
rect 308848 211898 309084 212134
rect 330917 212218 331153 212454
rect 330917 211898 331153 212134
rect 336848 212218 337084 212454
rect 336848 211898 337084 212134
rect 358917 212218 359153 212454
rect 358917 211898 359153 212134
rect 364848 212218 365084 212454
rect 364848 211898 365084 212134
rect 386917 212218 387153 212454
rect 386917 211898 387153 212134
rect 392848 212218 393084 212454
rect 392848 211898 393084 212134
rect 414917 212218 415153 212454
rect 414917 211898 415153 212134
rect 420848 212218 421084 212454
rect 420848 211898 421084 212134
rect 442917 212218 443153 212454
rect 442917 211898 443153 212134
rect 448848 212218 449084 212454
rect 448848 211898 449084 212134
rect 470917 212218 471153 212454
rect 470917 211898 471153 212134
rect 476848 212218 477084 212454
rect 476848 211898 477084 212134
rect 498917 212218 499153 212454
rect 498917 211898 499153 212134
rect 504848 212218 505084 212454
rect 504848 211898 505084 212134
rect 526917 212218 527153 212454
rect 526917 211898 527153 212134
rect 532848 212218 533084 212454
rect 532848 211898 533084 212134
rect 554917 212218 555153 212454
rect 554917 211898 555153 212134
rect 560848 212218 561084 212454
rect 560848 211898 561084 212134
rect -1974 188593 -1738 188829
rect -1654 188593 -1418 188829
rect -1974 188273 -1738 188509
rect -1654 188273 -1418 188509
rect 19952 188593 20188 188829
rect 19952 188273 20188 188509
rect 25882 188593 26118 188829
rect 25882 188273 26118 188509
rect 31813 188593 32049 188829
rect 31813 188273 32049 188509
rect 47952 188593 48188 188829
rect 47952 188273 48188 188509
rect 53882 188593 54118 188829
rect 53882 188273 54118 188509
rect 59813 188593 60049 188829
rect 59813 188273 60049 188509
rect 75952 188593 76188 188829
rect 75952 188273 76188 188509
rect 81882 188593 82118 188829
rect 81882 188273 82118 188509
rect 87813 188593 88049 188829
rect 87813 188273 88049 188509
rect 103952 188593 104188 188829
rect 103952 188273 104188 188509
rect 109882 188593 110118 188829
rect 109882 188273 110118 188509
rect 115813 188593 116049 188829
rect 115813 188273 116049 188509
rect 131952 188593 132188 188829
rect 131952 188273 132188 188509
rect 137882 188593 138118 188829
rect 137882 188273 138118 188509
rect 143813 188593 144049 188829
rect 143813 188273 144049 188509
rect 159952 188593 160188 188829
rect 159952 188273 160188 188509
rect 165882 188593 166118 188829
rect 165882 188273 166118 188509
rect 171813 188593 172049 188829
rect 171813 188273 172049 188509
rect 187952 188593 188188 188829
rect 187952 188273 188188 188509
rect 193882 188593 194118 188829
rect 193882 188273 194118 188509
rect 199813 188593 200049 188829
rect 199813 188273 200049 188509
rect 215952 188593 216188 188829
rect 215952 188273 216188 188509
rect 221882 188593 222118 188829
rect 221882 188273 222118 188509
rect 227813 188593 228049 188829
rect 227813 188273 228049 188509
rect 243952 188593 244188 188829
rect 243952 188273 244188 188509
rect 249882 188593 250118 188829
rect 249882 188273 250118 188509
rect 255813 188593 256049 188829
rect 255813 188273 256049 188509
rect 271952 188593 272188 188829
rect 271952 188273 272188 188509
rect 277882 188593 278118 188829
rect 277882 188273 278118 188509
rect 283813 188593 284049 188829
rect 283813 188273 284049 188509
rect 299952 188593 300188 188829
rect 299952 188273 300188 188509
rect 305882 188593 306118 188829
rect 305882 188273 306118 188509
rect 311813 188593 312049 188829
rect 311813 188273 312049 188509
rect 327952 188593 328188 188829
rect 327952 188273 328188 188509
rect 333882 188593 334118 188829
rect 333882 188273 334118 188509
rect 339813 188593 340049 188829
rect 339813 188273 340049 188509
rect 355952 188593 356188 188829
rect 355952 188273 356188 188509
rect 361882 188593 362118 188829
rect 361882 188273 362118 188509
rect 367813 188593 368049 188829
rect 367813 188273 368049 188509
rect 383952 188593 384188 188829
rect 383952 188273 384188 188509
rect 389882 188593 390118 188829
rect 389882 188273 390118 188509
rect 395813 188593 396049 188829
rect 395813 188273 396049 188509
rect 411952 188593 412188 188829
rect 411952 188273 412188 188509
rect 417882 188593 418118 188829
rect 417882 188273 418118 188509
rect 423813 188593 424049 188829
rect 423813 188273 424049 188509
rect 439952 188593 440188 188829
rect 439952 188273 440188 188509
rect 445882 188593 446118 188829
rect 445882 188273 446118 188509
rect 451813 188593 452049 188829
rect 451813 188273 452049 188509
rect 467952 188593 468188 188829
rect 467952 188273 468188 188509
rect 473882 188593 474118 188829
rect 473882 188273 474118 188509
rect 479813 188593 480049 188829
rect 479813 188273 480049 188509
rect 495952 188593 496188 188829
rect 495952 188273 496188 188509
rect 501882 188593 502118 188829
rect 501882 188273 502118 188509
rect 507813 188593 508049 188829
rect 507813 188273 508049 188509
rect 523952 188593 524188 188829
rect 523952 188273 524188 188509
rect 529882 188593 530118 188829
rect 529882 188273 530118 188509
rect 535813 188593 536049 188829
rect 535813 188273 536049 188509
rect 551952 188593 552188 188829
rect 551952 188273 552188 188509
rect 557882 188593 558118 188829
rect 557882 188273 558118 188509
rect 563813 188593 564049 188829
rect 563813 188273 564049 188509
rect 573526 188593 573762 188829
rect 573846 188593 574082 188829
rect 573526 188273 573762 188509
rect 573846 188273 574082 188509
rect 22916 185218 23152 185454
rect 22916 184898 23152 185134
rect 28847 185218 29083 185454
rect 28847 184898 29083 185134
rect 50916 185218 51152 185454
rect 50916 184898 51152 185134
rect 56847 185218 57083 185454
rect 56847 184898 57083 185134
rect 78916 185218 79152 185454
rect 78916 184898 79152 185134
rect 84847 185218 85083 185454
rect 84847 184898 85083 185134
rect 106916 185218 107152 185454
rect 106916 184898 107152 185134
rect 112847 185218 113083 185454
rect 112847 184898 113083 185134
rect 134916 185218 135152 185454
rect 134916 184898 135152 185134
rect 140847 185218 141083 185454
rect 140847 184898 141083 185134
rect 162916 185218 163152 185454
rect 162916 184898 163152 185134
rect 168847 185218 169083 185454
rect 168847 184898 169083 185134
rect 190916 185218 191152 185454
rect 190916 184898 191152 185134
rect 196847 185218 197083 185454
rect 196847 184898 197083 185134
rect 218916 185218 219152 185454
rect 218916 184898 219152 185134
rect 224847 185218 225083 185454
rect 224847 184898 225083 185134
rect 246916 185218 247152 185454
rect 246916 184898 247152 185134
rect 252847 185218 253083 185454
rect 252847 184898 253083 185134
rect 274916 185218 275152 185454
rect 274916 184898 275152 185134
rect 280847 185218 281083 185454
rect 280847 184898 281083 185134
rect 302916 185218 303152 185454
rect 302916 184898 303152 185134
rect 308847 185218 309083 185454
rect 308847 184898 309083 185134
rect 330916 185218 331152 185454
rect 330916 184898 331152 185134
rect 336847 185218 337083 185454
rect 336847 184898 337083 185134
rect 358916 185218 359152 185454
rect 358916 184898 359152 185134
rect 364847 185218 365083 185454
rect 364847 184898 365083 185134
rect 386916 185218 387152 185454
rect 386916 184898 387152 185134
rect 392847 185218 393083 185454
rect 392847 184898 393083 185134
rect 414916 185218 415152 185454
rect 414916 184898 415152 185134
rect 420847 185218 421083 185454
rect 420847 184898 421083 185134
rect 442916 185218 443152 185454
rect 442916 184898 443152 185134
rect 448847 185218 449083 185454
rect 448847 184898 449083 185134
rect 470916 185218 471152 185454
rect 470916 184898 471152 185134
rect 476847 185218 477083 185454
rect 476847 184898 477083 185134
rect 498916 185218 499152 185454
rect 498916 184898 499152 185134
rect 504847 185218 505083 185454
rect 504847 184898 505083 185134
rect 526916 185218 527152 185454
rect 526916 184898 527152 185134
rect 532847 185218 533083 185454
rect 532847 184898 533083 185134
rect 554916 185218 555152 185454
rect 554916 184898 555152 185134
rect 560847 185218 561083 185454
rect 560847 184898 561083 185134
rect -1974 161593 -1738 161829
rect -1654 161593 -1418 161829
rect -1974 161273 -1738 161509
rect -1654 161273 -1418 161509
rect 19951 161593 20187 161829
rect 19951 161273 20187 161509
rect 25882 161593 26118 161829
rect 25882 161273 26118 161509
rect 31812 161593 32048 161829
rect 31812 161273 32048 161509
rect 47951 161593 48187 161829
rect 47951 161273 48187 161509
rect 53882 161593 54118 161829
rect 53882 161273 54118 161509
rect 59812 161593 60048 161829
rect 59812 161273 60048 161509
rect 75951 161593 76187 161829
rect 75951 161273 76187 161509
rect 81882 161593 82118 161829
rect 81882 161273 82118 161509
rect 87812 161593 88048 161829
rect 87812 161273 88048 161509
rect 103951 161593 104187 161829
rect 103951 161273 104187 161509
rect 109882 161593 110118 161829
rect 109882 161273 110118 161509
rect 115812 161593 116048 161829
rect 115812 161273 116048 161509
rect 131951 161593 132187 161829
rect 131951 161273 132187 161509
rect 137882 161593 138118 161829
rect 137882 161273 138118 161509
rect 143812 161593 144048 161829
rect 143812 161273 144048 161509
rect 159951 161593 160187 161829
rect 159951 161273 160187 161509
rect 165882 161593 166118 161829
rect 165882 161273 166118 161509
rect 171812 161593 172048 161829
rect 171812 161273 172048 161509
rect 187951 161593 188187 161829
rect 187951 161273 188187 161509
rect 193882 161593 194118 161829
rect 193882 161273 194118 161509
rect 199812 161593 200048 161829
rect 199812 161273 200048 161509
rect 215951 161593 216187 161829
rect 215951 161273 216187 161509
rect 221882 161593 222118 161829
rect 221882 161273 222118 161509
rect 227812 161593 228048 161829
rect 227812 161273 228048 161509
rect 243951 161593 244187 161829
rect 243951 161273 244187 161509
rect 249882 161593 250118 161829
rect 249882 161273 250118 161509
rect 255812 161593 256048 161829
rect 255812 161273 256048 161509
rect 271951 161593 272187 161829
rect 271951 161273 272187 161509
rect 277882 161593 278118 161829
rect 277882 161273 278118 161509
rect 283812 161593 284048 161829
rect 283812 161273 284048 161509
rect 299951 161593 300187 161829
rect 299951 161273 300187 161509
rect 305882 161593 306118 161829
rect 305882 161273 306118 161509
rect 311812 161593 312048 161829
rect 311812 161273 312048 161509
rect 327951 161593 328187 161829
rect 327951 161273 328187 161509
rect 333882 161593 334118 161829
rect 333882 161273 334118 161509
rect 339812 161593 340048 161829
rect 339812 161273 340048 161509
rect 355951 161593 356187 161829
rect 355951 161273 356187 161509
rect 361882 161593 362118 161829
rect 361882 161273 362118 161509
rect 367812 161593 368048 161829
rect 367812 161273 368048 161509
rect 383951 161593 384187 161829
rect 383951 161273 384187 161509
rect 389882 161593 390118 161829
rect 389882 161273 390118 161509
rect 395812 161593 396048 161829
rect 395812 161273 396048 161509
rect 411951 161593 412187 161829
rect 411951 161273 412187 161509
rect 417882 161593 418118 161829
rect 417882 161273 418118 161509
rect 423812 161593 424048 161829
rect 423812 161273 424048 161509
rect 439951 161593 440187 161829
rect 439951 161273 440187 161509
rect 445882 161593 446118 161829
rect 445882 161273 446118 161509
rect 451812 161593 452048 161829
rect 451812 161273 452048 161509
rect 467951 161593 468187 161829
rect 467951 161273 468187 161509
rect 473882 161593 474118 161829
rect 473882 161273 474118 161509
rect 479812 161593 480048 161829
rect 479812 161273 480048 161509
rect 495951 161593 496187 161829
rect 495951 161273 496187 161509
rect 501882 161593 502118 161829
rect 501882 161273 502118 161509
rect 507812 161593 508048 161829
rect 507812 161273 508048 161509
rect 523951 161593 524187 161829
rect 523951 161273 524187 161509
rect 529882 161593 530118 161829
rect 529882 161273 530118 161509
rect 535812 161593 536048 161829
rect 535812 161273 536048 161509
rect 551951 161593 552187 161829
rect 551951 161273 552187 161509
rect 557882 161593 558118 161829
rect 557882 161273 558118 161509
rect 563812 161593 564048 161829
rect 563812 161273 564048 161509
rect 573526 161593 573762 161829
rect 573846 161593 574082 161829
rect 573526 161273 573762 161509
rect 573846 161273 574082 161509
rect 22917 158218 23153 158454
rect 22917 157898 23153 158134
rect 28848 158218 29084 158454
rect 28848 157898 29084 158134
rect 50917 158218 51153 158454
rect 50917 157898 51153 158134
rect 56848 158218 57084 158454
rect 56848 157898 57084 158134
rect 78917 158218 79153 158454
rect 78917 157898 79153 158134
rect 84848 158218 85084 158454
rect 84848 157898 85084 158134
rect 106917 158218 107153 158454
rect 106917 157898 107153 158134
rect 112848 158218 113084 158454
rect 112848 157898 113084 158134
rect 134917 158218 135153 158454
rect 134917 157898 135153 158134
rect 140848 158218 141084 158454
rect 140848 157898 141084 158134
rect 162917 158218 163153 158454
rect 162917 157898 163153 158134
rect 168848 158218 169084 158454
rect 168848 157898 169084 158134
rect 190917 158218 191153 158454
rect 190917 157898 191153 158134
rect 196848 158218 197084 158454
rect 196848 157898 197084 158134
rect 218917 158218 219153 158454
rect 218917 157898 219153 158134
rect 224848 158218 225084 158454
rect 224848 157898 225084 158134
rect 246917 158218 247153 158454
rect 246917 157898 247153 158134
rect 252848 158218 253084 158454
rect 252848 157898 253084 158134
rect 274917 158218 275153 158454
rect 274917 157898 275153 158134
rect 280848 158218 281084 158454
rect 280848 157898 281084 158134
rect 302917 158218 303153 158454
rect 302917 157898 303153 158134
rect 308848 158218 309084 158454
rect 308848 157898 309084 158134
rect 330917 158218 331153 158454
rect 330917 157898 331153 158134
rect 336848 158218 337084 158454
rect 336848 157898 337084 158134
rect 358917 158218 359153 158454
rect 358917 157898 359153 158134
rect 364848 158218 365084 158454
rect 364848 157898 365084 158134
rect 386917 158218 387153 158454
rect 386917 157898 387153 158134
rect 392848 158218 393084 158454
rect 392848 157898 393084 158134
rect 414917 158218 415153 158454
rect 414917 157898 415153 158134
rect 420848 158218 421084 158454
rect 420848 157898 421084 158134
rect 442917 158218 443153 158454
rect 442917 157898 443153 158134
rect 448848 158218 449084 158454
rect 448848 157898 449084 158134
rect 470917 158218 471153 158454
rect 470917 157898 471153 158134
rect 476848 158218 477084 158454
rect 476848 157898 477084 158134
rect 498917 158218 499153 158454
rect 498917 157898 499153 158134
rect 504848 158218 505084 158454
rect 504848 157898 505084 158134
rect 526917 158218 527153 158454
rect 526917 157898 527153 158134
rect 532848 158218 533084 158454
rect 532848 157898 533084 158134
rect 554917 158218 555153 158454
rect 554917 157898 555153 158134
rect 560848 158218 561084 158454
rect 560848 157898 561084 158134
rect -1974 134593 -1738 134829
rect -1654 134593 -1418 134829
rect -1974 134273 -1738 134509
rect -1654 134273 -1418 134509
rect 19952 134593 20188 134829
rect 19952 134273 20188 134509
rect 25882 134593 26118 134829
rect 25882 134273 26118 134509
rect 31813 134593 32049 134829
rect 31813 134273 32049 134509
rect 47952 134593 48188 134829
rect 47952 134273 48188 134509
rect 53882 134593 54118 134829
rect 53882 134273 54118 134509
rect 59813 134593 60049 134829
rect 59813 134273 60049 134509
rect 75952 134593 76188 134829
rect 75952 134273 76188 134509
rect 81882 134593 82118 134829
rect 81882 134273 82118 134509
rect 87813 134593 88049 134829
rect 87813 134273 88049 134509
rect 103952 134593 104188 134829
rect 103952 134273 104188 134509
rect 109882 134593 110118 134829
rect 109882 134273 110118 134509
rect 115813 134593 116049 134829
rect 115813 134273 116049 134509
rect 131952 134593 132188 134829
rect 131952 134273 132188 134509
rect 137882 134593 138118 134829
rect 137882 134273 138118 134509
rect 143813 134593 144049 134829
rect 143813 134273 144049 134509
rect 159952 134593 160188 134829
rect 159952 134273 160188 134509
rect 165882 134593 166118 134829
rect 165882 134273 166118 134509
rect 171813 134593 172049 134829
rect 171813 134273 172049 134509
rect 187952 134593 188188 134829
rect 187952 134273 188188 134509
rect 193882 134593 194118 134829
rect 193882 134273 194118 134509
rect 199813 134593 200049 134829
rect 199813 134273 200049 134509
rect 215952 134593 216188 134829
rect 215952 134273 216188 134509
rect 221882 134593 222118 134829
rect 221882 134273 222118 134509
rect 227813 134593 228049 134829
rect 227813 134273 228049 134509
rect 243952 134593 244188 134829
rect 243952 134273 244188 134509
rect 249882 134593 250118 134829
rect 249882 134273 250118 134509
rect 255813 134593 256049 134829
rect 255813 134273 256049 134509
rect 271952 134593 272188 134829
rect 271952 134273 272188 134509
rect 277882 134593 278118 134829
rect 277882 134273 278118 134509
rect 283813 134593 284049 134829
rect 283813 134273 284049 134509
rect 299952 134593 300188 134829
rect 299952 134273 300188 134509
rect 305882 134593 306118 134829
rect 305882 134273 306118 134509
rect 311813 134593 312049 134829
rect 311813 134273 312049 134509
rect 327952 134593 328188 134829
rect 327952 134273 328188 134509
rect 333882 134593 334118 134829
rect 333882 134273 334118 134509
rect 339813 134593 340049 134829
rect 339813 134273 340049 134509
rect 355952 134593 356188 134829
rect 355952 134273 356188 134509
rect 361882 134593 362118 134829
rect 361882 134273 362118 134509
rect 367813 134593 368049 134829
rect 367813 134273 368049 134509
rect 383952 134593 384188 134829
rect 383952 134273 384188 134509
rect 389882 134593 390118 134829
rect 389882 134273 390118 134509
rect 395813 134593 396049 134829
rect 395813 134273 396049 134509
rect 411952 134593 412188 134829
rect 411952 134273 412188 134509
rect 417882 134593 418118 134829
rect 417882 134273 418118 134509
rect 423813 134593 424049 134829
rect 423813 134273 424049 134509
rect 439952 134593 440188 134829
rect 439952 134273 440188 134509
rect 445882 134593 446118 134829
rect 445882 134273 446118 134509
rect 451813 134593 452049 134829
rect 451813 134273 452049 134509
rect 467952 134593 468188 134829
rect 467952 134273 468188 134509
rect 473882 134593 474118 134829
rect 473882 134273 474118 134509
rect 479813 134593 480049 134829
rect 479813 134273 480049 134509
rect 495952 134593 496188 134829
rect 495952 134273 496188 134509
rect 501882 134593 502118 134829
rect 501882 134273 502118 134509
rect 507813 134593 508049 134829
rect 507813 134273 508049 134509
rect 523952 134593 524188 134829
rect 523952 134273 524188 134509
rect 529882 134593 530118 134829
rect 529882 134273 530118 134509
rect 535813 134593 536049 134829
rect 535813 134273 536049 134509
rect 551952 134593 552188 134829
rect 551952 134273 552188 134509
rect 557882 134593 558118 134829
rect 557882 134273 558118 134509
rect 563813 134593 564049 134829
rect 563813 134273 564049 134509
rect 573526 134593 573762 134829
rect 573846 134593 574082 134829
rect 573526 134273 573762 134509
rect 573846 134273 574082 134509
rect 22916 131218 23152 131454
rect 22916 130898 23152 131134
rect 28847 131218 29083 131454
rect 28847 130898 29083 131134
rect 50916 131218 51152 131454
rect 50916 130898 51152 131134
rect 56847 131218 57083 131454
rect 56847 130898 57083 131134
rect 78916 131218 79152 131454
rect 78916 130898 79152 131134
rect 84847 131218 85083 131454
rect 84847 130898 85083 131134
rect 106916 131218 107152 131454
rect 106916 130898 107152 131134
rect 112847 131218 113083 131454
rect 112847 130898 113083 131134
rect 134916 131218 135152 131454
rect 134916 130898 135152 131134
rect 140847 131218 141083 131454
rect 140847 130898 141083 131134
rect 162916 131218 163152 131454
rect 162916 130898 163152 131134
rect 168847 131218 169083 131454
rect 168847 130898 169083 131134
rect 190916 131218 191152 131454
rect 190916 130898 191152 131134
rect 196847 131218 197083 131454
rect 196847 130898 197083 131134
rect 218916 131218 219152 131454
rect 218916 130898 219152 131134
rect 224847 131218 225083 131454
rect 224847 130898 225083 131134
rect 246916 131218 247152 131454
rect 246916 130898 247152 131134
rect 252847 131218 253083 131454
rect 252847 130898 253083 131134
rect 274916 131218 275152 131454
rect 274916 130898 275152 131134
rect 280847 131218 281083 131454
rect 280847 130898 281083 131134
rect 302916 131218 303152 131454
rect 302916 130898 303152 131134
rect 308847 131218 309083 131454
rect 308847 130898 309083 131134
rect 330916 131218 331152 131454
rect 330916 130898 331152 131134
rect 336847 131218 337083 131454
rect 336847 130898 337083 131134
rect 358916 131218 359152 131454
rect 358916 130898 359152 131134
rect 364847 131218 365083 131454
rect 364847 130898 365083 131134
rect 386916 131218 387152 131454
rect 386916 130898 387152 131134
rect 392847 131218 393083 131454
rect 392847 130898 393083 131134
rect 414916 131218 415152 131454
rect 414916 130898 415152 131134
rect 420847 131218 421083 131454
rect 420847 130898 421083 131134
rect 442916 131218 443152 131454
rect 442916 130898 443152 131134
rect 448847 131218 449083 131454
rect 448847 130898 449083 131134
rect 470916 131218 471152 131454
rect 470916 130898 471152 131134
rect 476847 131218 477083 131454
rect 476847 130898 477083 131134
rect 498916 131218 499152 131454
rect 498916 130898 499152 131134
rect 504847 131218 505083 131454
rect 504847 130898 505083 131134
rect 526916 131218 527152 131454
rect 526916 130898 527152 131134
rect 532847 131218 533083 131454
rect 532847 130898 533083 131134
rect 554916 131218 555152 131454
rect 554916 130898 555152 131134
rect 560847 131218 561083 131454
rect 560847 130898 561083 131134
rect -1974 107593 -1738 107829
rect -1654 107593 -1418 107829
rect -1974 107273 -1738 107509
rect -1654 107273 -1418 107509
rect 19951 107593 20187 107829
rect 19951 107273 20187 107509
rect 25882 107593 26118 107829
rect 25882 107273 26118 107509
rect 31812 107593 32048 107829
rect 31812 107273 32048 107509
rect 47951 107593 48187 107829
rect 47951 107273 48187 107509
rect 53882 107593 54118 107829
rect 53882 107273 54118 107509
rect 59812 107593 60048 107829
rect 59812 107273 60048 107509
rect 75951 107593 76187 107829
rect 75951 107273 76187 107509
rect 81882 107593 82118 107829
rect 81882 107273 82118 107509
rect 87812 107593 88048 107829
rect 87812 107273 88048 107509
rect 103951 107593 104187 107829
rect 103951 107273 104187 107509
rect 109882 107593 110118 107829
rect 109882 107273 110118 107509
rect 115812 107593 116048 107829
rect 115812 107273 116048 107509
rect 131210 107593 131446 107829
rect 131210 107273 131446 107509
rect 135658 107593 135894 107829
rect 135658 107273 135894 107509
rect 140106 107593 140342 107829
rect 140106 107273 140342 107509
rect 144554 107593 144790 107829
rect 144554 107273 144790 107509
rect 159951 107593 160187 107829
rect 159951 107273 160187 107509
rect 165882 107593 166118 107829
rect 165882 107273 166118 107509
rect 171812 107593 172048 107829
rect 171812 107273 172048 107509
rect 187951 107593 188187 107829
rect 187951 107273 188187 107509
rect 193882 107593 194118 107829
rect 193882 107273 194118 107509
rect 199812 107593 200048 107829
rect 199812 107273 200048 107509
rect 215210 107593 215446 107829
rect 215210 107273 215446 107509
rect 219658 107593 219894 107829
rect 219658 107273 219894 107509
rect 224106 107593 224342 107829
rect 224106 107273 224342 107509
rect 228554 107593 228790 107829
rect 228554 107273 228790 107509
rect 243951 107593 244187 107829
rect 243951 107273 244187 107509
rect 249882 107593 250118 107829
rect 249882 107273 250118 107509
rect 255812 107593 256048 107829
rect 255812 107273 256048 107509
rect 271951 107593 272187 107829
rect 271951 107273 272187 107509
rect 277882 107593 278118 107829
rect 277882 107273 278118 107509
rect 283812 107593 284048 107829
rect 283812 107273 284048 107509
rect 299951 107593 300187 107829
rect 299951 107273 300187 107509
rect 305882 107593 306118 107829
rect 305882 107273 306118 107509
rect 311812 107593 312048 107829
rect 311812 107273 312048 107509
rect 327951 107593 328187 107829
rect 327951 107273 328187 107509
rect 333882 107593 334118 107829
rect 333882 107273 334118 107509
rect 339812 107593 340048 107829
rect 339812 107273 340048 107509
rect 355951 107593 356187 107829
rect 355951 107273 356187 107509
rect 361882 107593 362118 107829
rect 361882 107273 362118 107509
rect 367812 107593 368048 107829
rect 367812 107273 368048 107509
rect 383951 107593 384187 107829
rect 383951 107273 384187 107509
rect 389882 107593 390118 107829
rect 389882 107273 390118 107509
rect 395812 107593 396048 107829
rect 395812 107273 396048 107509
rect 411951 107593 412187 107829
rect 411951 107273 412187 107509
rect 417882 107593 418118 107829
rect 417882 107273 418118 107509
rect 423812 107593 424048 107829
rect 423812 107273 424048 107509
rect 439951 107593 440187 107829
rect 439951 107273 440187 107509
rect 445882 107593 446118 107829
rect 445882 107273 446118 107509
rect 451812 107593 452048 107829
rect 451812 107273 452048 107509
rect 467951 107593 468187 107829
rect 467951 107273 468187 107509
rect 473882 107593 474118 107829
rect 473882 107273 474118 107509
rect 479812 107593 480048 107829
rect 479812 107273 480048 107509
rect 495951 107593 496187 107829
rect 495951 107273 496187 107509
rect 501882 107593 502118 107829
rect 501882 107273 502118 107509
rect 507812 107593 508048 107829
rect 507812 107273 508048 107509
rect 523951 107593 524187 107829
rect 523951 107273 524187 107509
rect 529882 107593 530118 107829
rect 529882 107273 530118 107509
rect 535812 107593 536048 107829
rect 535812 107273 536048 107509
rect 551951 107593 552187 107829
rect 551951 107273 552187 107509
rect 557882 107593 558118 107829
rect 557882 107273 558118 107509
rect 563812 107593 564048 107829
rect 563812 107273 564048 107509
rect 573526 107593 573762 107829
rect 573846 107593 574082 107829
rect 573526 107273 573762 107509
rect 573846 107273 574082 107509
rect 22917 104218 23153 104454
rect 22917 103898 23153 104134
rect 28848 104218 29084 104454
rect 28848 103898 29084 104134
rect 50917 104218 51153 104454
rect 50917 103898 51153 104134
rect 56848 104218 57084 104454
rect 56848 103898 57084 104134
rect 78917 104218 79153 104454
rect 78917 103898 79153 104134
rect 84848 104218 85084 104454
rect 84848 103898 85084 104134
rect 106917 104218 107153 104454
rect 106917 103898 107153 104134
rect 112848 104218 113084 104454
rect 112848 103898 113084 104134
rect 133434 104218 133670 104454
rect 133434 103898 133670 104134
rect 137882 104218 138118 104454
rect 137882 103898 138118 104134
rect 142330 104218 142566 104454
rect 142330 103898 142566 104134
rect 162917 104218 163153 104454
rect 162917 103898 163153 104134
rect 168848 104218 169084 104454
rect 168848 103898 169084 104134
rect 190917 104218 191153 104454
rect 190917 103898 191153 104134
rect 196848 104218 197084 104454
rect 196848 103898 197084 104134
rect 217434 104218 217670 104454
rect 217434 103898 217670 104134
rect 221882 104218 222118 104454
rect 221882 103898 222118 104134
rect 226330 104218 226566 104454
rect 226330 103898 226566 104134
rect 246917 104218 247153 104454
rect 246917 103898 247153 104134
rect 252848 104218 253084 104454
rect 252848 103898 253084 104134
rect 274917 104218 275153 104454
rect 274917 103898 275153 104134
rect 280848 104218 281084 104454
rect 280848 103898 281084 104134
rect 302917 104218 303153 104454
rect 302917 103898 303153 104134
rect 308848 104218 309084 104454
rect 308848 103898 309084 104134
rect 330917 104218 331153 104454
rect 330917 103898 331153 104134
rect 336848 104218 337084 104454
rect 336848 103898 337084 104134
rect 358917 104218 359153 104454
rect 358917 103898 359153 104134
rect 364848 104218 365084 104454
rect 364848 103898 365084 104134
rect 386917 104218 387153 104454
rect 386917 103898 387153 104134
rect 392848 104218 393084 104454
rect 392848 103898 393084 104134
rect 414917 104218 415153 104454
rect 414917 103898 415153 104134
rect 420848 104218 421084 104454
rect 420848 103898 421084 104134
rect 442917 104218 443153 104454
rect 442917 103898 443153 104134
rect 448848 104218 449084 104454
rect 448848 103898 449084 104134
rect 470917 104218 471153 104454
rect 470917 103898 471153 104134
rect 476848 104218 477084 104454
rect 476848 103898 477084 104134
rect 498917 104218 499153 104454
rect 498917 103898 499153 104134
rect 504848 104218 505084 104454
rect 504848 103898 505084 104134
rect 526917 104218 527153 104454
rect 526917 103898 527153 104134
rect 532848 104218 533084 104454
rect 532848 103898 533084 104134
rect 554917 104218 555153 104454
rect 554917 103898 555153 104134
rect 560848 104218 561084 104454
rect 560848 103898 561084 104134
rect -1974 80593 -1738 80829
rect -1654 80593 -1418 80829
rect -1974 80273 -1738 80509
rect -1654 80273 -1418 80509
rect 19952 80593 20188 80829
rect 19952 80273 20188 80509
rect 25882 80593 26118 80829
rect 25882 80273 26118 80509
rect 31813 80593 32049 80829
rect 31813 80273 32049 80509
rect 47952 80593 48188 80829
rect 47952 80273 48188 80509
rect 53882 80593 54118 80829
rect 53882 80273 54118 80509
rect 59813 80593 60049 80829
rect 59813 80273 60049 80509
rect 75952 80593 76188 80829
rect 75952 80273 76188 80509
rect 81882 80593 82118 80829
rect 81882 80273 82118 80509
rect 87813 80593 88049 80829
rect 87813 80273 88049 80509
rect 103952 80593 104188 80829
rect 103952 80273 104188 80509
rect 109882 80593 110118 80829
rect 109882 80273 110118 80509
rect 115813 80593 116049 80829
rect 115813 80273 116049 80509
rect 131952 80593 132188 80829
rect 131952 80273 132188 80509
rect 137882 80593 138118 80829
rect 137882 80273 138118 80509
rect 143813 80593 144049 80829
rect 143813 80273 144049 80509
rect 159952 80593 160188 80829
rect 159952 80273 160188 80509
rect 165882 80593 166118 80829
rect 165882 80273 166118 80509
rect 171813 80593 172049 80829
rect 171813 80273 172049 80509
rect 187952 80593 188188 80829
rect 187952 80273 188188 80509
rect 193882 80593 194118 80829
rect 193882 80273 194118 80509
rect 199813 80593 200049 80829
rect 199813 80273 200049 80509
rect 215952 80593 216188 80829
rect 215952 80273 216188 80509
rect 221882 80593 222118 80829
rect 221882 80273 222118 80509
rect 227813 80593 228049 80829
rect 227813 80273 228049 80509
rect 243952 80593 244188 80829
rect 243952 80273 244188 80509
rect 249882 80593 250118 80829
rect 249882 80273 250118 80509
rect 255813 80593 256049 80829
rect 255813 80273 256049 80509
rect 271952 80593 272188 80829
rect 271952 80273 272188 80509
rect 277882 80593 278118 80829
rect 277882 80273 278118 80509
rect 283813 80593 284049 80829
rect 283813 80273 284049 80509
rect 299952 80593 300188 80829
rect 299952 80273 300188 80509
rect 305882 80593 306118 80829
rect 305882 80273 306118 80509
rect 311813 80593 312049 80829
rect 311813 80273 312049 80509
rect 327952 80593 328188 80829
rect 327952 80273 328188 80509
rect 333882 80593 334118 80829
rect 333882 80273 334118 80509
rect 339813 80593 340049 80829
rect 339813 80273 340049 80509
rect 355952 80593 356188 80829
rect 355952 80273 356188 80509
rect 361882 80593 362118 80829
rect 361882 80273 362118 80509
rect 367813 80593 368049 80829
rect 367813 80273 368049 80509
rect 383952 80593 384188 80829
rect 383952 80273 384188 80509
rect 389882 80593 390118 80829
rect 389882 80273 390118 80509
rect 395813 80593 396049 80829
rect 395813 80273 396049 80509
rect 411952 80593 412188 80829
rect 411952 80273 412188 80509
rect 417882 80593 418118 80829
rect 417882 80273 418118 80509
rect 423813 80593 424049 80829
rect 423813 80273 424049 80509
rect 439952 80593 440188 80829
rect 439952 80273 440188 80509
rect 445882 80593 446118 80829
rect 445882 80273 446118 80509
rect 451813 80593 452049 80829
rect 451813 80273 452049 80509
rect 467952 80593 468188 80829
rect 467952 80273 468188 80509
rect 473882 80593 474118 80829
rect 473882 80273 474118 80509
rect 479813 80593 480049 80829
rect 479813 80273 480049 80509
rect 495952 80593 496188 80829
rect 495952 80273 496188 80509
rect 501882 80593 502118 80829
rect 501882 80273 502118 80509
rect 507813 80593 508049 80829
rect 507813 80273 508049 80509
rect 523952 80593 524188 80829
rect 523952 80273 524188 80509
rect 529882 80593 530118 80829
rect 529882 80273 530118 80509
rect 535813 80593 536049 80829
rect 535813 80273 536049 80509
rect 551952 80593 552188 80829
rect 551952 80273 552188 80509
rect 557882 80593 558118 80829
rect 557882 80273 558118 80509
rect 563813 80593 564049 80829
rect 563813 80273 564049 80509
rect 573526 80593 573762 80829
rect 573846 80593 574082 80829
rect 573526 80273 573762 80509
rect 573846 80273 574082 80509
rect 22916 77218 23152 77454
rect 22916 76898 23152 77134
rect 28847 77218 29083 77454
rect 28847 76898 29083 77134
rect 50916 77218 51152 77454
rect 50916 76898 51152 77134
rect 56847 77218 57083 77454
rect 56847 76898 57083 77134
rect 78916 77218 79152 77454
rect 78916 76898 79152 77134
rect 84847 77218 85083 77454
rect 84847 76898 85083 77134
rect 106916 77218 107152 77454
rect 106916 76898 107152 77134
rect 112847 77218 113083 77454
rect 112847 76898 113083 77134
rect 134916 77218 135152 77454
rect 134916 76898 135152 77134
rect 140847 77218 141083 77454
rect 140847 76898 141083 77134
rect 162916 77218 163152 77454
rect 162916 76898 163152 77134
rect 168847 77218 169083 77454
rect 168847 76898 169083 77134
rect 190916 77218 191152 77454
rect 190916 76898 191152 77134
rect 196847 77218 197083 77454
rect 196847 76898 197083 77134
rect 218916 77218 219152 77454
rect 218916 76898 219152 77134
rect 224847 77218 225083 77454
rect 224847 76898 225083 77134
rect 246916 77218 247152 77454
rect 246916 76898 247152 77134
rect 252847 77218 253083 77454
rect 252847 76898 253083 77134
rect 274916 77218 275152 77454
rect 274916 76898 275152 77134
rect 280847 77218 281083 77454
rect 280847 76898 281083 77134
rect 302916 77218 303152 77454
rect 302916 76898 303152 77134
rect 308847 77218 309083 77454
rect 308847 76898 309083 77134
rect 330916 77218 331152 77454
rect 330916 76898 331152 77134
rect 336847 77218 337083 77454
rect 336847 76898 337083 77134
rect 358916 77218 359152 77454
rect 358916 76898 359152 77134
rect 364847 77218 365083 77454
rect 364847 76898 365083 77134
rect 386916 77218 387152 77454
rect 386916 76898 387152 77134
rect 392847 77218 393083 77454
rect 392847 76898 393083 77134
rect 414916 77218 415152 77454
rect 414916 76898 415152 77134
rect 420847 77218 421083 77454
rect 420847 76898 421083 77134
rect 442916 77218 443152 77454
rect 442916 76898 443152 77134
rect 448847 77218 449083 77454
rect 448847 76898 449083 77134
rect 470916 77218 471152 77454
rect 470916 76898 471152 77134
rect 476847 77218 477083 77454
rect 476847 76898 477083 77134
rect 498916 77218 499152 77454
rect 498916 76898 499152 77134
rect 504847 77218 505083 77454
rect 504847 76898 505083 77134
rect 526916 77218 527152 77454
rect 526916 76898 527152 77134
rect 532847 77218 533083 77454
rect 532847 76898 533083 77134
rect 554916 77218 555152 77454
rect 554916 76898 555152 77134
rect 560847 77218 561083 77454
rect 560847 76898 561083 77134
rect -1974 53593 -1738 53829
rect -1654 53593 -1418 53829
rect -1974 53273 -1738 53509
rect -1654 53273 -1418 53509
rect 19951 53593 20187 53829
rect 19951 53273 20187 53509
rect 25882 53593 26118 53829
rect 25882 53273 26118 53509
rect 31812 53593 32048 53829
rect 31812 53273 32048 53509
rect 47951 53593 48187 53829
rect 47951 53273 48187 53509
rect 53882 53593 54118 53829
rect 53882 53273 54118 53509
rect 59812 53593 60048 53829
rect 59812 53273 60048 53509
rect 75951 53593 76187 53829
rect 75951 53273 76187 53509
rect 81882 53593 82118 53829
rect 81882 53273 82118 53509
rect 87812 53593 88048 53829
rect 87812 53273 88048 53509
rect 103951 53593 104187 53829
rect 103951 53273 104187 53509
rect 109882 53593 110118 53829
rect 109882 53273 110118 53509
rect 115812 53593 116048 53829
rect 115812 53273 116048 53509
rect 131951 53593 132187 53829
rect 131951 53273 132187 53509
rect 137882 53593 138118 53829
rect 137882 53273 138118 53509
rect 143812 53593 144048 53829
rect 143812 53273 144048 53509
rect 159951 53593 160187 53829
rect 159951 53273 160187 53509
rect 165882 53593 166118 53829
rect 165882 53273 166118 53509
rect 171812 53593 172048 53829
rect 171812 53273 172048 53509
rect 187951 53593 188187 53829
rect 187951 53273 188187 53509
rect 193882 53593 194118 53829
rect 193882 53273 194118 53509
rect 199812 53593 200048 53829
rect 199812 53273 200048 53509
rect 215951 53593 216187 53829
rect 215951 53273 216187 53509
rect 221882 53593 222118 53829
rect 221882 53273 222118 53509
rect 227812 53593 228048 53829
rect 227812 53273 228048 53509
rect 243951 53593 244187 53829
rect 243951 53273 244187 53509
rect 249882 53593 250118 53829
rect 249882 53273 250118 53509
rect 255812 53593 256048 53829
rect 255812 53273 256048 53509
rect 271951 53593 272187 53829
rect 271951 53273 272187 53509
rect 277882 53593 278118 53829
rect 277882 53273 278118 53509
rect 283812 53593 284048 53829
rect 283812 53273 284048 53509
rect 299951 53593 300187 53829
rect 299951 53273 300187 53509
rect 305882 53593 306118 53829
rect 305882 53273 306118 53509
rect 311812 53593 312048 53829
rect 311812 53273 312048 53509
rect 327951 53593 328187 53829
rect 327951 53273 328187 53509
rect 333882 53593 334118 53829
rect 333882 53273 334118 53509
rect 339812 53593 340048 53829
rect 339812 53273 340048 53509
rect 355951 53593 356187 53829
rect 355951 53273 356187 53509
rect 361882 53593 362118 53829
rect 361882 53273 362118 53509
rect 367812 53593 368048 53829
rect 367812 53273 368048 53509
rect 383951 53593 384187 53829
rect 383951 53273 384187 53509
rect 389882 53593 390118 53829
rect 389882 53273 390118 53509
rect 395812 53593 396048 53829
rect 395812 53273 396048 53509
rect 411951 53593 412187 53829
rect 411951 53273 412187 53509
rect 417882 53593 418118 53829
rect 417882 53273 418118 53509
rect 423812 53593 424048 53829
rect 423812 53273 424048 53509
rect 439951 53593 440187 53829
rect 439951 53273 440187 53509
rect 445882 53593 446118 53829
rect 445882 53273 446118 53509
rect 451812 53593 452048 53829
rect 451812 53273 452048 53509
rect 467951 53593 468187 53829
rect 467951 53273 468187 53509
rect 473882 53593 474118 53829
rect 473882 53273 474118 53509
rect 479812 53593 480048 53829
rect 479812 53273 480048 53509
rect 495951 53593 496187 53829
rect 495951 53273 496187 53509
rect 501882 53593 502118 53829
rect 501882 53273 502118 53509
rect 507812 53593 508048 53829
rect 507812 53273 508048 53509
rect 523951 53593 524187 53829
rect 523951 53273 524187 53509
rect 529882 53593 530118 53829
rect 529882 53273 530118 53509
rect 535812 53593 536048 53829
rect 535812 53273 536048 53509
rect 551951 53593 552187 53829
rect 551951 53273 552187 53509
rect 557882 53593 558118 53829
rect 557882 53273 558118 53509
rect 563812 53593 564048 53829
rect 563812 53273 564048 53509
rect 573526 53593 573762 53829
rect 573846 53593 574082 53829
rect 573526 53273 573762 53509
rect 573846 53273 574082 53509
rect 22917 50218 23153 50454
rect 22917 49898 23153 50134
rect 28848 50218 29084 50454
rect 28848 49898 29084 50134
rect 50917 50218 51153 50454
rect 50917 49898 51153 50134
rect 56848 50218 57084 50454
rect 56848 49898 57084 50134
rect 78917 50218 79153 50454
rect 78917 49898 79153 50134
rect 84848 50218 85084 50454
rect 84848 49898 85084 50134
rect 106917 50218 107153 50454
rect 106917 49898 107153 50134
rect 112848 50218 113084 50454
rect 112848 49898 113084 50134
rect 134917 50218 135153 50454
rect 134917 49898 135153 50134
rect 140848 50218 141084 50454
rect 140848 49898 141084 50134
rect 162917 50218 163153 50454
rect 162917 49898 163153 50134
rect 168848 50218 169084 50454
rect 168848 49898 169084 50134
rect 190917 50218 191153 50454
rect 190917 49898 191153 50134
rect 196848 50218 197084 50454
rect 196848 49898 197084 50134
rect 218917 50218 219153 50454
rect 218917 49898 219153 50134
rect 224848 50218 225084 50454
rect 224848 49898 225084 50134
rect 246917 50218 247153 50454
rect 246917 49898 247153 50134
rect 252848 50218 253084 50454
rect 252848 49898 253084 50134
rect 274917 50218 275153 50454
rect 274917 49898 275153 50134
rect 280848 50218 281084 50454
rect 280848 49898 281084 50134
rect 302917 50218 303153 50454
rect 302917 49898 303153 50134
rect 308848 50218 309084 50454
rect 308848 49898 309084 50134
rect 330917 50218 331153 50454
rect 330917 49898 331153 50134
rect 336848 50218 337084 50454
rect 336848 49898 337084 50134
rect 358917 50218 359153 50454
rect 358917 49898 359153 50134
rect 364848 50218 365084 50454
rect 364848 49898 365084 50134
rect 386917 50218 387153 50454
rect 386917 49898 387153 50134
rect 392848 50218 393084 50454
rect 392848 49898 393084 50134
rect 414917 50218 415153 50454
rect 414917 49898 415153 50134
rect 420848 50218 421084 50454
rect 420848 49898 421084 50134
rect 442917 50218 443153 50454
rect 442917 49898 443153 50134
rect 448848 50218 449084 50454
rect 448848 49898 449084 50134
rect 470917 50218 471153 50454
rect 470917 49898 471153 50134
rect 476848 50218 477084 50454
rect 476848 49898 477084 50134
rect 498917 50218 499153 50454
rect 498917 49898 499153 50134
rect 504848 50218 505084 50454
rect 504848 49898 505084 50134
rect 526917 50218 527153 50454
rect 526917 49898 527153 50134
rect 532848 50218 533084 50454
rect 532848 49898 533084 50134
rect 554917 50218 555153 50454
rect 554917 49898 555153 50134
rect 560848 50218 561084 50454
rect 560848 49898 561084 50134
rect -1974 26593 -1738 26829
rect -1654 26593 -1418 26829
rect -1974 26273 -1738 26509
rect -1654 26273 -1418 26509
rect 22460 26593 22696 26829
rect 22460 26273 22696 26509
rect 33408 26593 33644 26829
rect 33408 26273 33644 26509
rect 27934 23218 28170 23454
rect 27934 22898 28170 23134
rect 38882 23218 39118 23454
rect 38882 22898 39118 23134
rect 44356 26593 44592 26829
rect 44356 26273 44592 26509
rect 55304 26593 55540 26829
rect 55304 26273 55540 26509
rect 49830 23218 50066 23454
rect 49830 22898 50066 23134
rect 60778 23218 61014 23454
rect 60778 22898 61014 23134
rect 75952 26593 76188 26829
rect 75952 26273 76188 26509
rect 81882 26593 82118 26829
rect 81882 26273 82118 26509
rect 87813 26593 88049 26829
rect 87813 26273 88049 26509
rect 103952 26593 104188 26829
rect 103952 26273 104188 26509
rect 109882 26593 110118 26829
rect 109882 26273 110118 26509
rect 115813 26593 116049 26829
rect 115813 26273 116049 26509
rect 131952 26593 132188 26829
rect 131952 26273 132188 26509
rect 137882 26593 138118 26829
rect 137882 26273 138118 26509
rect 143813 26593 144049 26829
rect 143813 26273 144049 26509
rect 159952 26593 160188 26829
rect 159952 26273 160188 26509
rect 165882 26593 166118 26829
rect 165882 26273 166118 26509
rect 171813 26593 172049 26829
rect 171813 26273 172049 26509
rect 187952 26593 188188 26829
rect 187952 26273 188188 26509
rect 193882 26593 194118 26829
rect 193882 26273 194118 26509
rect 199813 26593 200049 26829
rect 199813 26273 200049 26509
rect 215952 26593 216188 26829
rect 215952 26273 216188 26509
rect 221882 26593 222118 26829
rect 221882 26273 222118 26509
rect 227813 26593 228049 26829
rect 227813 26273 228049 26509
rect 243952 26593 244188 26829
rect 243952 26273 244188 26509
rect 249882 26593 250118 26829
rect 249882 26273 250118 26509
rect 255813 26593 256049 26829
rect 255813 26273 256049 26509
rect 271952 26593 272188 26829
rect 271952 26273 272188 26509
rect 277882 26593 278118 26829
rect 277882 26273 278118 26509
rect 283813 26593 284049 26829
rect 283813 26273 284049 26509
rect 299952 26593 300188 26829
rect 299952 26273 300188 26509
rect 305882 26593 306118 26829
rect 305882 26273 306118 26509
rect 311813 26593 312049 26829
rect 311813 26273 312049 26509
rect 327952 26593 328188 26829
rect 327952 26273 328188 26509
rect 333882 26593 334118 26829
rect 333882 26273 334118 26509
rect 339813 26593 340049 26829
rect 339813 26273 340049 26509
rect 355952 26593 356188 26829
rect 355952 26273 356188 26509
rect 361882 26593 362118 26829
rect 361882 26273 362118 26509
rect 367813 26593 368049 26829
rect 367813 26273 368049 26509
rect 383952 26593 384188 26829
rect 383952 26273 384188 26509
rect 389882 26593 390118 26829
rect 389882 26273 390118 26509
rect 395813 26593 396049 26829
rect 395813 26273 396049 26509
rect 411952 26593 412188 26829
rect 411952 26273 412188 26509
rect 417882 26593 418118 26829
rect 417882 26273 418118 26509
rect 423813 26593 424049 26829
rect 423813 26273 424049 26509
rect 439952 26593 440188 26829
rect 439952 26273 440188 26509
rect 445882 26593 446118 26829
rect 445882 26273 446118 26509
rect 451813 26593 452049 26829
rect 451813 26273 452049 26509
rect 467952 26593 468188 26829
rect 467952 26273 468188 26509
rect 473882 26593 474118 26829
rect 473882 26273 474118 26509
rect 479813 26593 480049 26829
rect 479813 26273 480049 26509
rect 495952 26593 496188 26829
rect 495952 26273 496188 26509
rect 501882 26593 502118 26829
rect 501882 26273 502118 26509
rect 507813 26593 508049 26829
rect 507813 26273 508049 26509
rect 523952 26593 524188 26829
rect 523952 26273 524188 26509
rect 529882 26593 530118 26829
rect 529882 26273 530118 26509
rect 535813 26593 536049 26829
rect 535813 26273 536049 26509
rect 551952 26593 552188 26829
rect 551952 26273 552188 26509
rect 557882 26593 558118 26829
rect 557882 26273 558118 26509
rect 563813 26593 564049 26829
rect 563813 26273 564049 26509
rect 573526 26593 573762 26829
rect 573846 26593 574082 26829
rect 573526 26273 573762 26509
rect 573846 26273 574082 26509
rect 66026 23218 66262 23454
rect 66346 23218 66582 23454
rect 66026 22898 66262 23134
rect 66346 22898 66582 23134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 78916 23218 79152 23454
rect 78916 22898 79152 23134
rect 84847 23218 85083 23454
rect 84847 22898 85083 23134
rect 106916 23218 107152 23454
rect 106916 22898 107152 23134
rect 112847 23218 113083 23454
rect 112847 22898 113083 23134
rect 134916 23218 135152 23454
rect 134916 22898 135152 23134
rect 140847 23218 141083 23454
rect 140847 22898 141083 23134
rect 162916 23218 163152 23454
rect 162916 22898 163152 23134
rect 168847 23218 169083 23454
rect 168847 22898 169083 23134
rect 190916 23218 191152 23454
rect 190916 22898 191152 23134
rect 196847 23218 197083 23454
rect 196847 22898 197083 23134
rect 218916 23218 219152 23454
rect 218916 22898 219152 23134
rect 224847 23218 225083 23454
rect 224847 22898 225083 23134
rect 246916 23218 247152 23454
rect 246916 22898 247152 23134
rect 252847 23218 253083 23454
rect 252847 22898 253083 23134
rect 274916 23218 275152 23454
rect 274916 22898 275152 23134
rect 280847 23218 281083 23454
rect 280847 22898 281083 23134
rect 302916 23218 303152 23454
rect 302916 22898 303152 23134
rect 308847 23218 309083 23454
rect 308847 22898 309083 23134
rect 330916 23218 331152 23454
rect 330916 22898 331152 23134
rect 336847 23218 337083 23454
rect 336847 22898 337083 23134
rect 358916 23218 359152 23454
rect 358916 22898 359152 23134
rect 364847 23218 365083 23454
rect 364847 22898 365083 23134
rect 386916 23218 387152 23454
rect 386916 22898 387152 23134
rect 392847 23218 393083 23454
rect 392847 22898 393083 23134
rect 414916 23218 415152 23454
rect 414916 22898 415152 23134
rect 420847 23218 421083 23454
rect 420847 22898 421083 23134
rect 442916 23218 443152 23454
rect 442916 22898 443152 23134
rect 448847 23218 449083 23454
rect 448847 22898 449083 23134
rect 470916 23218 471152 23454
rect 470916 22898 471152 23134
rect 476847 23218 477083 23454
rect 476847 22898 477083 23134
rect 498916 23218 499152 23454
rect 498916 22898 499152 23134
rect 504847 23218 505083 23454
rect 504847 22898 505083 23134
rect 526916 23218 527152 23454
rect 526916 22898 527152 23134
rect 532847 23218 533083 23454
rect 532847 22898 533083 23134
rect 554916 23218 555152 23454
rect 554916 22898 555152 23134
rect 560847 23218 561083 23454
rect 560847 22898 561083 23134
rect 66026 -1542 66262 -1306
rect 66346 -1542 66582 -1306
rect 66026 -1862 66262 -1626
rect 66346 -1862 66582 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 585342 647593 585578 647829
rect 585662 647593 585898 647829
rect 585342 647273 585578 647509
rect 585662 647273 585898 647509
rect 585342 620593 585578 620829
rect 585662 620593 585898 620829
rect 585342 620273 585578 620509
rect 585662 620273 585898 620509
rect 585342 593593 585578 593829
rect 585662 593593 585898 593829
rect 585342 593273 585578 593509
rect 585662 593273 585898 593509
rect 585342 566593 585578 566829
rect 585662 566593 585898 566829
rect 585342 566273 585578 566509
rect 585662 566273 585898 566509
rect 585342 539593 585578 539829
rect 585662 539593 585898 539829
rect 585342 539273 585578 539509
rect 585662 539273 585898 539509
rect 585342 512593 585578 512829
rect 585662 512593 585898 512829
rect 585342 512273 585578 512509
rect 585662 512273 585898 512509
rect 585342 485593 585578 485829
rect 585662 485593 585898 485829
rect 585342 485273 585578 485509
rect 585662 485273 585898 485509
rect 585342 458593 585578 458829
rect 585662 458593 585898 458829
rect 585342 458273 585578 458509
rect 585662 458273 585898 458509
rect 585342 431593 585578 431829
rect 585662 431593 585898 431829
rect 585342 431273 585578 431509
rect 585662 431273 585898 431509
rect 585342 404593 585578 404829
rect 585662 404593 585898 404829
rect 585342 404273 585578 404509
rect 585662 404273 585898 404509
rect 585342 377593 585578 377829
rect 585662 377593 585898 377829
rect 585342 377273 585578 377509
rect 585662 377273 585898 377509
rect 585342 350593 585578 350829
rect 585662 350593 585898 350829
rect 585342 350273 585578 350509
rect 585662 350273 585898 350509
rect 585342 323593 585578 323829
rect 585662 323593 585898 323829
rect 585342 323273 585578 323509
rect 585662 323273 585898 323509
rect 585342 296593 585578 296829
rect 585662 296593 585898 296829
rect 585342 296273 585578 296509
rect 585662 296273 585898 296509
rect 585342 269593 585578 269829
rect 585662 269593 585898 269829
rect 585342 269273 585578 269509
rect 585662 269273 585898 269509
rect 585342 242593 585578 242829
rect 585662 242593 585898 242829
rect 585342 242273 585578 242509
rect 585662 242273 585898 242509
rect 585342 215593 585578 215829
rect 585662 215593 585898 215829
rect 585342 215273 585578 215509
rect 585662 215273 585898 215509
rect 585342 188593 585578 188829
rect 585662 188593 585898 188829
rect 585342 188273 585578 188509
rect 585662 188273 585898 188509
rect 585342 161593 585578 161829
rect 585662 161593 585898 161829
rect 585342 161273 585578 161509
rect 585662 161273 585898 161509
rect 585342 134593 585578 134829
rect 585662 134593 585898 134829
rect 585342 134273 585578 134509
rect 585662 134273 585898 134509
rect 585342 107593 585578 107829
rect 585662 107593 585898 107829
rect 585342 107273 585578 107509
rect 585662 107273 585898 107509
rect 585342 80593 585578 80829
rect 585662 80593 585898 80829
rect 585342 80273 585578 80509
rect 585662 80273 585898 80509
rect 585342 53593 585578 53829
rect 585662 53593 585898 53829
rect 585342 53273 585578 53509
rect 585662 53273 585898 53509
rect 585342 26593 585578 26829
rect 585662 26593 585898 26829
rect 585342 26273 585578 26509
rect 585662 26273 585898 26509
rect 573526 -582 573762 -346
rect 573846 -582 574082 -346
rect 573526 -902 573762 -666
rect 573846 -902 574082 -666
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 698218 586538 698454
rect 586622 698218 586858 698454
rect 586302 697898 586538 698134
rect 586622 697898 586858 698134
rect 586302 671218 586538 671454
rect 586622 671218 586858 671454
rect 586302 670898 586538 671134
rect 586622 670898 586858 671134
rect 586302 644218 586538 644454
rect 586622 644218 586858 644454
rect 586302 643898 586538 644134
rect 586622 643898 586858 644134
rect 586302 617218 586538 617454
rect 586622 617218 586858 617454
rect 586302 616898 586538 617134
rect 586622 616898 586858 617134
rect 586302 590218 586538 590454
rect 586622 590218 586858 590454
rect 586302 589898 586538 590134
rect 586622 589898 586858 590134
rect 586302 563218 586538 563454
rect 586622 563218 586858 563454
rect 586302 562898 586538 563134
rect 586622 562898 586858 563134
rect 586302 536218 586538 536454
rect 586622 536218 586858 536454
rect 586302 535898 586538 536134
rect 586622 535898 586858 536134
rect 586302 509218 586538 509454
rect 586622 509218 586858 509454
rect 586302 508898 586538 509134
rect 586622 508898 586858 509134
rect 586302 482218 586538 482454
rect 586622 482218 586858 482454
rect 586302 481898 586538 482134
rect 586622 481898 586858 482134
rect 586302 455218 586538 455454
rect 586622 455218 586858 455454
rect 586302 454898 586538 455134
rect 586622 454898 586858 455134
rect 586302 428218 586538 428454
rect 586622 428218 586858 428454
rect 586302 427898 586538 428134
rect 586622 427898 586858 428134
rect 586302 401218 586538 401454
rect 586622 401218 586858 401454
rect 586302 400898 586538 401134
rect 586622 400898 586858 401134
rect 586302 374218 586538 374454
rect 586622 374218 586858 374454
rect 586302 373898 586538 374134
rect 586622 373898 586858 374134
rect 586302 347218 586538 347454
rect 586622 347218 586858 347454
rect 586302 346898 586538 347134
rect 586622 346898 586858 347134
rect 586302 320218 586538 320454
rect 586622 320218 586858 320454
rect 586302 319898 586538 320134
rect 586622 319898 586858 320134
rect 586302 293218 586538 293454
rect 586622 293218 586858 293454
rect 586302 292898 586538 293134
rect 586622 292898 586858 293134
rect 586302 266218 586538 266454
rect 586622 266218 586858 266454
rect 586302 265898 586538 266134
rect 586622 265898 586858 266134
rect 586302 239218 586538 239454
rect 586622 239218 586858 239454
rect 586302 238898 586538 239134
rect 586622 238898 586858 239134
rect 586302 212218 586538 212454
rect 586622 212218 586858 212454
rect 586302 211898 586538 212134
rect 586622 211898 586858 212134
rect 586302 185218 586538 185454
rect 586622 185218 586858 185454
rect 586302 184898 586538 185134
rect 586622 184898 586858 185134
rect 586302 158218 586538 158454
rect 586622 158218 586858 158454
rect 586302 157898 586538 158134
rect 586622 157898 586858 158134
rect 586302 131218 586538 131454
rect 586622 131218 586858 131454
rect 586302 130898 586538 131134
rect 586622 130898 586858 131134
rect 586302 104218 586538 104454
rect 586622 104218 586858 104454
rect 586302 103898 586538 104134
rect 586622 103898 586858 104134
rect 586302 77218 586538 77454
rect 586622 77218 586858 77454
rect 586302 76898 586538 77134
rect 586622 76898 586858 77134
rect 586302 50218 586538 50454
rect 586622 50218 586858 50454
rect 586302 49898 586538 50134
rect 586622 49898 586858 50134
rect 586302 23218 586538 23454
rect 586622 23218 586858 23454
rect 586302 22898 586538 23134
rect 586622 22898 586858 23134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 38026 705798
rect 38262 705562 38346 705798
rect 38582 705562 66026 705798
rect 66262 705562 66346 705798
rect 66582 705562 94026 705798
rect 94262 705562 94346 705798
rect 94582 705562 122026 705798
rect 122262 705562 122346 705798
rect 122582 705562 150026 705798
rect 150262 705562 150346 705798
rect 150582 705562 178026 705798
rect 178262 705562 178346 705798
rect 178582 705562 206026 705798
rect 206262 705562 206346 705798
rect 206582 705562 234026 705798
rect 234262 705562 234346 705798
rect 234582 705562 262026 705798
rect 262262 705562 262346 705798
rect 262582 705562 290026 705798
rect 290262 705562 290346 705798
rect 290582 705562 318026 705798
rect 318262 705562 318346 705798
rect 318582 705562 346026 705798
rect 346262 705562 346346 705798
rect 346582 705562 374026 705798
rect 374262 705562 374346 705798
rect 374582 705562 402026 705798
rect 402262 705562 402346 705798
rect 402582 705562 430026 705798
rect 430262 705562 430346 705798
rect 430582 705562 458026 705798
rect 458262 705562 458346 705798
rect 458582 705562 486026 705798
rect 486262 705562 486346 705798
rect 486582 705562 514026 705798
rect 514262 705562 514346 705798
rect 514582 705562 542026 705798
rect 542262 705562 542346 705798
rect 542582 705562 570026 705798
rect 570262 705562 570346 705798
rect 570582 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 38026 705478
rect 38262 705242 38346 705478
rect 38582 705242 66026 705478
rect 66262 705242 66346 705478
rect 66582 705242 94026 705478
rect 94262 705242 94346 705478
rect 94582 705242 122026 705478
rect 122262 705242 122346 705478
rect 122582 705242 150026 705478
rect 150262 705242 150346 705478
rect 150582 705242 178026 705478
rect 178262 705242 178346 705478
rect 178582 705242 206026 705478
rect 206262 705242 206346 705478
rect 206582 705242 234026 705478
rect 234262 705242 234346 705478
rect 234582 705242 262026 705478
rect 262262 705242 262346 705478
rect 262582 705242 290026 705478
rect 290262 705242 290346 705478
rect 290582 705242 318026 705478
rect 318262 705242 318346 705478
rect 318582 705242 346026 705478
rect 346262 705242 346346 705478
rect 346582 705242 374026 705478
rect 374262 705242 374346 705478
rect 374582 705242 402026 705478
rect 402262 705242 402346 705478
rect 402582 705242 430026 705478
rect 430262 705242 430346 705478
rect 430582 705242 458026 705478
rect 458262 705242 458346 705478
rect 458582 705242 486026 705478
rect 486262 705242 486346 705478
rect 486582 705242 514026 705478
rect 514262 705242 514346 705478
rect 514582 705242 542026 705478
rect 542262 705242 542346 705478
rect 542582 705242 570026 705478
rect 570262 705242 570346 705478
rect 570582 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 41526 704838
rect 41762 704602 41846 704838
rect 42082 704602 69526 704838
rect 69762 704602 69846 704838
rect 70082 704602 97526 704838
rect 97762 704602 97846 704838
rect 98082 704602 125526 704838
rect 125762 704602 125846 704838
rect 126082 704602 153526 704838
rect 153762 704602 153846 704838
rect 154082 704602 181526 704838
rect 181762 704602 181846 704838
rect 182082 704602 209526 704838
rect 209762 704602 209846 704838
rect 210082 704602 237526 704838
rect 237762 704602 237846 704838
rect 238082 704602 265526 704838
rect 265762 704602 265846 704838
rect 266082 704602 293526 704838
rect 293762 704602 293846 704838
rect 294082 704602 321526 704838
rect 321762 704602 321846 704838
rect 322082 704602 349526 704838
rect 349762 704602 349846 704838
rect 350082 704602 377526 704838
rect 377762 704602 377846 704838
rect 378082 704602 405526 704838
rect 405762 704602 405846 704838
rect 406082 704602 433526 704838
rect 433762 704602 433846 704838
rect 434082 704602 461526 704838
rect 461762 704602 461846 704838
rect 462082 704602 489526 704838
rect 489762 704602 489846 704838
rect 490082 704602 517526 704838
rect 517762 704602 517846 704838
rect 518082 704602 545526 704838
rect 545762 704602 545846 704838
rect 546082 704602 573526 704838
rect 573762 704602 573846 704838
rect 574082 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 41526 704518
rect 41762 704282 41846 704518
rect 42082 704282 69526 704518
rect 69762 704282 69846 704518
rect 70082 704282 97526 704518
rect 97762 704282 97846 704518
rect 98082 704282 125526 704518
rect 125762 704282 125846 704518
rect 126082 704282 153526 704518
rect 153762 704282 153846 704518
rect 154082 704282 181526 704518
rect 181762 704282 181846 704518
rect 182082 704282 209526 704518
rect 209762 704282 209846 704518
rect 210082 704282 237526 704518
rect 237762 704282 237846 704518
rect 238082 704282 265526 704518
rect 265762 704282 265846 704518
rect 266082 704282 293526 704518
rect 293762 704282 293846 704518
rect 294082 704282 321526 704518
rect 321762 704282 321846 704518
rect 322082 704282 349526 704518
rect 349762 704282 349846 704518
rect 350082 704282 377526 704518
rect 377762 704282 377846 704518
rect 378082 704282 405526 704518
rect 405762 704282 405846 704518
rect 406082 704282 433526 704518
rect 433762 704282 433846 704518
rect 434082 704282 461526 704518
rect 461762 704282 461846 704518
rect 462082 704282 489526 704518
rect 489762 704282 489846 704518
rect 490082 704282 517526 704518
rect 517762 704282 517846 704518
rect 518082 704282 545526 704518
rect 545762 704282 545846 704518
rect 546082 704282 573526 704518
rect 573762 704282 573846 704518
rect 574082 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 701829 592650 701861
rect -8726 701593 -1974 701829
rect -1738 701593 -1654 701829
rect -1418 701593 41526 701829
rect 41762 701593 41846 701829
rect 42082 701593 69526 701829
rect 69762 701593 69846 701829
rect 70082 701593 97526 701829
rect 97762 701593 97846 701829
rect 98082 701593 125526 701829
rect 125762 701593 125846 701829
rect 126082 701593 153526 701829
rect 153762 701593 153846 701829
rect 154082 701593 181526 701829
rect 181762 701593 181846 701829
rect 182082 701593 209526 701829
rect 209762 701593 209846 701829
rect 210082 701593 237526 701829
rect 237762 701593 237846 701829
rect 238082 701593 265526 701829
rect 265762 701593 265846 701829
rect 266082 701593 293526 701829
rect 293762 701593 293846 701829
rect 294082 701593 321526 701829
rect 321762 701593 321846 701829
rect 322082 701593 349526 701829
rect 349762 701593 349846 701829
rect 350082 701593 377526 701829
rect 377762 701593 377846 701829
rect 378082 701593 405526 701829
rect 405762 701593 405846 701829
rect 406082 701593 433526 701829
rect 433762 701593 433846 701829
rect 434082 701593 461526 701829
rect 461762 701593 461846 701829
rect 462082 701593 489526 701829
rect 489762 701593 489846 701829
rect 490082 701593 517526 701829
rect 517762 701593 517846 701829
rect 518082 701593 545526 701829
rect 545762 701593 545846 701829
rect 546082 701593 573526 701829
rect 573762 701593 573846 701829
rect 574082 701593 585342 701829
rect 585578 701593 585662 701829
rect 585898 701593 592650 701829
rect -8726 701509 592650 701593
rect -8726 701273 -1974 701509
rect -1738 701273 -1654 701509
rect -1418 701273 41526 701509
rect 41762 701273 41846 701509
rect 42082 701273 69526 701509
rect 69762 701273 69846 701509
rect 70082 701273 97526 701509
rect 97762 701273 97846 701509
rect 98082 701273 125526 701509
rect 125762 701273 125846 701509
rect 126082 701273 153526 701509
rect 153762 701273 153846 701509
rect 154082 701273 181526 701509
rect 181762 701273 181846 701509
rect 182082 701273 209526 701509
rect 209762 701273 209846 701509
rect 210082 701273 237526 701509
rect 237762 701273 237846 701509
rect 238082 701273 265526 701509
rect 265762 701273 265846 701509
rect 266082 701273 293526 701509
rect 293762 701273 293846 701509
rect 294082 701273 321526 701509
rect 321762 701273 321846 701509
rect 322082 701273 349526 701509
rect 349762 701273 349846 701509
rect 350082 701273 377526 701509
rect 377762 701273 377846 701509
rect 378082 701273 405526 701509
rect 405762 701273 405846 701509
rect 406082 701273 433526 701509
rect 433762 701273 433846 701509
rect 434082 701273 461526 701509
rect 461762 701273 461846 701509
rect 462082 701273 489526 701509
rect 489762 701273 489846 701509
rect 490082 701273 517526 701509
rect 517762 701273 517846 701509
rect 518082 701273 545526 701509
rect 545762 701273 545846 701509
rect 546082 701273 573526 701509
rect 573762 701273 573846 701509
rect 574082 701273 585342 701509
rect 585578 701273 585662 701509
rect 585898 701273 592650 701509
rect -8726 701241 592650 701273
rect -8726 698454 592650 698486
rect -8726 698218 -2934 698454
rect -2698 698218 -2614 698454
rect -2378 698218 38026 698454
rect 38262 698218 38346 698454
rect 38582 698218 66026 698454
rect 66262 698218 66346 698454
rect 66582 698218 94026 698454
rect 94262 698218 94346 698454
rect 94582 698218 122026 698454
rect 122262 698218 122346 698454
rect 122582 698218 150026 698454
rect 150262 698218 150346 698454
rect 150582 698218 178026 698454
rect 178262 698218 178346 698454
rect 178582 698218 206026 698454
rect 206262 698218 206346 698454
rect 206582 698218 234026 698454
rect 234262 698218 234346 698454
rect 234582 698218 262026 698454
rect 262262 698218 262346 698454
rect 262582 698218 290026 698454
rect 290262 698218 290346 698454
rect 290582 698218 318026 698454
rect 318262 698218 318346 698454
rect 318582 698218 346026 698454
rect 346262 698218 346346 698454
rect 346582 698218 374026 698454
rect 374262 698218 374346 698454
rect 374582 698218 402026 698454
rect 402262 698218 402346 698454
rect 402582 698218 430026 698454
rect 430262 698218 430346 698454
rect 430582 698218 458026 698454
rect 458262 698218 458346 698454
rect 458582 698218 486026 698454
rect 486262 698218 486346 698454
rect 486582 698218 514026 698454
rect 514262 698218 514346 698454
rect 514582 698218 542026 698454
rect 542262 698218 542346 698454
rect 542582 698218 570026 698454
rect 570262 698218 570346 698454
rect 570582 698218 586302 698454
rect 586538 698218 586622 698454
rect 586858 698218 592650 698454
rect -8726 698134 592650 698218
rect -8726 697898 -2934 698134
rect -2698 697898 -2614 698134
rect -2378 697898 38026 698134
rect 38262 697898 38346 698134
rect 38582 697898 66026 698134
rect 66262 697898 66346 698134
rect 66582 697898 94026 698134
rect 94262 697898 94346 698134
rect 94582 697898 122026 698134
rect 122262 697898 122346 698134
rect 122582 697898 150026 698134
rect 150262 697898 150346 698134
rect 150582 697898 178026 698134
rect 178262 697898 178346 698134
rect 178582 697898 206026 698134
rect 206262 697898 206346 698134
rect 206582 697898 234026 698134
rect 234262 697898 234346 698134
rect 234582 697898 262026 698134
rect 262262 697898 262346 698134
rect 262582 697898 290026 698134
rect 290262 697898 290346 698134
rect 290582 697898 318026 698134
rect 318262 697898 318346 698134
rect 318582 697898 346026 698134
rect 346262 697898 346346 698134
rect 346582 697898 374026 698134
rect 374262 697898 374346 698134
rect 374582 697898 402026 698134
rect 402262 697898 402346 698134
rect 402582 697898 430026 698134
rect 430262 697898 430346 698134
rect 430582 697898 458026 698134
rect 458262 697898 458346 698134
rect 458582 697898 486026 698134
rect 486262 697898 486346 698134
rect 486582 697898 514026 698134
rect 514262 697898 514346 698134
rect 514582 697898 542026 698134
rect 542262 697898 542346 698134
rect 542582 697898 570026 698134
rect 570262 697898 570346 698134
rect 570582 697898 586302 698134
rect 586538 697898 586622 698134
rect 586858 697898 592650 698134
rect -8726 697866 592650 697898
rect -8726 674829 592650 674861
rect -8726 674593 -1974 674829
rect -1738 674593 -1654 674829
rect -1418 674593 19952 674829
rect 20188 674593 25882 674829
rect 26118 674593 31813 674829
rect 32049 674593 47952 674829
rect 48188 674593 53882 674829
rect 54118 674593 59813 674829
rect 60049 674593 75952 674829
rect 76188 674593 81882 674829
rect 82118 674593 87813 674829
rect 88049 674593 103952 674829
rect 104188 674593 109882 674829
rect 110118 674593 115813 674829
rect 116049 674593 131952 674829
rect 132188 674593 137882 674829
rect 138118 674593 143813 674829
rect 144049 674593 159952 674829
rect 160188 674593 165882 674829
rect 166118 674593 171813 674829
rect 172049 674593 187952 674829
rect 188188 674593 193882 674829
rect 194118 674593 199813 674829
rect 200049 674593 215952 674829
rect 216188 674593 221882 674829
rect 222118 674593 227813 674829
rect 228049 674593 243952 674829
rect 244188 674593 249882 674829
rect 250118 674593 255813 674829
rect 256049 674593 271952 674829
rect 272188 674593 277882 674829
rect 278118 674593 283813 674829
rect 284049 674593 299952 674829
rect 300188 674593 305882 674829
rect 306118 674593 311813 674829
rect 312049 674593 327952 674829
rect 328188 674593 333882 674829
rect 334118 674593 339813 674829
rect 340049 674593 355952 674829
rect 356188 674593 361882 674829
rect 362118 674593 367813 674829
rect 368049 674593 383952 674829
rect 384188 674593 389882 674829
rect 390118 674593 395813 674829
rect 396049 674593 411952 674829
rect 412188 674593 417882 674829
rect 418118 674593 423813 674829
rect 424049 674593 439952 674829
rect 440188 674593 445882 674829
rect 446118 674593 451813 674829
rect 452049 674593 467952 674829
rect 468188 674593 473882 674829
rect 474118 674593 479813 674829
rect 480049 674593 495952 674829
rect 496188 674593 501882 674829
rect 502118 674593 507813 674829
rect 508049 674593 523952 674829
rect 524188 674593 529882 674829
rect 530118 674593 535813 674829
rect 536049 674593 551952 674829
rect 552188 674593 557882 674829
rect 558118 674593 563813 674829
rect 564049 674593 573526 674829
rect 573762 674593 573846 674829
rect 574082 674593 585342 674829
rect 585578 674593 585662 674829
rect 585898 674593 592650 674829
rect -8726 674509 592650 674593
rect -8726 674273 -1974 674509
rect -1738 674273 -1654 674509
rect -1418 674273 19952 674509
rect 20188 674273 25882 674509
rect 26118 674273 31813 674509
rect 32049 674273 47952 674509
rect 48188 674273 53882 674509
rect 54118 674273 59813 674509
rect 60049 674273 75952 674509
rect 76188 674273 81882 674509
rect 82118 674273 87813 674509
rect 88049 674273 103952 674509
rect 104188 674273 109882 674509
rect 110118 674273 115813 674509
rect 116049 674273 131952 674509
rect 132188 674273 137882 674509
rect 138118 674273 143813 674509
rect 144049 674273 159952 674509
rect 160188 674273 165882 674509
rect 166118 674273 171813 674509
rect 172049 674273 187952 674509
rect 188188 674273 193882 674509
rect 194118 674273 199813 674509
rect 200049 674273 215952 674509
rect 216188 674273 221882 674509
rect 222118 674273 227813 674509
rect 228049 674273 243952 674509
rect 244188 674273 249882 674509
rect 250118 674273 255813 674509
rect 256049 674273 271952 674509
rect 272188 674273 277882 674509
rect 278118 674273 283813 674509
rect 284049 674273 299952 674509
rect 300188 674273 305882 674509
rect 306118 674273 311813 674509
rect 312049 674273 327952 674509
rect 328188 674273 333882 674509
rect 334118 674273 339813 674509
rect 340049 674273 355952 674509
rect 356188 674273 361882 674509
rect 362118 674273 367813 674509
rect 368049 674273 383952 674509
rect 384188 674273 389882 674509
rect 390118 674273 395813 674509
rect 396049 674273 411952 674509
rect 412188 674273 417882 674509
rect 418118 674273 423813 674509
rect 424049 674273 439952 674509
rect 440188 674273 445882 674509
rect 446118 674273 451813 674509
rect 452049 674273 467952 674509
rect 468188 674273 473882 674509
rect 474118 674273 479813 674509
rect 480049 674273 495952 674509
rect 496188 674273 501882 674509
rect 502118 674273 507813 674509
rect 508049 674273 523952 674509
rect 524188 674273 529882 674509
rect 530118 674273 535813 674509
rect 536049 674273 551952 674509
rect 552188 674273 557882 674509
rect 558118 674273 563813 674509
rect 564049 674273 573526 674509
rect 573762 674273 573846 674509
rect 574082 674273 585342 674509
rect 585578 674273 585662 674509
rect 585898 674273 592650 674509
rect -8726 674241 592650 674273
rect -8726 671454 592650 671486
rect -8726 671218 -2934 671454
rect -2698 671218 -2614 671454
rect -2378 671218 22916 671454
rect 23152 671218 28847 671454
rect 29083 671218 50916 671454
rect 51152 671218 56847 671454
rect 57083 671218 78916 671454
rect 79152 671218 84847 671454
rect 85083 671218 106916 671454
rect 107152 671218 112847 671454
rect 113083 671218 134916 671454
rect 135152 671218 140847 671454
rect 141083 671218 162916 671454
rect 163152 671218 168847 671454
rect 169083 671218 190916 671454
rect 191152 671218 196847 671454
rect 197083 671218 218916 671454
rect 219152 671218 224847 671454
rect 225083 671218 246916 671454
rect 247152 671218 252847 671454
rect 253083 671218 274916 671454
rect 275152 671218 280847 671454
rect 281083 671218 302916 671454
rect 303152 671218 308847 671454
rect 309083 671218 330916 671454
rect 331152 671218 336847 671454
rect 337083 671218 358916 671454
rect 359152 671218 364847 671454
rect 365083 671218 386916 671454
rect 387152 671218 392847 671454
rect 393083 671218 414916 671454
rect 415152 671218 420847 671454
rect 421083 671218 442916 671454
rect 443152 671218 448847 671454
rect 449083 671218 470916 671454
rect 471152 671218 476847 671454
rect 477083 671218 498916 671454
rect 499152 671218 504847 671454
rect 505083 671218 526916 671454
rect 527152 671218 532847 671454
rect 533083 671218 554916 671454
rect 555152 671218 560847 671454
rect 561083 671218 586302 671454
rect 586538 671218 586622 671454
rect 586858 671218 592650 671454
rect -8726 671134 592650 671218
rect -8726 670898 -2934 671134
rect -2698 670898 -2614 671134
rect -2378 670898 22916 671134
rect 23152 670898 28847 671134
rect 29083 670898 50916 671134
rect 51152 670898 56847 671134
rect 57083 670898 78916 671134
rect 79152 670898 84847 671134
rect 85083 670898 106916 671134
rect 107152 670898 112847 671134
rect 113083 670898 134916 671134
rect 135152 670898 140847 671134
rect 141083 670898 162916 671134
rect 163152 670898 168847 671134
rect 169083 670898 190916 671134
rect 191152 670898 196847 671134
rect 197083 670898 218916 671134
rect 219152 670898 224847 671134
rect 225083 670898 246916 671134
rect 247152 670898 252847 671134
rect 253083 670898 274916 671134
rect 275152 670898 280847 671134
rect 281083 670898 302916 671134
rect 303152 670898 308847 671134
rect 309083 670898 330916 671134
rect 331152 670898 336847 671134
rect 337083 670898 358916 671134
rect 359152 670898 364847 671134
rect 365083 670898 386916 671134
rect 387152 670898 392847 671134
rect 393083 670898 414916 671134
rect 415152 670898 420847 671134
rect 421083 670898 442916 671134
rect 443152 670898 448847 671134
rect 449083 670898 470916 671134
rect 471152 670898 476847 671134
rect 477083 670898 498916 671134
rect 499152 670898 504847 671134
rect 505083 670898 526916 671134
rect 527152 670898 532847 671134
rect 533083 670898 554916 671134
rect 555152 670898 560847 671134
rect 561083 670898 586302 671134
rect 586538 670898 586622 671134
rect 586858 670898 592650 671134
rect -8726 670866 592650 670898
rect -8726 647829 592650 647861
rect -8726 647593 -1974 647829
rect -1738 647593 -1654 647829
rect -1418 647593 19951 647829
rect 20187 647593 25882 647829
rect 26118 647593 31812 647829
rect 32048 647593 47951 647829
rect 48187 647593 53882 647829
rect 54118 647593 59812 647829
rect 60048 647593 75951 647829
rect 76187 647593 81882 647829
rect 82118 647593 87812 647829
rect 88048 647593 103951 647829
rect 104187 647593 109882 647829
rect 110118 647593 115812 647829
rect 116048 647593 131951 647829
rect 132187 647593 137882 647829
rect 138118 647593 143812 647829
rect 144048 647593 159951 647829
rect 160187 647593 165882 647829
rect 166118 647593 171812 647829
rect 172048 647593 187951 647829
rect 188187 647593 193882 647829
rect 194118 647593 199812 647829
rect 200048 647593 215951 647829
rect 216187 647593 221882 647829
rect 222118 647593 227812 647829
rect 228048 647593 243951 647829
rect 244187 647593 249882 647829
rect 250118 647593 255812 647829
rect 256048 647593 271951 647829
rect 272187 647593 277882 647829
rect 278118 647593 283812 647829
rect 284048 647593 299951 647829
rect 300187 647593 305882 647829
rect 306118 647593 311812 647829
rect 312048 647593 327951 647829
rect 328187 647593 333882 647829
rect 334118 647593 339812 647829
rect 340048 647593 355951 647829
rect 356187 647593 361882 647829
rect 362118 647593 367812 647829
rect 368048 647593 383951 647829
rect 384187 647593 389882 647829
rect 390118 647593 395812 647829
rect 396048 647593 411951 647829
rect 412187 647593 417882 647829
rect 418118 647593 423812 647829
rect 424048 647593 439951 647829
rect 440187 647593 445882 647829
rect 446118 647593 451812 647829
rect 452048 647593 467951 647829
rect 468187 647593 473882 647829
rect 474118 647593 479812 647829
rect 480048 647593 495951 647829
rect 496187 647593 501882 647829
rect 502118 647593 507812 647829
rect 508048 647593 523951 647829
rect 524187 647593 529882 647829
rect 530118 647593 535812 647829
rect 536048 647593 551951 647829
rect 552187 647593 557882 647829
rect 558118 647593 563812 647829
rect 564048 647593 573526 647829
rect 573762 647593 573846 647829
rect 574082 647593 585342 647829
rect 585578 647593 585662 647829
rect 585898 647593 592650 647829
rect -8726 647509 592650 647593
rect -8726 647273 -1974 647509
rect -1738 647273 -1654 647509
rect -1418 647273 19951 647509
rect 20187 647273 25882 647509
rect 26118 647273 31812 647509
rect 32048 647273 47951 647509
rect 48187 647273 53882 647509
rect 54118 647273 59812 647509
rect 60048 647273 75951 647509
rect 76187 647273 81882 647509
rect 82118 647273 87812 647509
rect 88048 647273 103951 647509
rect 104187 647273 109882 647509
rect 110118 647273 115812 647509
rect 116048 647273 131951 647509
rect 132187 647273 137882 647509
rect 138118 647273 143812 647509
rect 144048 647273 159951 647509
rect 160187 647273 165882 647509
rect 166118 647273 171812 647509
rect 172048 647273 187951 647509
rect 188187 647273 193882 647509
rect 194118 647273 199812 647509
rect 200048 647273 215951 647509
rect 216187 647273 221882 647509
rect 222118 647273 227812 647509
rect 228048 647273 243951 647509
rect 244187 647273 249882 647509
rect 250118 647273 255812 647509
rect 256048 647273 271951 647509
rect 272187 647273 277882 647509
rect 278118 647273 283812 647509
rect 284048 647273 299951 647509
rect 300187 647273 305882 647509
rect 306118 647273 311812 647509
rect 312048 647273 327951 647509
rect 328187 647273 333882 647509
rect 334118 647273 339812 647509
rect 340048 647273 355951 647509
rect 356187 647273 361882 647509
rect 362118 647273 367812 647509
rect 368048 647273 383951 647509
rect 384187 647273 389882 647509
rect 390118 647273 395812 647509
rect 396048 647273 411951 647509
rect 412187 647273 417882 647509
rect 418118 647273 423812 647509
rect 424048 647273 439951 647509
rect 440187 647273 445882 647509
rect 446118 647273 451812 647509
rect 452048 647273 467951 647509
rect 468187 647273 473882 647509
rect 474118 647273 479812 647509
rect 480048 647273 495951 647509
rect 496187 647273 501882 647509
rect 502118 647273 507812 647509
rect 508048 647273 523951 647509
rect 524187 647273 529882 647509
rect 530118 647273 535812 647509
rect 536048 647273 551951 647509
rect 552187 647273 557882 647509
rect 558118 647273 563812 647509
rect 564048 647273 573526 647509
rect 573762 647273 573846 647509
rect 574082 647273 585342 647509
rect 585578 647273 585662 647509
rect 585898 647273 592650 647509
rect -8726 647241 592650 647273
rect -8726 644454 592650 644486
rect -8726 644218 -2934 644454
rect -2698 644218 -2614 644454
rect -2378 644218 22917 644454
rect 23153 644218 28848 644454
rect 29084 644218 50917 644454
rect 51153 644218 56848 644454
rect 57084 644218 78917 644454
rect 79153 644218 84848 644454
rect 85084 644218 106917 644454
rect 107153 644218 112848 644454
rect 113084 644218 134917 644454
rect 135153 644218 140848 644454
rect 141084 644218 162917 644454
rect 163153 644218 168848 644454
rect 169084 644218 190917 644454
rect 191153 644218 196848 644454
rect 197084 644218 218917 644454
rect 219153 644218 224848 644454
rect 225084 644218 246917 644454
rect 247153 644218 252848 644454
rect 253084 644218 274917 644454
rect 275153 644218 280848 644454
rect 281084 644218 302917 644454
rect 303153 644218 308848 644454
rect 309084 644218 330917 644454
rect 331153 644218 336848 644454
rect 337084 644218 358917 644454
rect 359153 644218 364848 644454
rect 365084 644218 386917 644454
rect 387153 644218 392848 644454
rect 393084 644218 414917 644454
rect 415153 644218 420848 644454
rect 421084 644218 442917 644454
rect 443153 644218 448848 644454
rect 449084 644218 470917 644454
rect 471153 644218 476848 644454
rect 477084 644218 498917 644454
rect 499153 644218 504848 644454
rect 505084 644218 526917 644454
rect 527153 644218 532848 644454
rect 533084 644218 554917 644454
rect 555153 644218 560848 644454
rect 561084 644218 586302 644454
rect 586538 644218 586622 644454
rect 586858 644218 592650 644454
rect -8726 644134 592650 644218
rect -8726 643898 -2934 644134
rect -2698 643898 -2614 644134
rect -2378 643898 22917 644134
rect 23153 643898 28848 644134
rect 29084 643898 50917 644134
rect 51153 643898 56848 644134
rect 57084 643898 78917 644134
rect 79153 643898 84848 644134
rect 85084 643898 106917 644134
rect 107153 643898 112848 644134
rect 113084 643898 134917 644134
rect 135153 643898 140848 644134
rect 141084 643898 162917 644134
rect 163153 643898 168848 644134
rect 169084 643898 190917 644134
rect 191153 643898 196848 644134
rect 197084 643898 218917 644134
rect 219153 643898 224848 644134
rect 225084 643898 246917 644134
rect 247153 643898 252848 644134
rect 253084 643898 274917 644134
rect 275153 643898 280848 644134
rect 281084 643898 302917 644134
rect 303153 643898 308848 644134
rect 309084 643898 330917 644134
rect 331153 643898 336848 644134
rect 337084 643898 358917 644134
rect 359153 643898 364848 644134
rect 365084 643898 386917 644134
rect 387153 643898 392848 644134
rect 393084 643898 414917 644134
rect 415153 643898 420848 644134
rect 421084 643898 442917 644134
rect 443153 643898 448848 644134
rect 449084 643898 470917 644134
rect 471153 643898 476848 644134
rect 477084 643898 498917 644134
rect 499153 643898 504848 644134
rect 505084 643898 526917 644134
rect 527153 643898 532848 644134
rect 533084 643898 554917 644134
rect 555153 643898 560848 644134
rect 561084 643898 586302 644134
rect 586538 643898 586622 644134
rect 586858 643898 592650 644134
rect -8726 643866 592650 643898
rect -8726 620829 592650 620861
rect -8726 620593 -1974 620829
rect -1738 620593 -1654 620829
rect -1418 620593 19952 620829
rect 20188 620593 25882 620829
rect 26118 620593 31813 620829
rect 32049 620593 47952 620829
rect 48188 620593 53882 620829
rect 54118 620593 59813 620829
rect 60049 620593 75952 620829
rect 76188 620593 81882 620829
rect 82118 620593 87813 620829
rect 88049 620593 103952 620829
rect 104188 620593 109882 620829
rect 110118 620593 115813 620829
rect 116049 620593 131952 620829
rect 132188 620593 137882 620829
rect 138118 620593 143813 620829
rect 144049 620593 159952 620829
rect 160188 620593 165882 620829
rect 166118 620593 171813 620829
rect 172049 620593 187952 620829
rect 188188 620593 193882 620829
rect 194118 620593 199813 620829
rect 200049 620593 215952 620829
rect 216188 620593 221882 620829
rect 222118 620593 227813 620829
rect 228049 620593 243952 620829
rect 244188 620593 249882 620829
rect 250118 620593 255813 620829
rect 256049 620593 271952 620829
rect 272188 620593 277882 620829
rect 278118 620593 283813 620829
rect 284049 620593 299952 620829
rect 300188 620593 305882 620829
rect 306118 620593 311813 620829
rect 312049 620593 327952 620829
rect 328188 620593 333882 620829
rect 334118 620593 339813 620829
rect 340049 620593 355952 620829
rect 356188 620593 361882 620829
rect 362118 620593 367813 620829
rect 368049 620593 383952 620829
rect 384188 620593 389882 620829
rect 390118 620593 395813 620829
rect 396049 620593 411952 620829
rect 412188 620593 417882 620829
rect 418118 620593 423813 620829
rect 424049 620593 439952 620829
rect 440188 620593 445882 620829
rect 446118 620593 451813 620829
rect 452049 620593 467952 620829
rect 468188 620593 473882 620829
rect 474118 620593 479813 620829
rect 480049 620593 495952 620829
rect 496188 620593 501882 620829
rect 502118 620593 507813 620829
rect 508049 620593 523952 620829
rect 524188 620593 529882 620829
rect 530118 620593 535813 620829
rect 536049 620593 551952 620829
rect 552188 620593 557882 620829
rect 558118 620593 563813 620829
rect 564049 620593 573526 620829
rect 573762 620593 573846 620829
rect 574082 620593 585342 620829
rect 585578 620593 585662 620829
rect 585898 620593 592650 620829
rect -8726 620509 592650 620593
rect -8726 620273 -1974 620509
rect -1738 620273 -1654 620509
rect -1418 620273 19952 620509
rect 20188 620273 25882 620509
rect 26118 620273 31813 620509
rect 32049 620273 47952 620509
rect 48188 620273 53882 620509
rect 54118 620273 59813 620509
rect 60049 620273 75952 620509
rect 76188 620273 81882 620509
rect 82118 620273 87813 620509
rect 88049 620273 103952 620509
rect 104188 620273 109882 620509
rect 110118 620273 115813 620509
rect 116049 620273 131952 620509
rect 132188 620273 137882 620509
rect 138118 620273 143813 620509
rect 144049 620273 159952 620509
rect 160188 620273 165882 620509
rect 166118 620273 171813 620509
rect 172049 620273 187952 620509
rect 188188 620273 193882 620509
rect 194118 620273 199813 620509
rect 200049 620273 215952 620509
rect 216188 620273 221882 620509
rect 222118 620273 227813 620509
rect 228049 620273 243952 620509
rect 244188 620273 249882 620509
rect 250118 620273 255813 620509
rect 256049 620273 271952 620509
rect 272188 620273 277882 620509
rect 278118 620273 283813 620509
rect 284049 620273 299952 620509
rect 300188 620273 305882 620509
rect 306118 620273 311813 620509
rect 312049 620273 327952 620509
rect 328188 620273 333882 620509
rect 334118 620273 339813 620509
rect 340049 620273 355952 620509
rect 356188 620273 361882 620509
rect 362118 620273 367813 620509
rect 368049 620273 383952 620509
rect 384188 620273 389882 620509
rect 390118 620273 395813 620509
rect 396049 620273 411952 620509
rect 412188 620273 417882 620509
rect 418118 620273 423813 620509
rect 424049 620273 439952 620509
rect 440188 620273 445882 620509
rect 446118 620273 451813 620509
rect 452049 620273 467952 620509
rect 468188 620273 473882 620509
rect 474118 620273 479813 620509
rect 480049 620273 495952 620509
rect 496188 620273 501882 620509
rect 502118 620273 507813 620509
rect 508049 620273 523952 620509
rect 524188 620273 529882 620509
rect 530118 620273 535813 620509
rect 536049 620273 551952 620509
rect 552188 620273 557882 620509
rect 558118 620273 563813 620509
rect 564049 620273 573526 620509
rect 573762 620273 573846 620509
rect 574082 620273 585342 620509
rect 585578 620273 585662 620509
rect 585898 620273 592650 620509
rect -8726 620241 592650 620273
rect -8726 617454 592650 617486
rect -8726 617218 -2934 617454
rect -2698 617218 -2614 617454
rect -2378 617218 22916 617454
rect 23152 617218 28847 617454
rect 29083 617218 50916 617454
rect 51152 617218 56847 617454
rect 57083 617218 78916 617454
rect 79152 617218 84847 617454
rect 85083 617218 106916 617454
rect 107152 617218 112847 617454
rect 113083 617218 134916 617454
rect 135152 617218 140847 617454
rect 141083 617218 162916 617454
rect 163152 617218 168847 617454
rect 169083 617218 190916 617454
rect 191152 617218 196847 617454
rect 197083 617218 218916 617454
rect 219152 617218 224847 617454
rect 225083 617218 246916 617454
rect 247152 617218 252847 617454
rect 253083 617218 274916 617454
rect 275152 617218 280847 617454
rect 281083 617218 302916 617454
rect 303152 617218 308847 617454
rect 309083 617218 330916 617454
rect 331152 617218 336847 617454
rect 337083 617218 358916 617454
rect 359152 617218 364847 617454
rect 365083 617218 386916 617454
rect 387152 617218 392847 617454
rect 393083 617218 414916 617454
rect 415152 617218 420847 617454
rect 421083 617218 442916 617454
rect 443152 617218 448847 617454
rect 449083 617218 470916 617454
rect 471152 617218 476847 617454
rect 477083 617218 498916 617454
rect 499152 617218 504847 617454
rect 505083 617218 526916 617454
rect 527152 617218 532847 617454
rect 533083 617218 554916 617454
rect 555152 617218 560847 617454
rect 561083 617218 586302 617454
rect 586538 617218 586622 617454
rect 586858 617218 592650 617454
rect -8726 617134 592650 617218
rect -8726 616898 -2934 617134
rect -2698 616898 -2614 617134
rect -2378 616898 22916 617134
rect 23152 616898 28847 617134
rect 29083 616898 50916 617134
rect 51152 616898 56847 617134
rect 57083 616898 78916 617134
rect 79152 616898 84847 617134
rect 85083 616898 106916 617134
rect 107152 616898 112847 617134
rect 113083 616898 134916 617134
rect 135152 616898 140847 617134
rect 141083 616898 162916 617134
rect 163152 616898 168847 617134
rect 169083 616898 190916 617134
rect 191152 616898 196847 617134
rect 197083 616898 218916 617134
rect 219152 616898 224847 617134
rect 225083 616898 246916 617134
rect 247152 616898 252847 617134
rect 253083 616898 274916 617134
rect 275152 616898 280847 617134
rect 281083 616898 302916 617134
rect 303152 616898 308847 617134
rect 309083 616898 330916 617134
rect 331152 616898 336847 617134
rect 337083 616898 358916 617134
rect 359152 616898 364847 617134
rect 365083 616898 386916 617134
rect 387152 616898 392847 617134
rect 393083 616898 414916 617134
rect 415152 616898 420847 617134
rect 421083 616898 442916 617134
rect 443152 616898 448847 617134
rect 449083 616898 470916 617134
rect 471152 616898 476847 617134
rect 477083 616898 498916 617134
rect 499152 616898 504847 617134
rect 505083 616898 526916 617134
rect 527152 616898 532847 617134
rect 533083 616898 554916 617134
rect 555152 616898 560847 617134
rect 561083 616898 586302 617134
rect 586538 616898 586622 617134
rect 586858 616898 592650 617134
rect -8726 616866 592650 616898
rect -8726 593829 592650 593861
rect -8726 593593 -1974 593829
rect -1738 593593 -1654 593829
rect -1418 593593 19951 593829
rect 20187 593593 25882 593829
rect 26118 593593 31812 593829
rect 32048 593593 47951 593829
rect 48187 593593 53882 593829
rect 54118 593593 59812 593829
rect 60048 593593 75951 593829
rect 76187 593593 81882 593829
rect 82118 593593 87812 593829
rect 88048 593593 103951 593829
rect 104187 593593 109882 593829
rect 110118 593593 115812 593829
rect 116048 593593 131951 593829
rect 132187 593593 137882 593829
rect 138118 593593 143812 593829
rect 144048 593593 159951 593829
rect 160187 593593 165882 593829
rect 166118 593593 171812 593829
rect 172048 593593 187951 593829
rect 188187 593593 193882 593829
rect 194118 593593 199812 593829
rect 200048 593593 215951 593829
rect 216187 593593 221882 593829
rect 222118 593593 227812 593829
rect 228048 593593 243951 593829
rect 244187 593593 249882 593829
rect 250118 593593 255812 593829
rect 256048 593593 271951 593829
rect 272187 593593 277882 593829
rect 278118 593593 283812 593829
rect 284048 593593 299951 593829
rect 300187 593593 305882 593829
rect 306118 593593 311812 593829
rect 312048 593593 327951 593829
rect 328187 593593 333882 593829
rect 334118 593593 339812 593829
rect 340048 593593 355951 593829
rect 356187 593593 361882 593829
rect 362118 593593 367812 593829
rect 368048 593593 383951 593829
rect 384187 593593 389882 593829
rect 390118 593593 395812 593829
rect 396048 593593 411951 593829
rect 412187 593593 417882 593829
rect 418118 593593 423812 593829
rect 424048 593593 439951 593829
rect 440187 593593 445882 593829
rect 446118 593593 451812 593829
rect 452048 593593 467951 593829
rect 468187 593593 473882 593829
rect 474118 593593 479812 593829
rect 480048 593593 495951 593829
rect 496187 593593 501882 593829
rect 502118 593593 507812 593829
rect 508048 593593 523951 593829
rect 524187 593593 529882 593829
rect 530118 593593 535812 593829
rect 536048 593593 551951 593829
rect 552187 593593 557882 593829
rect 558118 593593 563812 593829
rect 564048 593593 573526 593829
rect 573762 593593 573846 593829
rect 574082 593593 585342 593829
rect 585578 593593 585662 593829
rect 585898 593593 592650 593829
rect -8726 593509 592650 593593
rect -8726 593273 -1974 593509
rect -1738 593273 -1654 593509
rect -1418 593273 19951 593509
rect 20187 593273 25882 593509
rect 26118 593273 31812 593509
rect 32048 593273 47951 593509
rect 48187 593273 53882 593509
rect 54118 593273 59812 593509
rect 60048 593273 75951 593509
rect 76187 593273 81882 593509
rect 82118 593273 87812 593509
rect 88048 593273 103951 593509
rect 104187 593273 109882 593509
rect 110118 593273 115812 593509
rect 116048 593273 131951 593509
rect 132187 593273 137882 593509
rect 138118 593273 143812 593509
rect 144048 593273 159951 593509
rect 160187 593273 165882 593509
rect 166118 593273 171812 593509
rect 172048 593273 187951 593509
rect 188187 593273 193882 593509
rect 194118 593273 199812 593509
rect 200048 593273 215951 593509
rect 216187 593273 221882 593509
rect 222118 593273 227812 593509
rect 228048 593273 243951 593509
rect 244187 593273 249882 593509
rect 250118 593273 255812 593509
rect 256048 593273 271951 593509
rect 272187 593273 277882 593509
rect 278118 593273 283812 593509
rect 284048 593273 299951 593509
rect 300187 593273 305882 593509
rect 306118 593273 311812 593509
rect 312048 593273 327951 593509
rect 328187 593273 333882 593509
rect 334118 593273 339812 593509
rect 340048 593273 355951 593509
rect 356187 593273 361882 593509
rect 362118 593273 367812 593509
rect 368048 593273 383951 593509
rect 384187 593273 389882 593509
rect 390118 593273 395812 593509
rect 396048 593273 411951 593509
rect 412187 593273 417882 593509
rect 418118 593273 423812 593509
rect 424048 593273 439951 593509
rect 440187 593273 445882 593509
rect 446118 593273 451812 593509
rect 452048 593273 467951 593509
rect 468187 593273 473882 593509
rect 474118 593273 479812 593509
rect 480048 593273 495951 593509
rect 496187 593273 501882 593509
rect 502118 593273 507812 593509
rect 508048 593273 523951 593509
rect 524187 593273 529882 593509
rect 530118 593273 535812 593509
rect 536048 593273 551951 593509
rect 552187 593273 557882 593509
rect 558118 593273 563812 593509
rect 564048 593273 573526 593509
rect 573762 593273 573846 593509
rect 574082 593273 585342 593509
rect 585578 593273 585662 593509
rect 585898 593273 592650 593509
rect -8726 593241 592650 593273
rect -8726 590454 592650 590486
rect -8726 590218 -2934 590454
rect -2698 590218 -2614 590454
rect -2378 590218 22917 590454
rect 23153 590218 28848 590454
rect 29084 590218 50917 590454
rect 51153 590218 56848 590454
rect 57084 590218 78917 590454
rect 79153 590218 84848 590454
rect 85084 590218 106917 590454
rect 107153 590218 112848 590454
rect 113084 590218 134917 590454
rect 135153 590218 140848 590454
rect 141084 590218 162917 590454
rect 163153 590218 168848 590454
rect 169084 590218 190917 590454
rect 191153 590218 196848 590454
rect 197084 590218 218917 590454
rect 219153 590218 224848 590454
rect 225084 590218 246917 590454
rect 247153 590218 252848 590454
rect 253084 590218 274917 590454
rect 275153 590218 280848 590454
rect 281084 590218 302917 590454
rect 303153 590218 308848 590454
rect 309084 590218 330917 590454
rect 331153 590218 336848 590454
rect 337084 590218 358917 590454
rect 359153 590218 364848 590454
rect 365084 590218 386917 590454
rect 387153 590218 392848 590454
rect 393084 590218 414917 590454
rect 415153 590218 420848 590454
rect 421084 590218 442917 590454
rect 443153 590218 448848 590454
rect 449084 590218 470917 590454
rect 471153 590218 476848 590454
rect 477084 590218 498917 590454
rect 499153 590218 504848 590454
rect 505084 590218 526917 590454
rect 527153 590218 532848 590454
rect 533084 590218 554917 590454
rect 555153 590218 560848 590454
rect 561084 590218 586302 590454
rect 586538 590218 586622 590454
rect 586858 590218 592650 590454
rect -8726 590134 592650 590218
rect -8726 589898 -2934 590134
rect -2698 589898 -2614 590134
rect -2378 589898 22917 590134
rect 23153 589898 28848 590134
rect 29084 589898 50917 590134
rect 51153 589898 56848 590134
rect 57084 589898 78917 590134
rect 79153 589898 84848 590134
rect 85084 589898 106917 590134
rect 107153 589898 112848 590134
rect 113084 589898 134917 590134
rect 135153 589898 140848 590134
rect 141084 589898 162917 590134
rect 163153 589898 168848 590134
rect 169084 589898 190917 590134
rect 191153 589898 196848 590134
rect 197084 589898 218917 590134
rect 219153 589898 224848 590134
rect 225084 589898 246917 590134
rect 247153 589898 252848 590134
rect 253084 589898 274917 590134
rect 275153 589898 280848 590134
rect 281084 589898 302917 590134
rect 303153 589898 308848 590134
rect 309084 589898 330917 590134
rect 331153 589898 336848 590134
rect 337084 589898 358917 590134
rect 359153 589898 364848 590134
rect 365084 589898 386917 590134
rect 387153 589898 392848 590134
rect 393084 589898 414917 590134
rect 415153 589898 420848 590134
rect 421084 589898 442917 590134
rect 443153 589898 448848 590134
rect 449084 589898 470917 590134
rect 471153 589898 476848 590134
rect 477084 589898 498917 590134
rect 499153 589898 504848 590134
rect 505084 589898 526917 590134
rect 527153 589898 532848 590134
rect 533084 589898 554917 590134
rect 555153 589898 560848 590134
rect 561084 589898 586302 590134
rect 586538 589898 586622 590134
rect 586858 589898 592650 590134
rect -8726 589866 592650 589898
rect -8726 566829 592650 566861
rect -8726 566593 -1974 566829
rect -1738 566593 -1654 566829
rect -1418 566593 19952 566829
rect 20188 566593 25882 566829
rect 26118 566593 31813 566829
rect 32049 566593 47952 566829
rect 48188 566593 53882 566829
rect 54118 566593 59813 566829
rect 60049 566593 75952 566829
rect 76188 566593 81882 566829
rect 82118 566593 87813 566829
rect 88049 566593 103952 566829
rect 104188 566593 109882 566829
rect 110118 566593 115813 566829
rect 116049 566593 131952 566829
rect 132188 566593 137882 566829
rect 138118 566593 143813 566829
rect 144049 566593 159952 566829
rect 160188 566593 165882 566829
rect 166118 566593 171813 566829
rect 172049 566593 187952 566829
rect 188188 566593 193882 566829
rect 194118 566593 199813 566829
rect 200049 566593 215952 566829
rect 216188 566593 221882 566829
rect 222118 566593 227813 566829
rect 228049 566593 243952 566829
rect 244188 566593 249882 566829
rect 250118 566593 255813 566829
rect 256049 566593 271952 566829
rect 272188 566593 277882 566829
rect 278118 566593 283813 566829
rect 284049 566593 299952 566829
rect 300188 566593 305882 566829
rect 306118 566593 311813 566829
rect 312049 566593 327952 566829
rect 328188 566593 333882 566829
rect 334118 566593 339813 566829
rect 340049 566593 355952 566829
rect 356188 566593 361882 566829
rect 362118 566593 367813 566829
rect 368049 566593 383952 566829
rect 384188 566593 389882 566829
rect 390118 566593 395813 566829
rect 396049 566593 411952 566829
rect 412188 566593 417882 566829
rect 418118 566593 423813 566829
rect 424049 566593 439952 566829
rect 440188 566593 445882 566829
rect 446118 566593 451813 566829
rect 452049 566593 467952 566829
rect 468188 566593 473882 566829
rect 474118 566593 479813 566829
rect 480049 566593 495952 566829
rect 496188 566593 501882 566829
rect 502118 566593 507813 566829
rect 508049 566593 523952 566829
rect 524188 566593 529882 566829
rect 530118 566593 535813 566829
rect 536049 566593 551952 566829
rect 552188 566593 557882 566829
rect 558118 566593 563813 566829
rect 564049 566593 573526 566829
rect 573762 566593 573846 566829
rect 574082 566593 585342 566829
rect 585578 566593 585662 566829
rect 585898 566593 592650 566829
rect -8726 566509 592650 566593
rect -8726 566273 -1974 566509
rect -1738 566273 -1654 566509
rect -1418 566273 19952 566509
rect 20188 566273 25882 566509
rect 26118 566273 31813 566509
rect 32049 566273 47952 566509
rect 48188 566273 53882 566509
rect 54118 566273 59813 566509
rect 60049 566273 75952 566509
rect 76188 566273 81882 566509
rect 82118 566273 87813 566509
rect 88049 566273 103952 566509
rect 104188 566273 109882 566509
rect 110118 566273 115813 566509
rect 116049 566273 131952 566509
rect 132188 566273 137882 566509
rect 138118 566273 143813 566509
rect 144049 566273 159952 566509
rect 160188 566273 165882 566509
rect 166118 566273 171813 566509
rect 172049 566273 187952 566509
rect 188188 566273 193882 566509
rect 194118 566273 199813 566509
rect 200049 566273 215952 566509
rect 216188 566273 221882 566509
rect 222118 566273 227813 566509
rect 228049 566273 243952 566509
rect 244188 566273 249882 566509
rect 250118 566273 255813 566509
rect 256049 566273 271952 566509
rect 272188 566273 277882 566509
rect 278118 566273 283813 566509
rect 284049 566273 299952 566509
rect 300188 566273 305882 566509
rect 306118 566273 311813 566509
rect 312049 566273 327952 566509
rect 328188 566273 333882 566509
rect 334118 566273 339813 566509
rect 340049 566273 355952 566509
rect 356188 566273 361882 566509
rect 362118 566273 367813 566509
rect 368049 566273 383952 566509
rect 384188 566273 389882 566509
rect 390118 566273 395813 566509
rect 396049 566273 411952 566509
rect 412188 566273 417882 566509
rect 418118 566273 423813 566509
rect 424049 566273 439952 566509
rect 440188 566273 445882 566509
rect 446118 566273 451813 566509
rect 452049 566273 467952 566509
rect 468188 566273 473882 566509
rect 474118 566273 479813 566509
rect 480049 566273 495952 566509
rect 496188 566273 501882 566509
rect 502118 566273 507813 566509
rect 508049 566273 523952 566509
rect 524188 566273 529882 566509
rect 530118 566273 535813 566509
rect 536049 566273 551952 566509
rect 552188 566273 557882 566509
rect 558118 566273 563813 566509
rect 564049 566273 573526 566509
rect 573762 566273 573846 566509
rect 574082 566273 585342 566509
rect 585578 566273 585662 566509
rect 585898 566273 592650 566509
rect -8726 566241 592650 566273
rect -8726 563454 592650 563486
rect -8726 563218 -2934 563454
rect -2698 563218 -2614 563454
rect -2378 563218 22916 563454
rect 23152 563218 28847 563454
rect 29083 563218 50916 563454
rect 51152 563218 56847 563454
rect 57083 563218 78916 563454
rect 79152 563218 84847 563454
rect 85083 563218 106916 563454
rect 107152 563218 112847 563454
rect 113083 563218 134916 563454
rect 135152 563218 140847 563454
rect 141083 563218 162916 563454
rect 163152 563218 168847 563454
rect 169083 563218 190916 563454
rect 191152 563218 196847 563454
rect 197083 563218 218916 563454
rect 219152 563218 224847 563454
rect 225083 563218 246916 563454
rect 247152 563218 252847 563454
rect 253083 563218 274916 563454
rect 275152 563218 280847 563454
rect 281083 563218 302916 563454
rect 303152 563218 308847 563454
rect 309083 563218 330916 563454
rect 331152 563218 336847 563454
rect 337083 563218 358916 563454
rect 359152 563218 364847 563454
rect 365083 563218 386916 563454
rect 387152 563218 392847 563454
rect 393083 563218 414916 563454
rect 415152 563218 420847 563454
rect 421083 563218 442916 563454
rect 443152 563218 448847 563454
rect 449083 563218 470916 563454
rect 471152 563218 476847 563454
rect 477083 563218 498916 563454
rect 499152 563218 504847 563454
rect 505083 563218 526916 563454
rect 527152 563218 532847 563454
rect 533083 563218 554916 563454
rect 555152 563218 560847 563454
rect 561083 563218 586302 563454
rect 586538 563218 586622 563454
rect 586858 563218 592650 563454
rect -8726 563134 592650 563218
rect -8726 562898 -2934 563134
rect -2698 562898 -2614 563134
rect -2378 562898 22916 563134
rect 23152 562898 28847 563134
rect 29083 562898 50916 563134
rect 51152 562898 56847 563134
rect 57083 562898 78916 563134
rect 79152 562898 84847 563134
rect 85083 562898 106916 563134
rect 107152 562898 112847 563134
rect 113083 562898 134916 563134
rect 135152 562898 140847 563134
rect 141083 562898 162916 563134
rect 163152 562898 168847 563134
rect 169083 562898 190916 563134
rect 191152 562898 196847 563134
rect 197083 562898 218916 563134
rect 219152 562898 224847 563134
rect 225083 562898 246916 563134
rect 247152 562898 252847 563134
rect 253083 562898 274916 563134
rect 275152 562898 280847 563134
rect 281083 562898 302916 563134
rect 303152 562898 308847 563134
rect 309083 562898 330916 563134
rect 331152 562898 336847 563134
rect 337083 562898 358916 563134
rect 359152 562898 364847 563134
rect 365083 562898 386916 563134
rect 387152 562898 392847 563134
rect 393083 562898 414916 563134
rect 415152 562898 420847 563134
rect 421083 562898 442916 563134
rect 443152 562898 448847 563134
rect 449083 562898 470916 563134
rect 471152 562898 476847 563134
rect 477083 562898 498916 563134
rect 499152 562898 504847 563134
rect 505083 562898 526916 563134
rect 527152 562898 532847 563134
rect 533083 562898 554916 563134
rect 555152 562898 560847 563134
rect 561083 562898 586302 563134
rect 586538 562898 586622 563134
rect 586858 562898 592650 563134
rect -8726 562866 592650 562898
rect -8726 539829 592650 539861
rect -8726 539593 -1974 539829
rect -1738 539593 -1654 539829
rect -1418 539593 19951 539829
rect 20187 539593 25882 539829
rect 26118 539593 31812 539829
rect 32048 539593 47951 539829
rect 48187 539593 53882 539829
rect 54118 539593 59812 539829
rect 60048 539593 75951 539829
rect 76187 539593 81882 539829
rect 82118 539593 87812 539829
rect 88048 539593 103951 539829
rect 104187 539593 109882 539829
rect 110118 539593 115812 539829
rect 116048 539593 131951 539829
rect 132187 539593 137882 539829
rect 138118 539593 143812 539829
rect 144048 539593 159951 539829
rect 160187 539593 165882 539829
rect 166118 539593 171812 539829
rect 172048 539593 187951 539829
rect 188187 539593 193882 539829
rect 194118 539593 199812 539829
rect 200048 539593 215951 539829
rect 216187 539593 221882 539829
rect 222118 539593 227812 539829
rect 228048 539593 243951 539829
rect 244187 539593 249882 539829
rect 250118 539593 255812 539829
rect 256048 539593 271951 539829
rect 272187 539593 277882 539829
rect 278118 539593 283812 539829
rect 284048 539593 299951 539829
rect 300187 539593 305882 539829
rect 306118 539593 311812 539829
rect 312048 539593 327951 539829
rect 328187 539593 333882 539829
rect 334118 539593 339812 539829
rect 340048 539593 355951 539829
rect 356187 539593 361882 539829
rect 362118 539593 367812 539829
rect 368048 539593 383951 539829
rect 384187 539593 389882 539829
rect 390118 539593 395812 539829
rect 396048 539593 411951 539829
rect 412187 539593 417882 539829
rect 418118 539593 423812 539829
rect 424048 539593 439951 539829
rect 440187 539593 445882 539829
rect 446118 539593 451812 539829
rect 452048 539593 467951 539829
rect 468187 539593 473882 539829
rect 474118 539593 479812 539829
rect 480048 539593 495951 539829
rect 496187 539593 501882 539829
rect 502118 539593 507812 539829
rect 508048 539593 523951 539829
rect 524187 539593 529882 539829
rect 530118 539593 535812 539829
rect 536048 539593 551951 539829
rect 552187 539593 557882 539829
rect 558118 539593 563812 539829
rect 564048 539593 573526 539829
rect 573762 539593 573846 539829
rect 574082 539593 585342 539829
rect 585578 539593 585662 539829
rect 585898 539593 592650 539829
rect -8726 539509 592650 539593
rect -8726 539273 -1974 539509
rect -1738 539273 -1654 539509
rect -1418 539273 19951 539509
rect 20187 539273 25882 539509
rect 26118 539273 31812 539509
rect 32048 539273 47951 539509
rect 48187 539273 53882 539509
rect 54118 539273 59812 539509
rect 60048 539273 75951 539509
rect 76187 539273 81882 539509
rect 82118 539273 87812 539509
rect 88048 539273 103951 539509
rect 104187 539273 109882 539509
rect 110118 539273 115812 539509
rect 116048 539273 131951 539509
rect 132187 539273 137882 539509
rect 138118 539273 143812 539509
rect 144048 539273 159951 539509
rect 160187 539273 165882 539509
rect 166118 539273 171812 539509
rect 172048 539273 187951 539509
rect 188187 539273 193882 539509
rect 194118 539273 199812 539509
rect 200048 539273 215951 539509
rect 216187 539273 221882 539509
rect 222118 539273 227812 539509
rect 228048 539273 243951 539509
rect 244187 539273 249882 539509
rect 250118 539273 255812 539509
rect 256048 539273 271951 539509
rect 272187 539273 277882 539509
rect 278118 539273 283812 539509
rect 284048 539273 299951 539509
rect 300187 539273 305882 539509
rect 306118 539273 311812 539509
rect 312048 539273 327951 539509
rect 328187 539273 333882 539509
rect 334118 539273 339812 539509
rect 340048 539273 355951 539509
rect 356187 539273 361882 539509
rect 362118 539273 367812 539509
rect 368048 539273 383951 539509
rect 384187 539273 389882 539509
rect 390118 539273 395812 539509
rect 396048 539273 411951 539509
rect 412187 539273 417882 539509
rect 418118 539273 423812 539509
rect 424048 539273 439951 539509
rect 440187 539273 445882 539509
rect 446118 539273 451812 539509
rect 452048 539273 467951 539509
rect 468187 539273 473882 539509
rect 474118 539273 479812 539509
rect 480048 539273 495951 539509
rect 496187 539273 501882 539509
rect 502118 539273 507812 539509
rect 508048 539273 523951 539509
rect 524187 539273 529882 539509
rect 530118 539273 535812 539509
rect 536048 539273 551951 539509
rect 552187 539273 557882 539509
rect 558118 539273 563812 539509
rect 564048 539273 573526 539509
rect 573762 539273 573846 539509
rect 574082 539273 585342 539509
rect 585578 539273 585662 539509
rect 585898 539273 592650 539509
rect -8726 539241 592650 539273
rect -8726 536454 592650 536486
rect -8726 536218 -2934 536454
rect -2698 536218 -2614 536454
rect -2378 536218 22917 536454
rect 23153 536218 28848 536454
rect 29084 536218 50917 536454
rect 51153 536218 56848 536454
rect 57084 536218 78917 536454
rect 79153 536218 84848 536454
rect 85084 536218 106917 536454
rect 107153 536218 112848 536454
rect 113084 536218 134917 536454
rect 135153 536218 140848 536454
rect 141084 536218 162917 536454
rect 163153 536218 168848 536454
rect 169084 536218 190917 536454
rect 191153 536218 196848 536454
rect 197084 536218 218917 536454
rect 219153 536218 224848 536454
rect 225084 536218 246917 536454
rect 247153 536218 252848 536454
rect 253084 536218 274917 536454
rect 275153 536218 280848 536454
rect 281084 536218 302917 536454
rect 303153 536218 308848 536454
rect 309084 536218 330917 536454
rect 331153 536218 336848 536454
rect 337084 536218 358917 536454
rect 359153 536218 364848 536454
rect 365084 536218 386917 536454
rect 387153 536218 392848 536454
rect 393084 536218 414917 536454
rect 415153 536218 420848 536454
rect 421084 536218 442917 536454
rect 443153 536218 448848 536454
rect 449084 536218 470917 536454
rect 471153 536218 476848 536454
rect 477084 536218 498917 536454
rect 499153 536218 504848 536454
rect 505084 536218 526917 536454
rect 527153 536218 532848 536454
rect 533084 536218 554917 536454
rect 555153 536218 560848 536454
rect 561084 536218 586302 536454
rect 586538 536218 586622 536454
rect 586858 536218 592650 536454
rect -8726 536134 592650 536218
rect -8726 535898 -2934 536134
rect -2698 535898 -2614 536134
rect -2378 535898 22917 536134
rect 23153 535898 28848 536134
rect 29084 535898 50917 536134
rect 51153 535898 56848 536134
rect 57084 535898 78917 536134
rect 79153 535898 84848 536134
rect 85084 535898 106917 536134
rect 107153 535898 112848 536134
rect 113084 535898 134917 536134
rect 135153 535898 140848 536134
rect 141084 535898 162917 536134
rect 163153 535898 168848 536134
rect 169084 535898 190917 536134
rect 191153 535898 196848 536134
rect 197084 535898 218917 536134
rect 219153 535898 224848 536134
rect 225084 535898 246917 536134
rect 247153 535898 252848 536134
rect 253084 535898 274917 536134
rect 275153 535898 280848 536134
rect 281084 535898 302917 536134
rect 303153 535898 308848 536134
rect 309084 535898 330917 536134
rect 331153 535898 336848 536134
rect 337084 535898 358917 536134
rect 359153 535898 364848 536134
rect 365084 535898 386917 536134
rect 387153 535898 392848 536134
rect 393084 535898 414917 536134
rect 415153 535898 420848 536134
rect 421084 535898 442917 536134
rect 443153 535898 448848 536134
rect 449084 535898 470917 536134
rect 471153 535898 476848 536134
rect 477084 535898 498917 536134
rect 499153 535898 504848 536134
rect 505084 535898 526917 536134
rect 527153 535898 532848 536134
rect 533084 535898 554917 536134
rect 555153 535898 560848 536134
rect 561084 535898 586302 536134
rect 586538 535898 586622 536134
rect 586858 535898 592650 536134
rect -8726 535866 592650 535898
rect -8726 512829 592650 512861
rect -8726 512593 -1974 512829
rect -1738 512593 -1654 512829
rect -1418 512593 19952 512829
rect 20188 512593 25882 512829
rect 26118 512593 31813 512829
rect 32049 512593 47952 512829
rect 48188 512593 53882 512829
rect 54118 512593 59813 512829
rect 60049 512593 75952 512829
rect 76188 512593 81882 512829
rect 82118 512593 87813 512829
rect 88049 512593 103952 512829
rect 104188 512593 109882 512829
rect 110118 512593 115813 512829
rect 116049 512593 131952 512829
rect 132188 512593 137882 512829
rect 138118 512593 143813 512829
rect 144049 512593 159952 512829
rect 160188 512593 165882 512829
rect 166118 512593 171813 512829
rect 172049 512593 187952 512829
rect 188188 512593 193882 512829
rect 194118 512593 199813 512829
rect 200049 512593 215952 512829
rect 216188 512593 221882 512829
rect 222118 512593 227813 512829
rect 228049 512593 243952 512829
rect 244188 512593 249882 512829
rect 250118 512593 255813 512829
rect 256049 512593 271952 512829
rect 272188 512593 277882 512829
rect 278118 512593 283813 512829
rect 284049 512593 299952 512829
rect 300188 512593 305882 512829
rect 306118 512593 311813 512829
rect 312049 512593 327952 512829
rect 328188 512593 333882 512829
rect 334118 512593 339813 512829
rect 340049 512593 355952 512829
rect 356188 512593 361882 512829
rect 362118 512593 367813 512829
rect 368049 512593 383952 512829
rect 384188 512593 389882 512829
rect 390118 512593 395813 512829
rect 396049 512593 411952 512829
rect 412188 512593 417882 512829
rect 418118 512593 423813 512829
rect 424049 512593 439952 512829
rect 440188 512593 445882 512829
rect 446118 512593 451813 512829
rect 452049 512593 467952 512829
rect 468188 512593 473882 512829
rect 474118 512593 479813 512829
rect 480049 512593 495952 512829
rect 496188 512593 501882 512829
rect 502118 512593 507813 512829
rect 508049 512593 523952 512829
rect 524188 512593 529882 512829
rect 530118 512593 535813 512829
rect 536049 512593 551952 512829
rect 552188 512593 557882 512829
rect 558118 512593 563813 512829
rect 564049 512593 573526 512829
rect 573762 512593 573846 512829
rect 574082 512593 585342 512829
rect 585578 512593 585662 512829
rect 585898 512593 592650 512829
rect -8726 512509 592650 512593
rect -8726 512273 -1974 512509
rect -1738 512273 -1654 512509
rect -1418 512273 19952 512509
rect 20188 512273 25882 512509
rect 26118 512273 31813 512509
rect 32049 512273 47952 512509
rect 48188 512273 53882 512509
rect 54118 512273 59813 512509
rect 60049 512273 75952 512509
rect 76188 512273 81882 512509
rect 82118 512273 87813 512509
rect 88049 512273 103952 512509
rect 104188 512273 109882 512509
rect 110118 512273 115813 512509
rect 116049 512273 131952 512509
rect 132188 512273 137882 512509
rect 138118 512273 143813 512509
rect 144049 512273 159952 512509
rect 160188 512273 165882 512509
rect 166118 512273 171813 512509
rect 172049 512273 187952 512509
rect 188188 512273 193882 512509
rect 194118 512273 199813 512509
rect 200049 512273 215952 512509
rect 216188 512273 221882 512509
rect 222118 512273 227813 512509
rect 228049 512273 243952 512509
rect 244188 512273 249882 512509
rect 250118 512273 255813 512509
rect 256049 512273 271952 512509
rect 272188 512273 277882 512509
rect 278118 512273 283813 512509
rect 284049 512273 299952 512509
rect 300188 512273 305882 512509
rect 306118 512273 311813 512509
rect 312049 512273 327952 512509
rect 328188 512273 333882 512509
rect 334118 512273 339813 512509
rect 340049 512273 355952 512509
rect 356188 512273 361882 512509
rect 362118 512273 367813 512509
rect 368049 512273 383952 512509
rect 384188 512273 389882 512509
rect 390118 512273 395813 512509
rect 396049 512273 411952 512509
rect 412188 512273 417882 512509
rect 418118 512273 423813 512509
rect 424049 512273 439952 512509
rect 440188 512273 445882 512509
rect 446118 512273 451813 512509
rect 452049 512273 467952 512509
rect 468188 512273 473882 512509
rect 474118 512273 479813 512509
rect 480049 512273 495952 512509
rect 496188 512273 501882 512509
rect 502118 512273 507813 512509
rect 508049 512273 523952 512509
rect 524188 512273 529882 512509
rect 530118 512273 535813 512509
rect 536049 512273 551952 512509
rect 552188 512273 557882 512509
rect 558118 512273 563813 512509
rect 564049 512273 573526 512509
rect 573762 512273 573846 512509
rect 574082 512273 585342 512509
rect 585578 512273 585662 512509
rect 585898 512273 592650 512509
rect -8726 512241 592650 512273
rect -8726 509454 592650 509486
rect -8726 509218 -2934 509454
rect -2698 509218 -2614 509454
rect -2378 509218 22916 509454
rect 23152 509218 28847 509454
rect 29083 509218 50916 509454
rect 51152 509218 56847 509454
rect 57083 509218 78916 509454
rect 79152 509218 84847 509454
rect 85083 509218 106916 509454
rect 107152 509218 112847 509454
rect 113083 509218 134916 509454
rect 135152 509218 140847 509454
rect 141083 509218 162916 509454
rect 163152 509218 168847 509454
rect 169083 509218 190916 509454
rect 191152 509218 196847 509454
rect 197083 509218 218916 509454
rect 219152 509218 224847 509454
rect 225083 509218 246916 509454
rect 247152 509218 252847 509454
rect 253083 509218 274916 509454
rect 275152 509218 280847 509454
rect 281083 509218 302916 509454
rect 303152 509218 308847 509454
rect 309083 509218 330916 509454
rect 331152 509218 336847 509454
rect 337083 509218 358916 509454
rect 359152 509218 364847 509454
rect 365083 509218 386916 509454
rect 387152 509218 392847 509454
rect 393083 509218 414916 509454
rect 415152 509218 420847 509454
rect 421083 509218 442916 509454
rect 443152 509218 448847 509454
rect 449083 509218 470916 509454
rect 471152 509218 476847 509454
rect 477083 509218 498916 509454
rect 499152 509218 504847 509454
rect 505083 509218 526916 509454
rect 527152 509218 532847 509454
rect 533083 509218 554916 509454
rect 555152 509218 560847 509454
rect 561083 509218 586302 509454
rect 586538 509218 586622 509454
rect 586858 509218 592650 509454
rect -8726 509134 592650 509218
rect -8726 508898 -2934 509134
rect -2698 508898 -2614 509134
rect -2378 508898 22916 509134
rect 23152 508898 28847 509134
rect 29083 508898 50916 509134
rect 51152 508898 56847 509134
rect 57083 508898 78916 509134
rect 79152 508898 84847 509134
rect 85083 508898 106916 509134
rect 107152 508898 112847 509134
rect 113083 508898 134916 509134
rect 135152 508898 140847 509134
rect 141083 508898 162916 509134
rect 163152 508898 168847 509134
rect 169083 508898 190916 509134
rect 191152 508898 196847 509134
rect 197083 508898 218916 509134
rect 219152 508898 224847 509134
rect 225083 508898 246916 509134
rect 247152 508898 252847 509134
rect 253083 508898 274916 509134
rect 275152 508898 280847 509134
rect 281083 508898 302916 509134
rect 303152 508898 308847 509134
rect 309083 508898 330916 509134
rect 331152 508898 336847 509134
rect 337083 508898 358916 509134
rect 359152 508898 364847 509134
rect 365083 508898 386916 509134
rect 387152 508898 392847 509134
rect 393083 508898 414916 509134
rect 415152 508898 420847 509134
rect 421083 508898 442916 509134
rect 443152 508898 448847 509134
rect 449083 508898 470916 509134
rect 471152 508898 476847 509134
rect 477083 508898 498916 509134
rect 499152 508898 504847 509134
rect 505083 508898 526916 509134
rect 527152 508898 532847 509134
rect 533083 508898 554916 509134
rect 555152 508898 560847 509134
rect 561083 508898 586302 509134
rect 586538 508898 586622 509134
rect 586858 508898 592650 509134
rect -8726 508866 592650 508898
rect -8726 485829 592650 485861
rect -8726 485593 -1974 485829
rect -1738 485593 -1654 485829
rect -1418 485593 19951 485829
rect 20187 485593 25882 485829
rect 26118 485593 31812 485829
rect 32048 485593 47951 485829
rect 48187 485593 53882 485829
rect 54118 485593 59812 485829
rect 60048 485593 75951 485829
rect 76187 485593 81882 485829
rect 82118 485593 87812 485829
rect 88048 485593 103951 485829
rect 104187 485593 109882 485829
rect 110118 485593 115812 485829
rect 116048 485593 131951 485829
rect 132187 485593 137882 485829
rect 138118 485593 143812 485829
rect 144048 485593 159951 485829
rect 160187 485593 165882 485829
rect 166118 485593 171812 485829
rect 172048 485593 187951 485829
rect 188187 485593 193882 485829
rect 194118 485593 199812 485829
rect 200048 485593 215951 485829
rect 216187 485593 221882 485829
rect 222118 485593 227812 485829
rect 228048 485593 243951 485829
rect 244187 485593 249882 485829
rect 250118 485593 255812 485829
rect 256048 485593 271951 485829
rect 272187 485593 277882 485829
rect 278118 485593 283812 485829
rect 284048 485593 299951 485829
rect 300187 485593 305882 485829
rect 306118 485593 311812 485829
rect 312048 485593 327951 485829
rect 328187 485593 333882 485829
rect 334118 485593 339812 485829
rect 340048 485593 355951 485829
rect 356187 485593 361882 485829
rect 362118 485593 367812 485829
rect 368048 485593 383951 485829
rect 384187 485593 389882 485829
rect 390118 485593 395812 485829
rect 396048 485593 411951 485829
rect 412187 485593 417882 485829
rect 418118 485593 423812 485829
rect 424048 485593 439951 485829
rect 440187 485593 445882 485829
rect 446118 485593 451812 485829
rect 452048 485593 467951 485829
rect 468187 485593 473882 485829
rect 474118 485593 479812 485829
rect 480048 485593 495951 485829
rect 496187 485593 501882 485829
rect 502118 485593 507812 485829
rect 508048 485593 523951 485829
rect 524187 485593 529882 485829
rect 530118 485593 535812 485829
rect 536048 485593 551951 485829
rect 552187 485593 557882 485829
rect 558118 485593 563812 485829
rect 564048 485593 573526 485829
rect 573762 485593 573846 485829
rect 574082 485593 585342 485829
rect 585578 485593 585662 485829
rect 585898 485593 592650 485829
rect -8726 485509 592650 485593
rect -8726 485273 -1974 485509
rect -1738 485273 -1654 485509
rect -1418 485273 19951 485509
rect 20187 485273 25882 485509
rect 26118 485273 31812 485509
rect 32048 485273 47951 485509
rect 48187 485273 53882 485509
rect 54118 485273 59812 485509
rect 60048 485273 75951 485509
rect 76187 485273 81882 485509
rect 82118 485273 87812 485509
rect 88048 485273 103951 485509
rect 104187 485273 109882 485509
rect 110118 485273 115812 485509
rect 116048 485273 131951 485509
rect 132187 485273 137882 485509
rect 138118 485273 143812 485509
rect 144048 485273 159951 485509
rect 160187 485273 165882 485509
rect 166118 485273 171812 485509
rect 172048 485273 187951 485509
rect 188187 485273 193882 485509
rect 194118 485273 199812 485509
rect 200048 485273 215951 485509
rect 216187 485273 221882 485509
rect 222118 485273 227812 485509
rect 228048 485273 243951 485509
rect 244187 485273 249882 485509
rect 250118 485273 255812 485509
rect 256048 485273 271951 485509
rect 272187 485273 277882 485509
rect 278118 485273 283812 485509
rect 284048 485273 299951 485509
rect 300187 485273 305882 485509
rect 306118 485273 311812 485509
rect 312048 485273 327951 485509
rect 328187 485273 333882 485509
rect 334118 485273 339812 485509
rect 340048 485273 355951 485509
rect 356187 485273 361882 485509
rect 362118 485273 367812 485509
rect 368048 485273 383951 485509
rect 384187 485273 389882 485509
rect 390118 485273 395812 485509
rect 396048 485273 411951 485509
rect 412187 485273 417882 485509
rect 418118 485273 423812 485509
rect 424048 485273 439951 485509
rect 440187 485273 445882 485509
rect 446118 485273 451812 485509
rect 452048 485273 467951 485509
rect 468187 485273 473882 485509
rect 474118 485273 479812 485509
rect 480048 485273 495951 485509
rect 496187 485273 501882 485509
rect 502118 485273 507812 485509
rect 508048 485273 523951 485509
rect 524187 485273 529882 485509
rect 530118 485273 535812 485509
rect 536048 485273 551951 485509
rect 552187 485273 557882 485509
rect 558118 485273 563812 485509
rect 564048 485273 573526 485509
rect 573762 485273 573846 485509
rect 574082 485273 585342 485509
rect 585578 485273 585662 485509
rect 585898 485273 592650 485509
rect -8726 485241 592650 485273
rect -8726 482454 592650 482486
rect -8726 482218 -2934 482454
rect -2698 482218 -2614 482454
rect -2378 482218 22917 482454
rect 23153 482218 28848 482454
rect 29084 482218 50917 482454
rect 51153 482218 56848 482454
rect 57084 482218 78917 482454
rect 79153 482218 84848 482454
rect 85084 482218 106917 482454
rect 107153 482218 112848 482454
rect 113084 482218 134917 482454
rect 135153 482218 140848 482454
rect 141084 482218 162917 482454
rect 163153 482218 168848 482454
rect 169084 482218 190917 482454
rect 191153 482218 196848 482454
rect 197084 482218 218917 482454
rect 219153 482218 224848 482454
rect 225084 482218 246917 482454
rect 247153 482218 252848 482454
rect 253084 482218 274917 482454
rect 275153 482218 280848 482454
rect 281084 482218 302917 482454
rect 303153 482218 308848 482454
rect 309084 482218 330917 482454
rect 331153 482218 336848 482454
rect 337084 482218 358917 482454
rect 359153 482218 364848 482454
rect 365084 482218 386917 482454
rect 387153 482218 392848 482454
rect 393084 482218 414917 482454
rect 415153 482218 420848 482454
rect 421084 482218 442917 482454
rect 443153 482218 448848 482454
rect 449084 482218 470917 482454
rect 471153 482218 476848 482454
rect 477084 482218 498917 482454
rect 499153 482218 504848 482454
rect 505084 482218 526917 482454
rect 527153 482218 532848 482454
rect 533084 482218 554917 482454
rect 555153 482218 560848 482454
rect 561084 482218 586302 482454
rect 586538 482218 586622 482454
rect 586858 482218 592650 482454
rect -8726 482134 592650 482218
rect -8726 481898 -2934 482134
rect -2698 481898 -2614 482134
rect -2378 481898 22917 482134
rect 23153 481898 28848 482134
rect 29084 481898 50917 482134
rect 51153 481898 56848 482134
rect 57084 481898 78917 482134
rect 79153 481898 84848 482134
rect 85084 481898 106917 482134
rect 107153 481898 112848 482134
rect 113084 481898 134917 482134
rect 135153 481898 140848 482134
rect 141084 481898 162917 482134
rect 163153 481898 168848 482134
rect 169084 481898 190917 482134
rect 191153 481898 196848 482134
rect 197084 481898 218917 482134
rect 219153 481898 224848 482134
rect 225084 481898 246917 482134
rect 247153 481898 252848 482134
rect 253084 481898 274917 482134
rect 275153 481898 280848 482134
rect 281084 481898 302917 482134
rect 303153 481898 308848 482134
rect 309084 481898 330917 482134
rect 331153 481898 336848 482134
rect 337084 481898 358917 482134
rect 359153 481898 364848 482134
rect 365084 481898 386917 482134
rect 387153 481898 392848 482134
rect 393084 481898 414917 482134
rect 415153 481898 420848 482134
rect 421084 481898 442917 482134
rect 443153 481898 448848 482134
rect 449084 481898 470917 482134
rect 471153 481898 476848 482134
rect 477084 481898 498917 482134
rect 499153 481898 504848 482134
rect 505084 481898 526917 482134
rect 527153 481898 532848 482134
rect 533084 481898 554917 482134
rect 555153 481898 560848 482134
rect 561084 481898 586302 482134
rect 586538 481898 586622 482134
rect 586858 481898 592650 482134
rect -8726 481866 592650 481898
rect -8726 458829 592650 458861
rect -8726 458593 -1974 458829
rect -1738 458593 -1654 458829
rect -1418 458593 19952 458829
rect 20188 458593 25882 458829
rect 26118 458593 31813 458829
rect 32049 458593 47952 458829
rect 48188 458593 53882 458829
rect 54118 458593 59813 458829
rect 60049 458593 75952 458829
rect 76188 458593 81882 458829
rect 82118 458593 87813 458829
rect 88049 458593 103952 458829
rect 104188 458593 109882 458829
rect 110118 458593 115813 458829
rect 116049 458593 131952 458829
rect 132188 458593 137882 458829
rect 138118 458593 143813 458829
rect 144049 458593 159952 458829
rect 160188 458593 165882 458829
rect 166118 458593 171813 458829
rect 172049 458593 187952 458829
rect 188188 458593 193882 458829
rect 194118 458593 199813 458829
rect 200049 458593 215952 458829
rect 216188 458593 221882 458829
rect 222118 458593 227813 458829
rect 228049 458593 243952 458829
rect 244188 458593 249882 458829
rect 250118 458593 255813 458829
rect 256049 458593 271952 458829
rect 272188 458593 277882 458829
rect 278118 458593 283813 458829
rect 284049 458593 299952 458829
rect 300188 458593 305882 458829
rect 306118 458593 311813 458829
rect 312049 458593 327952 458829
rect 328188 458593 333882 458829
rect 334118 458593 339813 458829
rect 340049 458593 355952 458829
rect 356188 458593 361882 458829
rect 362118 458593 367813 458829
rect 368049 458593 383952 458829
rect 384188 458593 389882 458829
rect 390118 458593 395813 458829
rect 396049 458593 411952 458829
rect 412188 458593 417882 458829
rect 418118 458593 423813 458829
rect 424049 458593 439952 458829
rect 440188 458593 445882 458829
rect 446118 458593 451813 458829
rect 452049 458593 467952 458829
rect 468188 458593 473882 458829
rect 474118 458593 479813 458829
rect 480049 458593 495952 458829
rect 496188 458593 501882 458829
rect 502118 458593 507813 458829
rect 508049 458593 523952 458829
rect 524188 458593 529882 458829
rect 530118 458593 535813 458829
rect 536049 458593 551952 458829
rect 552188 458593 557882 458829
rect 558118 458593 563813 458829
rect 564049 458593 573526 458829
rect 573762 458593 573846 458829
rect 574082 458593 585342 458829
rect 585578 458593 585662 458829
rect 585898 458593 592650 458829
rect -8726 458509 592650 458593
rect -8726 458273 -1974 458509
rect -1738 458273 -1654 458509
rect -1418 458273 19952 458509
rect 20188 458273 25882 458509
rect 26118 458273 31813 458509
rect 32049 458273 47952 458509
rect 48188 458273 53882 458509
rect 54118 458273 59813 458509
rect 60049 458273 75952 458509
rect 76188 458273 81882 458509
rect 82118 458273 87813 458509
rect 88049 458273 103952 458509
rect 104188 458273 109882 458509
rect 110118 458273 115813 458509
rect 116049 458273 131952 458509
rect 132188 458273 137882 458509
rect 138118 458273 143813 458509
rect 144049 458273 159952 458509
rect 160188 458273 165882 458509
rect 166118 458273 171813 458509
rect 172049 458273 187952 458509
rect 188188 458273 193882 458509
rect 194118 458273 199813 458509
rect 200049 458273 215952 458509
rect 216188 458273 221882 458509
rect 222118 458273 227813 458509
rect 228049 458273 243952 458509
rect 244188 458273 249882 458509
rect 250118 458273 255813 458509
rect 256049 458273 271952 458509
rect 272188 458273 277882 458509
rect 278118 458273 283813 458509
rect 284049 458273 299952 458509
rect 300188 458273 305882 458509
rect 306118 458273 311813 458509
rect 312049 458273 327952 458509
rect 328188 458273 333882 458509
rect 334118 458273 339813 458509
rect 340049 458273 355952 458509
rect 356188 458273 361882 458509
rect 362118 458273 367813 458509
rect 368049 458273 383952 458509
rect 384188 458273 389882 458509
rect 390118 458273 395813 458509
rect 396049 458273 411952 458509
rect 412188 458273 417882 458509
rect 418118 458273 423813 458509
rect 424049 458273 439952 458509
rect 440188 458273 445882 458509
rect 446118 458273 451813 458509
rect 452049 458273 467952 458509
rect 468188 458273 473882 458509
rect 474118 458273 479813 458509
rect 480049 458273 495952 458509
rect 496188 458273 501882 458509
rect 502118 458273 507813 458509
rect 508049 458273 523952 458509
rect 524188 458273 529882 458509
rect 530118 458273 535813 458509
rect 536049 458273 551952 458509
rect 552188 458273 557882 458509
rect 558118 458273 563813 458509
rect 564049 458273 573526 458509
rect 573762 458273 573846 458509
rect 574082 458273 585342 458509
rect 585578 458273 585662 458509
rect 585898 458273 592650 458509
rect -8726 458241 592650 458273
rect -8726 455454 592650 455486
rect -8726 455218 -2934 455454
rect -2698 455218 -2614 455454
rect -2378 455218 22916 455454
rect 23152 455218 28847 455454
rect 29083 455218 50916 455454
rect 51152 455218 56847 455454
rect 57083 455218 78916 455454
rect 79152 455218 84847 455454
rect 85083 455218 106916 455454
rect 107152 455218 112847 455454
rect 113083 455218 134916 455454
rect 135152 455218 140847 455454
rect 141083 455218 162916 455454
rect 163152 455218 168847 455454
rect 169083 455218 190916 455454
rect 191152 455218 196847 455454
rect 197083 455218 218916 455454
rect 219152 455218 224847 455454
rect 225083 455218 246916 455454
rect 247152 455218 252847 455454
rect 253083 455218 274916 455454
rect 275152 455218 280847 455454
rect 281083 455218 302916 455454
rect 303152 455218 308847 455454
rect 309083 455218 330916 455454
rect 331152 455218 336847 455454
rect 337083 455218 358916 455454
rect 359152 455218 364847 455454
rect 365083 455218 386916 455454
rect 387152 455218 392847 455454
rect 393083 455218 414916 455454
rect 415152 455218 420847 455454
rect 421083 455218 442916 455454
rect 443152 455218 448847 455454
rect 449083 455218 470916 455454
rect 471152 455218 476847 455454
rect 477083 455218 498916 455454
rect 499152 455218 504847 455454
rect 505083 455218 526916 455454
rect 527152 455218 532847 455454
rect 533083 455218 554916 455454
rect 555152 455218 560847 455454
rect 561083 455218 586302 455454
rect 586538 455218 586622 455454
rect 586858 455218 592650 455454
rect -8726 455134 592650 455218
rect -8726 454898 -2934 455134
rect -2698 454898 -2614 455134
rect -2378 454898 22916 455134
rect 23152 454898 28847 455134
rect 29083 454898 50916 455134
rect 51152 454898 56847 455134
rect 57083 454898 78916 455134
rect 79152 454898 84847 455134
rect 85083 454898 106916 455134
rect 107152 454898 112847 455134
rect 113083 454898 134916 455134
rect 135152 454898 140847 455134
rect 141083 454898 162916 455134
rect 163152 454898 168847 455134
rect 169083 454898 190916 455134
rect 191152 454898 196847 455134
rect 197083 454898 218916 455134
rect 219152 454898 224847 455134
rect 225083 454898 246916 455134
rect 247152 454898 252847 455134
rect 253083 454898 274916 455134
rect 275152 454898 280847 455134
rect 281083 454898 302916 455134
rect 303152 454898 308847 455134
rect 309083 454898 330916 455134
rect 331152 454898 336847 455134
rect 337083 454898 358916 455134
rect 359152 454898 364847 455134
rect 365083 454898 386916 455134
rect 387152 454898 392847 455134
rect 393083 454898 414916 455134
rect 415152 454898 420847 455134
rect 421083 454898 442916 455134
rect 443152 454898 448847 455134
rect 449083 454898 470916 455134
rect 471152 454898 476847 455134
rect 477083 454898 498916 455134
rect 499152 454898 504847 455134
rect 505083 454898 526916 455134
rect 527152 454898 532847 455134
rect 533083 454898 554916 455134
rect 555152 454898 560847 455134
rect 561083 454898 586302 455134
rect 586538 454898 586622 455134
rect 586858 454898 592650 455134
rect -8726 454866 592650 454898
rect -8726 431829 592650 431861
rect -8726 431593 -1974 431829
rect -1738 431593 -1654 431829
rect -1418 431593 19951 431829
rect 20187 431593 25882 431829
rect 26118 431593 31812 431829
rect 32048 431593 47951 431829
rect 48187 431593 53882 431829
rect 54118 431593 59812 431829
rect 60048 431593 75951 431829
rect 76187 431593 81882 431829
rect 82118 431593 87812 431829
rect 88048 431593 103951 431829
rect 104187 431593 109882 431829
rect 110118 431593 115812 431829
rect 116048 431593 131951 431829
rect 132187 431593 137882 431829
rect 138118 431593 143812 431829
rect 144048 431593 159951 431829
rect 160187 431593 165882 431829
rect 166118 431593 171812 431829
rect 172048 431593 187951 431829
rect 188187 431593 193882 431829
rect 194118 431593 199812 431829
rect 200048 431593 215951 431829
rect 216187 431593 221882 431829
rect 222118 431593 227812 431829
rect 228048 431593 243951 431829
rect 244187 431593 249882 431829
rect 250118 431593 255812 431829
rect 256048 431593 271951 431829
rect 272187 431593 277882 431829
rect 278118 431593 283812 431829
rect 284048 431593 299951 431829
rect 300187 431593 305882 431829
rect 306118 431593 311812 431829
rect 312048 431593 327951 431829
rect 328187 431593 333882 431829
rect 334118 431593 339812 431829
rect 340048 431593 355951 431829
rect 356187 431593 361882 431829
rect 362118 431593 367812 431829
rect 368048 431593 383951 431829
rect 384187 431593 389882 431829
rect 390118 431593 395812 431829
rect 396048 431593 411951 431829
rect 412187 431593 417882 431829
rect 418118 431593 423812 431829
rect 424048 431593 439951 431829
rect 440187 431593 445882 431829
rect 446118 431593 451812 431829
rect 452048 431593 467951 431829
rect 468187 431593 473882 431829
rect 474118 431593 479812 431829
rect 480048 431593 495951 431829
rect 496187 431593 501882 431829
rect 502118 431593 507812 431829
rect 508048 431593 523951 431829
rect 524187 431593 529882 431829
rect 530118 431593 535812 431829
rect 536048 431593 551951 431829
rect 552187 431593 557882 431829
rect 558118 431593 563812 431829
rect 564048 431593 573526 431829
rect 573762 431593 573846 431829
rect 574082 431593 585342 431829
rect 585578 431593 585662 431829
rect 585898 431593 592650 431829
rect -8726 431509 592650 431593
rect -8726 431273 -1974 431509
rect -1738 431273 -1654 431509
rect -1418 431273 19951 431509
rect 20187 431273 25882 431509
rect 26118 431273 31812 431509
rect 32048 431273 47951 431509
rect 48187 431273 53882 431509
rect 54118 431273 59812 431509
rect 60048 431273 75951 431509
rect 76187 431273 81882 431509
rect 82118 431273 87812 431509
rect 88048 431273 103951 431509
rect 104187 431273 109882 431509
rect 110118 431273 115812 431509
rect 116048 431273 131951 431509
rect 132187 431273 137882 431509
rect 138118 431273 143812 431509
rect 144048 431273 159951 431509
rect 160187 431273 165882 431509
rect 166118 431273 171812 431509
rect 172048 431273 187951 431509
rect 188187 431273 193882 431509
rect 194118 431273 199812 431509
rect 200048 431273 215951 431509
rect 216187 431273 221882 431509
rect 222118 431273 227812 431509
rect 228048 431273 243951 431509
rect 244187 431273 249882 431509
rect 250118 431273 255812 431509
rect 256048 431273 271951 431509
rect 272187 431273 277882 431509
rect 278118 431273 283812 431509
rect 284048 431273 299951 431509
rect 300187 431273 305882 431509
rect 306118 431273 311812 431509
rect 312048 431273 327951 431509
rect 328187 431273 333882 431509
rect 334118 431273 339812 431509
rect 340048 431273 355951 431509
rect 356187 431273 361882 431509
rect 362118 431273 367812 431509
rect 368048 431273 383951 431509
rect 384187 431273 389882 431509
rect 390118 431273 395812 431509
rect 396048 431273 411951 431509
rect 412187 431273 417882 431509
rect 418118 431273 423812 431509
rect 424048 431273 439951 431509
rect 440187 431273 445882 431509
rect 446118 431273 451812 431509
rect 452048 431273 467951 431509
rect 468187 431273 473882 431509
rect 474118 431273 479812 431509
rect 480048 431273 495951 431509
rect 496187 431273 501882 431509
rect 502118 431273 507812 431509
rect 508048 431273 523951 431509
rect 524187 431273 529882 431509
rect 530118 431273 535812 431509
rect 536048 431273 551951 431509
rect 552187 431273 557882 431509
rect 558118 431273 563812 431509
rect 564048 431273 573526 431509
rect 573762 431273 573846 431509
rect 574082 431273 585342 431509
rect 585578 431273 585662 431509
rect 585898 431273 592650 431509
rect -8726 431241 592650 431273
rect -8726 428454 592650 428486
rect -8726 428218 -2934 428454
rect -2698 428218 -2614 428454
rect -2378 428218 22917 428454
rect 23153 428218 28848 428454
rect 29084 428218 50917 428454
rect 51153 428218 56848 428454
rect 57084 428218 78917 428454
rect 79153 428218 84848 428454
rect 85084 428218 106917 428454
rect 107153 428218 112848 428454
rect 113084 428218 134917 428454
rect 135153 428218 140848 428454
rect 141084 428218 162917 428454
rect 163153 428218 168848 428454
rect 169084 428218 190917 428454
rect 191153 428218 196848 428454
rect 197084 428218 218917 428454
rect 219153 428218 224848 428454
rect 225084 428218 246917 428454
rect 247153 428218 252848 428454
rect 253084 428218 274917 428454
rect 275153 428218 280848 428454
rect 281084 428218 302917 428454
rect 303153 428218 308848 428454
rect 309084 428218 330917 428454
rect 331153 428218 336848 428454
rect 337084 428218 358917 428454
rect 359153 428218 364848 428454
rect 365084 428218 386917 428454
rect 387153 428218 392848 428454
rect 393084 428218 414917 428454
rect 415153 428218 420848 428454
rect 421084 428218 442917 428454
rect 443153 428218 448848 428454
rect 449084 428218 470917 428454
rect 471153 428218 476848 428454
rect 477084 428218 498917 428454
rect 499153 428218 504848 428454
rect 505084 428218 526917 428454
rect 527153 428218 532848 428454
rect 533084 428218 554917 428454
rect 555153 428218 560848 428454
rect 561084 428218 586302 428454
rect 586538 428218 586622 428454
rect 586858 428218 592650 428454
rect -8726 428134 592650 428218
rect -8726 427898 -2934 428134
rect -2698 427898 -2614 428134
rect -2378 427898 22917 428134
rect 23153 427898 28848 428134
rect 29084 427898 50917 428134
rect 51153 427898 56848 428134
rect 57084 427898 78917 428134
rect 79153 427898 84848 428134
rect 85084 427898 106917 428134
rect 107153 427898 112848 428134
rect 113084 427898 134917 428134
rect 135153 427898 140848 428134
rect 141084 427898 162917 428134
rect 163153 427898 168848 428134
rect 169084 427898 190917 428134
rect 191153 427898 196848 428134
rect 197084 427898 218917 428134
rect 219153 427898 224848 428134
rect 225084 427898 246917 428134
rect 247153 427898 252848 428134
rect 253084 427898 274917 428134
rect 275153 427898 280848 428134
rect 281084 427898 302917 428134
rect 303153 427898 308848 428134
rect 309084 427898 330917 428134
rect 331153 427898 336848 428134
rect 337084 427898 358917 428134
rect 359153 427898 364848 428134
rect 365084 427898 386917 428134
rect 387153 427898 392848 428134
rect 393084 427898 414917 428134
rect 415153 427898 420848 428134
rect 421084 427898 442917 428134
rect 443153 427898 448848 428134
rect 449084 427898 470917 428134
rect 471153 427898 476848 428134
rect 477084 427898 498917 428134
rect 499153 427898 504848 428134
rect 505084 427898 526917 428134
rect 527153 427898 532848 428134
rect 533084 427898 554917 428134
rect 555153 427898 560848 428134
rect 561084 427898 586302 428134
rect 586538 427898 586622 428134
rect 586858 427898 592650 428134
rect -8726 427866 592650 427898
rect -8726 404829 592650 404861
rect -8726 404593 -1974 404829
rect -1738 404593 -1654 404829
rect -1418 404593 19952 404829
rect 20188 404593 25882 404829
rect 26118 404593 31813 404829
rect 32049 404593 47952 404829
rect 48188 404593 53882 404829
rect 54118 404593 59813 404829
rect 60049 404593 75952 404829
rect 76188 404593 81882 404829
rect 82118 404593 87813 404829
rect 88049 404593 103952 404829
rect 104188 404593 109882 404829
rect 110118 404593 115813 404829
rect 116049 404593 131952 404829
rect 132188 404593 137882 404829
rect 138118 404593 143813 404829
rect 144049 404593 159952 404829
rect 160188 404593 165882 404829
rect 166118 404593 171813 404829
rect 172049 404593 187952 404829
rect 188188 404593 193882 404829
rect 194118 404593 199813 404829
rect 200049 404593 215952 404829
rect 216188 404593 221882 404829
rect 222118 404593 227813 404829
rect 228049 404593 243952 404829
rect 244188 404593 249882 404829
rect 250118 404593 255813 404829
rect 256049 404593 271952 404829
rect 272188 404593 277882 404829
rect 278118 404593 283813 404829
rect 284049 404593 299952 404829
rect 300188 404593 305882 404829
rect 306118 404593 311813 404829
rect 312049 404593 327952 404829
rect 328188 404593 333882 404829
rect 334118 404593 339813 404829
rect 340049 404593 355952 404829
rect 356188 404593 361882 404829
rect 362118 404593 367813 404829
rect 368049 404593 383952 404829
rect 384188 404593 389882 404829
rect 390118 404593 395813 404829
rect 396049 404593 411952 404829
rect 412188 404593 417882 404829
rect 418118 404593 423813 404829
rect 424049 404593 439952 404829
rect 440188 404593 445882 404829
rect 446118 404593 451813 404829
rect 452049 404593 467952 404829
rect 468188 404593 473882 404829
rect 474118 404593 479813 404829
rect 480049 404593 495952 404829
rect 496188 404593 501882 404829
rect 502118 404593 507813 404829
rect 508049 404593 523952 404829
rect 524188 404593 529882 404829
rect 530118 404593 535813 404829
rect 536049 404593 551952 404829
rect 552188 404593 557882 404829
rect 558118 404593 563813 404829
rect 564049 404593 573526 404829
rect 573762 404593 573846 404829
rect 574082 404593 585342 404829
rect 585578 404593 585662 404829
rect 585898 404593 592650 404829
rect -8726 404509 592650 404593
rect -8726 404273 -1974 404509
rect -1738 404273 -1654 404509
rect -1418 404273 19952 404509
rect 20188 404273 25882 404509
rect 26118 404273 31813 404509
rect 32049 404273 47952 404509
rect 48188 404273 53882 404509
rect 54118 404273 59813 404509
rect 60049 404273 75952 404509
rect 76188 404273 81882 404509
rect 82118 404273 87813 404509
rect 88049 404273 103952 404509
rect 104188 404273 109882 404509
rect 110118 404273 115813 404509
rect 116049 404273 131952 404509
rect 132188 404273 137882 404509
rect 138118 404273 143813 404509
rect 144049 404273 159952 404509
rect 160188 404273 165882 404509
rect 166118 404273 171813 404509
rect 172049 404273 187952 404509
rect 188188 404273 193882 404509
rect 194118 404273 199813 404509
rect 200049 404273 215952 404509
rect 216188 404273 221882 404509
rect 222118 404273 227813 404509
rect 228049 404273 243952 404509
rect 244188 404273 249882 404509
rect 250118 404273 255813 404509
rect 256049 404273 271952 404509
rect 272188 404273 277882 404509
rect 278118 404273 283813 404509
rect 284049 404273 299952 404509
rect 300188 404273 305882 404509
rect 306118 404273 311813 404509
rect 312049 404273 327952 404509
rect 328188 404273 333882 404509
rect 334118 404273 339813 404509
rect 340049 404273 355952 404509
rect 356188 404273 361882 404509
rect 362118 404273 367813 404509
rect 368049 404273 383952 404509
rect 384188 404273 389882 404509
rect 390118 404273 395813 404509
rect 396049 404273 411952 404509
rect 412188 404273 417882 404509
rect 418118 404273 423813 404509
rect 424049 404273 439952 404509
rect 440188 404273 445882 404509
rect 446118 404273 451813 404509
rect 452049 404273 467952 404509
rect 468188 404273 473882 404509
rect 474118 404273 479813 404509
rect 480049 404273 495952 404509
rect 496188 404273 501882 404509
rect 502118 404273 507813 404509
rect 508049 404273 523952 404509
rect 524188 404273 529882 404509
rect 530118 404273 535813 404509
rect 536049 404273 551952 404509
rect 552188 404273 557882 404509
rect 558118 404273 563813 404509
rect 564049 404273 573526 404509
rect 573762 404273 573846 404509
rect 574082 404273 585342 404509
rect 585578 404273 585662 404509
rect 585898 404273 592650 404509
rect -8726 404241 592650 404273
rect -8726 401454 592650 401486
rect -8726 401218 -2934 401454
rect -2698 401218 -2614 401454
rect -2378 401218 22916 401454
rect 23152 401218 28847 401454
rect 29083 401218 50916 401454
rect 51152 401218 56847 401454
rect 57083 401218 78916 401454
rect 79152 401218 84847 401454
rect 85083 401218 106916 401454
rect 107152 401218 112847 401454
rect 113083 401218 134916 401454
rect 135152 401218 140847 401454
rect 141083 401218 162916 401454
rect 163152 401218 168847 401454
rect 169083 401218 190916 401454
rect 191152 401218 196847 401454
rect 197083 401218 218916 401454
rect 219152 401218 224847 401454
rect 225083 401218 246916 401454
rect 247152 401218 252847 401454
rect 253083 401218 274916 401454
rect 275152 401218 280847 401454
rect 281083 401218 302916 401454
rect 303152 401218 308847 401454
rect 309083 401218 330916 401454
rect 331152 401218 336847 401454
rect 337083 401218 358916 401454
rect 359152 401218 364847 401454
rect 365083 401218 386916 401454
rect 387152 401218 392847 401454
rect 393083 401218 414916 401454
rect 415152 401218 420847 401454
rect 421083 401218 442916 401454
rect 443152 401218 448847 401454
rect 449083 401218 470916 401454
rect 471152 401218 476847 401454
rect 477083 401218 498916 401454
rect 499152 401218 504847 401454
rect 505083 401218 526916 401454
rect 527152 401218 532847 401454
rect 533083 401218 554916 401454
rect 555152 401218 560847 401454
rect 561083 401218 586302 401454
rect 586538 401218 586622 401454
rect 586858 401218 592650 401454
rect -8726 401134 592650 401218
rect -8726 400898 -2934 401134
rect -2698 400898 -2614 401134
rect -2378 400898 22916 401134
rect 23152 400898 28847 401134
rect 29083 400898 50916 401134
rect 51152 400898 56847 401134
rect 57083 400898 78916 401134
rect 79152 400898 84847 401134
rect 85083 400898 106916 401134
rect 107152 400898 112847 401134
rect 113083 400898 134916 401134
rect 135152 400898 140847 401134
rect 141083 400898 162916 401134
rect 163152 400898 168847 401134
rect 169083 400898 190916 401134
rect 191152 400898 196847 401134
rect 197083 400898 218916 401134
rect 219152 400898 224847 401134
rect 225083 400898 246916 401134
rect 247152 400898 252847 401134
rect 253083 400898 274916 401134
rect 275152 400898 280847 401134
rect 281083 400898 302916 401134
rect 303152 400898 308847 401134
rect 309083 400898 330916 401134
rect 331152 400898 336847 401134
rect 337083 400898 358916 401134
rect 359152 400898 364847 401134
rect 365083 400898 386916 401134
rect 387152 400898 392847 401134
rect 393083 400898 414916 401134
rect 415152 400898 420847 401134
rect 421083 400898 442916 401134
rect 443152 400898 448847 401134
rect 449083 400898 470916 401134
rect 471152 400898 476847 401134
rect 477083 400898 498916 401134
rect 499152 400898 504847 401134
rect 505083 400898 526916 401134
rect 527152 400898 532847 401134
rect 533083 400898 554916 401134
rect 555152 400898 560847 401134
rect 561083 400898 586302 401134
rect 586538 400898 586622 401134
rect 586858 400898 592650 401134
rect -8726 400866 592650 400898
rect -8726 377829 592650 377861
rect -8726 377593 -1974 377829
rect -1738 377593 -1654 377829
rect -1418 377593 19951 377829
rect 20187 377593 25882 377829
rect 26118 377593 31812 377829
rect 32048 377593 47951 377829
rect 48187 377593 53882 377829
rect 54118 377593 59812 377829
rect 60048 377593 75951 377829
rect 76187 377593 81882 377829
rect 82118 377593 87812 377829
rect 88048 377593 103951 377829
rect 104187 377593 109882 377829
rect 110118 377593 115812 377829
rect 116048 377593 131951 377829
rect 132187 377593 137882 377829
rect 138118 377593 143812 377829
rect 144048 377593 159951 377829
rect 160187 377593 165882 377829
rect 166118 377593 171812 377829
rect 172048 377593 187951 377829
rect 188187 377593 193882 377829
rect 194118 377593 199812 377829
rect 200048 377593 215951 377829
rect 216187 377593 221882 377829
rect 222118 377593 227812 377829
rect 228048 377593 243951 377829
rect 244187 377593 249882 377829
rect 250118 377593 255812 377829
rect 256048 377593 271951 377829
rect 272187 377593 277882 377829
rect 278118 377593 283812 377829
rect 284048 377593 299951 377829
rect 300187 377593 305882 377829
rect 306118 377593 311812 377829
rect 312048 377593 327951 377829
rect 328187 377593 333882 377829
rect 334118 377593 339812 377829
rect 340048 377593 355951 377829
rect 356187 377593 361882 377829
rect 362118 377593 367812 377829
rect 368048 377593 383951 377829
rect 384187 377593 389882 377829
rect 390118 377593 395812 377829
rect 396048 377593 411951 377829
rect 412187 377593 417882 377829
rect 418118 377593 423812 377829
rect 424048 377593 439951 377829
rect 440187 377593 445882 377829
rect 446118 377593 451812 377829
rect 452048 377593 467951 377829
rect 468187 377593 473882 377829
rect 474118 377593 479812 377829
rect 480048 377593 495951 377829
rect 496187 377593 501882 377829
rect 502118 377593 507812 377829
rect 508048 377593 523951 377829
rect 524187 377593 529882 377829
rect 530118 377593 535812 377829
rect 536048 377593 551951 377829
rect 552187 377593 557882 377829
rect 558118 377593 563812 377829
rect 564048 377593 573526 377829
rect 573762 377593 573846 377829
rect 574082 377593 585342 377829
rect 585578 377593 585662 377829
rect 585898 377593 592650 377829
rect -8726 377509 592650 377593
rect -8726 377273 -1974 377509
rect -1738 377273 -1654 377509
rect -1418 377273 19951 377509
rect 20187 377273 25882 377509
rect 26118 377273 31812 377509
rect 32048 377273 47951 377509
rect 48187 377273 53882 377509
rect 54118 377273 59812 377509
rect 60048 377273 75951 377509
rect 76187 377273 81882 377509
rect 82118 377273 87812 377509
rect 88048 377273 103951 377509
rect 104187 377273 109882 377509
rect 110118 377273 115812 377509
rect 116048 377273 131951 377509
rect 132187 377273 137882 377509
rect 138118 377273 143812 377509
rect 144048 377273 159951 377509
rect 160187 377273 165882 377509
rect 166118 377273 171812 377509
rect 172048 377273 187951 377509
rect 188187 377273 193882 377509
rect 194118 377273 199812 377509
rect 200048 377273 215951 377509
rect 216187 377273 221882 377509
rect 222118 377273 227812 377509
rect 228048 377273 243951 377509
rect 244187 377273 249882 377509
rect 250118 377273 255812 377509
rect 256048 377273 271951 377509
rect 272187 377273 277882 377509
rect 278118 377273 283812 377509
rect 284048 377273 299951 377509
rect 300187 377273 305882 377509
rect 306118 377273 311812 377509
rect 312048 377273 327951 377509
rect 328187 377273 333882 377509
rect 334118 377273 339812 377509
rect 340048 377273 355951 377509
rect 356187 377273 361882 377509
rect 362118 377273 367812 377509
rect 368048 377273 383951 377509
rect 384187 377273 389882 377509
rect 390118 377273 395812 377509
rect 396048 377273 411951 377509
rect 412187 377273 417882 377509
rect 418118 377273 423812 377509
rect 424048 377273 439951 377509
rect 440187 377273 445882 377509
rect 446118 377273 451812 377509
rect 452048 377273 467951 377509
rect 468187 377273 473882 377509
rect 474118 377273 479812 377509
rect 480048 377273 495951 377509
rect 496187 377273 501882 377509
rect 502118 377273 507812 377509
rect 508048 377273 523951 377509
rect 524187 377273 529882 377509
rect 530118 377273 535812 377509
rect 536048 377273 551951 377509
rect 552187 377273 557882 377509
rect 558118 377273 563812 377509
rect 564048 377273 573526 377509
rect 573762 377273 573846 377509
rect 574082 377273 585342 377509
rect 585578 377273 585662 377509
rect 585898 377273 592650 377509
rect -8726 377241 592650 377273
rect -8726 374454 592650 374486
rect -8726 374218 -2934 374454
rect -2698 374218 -2614 374454
rect -2378 374218 22917 374454
rect 23153 374218 28848 374454
rect 29084 374218 50917 374454
rect 51153 374218 56848 374454
rect 57084 374218 78917 374454
rect 79153 374218 84848 374454
rect 85084 374218 106917 374454
rect 107153 374218 112848 374454
rect 113084 374218 134917 374454
rect 135153 374218 140848 374454
rect 141084 374218 162917 374454
rect 163153 374218 168848 374454
rect 169084 374218 190917 374454
rect 191153 374218 196848 374454
rect 197084 374218 218917 374454
rect 219153 374218 224848 374454
rect 225084 374218 246917 374454
rect 247153 374218 252848 374454
rect 253084 374218 274917 374454
rect 275153 374218 280848 374454
rect 281084 374218 302917 374454
rect 303153 374218 308848 374454
rect 309084 374218 330917 374454
rect 331153 374218 336848 374454
rect 337084 374218 358917 374454
rect 359153 374218 364848 374454
rect 365084 374218 386917 374454
rect 387153 374218 392848 374454
rect 393084 374218 414917 374454
rect 415153 374218 420848 374454
rect 421084 374218 442917 374454
rect 443153 374218 448848 374454
rect 449084 374218 470917 374454
rect 471153 374218 476848 374454
rect 477084 374218 498917 374454
rect 499153 374218 504848 374454
rect 505084 374218 526917 374454
rect 527153 374218 532848 374454
rect 533084 374218 554917 374454
rect 555153 374218 560848 374454
rect 561084 374218 586302 374454
rect 586538 374218 586622 374454
rect 586858 374218 592650 374454
rect -8726 374134 592650 374218
rect -8726 373898 -2934 374134
rect -2698 373898 -2614 374134
rect -2378 373898 22917 374134
rect 23153 373898 28848 374134
rect 29084 373898 50917 374134
rect 51153 373898 56848 374134
rect 57084 373898 78917 374134
rect 79153 373898 84848 374134
rect 85084 373898 106917 374134
rect 107153 373898 112848 374134
rect 113084 373898 134917 374134
rect 135153 373898 140848 374134
rect 141084 373898 162917 374134
rect 163153 373898 168848 374134
rect 169084 373898 190917 374134
rect 191153 373898 196848 374134
rect 197084 373898 218917 374134
rect 219153 373898 224848 374134
rect 225084 373898 246917 374134
rect 247153 373898 252848 374134
rect 253084 373898 274917 374134
rect 275153 373898 280848 374134
rect 281084 373898 302917 374134
rect 303153 373898 308848 374134
rect 309084 373898 330917 374134
rect 331153 373898 336848 374134
rect 337084 373898 358917 374134
rect 359153 373898 364848 374134
rect 365084 373898 386917 374134
rect 387153 373898 392848 374134
rect 393084 373898 414917 374134
rect 415153 373898 420848 374134
rect 421084 373898 442917 374134
rect 443153 373898 448848 374134
rect 449084 373898 470917 374134
rect 471153 373898 476848 374134
rect 477084 373898 498917 374134
rect 499153 373898 504848 374134
rect 505084 373898 526917 374134
rect 527153 373898 532848 374134
rect 533084 373898 554917 374134
rect 555153 373898 560848 374134
rect 561084 373898 586302 374134
rect 586538 373898 586622 374134
rect 586858 373898 592650 374134
rect -8726 373866 592650 373898
rect -8726 350829 592650 350861
rect -8726 350593 -1974 350829
rect -1738 350593 -1654 350829
rect -1418 350593 19952 350829
rect 20188 350593 25882 350829
rect 26118 350593 31813 350829
rect 32049 350593 47952 350829
rect 48188 350593 53882 350829
rect 54118 350593 59813 350829
rect 60049 350593 75952 350829
rect 76188 350593 81882 350829
rect 82118 350593 87813 350829
rect 88049 350593 103952 350829
rect 104188 350593 109882 350829
rect 110118 350593 115813 350829
rect 116049 350593 131952 350829
rect 132188 350593 137882 350829
rect 138118 350593 143813 350829
rect 144049 350593 159952 350829
rect 160188 350593 165882 350829
rect 166118 350593 171813 350829
rect 172049 350593 187952 350829
rect 188188 350593 193882 350829
rect 194118 350593 199813 350829
rect 200049 350593 215952 350829
rect 216188 350593 221882 350829
rect 222118 350593 227813 350829
rect 228049 350593 243952 350829
rect 244188 350593 249882 350829
rect 250118 350593 255813 350829
rect 256049 350593 271952 350829
rect 272188 350593 277882 350829
rect 278118 350593 283813 350829
rect 284049 350593 299952 350829
rect 300188 350593 305882 350829
rect 306118 350593 311813 350829
rect 312049 350593 327952 350829
rect 328188 350593 333882 350829
rect 334118 350593 339813 350829
rect 340049 350593 355952 350829
rect 356188 350593 361882 350829
rect 362118 350593 367813 350829
rect 368049 350593 383952 350829
rect 384188 350593 389882 350829
rect 390118 350593 395813 350829
rect 396049 350593 411952 350829
rect 412188 350593 417882 350829
rect 418118 350593 423813 350829
rect 424049 350593 439952 350829
rect 440188 350593 445882 350829
rect 446118 350593 451813 350829
rect 452049 350593 467952 350829
rect 468188 350593 473882 350829
rect 474118 350593 479813 350829
rect 480049 350593 495952 350829
rect 496188 350593 501882 350829
rect 502118 350593 507813 350829
rect 508049 350593 523952 350829
rect 524188 350593 529882 350829
rect 530118 350593 535813 350829
rect 536049 350593 551952 350829
rect 552188 350593 557882 350829
rect 558118 350593 563813 350829
rect 564049 350593 573526 350829
rect 573762 350593 573846 350829
rect 574082 350593 585342 350829
rect 585578 350593 585662 350829
rect 585898 350593 592650 350829
rect -8726 350509 592650 350593
rect -8726 350273 -1974 350509
rect -1738 350273 -1654 350509
rect -1418 350273 19952 350509
rect 20188 350273 25882 350509
rect 26118 350273 31813 350509
rect 32049 350273 47952 350509
rect 48188 350273 53882 350509
rect 54118 350273 59813 350509
rect 60049 350273 75952 350509
rect 76188 350273 81882 350509
rect 82118 350273 87813 350509
rect 88049 350273 103952 350509
rect 104188 350273 109882 350509
rect 110118 350273 115813 350509
rect 116049 350273 131952 350509
rect 132188 350273 137882 350509
rect 138118 350273 143813 350509
rect 144049 350273 159952 350509
rect 160188 350273 165882 350509
rect 166118 350273 171813 350509
rect 172049 350273 187952 350509
rect 188188 350273 193882 350509
rect 194118 350273 199813 350509
rect 200049 350273 215952 350509
rect 216188 350273 221882 350509
rect 222118 350273 227813 350509
rect 228049 350273 243952 350509
rect 244188 350273 249882 350509
rect 250118 350273 255813 350509
rect 256049 350273 271952 350509
rect 272188 350273 277882 350509
rect 278118 350273 283813 350509
rect 284049 350273 299952 350509
rect 300188 350273 305882 350509
rect 306118 350273 311813 350509
rect 312049 350273 327952 350509
rect 328188 350273 333882 350509
rect 334118 350273 339813 350509
rect 340049 350273 355952 350509
rect 356188 350273 361882 350509
rect 362118 350273 367813 350509
rect 368049 350273 383952 350509
rect 384188 350273 389882 350509
rect 390118 350273 395813 350509
rect 396049 350273 411952 350509
rect 412188 350273 417882 350509
rect 418118 350273 423813 350509
rect 424049 350273 439952 350509
rect 440188 350273 445882 350509
rect 446118 350273 451813 350509
rect 452049 350273 467952 350509
rect 468188 350273 473882 350509
rect 474118 350273 479813 350509
rect 480049 350273 495952 350509
rect 496188 350273 501882 350509
rect 502118 350273 507813 350509
rect 508049 350273 523952 350509
rect 524188 350273 529882 350509
rect 530118 350273 535813 350509
rect 536049 350273 551952 350509
rect 552188 350273 557882 350509
rect 558118 350273 563813 350509
rect 564049 350273 573526 350509
rect 573762 350273 573846 350509
rect 574082 350273 585342 350509
rect 585578 350273 585662 350509
rect 585898 350273 592650 350509
rect -8726 350241 592650 350273
rect -8726 347454 592650 347486
rect -8726 347218 -2934 347454
rect -2698 347218 -2614 347454
rect -2378 347218 22916 347454
rect 23152 347218 28847 347454
rect 29083 347218 50916 347454
rect 51152 347218 56847 347454
rect 57083 347218 78916 347454
rect 79152 347218 84847 347454
rect 85083 347218 106916 347454
rect 107152 347218 112847 347454
rect 113083 347218 134916 347454
rect 135152 347218 140847 347454
rect 141083 347218 162916 347454
rect 163152 347218 168847 347454
rect 169083 347218 190916 347454
rect 191152 347218 196847 347454
rect 197083 347218 218916 347454
rect 219152 347218 224847 347454
rect 225083 347218 246916 347454
rect 247152 347218 252847 347454
rect 253083 347218 274916 347454
rect 275152 347218 280847 347454
rect 281083 347218 302916 347454
rect 303152 347218 308847 347454
rect 309083 347218 330916 347454
rect 331152 347218 336847 347454
rect 337083 347218 358916 347454
rect 359152 347218 364847 347454
rect 365083 347218 386916 347454
rect 387152 347218 392847 347454
rect 393083 347218 414916 347454
rect 415152 347218 420847 347454
rect 421083 347218 442916 347454
rect 443152 347218 448847 347454
rect 449083 347218 470916 347454
rect 471152 347218 476847 347454
rect 477083 347218 498916 347454
rect 499152 347218 504847 347454
rect 505083 347218 526916 347454
rect 527152 347218 532847 347454
rect 533083 347218 554916 347454
rect 555152 347218 560847 347454
rect 561083 347218 586302 347454
rect 586538 347218 586622 347454
rect 586858 347218 592650 347454
rect -8726 347134 592650 347218
rect -8726 346898 -2934 347134
rect -2698 346898 -2614 347134
rect -2378 346898 22916 347134
rect 23152 346898 28847 347134
rect 29083 346898 50916 347134
rect 51152 346898 56847 347134
rect 57083 346898 78916 347134
rect 79152 346898 84847 347134
rect 85083 346898 106916 347134
rect 107152 346898 112847 347134
rect 113083 346898 134916 347134
rect 135152 346898 140847 347134
rect 141083 346898 162916 347134
rect 163152 346898 168847 347134
rect 169083 346898 190916 347134
rect 191152 346898 196847 347134
rect 197083 346898 218916 347134
rect 219152 346898 224847 347134
rect 225083 346898 246916 347134
rect 247152 346898 252847 347134
rect 253083 346898 274916 347134
rect 275152 346898 280847 347134
rect 281083 346898 302916 347134
rect 303152 346898 308847 347134
rect 309083 346898 330916 347134
rect 331152 346898 336847 347134
rect 337083 346898 358916 347134
rect 359152 346898 364847 347134
rect 365083 346898 386916 347134
rect 387152 346898 392847 347134
rect 393083 346898 414916 347134
rect 415152 346898 420847 347134
rect 421083 346898 442916 347134
rect 443152 346898 448847 347134
rect 449083 346898 470916 347134
rect 471152 346898 476847 347134
rect 477083 346898 498916 347134
rect 499152 346898 504847 347134
rect 505083 346898 526916 347134
rect 527152 346898 532847 347134
rect 533083 346898 554916 347134
rect 555152 346898 560847 347134
rect 561083 346898 586302 347134
rect 586538 346898 586622 347134
rect 586858 346898 592650 347134
rect -8726 346866 592650 346898
rect -8726 323829 592650 323861
rect -8726 323593 -1974 323829
rect -1738 323593 -1654 323829
rect -1418 323593 19951 323829
rect 20187 323593 25882 323829
rect 26118 323593 31812 323829
rect 32048 323593 47951 323829
rect 48187 323593 53882 323829
rect 54118 323593 59812 323829
rect 60048 323593 75951 323829
rect 76187 323593 81882 323829
rect 82118 323593 87812 323829
rect 88048 323593 103951 323829
rect 104187 323593 109882 323829
rect 110118 323593 115812 323829
rect 116048 323593 131951 323829
rect 132187 323593 137882 323829
rect 138118 323593 143812 323829
rect 144048 323593 159951 323829
rect 160187 323593 165882 323829
rect 166118 323593 171812 323829
rect 172048 323593 187951 323829
rect 188187 323593 193882 323829
rect 194118 323593 199812 323829
rect 200048 323593 215951 323829
rect 216187 323593 221882 323829
rect 222118 323593 227812 323829
rect 228048 323593 243951 323829
rect 244187 323593 249882 323829
rect 250118 323593 255812 323829
rect 256048 323593 271951 323829
rect 272187 323593 277882 323829
rect 278118 323593 283812 323829
rect 284048 323593 299951 323829
rect 300187 323593 305882 323829
rect 306118 323593 311812 323829
rect 312048 323593 327951 323829
rect 328187 323593 333882 323829
rect 334118 323593 339812 323829
rect 340048 323593 355951 323829
rect 356187 323593 361882 323829
rect 362118 323593 367812 323829
rect 368048 323593 383951 323829
rect 384187 323593 389882 323829
rect 390118 323593 395812 323829
rect 396048 323593 411951 323829
rect 412187 323593 417882 323829
rect 418118 323593 423812 323829
rect 424048 323593 439951 323829
rect 440187 323593 445882 323829
rect 446118 323593 451812 323829
rect 452048 323593 467951 323829
rect 468187 323593 473882 323829
rect 474118 323593 479812 323829
rect 480048 323593 495951 323829
rect 496187 323593 501882 323829
rect 502118 323593 507812 323829
rect 508048 323593 523951 323829
rect 524187 323593 529882 323829
rect 530118 323593 535812 323829
rect 536048 323593 551951 323829
rect 552187 323593 557882 323829
rect 558118 323593 563812 323829
rect 564048 323593 573526 323829
rect 573762 323593 573846 323829
rect 574082 323593 585342 323829
rect 585578 323593 585662 323829
rect 585898 323593 592650 323829
rect -8726 323509 592650 323593
rect -8726 323273 -1974 323509
rect -1738 323273 -1654 323509
rect -1418 323273 19951 323509
rect 20187 323273 25882 323509
rect 26118 323273 31812 323509
rect 32048 323273 47951 323509
rect 48187 323273 53882 323509
rect 54118 323273 59812 323509
rect 60048 323273 75951 323509
rect 76187 323273 81882 323509
rect 82118 323273 87812 323509
rect 88048 323273 103951 323509
rect 104187 323273 109882 323509
rect 110118 323273 115812 323509
rect 116048 323273 131951 323509
rect 132187 323273 137882 323509
rect 138118 323273 143812 323509
rect 144048 323273 159951 323509
rect 160187 323273 165882 323509
rect 166118 323273 171812 323509
rect 172048 323273 187951 323509
rect 188187 323273 193882 323509
rect 194118 323273 199812 323509
rect 200048 323273 215951 323509
rect 216187 323273 221882 323509
rect 222118 323273 227812 323509
rect 228048 323273 243951 323509
rect 244187 323273 249882 323509
rect 250118 323273 255812 323509
rect 256048 323273 271951 323509
rect 272187 323273 277882 323509
rect 278118 323273 283812 323509
rect 284048 323273 299951 323509
rect 300187 323273 305882 323509
rect 306118 323273 311812 323509
rect 312048 323273 327951 323509
rect 328187 323273 333882 323509
rect 334118 323273 339812 323509
rect 340048 323273 355951 323509
rect 356187 323273 361882 323509
rect 362118 323273 367812 323509
rect 368048 323273 383951 323509
rect 384187 323273 389882 323509
rect 390118 323273 395812 323509
rect 396048 323273 411951 323509
rect 412187 323273 417882 323509
rect 418118 323273 423812 323509
rect 424048 323273 439951 323509
rect 440187 323273 445882 323509
rect 446118 323273 451812 323509
rect 452048 323273 467951 323509
rect 468187 323273 473882 323509
rect 474118 323273 479812 323509
rect 480048 323273 495951 323509
rect 496187 323273 501882 323509
rect 502118 323273 507812 323509
rect 508048 323273 523951 323509
rect 524187 323273 529882 323509
rect 530118 323273 535812 323509
rect 536048 323273 551951 323509
rect 552187 323273 557882 323509
rect 558118 323273 563812 323509
rect 564048 323273 573526 323509
rect 573762 323273 573846 323509
rect 574082 323273 585342 323509
rect 585578 323273 585662 323509
rect 585898 323273 592650 323509
rect -8726 323241 592650 323273
rect -8726 320454 592650 320486
rect -8726 320218 -2934 320454
rect -2698 320218 -2614 320454
rect -2378 320218 22917 320454
rect 23153 320218 28848 320454
rect 29084 320218 50917 320454
rect 51153 320218 56848 320454
rect 57084 320218 78917 320454
rect 79153 320218 84848 320454
rect 85084 320218 106917 320454
rect 107153 320218 112848 320454
rect 113084 320218 134917 320454
rect 135153 320218 140848 320454
rect 141084 320218 162917 320454
rect 163153 320218 168848 320454
rect 169084 320218 190917 320454
rect 191153 320218 196848 320454
rect 197084 320218 218917 320454
rect 219153 320218 224848 320454
rect 225084 320218 246917 320454
rect 247153 320218 252848 320454
rect 253084 320218 274917 320454
rect 275153 320218 280848 320454
rect 281084 320218 302917 320454
rect 303153 320218 308848 320454
rect 309084 320218 330917 320454
rect 331153 320218 336848 320454
rect 337084 320218 358917 320454
rect 359153 320218 364848 320454
rect 365084 320218 386917 320454
rect 387153 320218 392848 320454
rect 393084 320218 414917 320454
rect 415153 320218 420848 320454
rect 421084 320218 442917 320454
rect 443153 320218 448848 320454
rect 449084 320218 470917 320454
rect 471153 320218 476848 320454
rect 477084 320218 498917 320454
rect 499153 320218 504848 320454
rect 505084 320218 526917 320454
rect 527153 320218 532848 320454
rect 533084 320218 554917 320454
rect 555153 320218 560848 320454
rect 561084 320218 586302 320454
rect 586538 320218 586622 320454
rect 586858 320218 592650 320454
rect -8726 320134 592650 320218
rect -8726 319898 -2934 320134
rect -2698 319898 -2614 320134
rect -2378 319898 22917 320134
rect 23153 319898 28848 320134
rect 29084 319898 50917 320134
rect 51153 319898 56848 320134
rect 57084 319898 78917 320134
rect 79153 319898 84848 320134
rect 85084 319898 106917 320134
rect 107153 319898 112848 320134
rect 113084 319898 134917 320134
rect 135153 319898 140848 320134
rect 141084 319898 162917 320134
rect 163153 319898 168848 320134
rect 169084 319898 190917 320134
rect 191153 319898 196848 320134
rect 197084 319898 218917 320134
rect 219153 319898 224848 320134
rect 225084 319898 246917 320134
rect 247153 319898 252848 320134
rect 253084 319898 274917 320134
rect 275153 319898 280848 320134
rect 281084 319898 302917 320134
rect 303153 319898 308848 320134
rect 309084 319898 330917 320134
rect 331153 319898 336848 320134
rect 337084 319898 358917 320134
rect 359153 319898 364848 320134
rect 365084 319898 386917 320134
rect 387153 319898 392848 320134
rect 393084 319898 414917 320134
rect 415153 319898 420848 320134
rect 421084 319898 442917 320134
rect 443153 319898 448848 320134
rect 449084 319898 470917 320134
rect 471153 319898 476848 320134
rect 477084 319898 498917 320134
rect 499153 319898 504848 320134
rect 505084 319898 526917 320134
rect 527153 319898 532848 320134
rect 533084 319898 554917 320134
rect 555153 319898 560848 320134
rect 561084 319898 586302 320134
rect 586538 319898 586622 320134
rect 586858 319898 592650 320134
rect -8726 319866 592650 319898
rect -8726 296829 592650 296861
rect -8726 296593 -1974 296829
rect -1738 296593 -1654 296829
rect -1418 296593 19952 296829
rect 20188 296593 25882 296829
rect 26118 296593 31813 296829
rect 32049 296593 47952 296829
rect 48188 296593 53882 296829
rect 54118 296593 59813 296829
rect 60049 296593 75952 296829
rect 76188 296593 81882 296829
rect 82118 296593 87813 296829
rect 88049 296593 103952 296829
rect 104188 296593 109882 296829
rect 110118 296593 115813 296829
rect 116049 296593 131952 296829
rect 132188 296593 137882 296829
rect 138118 296593 143813 296829
rect 144049 296593 159952 296829
rect 160188 296593 165882 296829
rect 166118 296593 171813 296829
rect 172049 296593 187952 296829
rect 188188 296593 193882 296829
rect 194118 296593 199813 296829
rect 200049 296593 215952 296829
rect 216188 296593 221882 296829
rect 222118 296593 227813 296829
rect 228049 296593 243952 296829
rect 244188 296593 249882 296829
rect 250118 296593 255813 296829
rect 256049 296593 271952 296829
rect 272188 296593 277882 296829
rect 278118 296593 283813 296829
rect 284049 296593 299952 296829
rect 300188 296593 305882 296829
rect 306118 296593 311813 296829
rect 312049 296593 327952 296829
rect 328188 296593 333882 296829
rect 334118 296593 339813 296829
rect 340049 296593 355952 296829
rect 356188 296593 361882 296829
rect 362118 296593 367813 296829
rect 368049 296593 383952 296829
rect 384188 296593 389882 296829
rect 390118 296593 395813 296829
rect 396049 296593 411952 296829
rect 412188 296593 417882 296829
rect 418118 296593 423813 296829
rect 424049 296593 439952 296829
rect 440188 296593 445882 296829
rect 446118 296593 451813 296829
rect 452049 296593 467952 296829
rect 468188 296593 473882 296829
rect 474118 296593 479813 296829
rect 480049 296593 495952 296829
rect 496188 296593 501882 296829
rect 502118 296593 507813 296829
rect 508049 296593 523952 296829
rect 524188 296593 529882 296829
rect 530118 296593 535813 296829
rect 536049 296593 551952 296829
rect 552188 296593 557882 296829
rect 558118 296593 563813 296829
rect 564049 296593 573526 296829
rect 573762 296593 573846 296829
rect 574082 296593 585342 296829
rect 585578 296593 585662 296829
rect 585898 296593 592650 296829
rect -8726 296509 592650 296593
rect -8726 296273 -1974 296509
rect -1738 296273 -1654 296509
rect -1418 296273 19952 296509
rect 20188 296273 25882 296509
rect 26118 296273 31813 296509
rect 32049 296273 47952 296509
rect 48188 296273 53882 296509
rect 54118 296273 59813 296509
rect 60049 296273 75952 296509
rect 76188 296273 81882 296509
rect 82118 296273 87813 296509
rect 88049 296273 103952 296509
rect 104188 296273 109882 296509
rect 110118 296273 115813 296509
rect 116049 296273 131952 296509
rect 132188 296273 137882 296509
rect 138118 296273 143813 296509
rect 144049 296273 159952 296509
rect 160188 296273 165882 296509
rect 166118 296273 171813 296509
rect 172049 296273 187952 296509
rect 188188 296273 193882 296509
rect 194118 296273 199813 296509
rect 200049 296273 215952 296509
rect 216188 296273 221882 296509
rect 222118 296273 227813 296509
rect 228049 296273 243952 296509
rect 244188 296273 249882 296509
rect 250118 296273 255813 296509
rect 256049 296273 271952 296509
rect 272188 296273 277882 296509
rect 278118 296273 283813 296509
rect 284049 296273 299952 296509
rect 300188 296273 305882 296509
rect 306118 296273 311813 296509
rect 312049 296273 327952 296509
rect 328188 296273 333882 296509
rect 334118 296273 339813 296509
rect 340049 296273 355952 296509
rect 356188 296273 361882 296509
rect 362118 296273 367813 296509
rect 368049 296273 383952 296509
rect 384188 296273 389882 296509
rect 390118 296273 395813 296509
rect 396049 296273 411952 296509
rect 412188 296273 417882 296509
rect 418118 296273 423813 296509
rect 424049 296273 439952 296509
rect 440188 296273 445882 296509
rect 446118 296273 451813 296509
rect 452049 296273 467952 296509
rect 468188 296273 473882 296509
rect 474118 296273 479813 296509
rect 480049 296273 495952 296509
rect 496188 296273 501882 296509
rect 502118 296273 507813 296509
rect 508049 296273 523952 296509
rect 524188 296273 529882 296509
rect 530118 296273 535813 296509
rect 536049 296273 551952 296509
rect 552188 296273 557882 296509
rect 558118 296273 563813 296509
rect 564049 296273 573526 296509
rect 573762 296273 573846 296509
rect 574082 296273 585342 296509
rect 585578 296273 585662 296509
rect 585898 296273 592650 296509
rect -8726 296241 592650 296273
rect -8726 293454 592650 293486
rect -8726 293218 -2934 293454
rect -2698 293218 -2614 293454
rect -2378 293218 22916 293454
rect 23152 293218 28847 293454
rect 29083 293218 50916 293454
rect 51152 293218 56847 293454
rect 57083 293218 78916 293454
rect 79152 293218 84847 293454
rect 85083 293218 106916 293454
rect 107152 293218 112847 293454
rect 113083 293218 134916 293454
rect 135152 293218 140847 293454
rect 141083 293218 162916 293454
rect 163152 293218 168847 293454
rect 169083 293218 190916 293454
rect 191152 293218 196847 293454
rect 197083 293218 218916 293454
rect 219152 293218 224847 293454
rect 225083 293218 246916 293454
rect 247152 293218 252847 293454
rect 253083 293218 274916 293454
rect 275152 293218 280847 293454
rect 281083 293218 302916 293454
rect 303152 293218 308847 293454
rect 309083 293218 330916 293454
rect 331152 293218 336847 293454
rect 337083 293218 358916 293454
rect 359152 293218 364847 293454
rect 365083 293218 386916 293454
rect 387152 293218 392847 293454
rect 393083 293218 414916 293454
rect 415152 293218 420847 293454
rect 421083 293218 442916 293454
rect 443152 293218 448847 293454
rect 449083 293218 470916 293454
rect 471152 293218 476847 293454
rect 477083 293218 498916 293454
rect 499152 293218 504847 293454
rect 505083 293218 526916 293454
rect 527152 293218 532847 293454
rect 533083 293218 554916 293454
rect 555152 293218 560847 293454
rect 561083 293218 586302 293454
rect 586538 293218 586622 293454
rect 586858 293218 592650 293454
rect -8726 293134 592650 293218
rect -8726 292898 -2934 293134
rect -2698 292898 -2614 293134
rect -2378 292898 22916 293134
rect 23152 292898 28847 293134
rect 29083 292898 50916 293134
rect 51152 292898 56847 293134
rect 57083 292898 78916 293134
rect 79152 292898 84847 293134
rect 85083 292898 106916 293134
rect 107152 292898 112847 293134
rect 113083 292898 134916 293134
rect 135152 292898 140847 293134
rect 141083 292898 162916 293134
rect 163152 292898 168847 293134
rect 169083 292898 190916 293134
rect 191152 292898 196847 293134
rect 197083 292898 218916 293134
rect 219152 292898 224847 293134
rect 225083 292898 246916 293134
rect 247152 292898 252847 293134
rect 253083 292898 274916 293134
rect 275152 292898 280847 293134
rect 281083 292898 302916 293134
rect 303152 292898 308847 293134
rect 309083 292898 330916 293134
rect 331152 292898 336847 293134
rect 337083 292898 358916 293134
rect 359152 292898 364847 293134
rect 365083 292898 386916 293134
rect 387152 292898 392847 293134
rect 393083 292898 414916 293134
rect 415152 292898 420847 293134
rect 421083 292898 442916 293134
rect 443152 292898 448847 293134
rect 449083 292898 470916 293134
rect 471152 292898 476847 293134
rect 477083 292898 498916 293134
rect 499152 292898 504847 293134
rect 505083 292898 526916 293134
rect 527152 292898 532847 293134
rect 533083 292898 554916 293134
rect 555152 292898 560847 293134
rect 561083 292898 586302 293134
rect 586538 292898 586622 293134
rect 586858 292898 592650 293134
rect -8726 292866 592650 292898
rect -8726 269829 592650 269861
rect -8726 269593 -1974 269829
rect -1738 269593 -1654 269829
rect -1418 269593 19951 269829
rect 20187 269593 25882 269829
rect 26118 269593 31812 269829
rect 32048 269593 47951 269829
rect 48187 269593 53882 269829
rect 54118 269593 59812 269829
rect 60048 269593 75951 269829
rect 76187 269593 81882 269829
rect 82118 269593 87812 269829
rect 88048 269593 103951 269829
rect 104187 269593 109882 269829
rect 110118 269593 115812 269829
rect 116048 269593 131951 269829
rect 132187 269593 137882 269829
rect 138118 269593 143812 269829
rect 144048 269593 159951 269829
rect 160187 269593 165882 269829
rect 166118 269593 171812 269829
rect 172048 269593 187951 269829
rect 188187 269593 193882 269829
rect 194118 269593 199812 269829
rect 200048 269593 215951 269829
rect 216187 269593 221882 269829
rect 222118 269593 227812 269829
rect 228048 269593 243951 269829
rect 244187 269593 249882 269829
rect 250118 269593 255812 269829
rect 256048 269593 271951 269829
rect 272187 269593 277882 269829
rect 278118 269593 283812 269829
rect 284048 269593 299951 269829
rect 300187 269593 305882 269829
rect 306118 269593 311812 269829
rect 312048 269593 327951 269829
rect 328187 269593 333882 269829
rect 334118 269593 339812 269829
rect 340048 269593 355951 269829
rect 356187 269593 361882 269829
rect 362118 269593 367812 269829
rect 368048 269593 383951 269829
rect 384187 269593 389882 269829
rect 390118 269593 395812 269829
rect 396048 269593 411951 269829
rect 412187 269593 417882 269829
rect 418118 269593 423812 269829
rect 424048 269593 439951 269829
rect 440187 269593 445882 269829
rect 446118 269593 451812 269829
rect 452048 269593 467951 269829
rect 468187 269593 473882 269829
rect 474118 269593 479812 269829
rect 480048 269593 495951 269829
rect 496187 269593 501882 269829
rect 502118 269593 507812 269829
rect 508048 269593 523951 269829
rect 524187 269593 529882 269829
rect 530118 269593 535812 269829
rect 536048 269593 551951 269829
rect 552187 269593 557882 269829
rect 558118 269593 563812 269829
rect 564048 269593 573526 269829
rect 573762 269593 573846 269829
rect 574082 269593 585342 269829
rect 585578 269593 585662 269829
rect 585898 269593 592650 269829
rect -8726 269509 592650 269593
rect -8726 269273 -1974 269509
rect -1738 269273 -1654 269509
rect -1418 269273 19951 269509
rect 20187 269273 25882 269509
rect 26118 269273 31812 269509
rect 32048 269273 47951 269509
rect 48187 269273 53882 269509
rect 54118 269273 59812 269509
rect 60048 269273 75951 269509
rect 76187 269273 81882 269509
rect 82118 269273 87812 269509
rect 88048 269273 103951 269509
rect 104187 269273 109882 269509
rect 110118 269273 115812 269509
rect 116048 269273 131951 269509
rect 132187 269273 137882 269509
rect 138118 269273 143812 269509
rect 144048 269273 159951 269509
rect 160187 269273 165882 269509
rect 166118 269273 171812 269509
rect 172048 269273 187951 269509
rect 188187 269273 193882 269509
rect 194118 269273 199812 269509
rect 200048 269273 215951 269509
rect 216187 269273 221882 269509
rect 222118 269273 227812 269509
rect 228048 269273 243951 269509
rect 244187 269273 249882 269509
rect 250118 269273 255812 269509
rect 256048 269273 271951 269509
rect 272187 269273 277882 269509
rect 278118 269273 283812 269509
rect 284048 269273 299951 269509
rect 300187 269273 305882 269509
rect 306118 269273 311812 269509
rect 312048 269273 327951 269509
rect 328187 269273 333882 269509
rect 334118 269273 339812 269509
rect 340048 269273 355951 269509
rect 356187 269273 361882 269509
rect 362118 269273 367812 269509
rect 368048 269273 383951 269509
rect 384187 269273 389882 269509
rect 390118 269273 395812 269509
rect 396048 269273 411951 269509
rect 412187 269273 417882 269509
rect 418118 269273 423812 269509
rect 424048 269273 439951 269509
rect 440187 269273 445882 269509
rect 446118 269273 451812 269509
rect 452048 269273 467951 269509
rect 468187 269273 473882 269509
rect 474118 269273 479812 269509
rect 480048 269273 495951 269509
rect 496187 269273 501882 269509
rect 502118 269273 507812 269509
rect 508048 269273 523951 269509
rect 524187 269273 529882 269509
rect 530118 269273 535812 269509
rect 536048 269273 551951 269509
rect 552187 269273 557882 269509
rect 558118 269273 563812 269509
rect 564048 269273 573526 269509
rect 573762 269273 573846 269509
rect 574082 269273 585342 269509
rect 585578 269273 585662 269509
rect 585898 269273 592650 269509
rect -8726 269241 592650 269273
rect -8726 266454 592650 266486
rect -8726 266218 -2934 266454
rect -2698 266218 -2614 266454
rect -2378 266218 22917 266454
rect 23153 266218 28848 266454
rect 29084 266218 50917 266454
rect 51153 266218 56848 266454
rect 57084 266218 78917 266454
rect 79153 266218 84848 266454
rect 85084 266218 106917 266454
rect 107153 266218 112848 266454
rect 113084 266218 134917 266454
rect 135153 266218 140848 266454
rect 141084 266218 162917 266454
rect 163153 266218 168848 266454
rect 169084 266218 190917 266454
rect 191153 266218 196848 266454
rect 197084 266218 218917 266454
rect 219153 266218 224848 266454
rect 225084 266218 246917 266454
rect 247153 266218 252848 266454
rect 253084 266218 274917 266454
rect 275153 266218 280848 266454
rect 281084 266218 302917 266454
rect 303153 266218 308848 266454
rect 309084 266218 330917 266454
rect 331153 266218 336848 266454
rect 337084 266218 358917 266454
rect 359153 266218 364848 266454
rect 365084 266218 386917 266454
rect 387153 266218 392848 266454
rect 393084 266218 414917 266454
rect 415153 266218 420848 266454
rect 421084 266218 442917 266454
rect 443153 266218 448848 266454
rect 449084 266218 470917 266454
rect 471153 266218 476848 266454
rect 477084 266218 498917 266454
rect 499153 266218 504848 266454
rect 505084 266218 526917 266454
rect 527153 266218 532848 266454
rect 533084 266218 554917 266454
rect 555153 266218 560848 266454
rect 561084 266218 586302 266454
rect 586538 266218 586622 266454
rect 586858 266218 592650 266454
rect -8726 266134 592650 266218
rect -8726 265898 -2934 266134
rect -2698 265898 -2614 266134
rect -2378 265898 22917 266134
rect 23153 265898 28848 266134
rect 29084 265898 50917 266134
rect 51153 265898 56848 266134
rect 57084 265898 78917 266134
rect 79153 265898 84848 266134
rect 85084 265898 106917 266134
rect 107153 265898 112848 266134
rect 113084 265898 134917 266134
rect 135153 265898 140848 266134
rect 141084 265898 162917 266134
rect 163153 265898 168848 266134
rect 169084 265898 190917 266134
rect 191153 265898 196848 266134
rect 197084 265898 218917 266134
rect 219153 265898 224848 266134
rect 225084 265898 246917 266134
rect 247153 265898 252848 266134
rect 253084 265898 274917 266134
rect 275153 265898 280848 266134
rect 281084 265898 302917 266134
rect 303153 265898 308848 266134
rect 309084 265898 330917 266134
rect 331153 265898 336848 266134
rect 337084 265898 358917 266134
rect 359153 265898 364848 266134
rect 365084 265898 386917 266134
rect 387153 265898 392848 266134
rect 393084 265898 414917 266134
rect 415153 265898 420848 266134
rect 421084 265898 442917 266134
rect 443153 265898 448848 266134
rect 449084 265898 470917 266134
rect 471153 265898 476848 266134
rect 477084 265898 498917 266134
rect 499153 265898 504848 266134
rect 505084 265898 526917 266134
rect 527153 265898 532848 266134
rect 533084 265898 554917 266134
rect 555153 265898 560848 266134
rect 561084 265898 586302 266134
rect 586538 265898 586622 266134
rect 586858 265898 592650 266134
rect -8726 265866 592650 265898
rect -8726 242829 592650 242861
rect -8726 242593 -1974 242829
rect -1738 242593 -1654 242829
rect -1418 242593 19952 242829
rect 20188 242593 25882 242829
rect 26118 242593 31813 242829
rect 32049 242593 47952 242829
rect 48188 242593 53882 242829
rect 54118 242593 59813 242829
rect 60049 242593 75952 242829
rect 76188 242593 81882 242829
rect 82118 242593 87813 242829
rect 88049 242593 103952 242829
rect 104188 242593 109882 242829
rect 110118 242593 115813 242829
rect 116049 242593 131952 242829
rect 132188 242593 137882 242829
rect 138118 242593 143813 242829
rect 144049 242593 159952 242829
rect 160188 242593 165882 242829
rect 166118 242593 171813 242829
rect 172049 242593 187952 242829
rect 188188 242593 193882 242829
rect 194118 242593 199813 242829
rect 200049 242593 215952 242829
rect 216188 242593 221882 242829
rect 222118 242593 227813 242829
rect 228049 242593 243952 242829
rect 244188 242593 249882 242829
rect 250118 242593 255813 242829
rect 256049 242593 271952 242829
rect 272188 242593 277882 242829
rect 278118 242593 283813 242829
rect 284049 242593 299952 242829
rect 300188 242593 305882 242829
rect 306118 242593 311813 242829
rect 312049 242593 327952 242829
rect 328188 242593 333882 242829
rect 334118 242593 339813 242829
rect 340049 242593 355952 242829
rect 356188 242593 361882 242829
rect 362118 242593 367813 242829
rect 368049 242593 383952 242829
rect 384188 242593 389882 242829
rect 390118 242593 395813 242829
rect 396049 242593 411952 242829
rect 412188 242593 417882 242829
rect 418118 242593 423813 242829
rect 424049 242593 439952 242829
rect 440188 242593 445882 242829
rect 446118 242593 451813 242829
rect 452049 242593 467952 242829
rect 468188 242593 473882 242829
rect 474118 242593 479813 242829
rect 480049 242593 495952 242829
rect 496188 242593 501882 242829
rect 502118 242593 507813 242829
rect 508049 242593 523952 242829
rect 524188 242593 529882 242829
rect 530118 242593 535813 242829
rect 536049 242593 551952 242829
rect 552188 242593 557882 242829
rect 558118 242593 563813 242829
rect 564049 242593 573526 242829
rect 573762 242593 573846 242829
rect 574082 242593 585342 242829
rect 585578 242593 585662 242829
rect 585898 242593 592650 242829
rect -8726 242509 592650 242593
rect -8726 242273 -1974 242509
rect -1738 242273 -1654 242509
rect -1418 242273 19952 242509
rect 20188 242273 25882 242509
rect 26118 242273 31813 242509
rect 32049 242273 47952 242509
rect 48188 242273 53882 242509
rect 54118 242273 59813 242509
rect 60049 242273 75952 242509
rect 76188 242273 81882 242509
rect 82118 242273 87813 242509
rect 88049 242273 103952 242509
rect 104188 242273 109882 242509
rect 110118 242273 115813 242509
rect 116049 242273 131952 242509
rect 132188 242273 137882 242509
rect 138118 242273 143813 242509
rect 144049 242273 159952 242509
rect 160188 242273 165882 242509
rect 166118 242273 171813 242509
rect 172049 242273 187952 242509
rect 188188 242273 193882 242509
rect 194118 242273 199813 242509
rect 200049 242273 215952 242509
rect 216188 242273 221882 242509
rect 222118 242273 227813 242509
rect 228049 242273 243952 242509
rect 244188 242273 249882 242509
rect 250118 242273 255813 242509
rect 256049 242273 271952 242509
rect 272188 242273 277882 242509
rect 278118 242273 283813 242509
rect 284049 242273 299952 242509
rect 300188 242273 305882 242509
rect 306118 242273 311813 242509
rect 312049 242273 327952 242509
rect 328188 242273 333882 242509
rect 334118 242273 339813 242509
rect 340049 242273 355952 242509
rect 356188 242273 361882 242509
rect 362118 242273 367813 242509
rect 368049 242273 383952 242509
rect 384188 242273 389882 242509
rect 390118 242273 395813 242509
rect 396049 242273 411952 242509
rect 412188 242273 417882 242509
rect 418118 242273 423813 242509
rect 424049 242273 439952 242509
rect 440188 242273 445882 242509
rect 446118 242273 451813 242509
rect 452049 242273 467952 242509
rect 468188 242273 473882 242509
rect 474118 242273 479813 242509
rect 480049 242273 495952 242509
rect 496188 242273 501882 242509
rect 502118 242273 507813 242509
rect 508049 242273 523952 242509
rect 524188 242273 529882 242509
rect 530118 242273 535813 242509
rect 536049 242273 551952 242509
rect 552188 242273 557882 242509
rect 558118 242273 563813 242509
rect 564049 242273 573526 242509
rect 573762 242273 573846 242509
rect 574082 242273 585342 242509
rect 585578 242273 585662 242509
rect 585898 242273 592650 242509
rect -8726 242241 592650 242273
rect -8726 239454 592650 239486
rect -8726 239218 -2934 239454
rect -2698 239218 -2614 239454
rect -2378 239218 22916 239454
rect 23152 239218 28847 239454
rect 29083 239218 50916 239454
rect 51152 239218 56847 239454
rect 57083 239218 78916 239454
rect 79152 239218 84847 239454
rect 85083 239218 106916 239454
rect 107152 239218 112847 239454
rect 113083 239218 134916 239454
rect 135152 239218 140847 239454
rect 141083 239218 162916 239454
rect 163152 239218 168847 239454
rect 169083 239218 190916 239454
rect 191152 239218 196847 239454
rect 197083 239218 218916 239454
rect 219152 239218 224847 239454
rect 225083 239218 246916 239454
rect 247152 239218 252847 239454
rect 253083 239218 274916 239454
rect 275152 239218 280847 239454
rect 281083 239218 302916 239454
rect 303152 239218 308847 239454
rect 309083 239218 330916 239454
rect 331152 239218 336847 239454
rect 337083 239218 358916 239454
rect 359152 239218 364847 239454
rect 365083 239218 386916 239454
rect 387152 239218 392847 239454
rect 393083 239218 414916 239454
rect 415152 239218 420847 239454
rect 421083 239218 442916 239454
rect 443152 239218 448847 239454
rect 449083 239218 470916 239454
rect 471152 239218 476847 239454
rect 477083 239218 498916 239454
rect 499152 239218 504847 239454
rect 505083 239218 526916 239454
rect 527152 239218 532847 239454
rect 533083 239218 554916 239454
rect 555152 239218 560847 239454
rect 561083 239218 586302 239454
rect 586538 239218 586622 239454
rect 586858 239218 592650 239454
rect -8726 239134 592650 239218
rect -8726 238898 -2934 239134
rect -2698 238898 -2614 239134
rect -2378 238898 22916 239134
rect 23152 238898 28847 239134
rect 29083 238898 50916 239134
rect 51152 238898 56847 239134
rect 57083 238898 78916 239134
rect 79152 238898 84847 239134
rect 85083 238898 106916 239134
rect 107152 238898 112847 239134
rect 113083 238898 134916 239134
rect 135152 238898 140847 239134
rect 141083 238898 162916 239134
rect 163152 238898 168847 239134
rect 169083 238898 190916 239134
rect 191152 238898 196847 239134
rect 197083 238898 218916 239134
rect 219152 238898 224847 239134
rect 225083 238898 246916 239134
rect 247152 238898 252847 239134
rect 253083 238898 274916 239134
rect 275152 238898 280847 239134
rect 281083 238898 302916 239134
rect 303152 238898 308847 239134
rect 309083 238898 330916 239134
rect 331152 238898 336847 239134
rect 337083 238898 358916 239134
rect 359152 238898 364847 239134
rect 365083 238898 386916 239134
rect 387152 238898 392847 239134
rect 393083 238898 414916 239134
rect 415152 238898 420847 239134
rect 421083 238898 442916 239134
rect 443152 238898 448847 239134
rect 449083 238898 470916 239134
rect 471152 238898 476847 239134
rect 477083 238898 498916 239134
rect 499152 238898 504847 239134
rect 505083 238898 526916 239134
rect 527152 238898 532847 239134
rect 533083 238898 554916 239134
rect 555152 238898 560847 239134
rect 561083 238898 586302 239134
rect 586538 238898 586622 239134
rect 586858 238898 592650 239134
rect -8726 238866 592650 238898
rect -8726 215829 592650 215861
rect -8726 215593 -1974 215829
rect -1738 215593 -1654 215829
rect -1418 215593 19951 215829
rect 20187 215593 25882 215829
rect 26118 215593 31812 215829
rect 32048 215593 47951 215829
rect 48187 215593 53882 215829
rect 54118 215593 59812 215829
rect 60048 215593 75951 215829
rect 76187 215593 81882 215829
rect 82118 215593 87812 215829
rect 88048 215593 103951 215829
rect 104187 215593 109882 215829
rect 110118 215593 115812 215829
rect 116048 215593 131951 215829
rect 132187 215593 137882 215829
rect 138118 215593 143812 215829
rect 144048 215593 159951 215829
rect 160187 215593 165882 215829
rect 166118 215593 171812 215829
rect 172048 215593 187951 215829
rect 188187 215593 193882 215829
rect 194118 215593 199812 215829
rect 200048 215593 215951 215829
rect 216187 215593 221882 215829
rect 222118 215593 227812 215829
rect 228048 215593 243951 215829
rect 244187 215593 249882 215829
rect 250118 215593 255812 215829
rect 256048 215593 271951 215829
rect 272187 215593 277882 215829
rect 278118 215593 283812 215829
rect 284048 215593 299951 215829
rect 300187 215593 305882 215829
rect 306118 215593 311812 215829
rect 312048 215593 327951 215829
rect 328187 215593 333882 215829
rect 334118 215593 339812 215829
rect 340048 215593 355951 215829
rect 356187 215593 361882 215829
rect 362118 215593 367812 215829
rect 368048 215593 383951 215829
rect 384187 215593 389882 215829
rect 390118 215593 395812 215829
rect 396048 215593 411951 215829
rect 412187 215593 417882 215829
rect 418118 215593 423812 215829
rect 424048 215593 439951 215829
rect 440187 215593 445882 215829
rect 446118 215593 451812 215829
rect 452048 215593 467951 215829
rect 468187 215593 473882 215829
rect 474118 215593 479812 215829
rect 480048 215593 495951 215829
rect 496187 215593 501882 215829
rect 502118 215593 507812 215829
rect 508048 215593 523951 215829
rect 524187 215593 529882 215829
rect 530118 215593 535812 215829
rect 536048 215593 551951 215829
rect 552187 215593 557882 215829
rect 558118 215593 563812 215829
rect 564048 215593 573526 215829
rect 573762 215593 573846 215829
rect 574082 215593 585342 215829
rect 585578 215593 585662 215829
rect 585898 215593 592650 215829
rect -8726 215509 592650 215593
rect -8726 215273 -1974 215509
rect -1738 215273 -1654 215509
rect -1418 215273 19951 215509
rect 20187 215273 25882 215509
rect 26118 215273 31812 215509
rect 32048 215273 47951 215509
rect 48187 215273 53882 215509
rect 54118 215273 59812 215509
rect 60048 215273 75951 215509
rect 76187 215273 81882 215509
rect 82118 215273 87812 215509
rect 88048 215273 103951 215509
rect 104187 215273 109882 215509
rect 110118 215273 115812 215509
rect 116048 215273 131951 215509
rect 132187 215273 137882 215509
rect 138118 215273 143812 215509
rect 144048 215273 159951 215509
rect 160187 215273 165882 215509
rect 166118 215273 171812 215509
rect 172048 215273 187951 215509
rect 188187 215273 193882 215509
rect 194118 215273 199812 215509
rect 200048 215273 215951 215509
rect 216187 215273 221882 215509
rect 222118 215273 227812 215509
rect 228048 215273 243951 215509
rect 244187 215273 249882 215509
rect 250118 215273 255812 215509
rect 256048 215273 271951 215509
rect 272187 215273 277882 215509
rect 278118 215273 283812 215509
rect 284048 215273 299951 215509
rect 300187 215273 305882 215509
rect 306118 215273 311812 215509
rect 312048 215273 327951 215509
rect 328187 215273 333882 215509
rect 334118 215273 339812 215509
rect 340048 215273 355951 215509
rect 356187 215273 361882 215509
rect 362118 215273 367812 215509
rect 368048 215273 383951 215509
rect 384187 215273 389882 215509
rect 390118 215273 395812 215509
rect 396048 215273 411951 215509
rect 412187 215273 417882 215509
rect 418118 215273 423812 215509
rect 424048 215273 439951 215509
rect 440187 215273 445882 215509
rect 446118 215273 451812 215509
rect 452048 215273 467951 215509
rect 468187 215273 473882 215509
rect 474118 215273 479812 215509
rect 480048 215273 495951 215509
rect 496187 215273 501882 215509
rect 502118 215273 507812 215509
rect 508048 215273 523951 215509
rect 524187 215273 529882 215509
rect 530118 215273 535812 215509
rect 536048 215273 551951 215509
rect 552187 215273 557882 215509
rect 558118 215273 563812 215509
rect 564048 215273 573526 215509
rect 573762 215273 573846 215509
rect 574082 215273 585342 215509
rect 585578 215273 585662 215509
rect 585898 215273 592650 215509
rect -8726 215241 592650 215273
rect -8726 212454 592650 212486
rect -8726 212218 -2934 212454
rect -2698 212218 -2614 212454
rect -2378 212218 22917 212454
rect 23153 212218 28848 212454
rect 29084 212218 50917 212454
rect 51153 212218 56848 212454
rect 57084 212218 78917 212454
rect 79153 212218 84848 212454
rect 85084 212218 106917 212454
rect 107153 212218 112848 212454
rect 113084 212218 134917 212454
rect 135153 212218 140848 212454
rect 141084 212218 162917 212454
rect 163153 212218 168848 212454
rect 169084 212218 190917 212454
rect 191153 212218 196848 212454
rect 197084 212218 218917 212454
rect 219153 212218 224848 212454
rect 225084 212218 246917 212454
rect 247153 212218 252848 212454
rect 253084 212218 274917 212454
rect 275153 212218 280848 212454
rect 281084 212218 302917 212454
rect 303153 212218 308848 212454
rect 309084 212218 330917 212454
rect 331153 212218 336848 212454
rect 337084 212218 358917 212454
rect 359153 212218 364848 212454
rect 365084 212218 386917 212454
rect 387153 212218 392848 212454
rect 393084 212218 414917 212454
rect 415153 212218 420848 212454
rect 421084 212218 442917 212454
rect 443153 212218 448848 212454
rect 449084 212218 470917 212454
rect 471153 212218 476848 212454
rect 477084 212218 498917 212454
rect 499153 212218 504848 212454
rect 505084 212218 526917 212454
rect 527153 212218 532848 212454
rect 533084 212218 554917 212454
rect 555153 212218 560848 212454
rect 561084 212218 586302 212454
rect 586538 212218 586622 212454
rect 586858 212218 592650 212454
rect -8726 212134 592650 212218
rect -8726 211898 -2934 212134
rect -2698 211898 -2614 212134
rect -2378 211898 22917 212134
rect 23153 211898 28848 212134
rect 29084 211898 50917 212134
rect 51153 211898 56848 212134
rect 57084 211898 78917 212134
rect 79153 211898 84848 212134
rect 85084 211898 106917 212134
rect 107153 211898 112848 212134
rect 113084 211898 134917 212134
rect 135153 211898 140848 212134
rect 141084 211898 162917 212134
rect 163153 211898 168848 212134
rect 169084 211898 190917 212134
rect 191153 211898 196848 212134
rect 197084 211898 218917 212134
rect 219153 211898 224848 212134
rect 225084 211898 246917 212134
rect 247153 211898 252848 212134
rect 253084 211898 274917 212134
rect 275153 211898 280848 212134
rect 281084 211898 302917 212134
rect 303153 211898 308848 212134
rect 309084 211898 330917 212134
rect 331153 211898 336848 212134
rect 337084 211898 358917 212134
rect 359153 211898 364848 212134
rect 365084 211898 386917 212134
rect 387153 211898 392848 212134
rect 393084 211898 414917 212134
rect 415153 211898 420848 212134
rect 421084 211898 442917 212134
rect 443153 211898 448848 212134
rect 449084 211898 470917 212134
rect 471153 211898 476848 212134
rect 477084 211898 498917 212134
rect 499153 211898 504848 212134
rect 505084 211898 526917 212134
rect 527153 211898 532848 212134
rect 533084 211898 554917 212134
rect 555153 211898 560848 212134
rect 561084 211898 586302 212134
rect 586538 211898 586622 212134
rect 586858 211898 592650 212134
rect -8726 211866 592650 211898
rect -8726 188829 592650 188861
rect -8726 188593 -1974 188829
rect -1738 188593 -1654 188829
rect -1418 188593 19952 188829
rect 20188 188593 25882 188829
rect 26118 188593 31813 188829
rect 32049 188593 47952 188829
rect 48188 188593 53882 188829
rect 54118 188593 59813 188829
rect 60049 188593 75952 188829
rect 76188 188593 81882 188829
rect 82118 188593 87813 188829
rect 88049 188593 103952 188829
rect 104188 188593 109882 188829
rect 110118 188593 115813 188829
rect 116049 188593 131952 188829
rect 132188 188593 137882 188829
rect 138118 188593 143813 188829
rect 144049 188593 159952 188829
rect 160188 188593 165882 188829
rect 166118 188593 171813 188829
rect 172049 188593 187952 188829
rect 188188 188593 193882 188829
rect 194118 188593 199813 188829
rect 200049 188593 215952 188829
rect 216188 188593 221882 188829
rect 222118 188593 227813 188829
rect 228049 188593 243952 188829
rect 244188 188593 249882 188829
rect 250118 188593 255813 188829
rect 256049 188593 271952 188829
rect 272188 188593 277882 188829
rect 278118 188593 283813 188829
rect 284049 188593 299952 188829
rect 300188 188593 305882 188829
rect 306118 188593 311813 188829
rect 312049 188593 327952 188829
rect 328188 188593 333882 188829
rect 334118 188593 339813 188829
rect 340049 188593 355952 188829
rect 356188 188593 361882 188829
rect 362118 188593 367813 188829
rect 368049 188593 383952 188829
rect 384188 188593 389882 188829
rect 390118 188593 395813 188829
rect 396049 188593 411952 188829
rect 412188 188593 417882 188829
rect 418118 188593 423813 188829
rect 424049 188593 439952 188829
rect 440188 188593 445882 188829
rect 446118 188593 451813 188829
rect 452049 188593 467952 188829
rect 468188 188593 473882 188829
rect 474118 188593 479813 188829
rect 480049 188593 495952 188829
rect 496188 188593 501882 188829
rect 502118 188593 507813 188829
rect 508049 188593 523952 188829
rect 524188 188593 529882 188829
rect 530118 188593 535813 188829
rect 536049 188593 551952 188829
rect 552188 188593 557882 188829
rect 558118 188593 563813 188829
rect 564049 188593 573526 188829
rect 573762 188593 573846 188829
rect 574082 188593 585342 188829
rect 585578 188593 585662 188829
rect 585898 188593 592650 188829
rect -8726 188509 592650 188593
rect -8726 188273 -1974 188509
rect -1738 188273 -1654 188509
rect -1418 188273 19952 188509
rect 20188 188273 25882 188509
rect 26118 188273 31813 188509
rect 32049 188273 47952 188509
rect 48188 188273 53882 188509
rect 54118 188273 59813 188509
rect 60049 188273 75952 188509
rect 76188 188273 81882 188509
rect 82118 188273 87813 188509
rect 88049 188273 103952 188509
rect 104188 188273 109882 188509
rect 110118 188273 115813 188509
rect 116049 188273 131952 188509
rect 132188 188273 137882 188509
rect 138118 188273 143813 188509
rect 144049 188273 159952 188509
rect 160188 188273 165882 188509
rect 166118 188273 171813 188509
rect 172049 188273 187952 188509
rect 188188 188273 193882 188509
rect 194118 188273 199813 188509
rect 200049 188273 215952 188509
rect 216188 188273 221882 188509
rect 222118 188273 227813 188509
rect 228049 188273 243952 188509
rect 244188 188273 249882 188509
rect 250118 188273 255813 188509
rect 256049 188273 271952 188509
rect 272188 188273 277882 188509
rect 278118 188273 283813 188509
rect 284049 188273 299952 188509
rect 300188 188273 305882 188509
rect 306118 188273 311813 188509
rect 312049 188273 327952 188509
rect 328188 188273 333882 188509
rect 334118 188273 339813 188509
rect 340049 188273 355952 188509
rect 356188 188273 361882 188509
rect 362118 188273 367813 188509
rect 368049 188273 383952 188509
rect 384188 188273 389882 188509
rect 390118 188273 395813 188509
rect 396049 188273 411952 188509
rect 412188 188273 417882 188509
rect 418118 188273 423813 188509
rect 424049 188273 439952 188509
rect 440188 188273 445882 188509
rect 446118 188273 451813 188509
rect 452049 188273 467952 188509
rect 468188 188273 473882 188509
rect 474118 188273 479813 188509
rect 480049 188273 495952 188509
rect 496188 188273 501882 188509
rect 502118 188273 507813 188509
rect 508049 188273 523952 188509
rect 524188 188273 529882 188509
rect 530118 188273 535813 188509
rect 536049 188273 551952 188509
rect 552188 188273 557882 188509
rect 558118 188273 563813 188509
rect 564049 188273 573526 188509
rect 573762 188273 573846 188509
rect 574082 188273 585342 188509
rect 585578 188273 585662 188509
rect 585898 188273 592650 188509
rect -8726 188241 592650 188273
rect -8726 185454 592650 185486
rect -8726 185218 -2934 185454
rect -2698 185218 -2614 185454
rect -2378 185218 22916 185454
rect 23152 185218 28847 185454
rect 29083 185218 50916 185454
rect 51152 185218 56847 185454
rect 57083 185218 78916 185454
rect 79152 185218 84847 185454
rect 85083 185218 106916 185454
rect 107152 185218 112847 185454
rect 113083 185218 134916 185454
rect 135152 185218 140847 185454
rect 141083 185218 162916 185454
rect 163152 185218 168847 185454
rect 169083 185218 190916 185454
rect 191152 185218 196847 185454
rect 197083 185218 218916 185454
rect 219152 185218 224847 185454
rect 225083 185218 246916 185454
rect 247152 185218 252847 185454
rect 253083 185218 274916 185454
rect 275152 185218 280847 185454
rect 281083 185218 302916 185454
rect 303152 185218 308847 185454
rect 309083 185218 330916 185454
rect 331152 185218 336847 185454
rect 337083 185218 358916 185454
rect 359152 185218 364847 185454
rect 365083 185218 386916 185454
rect 387152 185218 392847 185454
rect 393083 185218 414916 185454
rect 415152 185218 420847 185454
rect 421083 185218 442916 185454
rect 443152 185218 448847 185454
rect 449083 185218 470916 185454
rect 471152 185218 476847 185454
rect 477083 185218 498916 185454
rect 499152 185218 504847 185454
rect 505083 185218 526916 185454
rect 527152 185218 532847 185454
rect 533083 185218 554916 185454
rect 555152 185218 560847 185454
rect 561083 185218 586302 185454
rect 586538 185218 586622 185454
rect 586858 185218 592650 185454
rect -8726 185134 592650 185218
rect -8726 184898 -2934 185134
rect -2698 184898 -2614 185134
rect -2378 184898 22916 185134
rect 23152 184898 28847 185134
rect 29083 184898 50916 185134
rect 51152 184898 56847 185134
rect 57083 184898 78916 185134
rect 79152 184898 84847 185134
rect 85083 184898 106916 185134
rect 107152 184898 112847 185134
rect 113083 184898 134916 185134
rect 135152 184898 140847 185134
rect 141083 184898 162916 185134
rect 163152 184898 168847 185134
rect 169083 184898 190916 185134
rect 191152 184898 196847 185134
rect 197083 184898 218916 185134
rect 219152 184898 224847 185134
rect 225083 184898 246916 185134
rect 247152 184898 252847 185134
rect 253083 184898 274916 185134
rect 275152 184898 280847 185134
rect 281083 184898 302916 185134
rect 303152 184898 308847 185134
rect 309083 184898 330916 185134
rect 331152 184898 336847 185134
rect 337083 184898 358916 185134
rect 359152 184898 364847 185134
rect 365083 184898 386916 185134
rect 387152 184898 392847 185134
rect 393083 184898 414916 185134
rect 415152 184898 420847 185134
rect 421083 184898 442916 185134
rect 443152 184898 448847 185134
rect 449083 184898 470916 185134
rect 471152 184898 476847 185134
rect 477083 184898 498916 185134
rect 499152 184898 504847 185134
rect 505083 184898 526916 185134
rect 527152 184898 532847 185134
rect 533083 184898 554916 185134
rect 555152 184898 560847 185134
rect 561083 184898 586302 185134
rect 586538 184898 586622 185134
rect 586858 184898 592650 185134
rect -8726 184866 592650 184898
rect -8726 161829 592650 161861
rect -8726 161593 -1974 161829
rect -1738 161593 -1654 161829
rect -1418 161593 19951 161829
rect 20187 161593 25882 161829
rect 26118 161593 31812 161829
rect 32048 161593 47951 161829
rect 48187 161593 53882 161829
rect 54118 161593 59812 161829
rect 60048 161593 75951 161829
rect 76187 161593 81882 161829
rect 82118 161593 87812 161829
rect 88048 161593 103951 161829
rect 104187 161593 109882 161829
rect 110118 161593 115812 161829
rect 116048 161593 131951 161829
rect 132187 161593 137882 161829
rect 138118 161593 143812 161829
rect 144048 161593 159951 161829
rect 160187 161593 165882 161829
rect 166118 161593 171812 161829
rect 172048 161593 187951 161829
rect 188187 161593 193882 161829
rect 194118 161593 199812 161829
rect 200048 161593 215951 161829
rect 216187 161593 221882 161829
rect 222118 161593 227812 161829
rect 228048 161593 243951 161829
rect 244187 161593 249882 161829
rect 250118 161593 255812 161829
rect 256048 161593 271951 161829
rect 272187 161593 277882 161829
rect 278118 161593 283812 161829
rect 284048 161593 299951 161829
rect 300187 161593 305882 161829
rect 306118 161593 311812 161829
rect 312048 161593 327951 161829
rect 328187 161593 333882 161829
rect 334118 161593 339812 161829
rect 340048 161593 355951 161829
rect 356187 161593 361882 161829
rect 362118 161593 367812 161829
rect 368048 161593 383951 161829
rect 384187 161593 389882 161829
rect 390118 161593 395812 161829
rect 396048 161593 411951 161829
rect 412187 161593 417882 161829
rect 418118 161593 423812 161829
rect 424048 161593 439951 161829
rect 440187 161593 445882 161829
rect 446118 161593 451812 161829
rect 452048 161593 467951 161829
rect 468187 161593 473882 161829
rect 474118 161593 479812 161829
rect 480048 161593 495951 161829
rect 496187 161593 501882 161829
rect 502118 161593 507812 161829
rect 508048 161593 523951 161829
rect 524187 161593 529882 161829
rect 530118 161593 535812 161829
rect 536048 161593 551951 161829
rect 552187 161593 557882 161829
rect 558118 161593 563812 161829
rect 564048 161593 573526 161829
rect 573762 161593 573846 161829
rect 574082 161593 585342 161829
rect 585578 161593 585662 161829
rect 585898 161593 592650 161829
rect -8726 161509 592650 161593
rect -8726 161273 -1974 161509
rect -1738 161273 -1654 161509
rect -1418 161273 19951 161509
rect 20187 161273 25882 161509
rect 26118 161273 31812 161509
rect 32048 161273 47951 161509
rect 48187 161273 53882 161509
rect 54118 161273 59812 161509
rect 60048 161273 75951 161509
rect 76187 161273 81882 161509
rect 82118 161273 87812 161509
rect 88048 161273 103951 161509
rect 104187 161273 109882 161509
rect 110118 161273 115812 161509
rect 116048 161273 131951 161509
rect 132187 161273 137882 161509
rect 138118 161273 143812 161509
rect 144048 161273 159951 161509
rect 160187 161273 165882 161509
rect 166118 161273 171812 161509
rect 172048 161273 187951 161509
rect 188187 161273 193882 161509
rect 194118 161273 199812 161509
rect 200048 161273 215951 161509
rect 216187 161273 221882 161509
rect 222118 161273 227812 161509
rect 228048 161273 243951 161509
rect 244187 161273 249882 161509
rect 250118 161273 255812 161509
rect 256048 161273 271951 161509
rect 272187 161273 277882 161509
rect 278118 161273 283812 161509
rect 284048 161273 299951 161509
rect 300187 161273 305882 161509
rect 306118 161273 311812 161509
rect 312048 161273 327951 161509
rect 328187 161273 333882 161509
rect 334118 161273 339812 161509
rect 340048 161273 355951 161509
rect 356187 161273 361882 161509
rect 362118 161273 367812 161509
rect 368048 161273 383951 161509
rect 384187 161273 389882 161509
rect 390118 161273 395812 161509
rect 396048 161273 411951 161509
rect 412187 161273 417882 161509
rect 418118 161273 423812 161509
rect 424048 161273 439951 161509
rect 440187 161273 445882 161509
rect 446118 161273 451812 161509
rect 452048 161273 467951 161509
rect 468187 161273 473882 161509
rect 474118 161273 479812 161509
rect 480048 161273 495951 161509
rect 496187 161273 501882 161509
rect 502118 161273 507812 161509
rect 508048 161273 523951 161509
rect 524187 161273 529882 161509
rect 530118 161273 535812 161509
rect 536048 161273 551951 161509
rect 552187 161273 557882 161509
rect 558118 161273 563812 161509
rect 564048 161273 573526 161509
rect 573762 161273 573846 161509
rect 574082 161273 585342 161509
rect 585578 161273 585662 161509
rect 585898 161273 592650 161509
rect -8726 161241 592650 161273
rect -8726 158454 592650 158486
rect -8726 158218 -2934 158454
rect -2698 158218 -2614 158454
rect -2378 158218 22917 158454
rect 23153 158218 28848 158454
rect 29084 158218 50917 158454
rect 51153 158218 56848 158454
rect 57084 158218 78917 158454
rect 79153 158218 84848 158454
rect 85084 158218 106917 158454
rect 107153 158218 112848 158454
rect 113084 158218 134917 158454
rect 135153 158218 140848 158454
rect 141084 158218 162917 158454
rect 163153 158218 168848 158454
rect 169084 158218 190917 158454
rect 191153 158218 196848 158454
rect 197084 158218 218917 158454
rect 219153 158218 224848 158454
rect 225084 158218 246917 158454
rect 247153 158218 252848 158454
rect 253084 158218 274917 158454
rect 275153 158218 280848 158454
rect 281084 158218 302917 158454
rect 303153 158218 308848 158454
rect 309084 158218 330917 158454
rect 331153 158218 336848 158454
rect 337084 158218 358917 158454
rect 359153 158218 364848 158454
rect 365084 158218 386917 158454
rect 387153 158218 392848 158454
rect 393084 158218 414917 158454
rect 415153 158218 420848 158454
rect 421084 158218 442917 158454
rect 443153 158218 448848 158454
rect 449084 158218 470917 158454
rect 471153 158218 476848 158454
rect 477084 158218 498917 158454
rect 499153 158218 504848 158454
rect 505084 158218 526917 158454
rect 527153 158218 532848 158454
rect 533084 158218 554917 158454
rect 555153 158218 560848 158454
rect 561084 158218 586302 158454
rect 586538 158218 586622 158454
rect 586858 158218 592650 158454
rect -8726 158134 592650 158218
rect -8726 157898 -2934 158134
rect -2698 157898 -2614 158134
rect -2378 157898 22917 158134
rect 23153 157898 28848 158134
rect 29084 157898 50917 158134
rect 51153 157898 56848 158134
rect 57084 157898 78917 158134
rect 79153 157898 84848 158134
rect 85084 157898 106917 158134
rect 107153 157898 112848 158134
rect 113084 157898 134917 158134
rect 135153 157898 140848 158134
rect 141084 157898 162917 158134
rect 163153 157898 168848 158134
rect 169084 157898 190917 158134
rect 191153 157898 196848 158134
rect 197084 157898 218917 158134
rect 219153 157898 224848 158134
rect 225084 157898 246917 158134
rect 247153 157898 252848 158134
rect 253084 157898 274917 158134
rect 275153 157898 280848 158134
rect 281084 157898 302917 158134
rect 303153 157898 308848 158134
rect 309084 157898 330917 158134
rect 331153 157898 336848 158134
rect 337084 157898 358917 158134
rect 359153 157898 364848 158134
rect 365084 157898 386917 158134
rect 387153 157898 392848 158134
rect 393084 157898 414917 158134
rect 415153 157898 420848 158134
rect 421084 157898 442917 158134
rect 443153 157898 448848 158134
rect 449084 157898 470917 158134
rect 471153 157898 476848 158134
rect 477084 157898 498917 158134
rect 499153 157898 504848 158134
rect 505084 157898 526917 158134
rect 527153 157898 532848 158134
rect 533084 157898 554917 158134
rect 555153 157898 560848 158134
rect 561084 157898 586302 158134
rect 586538 157898 586622 158134
rect 586858 157898 592650 158134
rect -8726 157866 592650 157898
rect -8726 134829 592650 134861
rect -8726 134593 -1974 134829
rect -1738 134593 -1654 134829
rect -1418 134593 19952 134829
rect 20188 134593 25882 134829
rect 26118 134593 31813 134829
rect 32049 134593 47952 134829
rect 48188 134593 53882 134829
rect 54118 134593 59813 134829
rect 60049 134593 75952 134829
rect 76188 134593 81882 134829
rect 82118 134593 87813 134829
rect 88049 134593 103952 134829
rect 104188 134593 109882 134829
rect 110118 134593 115813 134829
rect 116049 134593 131952 134829
rect 132188 134593 137882 134829
rect 138118 134593 143813 134829
rect 144049 134593 159952 134829
rect 160188 134593 165882 134829
rect 166118 134593 171813 134829
rect 172049 134593 187952 134829
rect 188188 134593 193882 134829
rect 194118 134593 199813 134829
rect 200049 134593 215952 134829
rect 216188 134593 221882 134829
rect 222118 134593 227813 134829
rect 228049 134593 243952 134829
rect 244188 134593 249882 134829
rect 250118 134593 255813 134829
rect 256049 134593 271952 134829
rect 272188 134593 277882 134829
rect 278118 134593 283813 134829
rect 284049 134593 299952 134829
rect 300188 134593 305882 134829
rect 306118 134593 311813 134829
rect 312049 134593 327952 134829
rect 328188 134593 333882 134829
rect 334118 134593 339813 134829
rect 340049 134593 355952 134829
rect 356188 134593 361882 134829
rect 362118 134593 367813 134829
rect 368049 134593 383952 134829
rect 384188 134593 389882 134829
rect 390118 134593 395813 134829
rect 396049 134593 411952 134829
rect 412188 134593 417882 134829
rect 418118 134593 423813 134829
rect 424049 134593 439952 134829
rect 440188 134593 445882 134829
rect 446118 134593 451813 134829
rect 452049 134593 467952 134829
rect 468188 134593 473882 134829
rect 474118 134593 479813 134829
rect 480049 134593 495952 134829
rect 496188 134593 501882 134829
rect 502118 134593 507813 134829
rect 508049 134593 523952 134829
rect 524188 134593 529882 134829
rect 530118 134593 535813 134829
rect 536049 134593 551952 134829
rect 552188 134593 557882 134829
rect 558118 134593 563813 134829
rect 564049 134593 573526 134829
rect 573762 134593 573846 134829
rect 574082 134593 585342 134829
rect 585578 134593 585662 134829
rect 585898 134593 592650 134829
rect -8726 134509 592650 134593
rect -8726 134273 -1974 134509
rect -1738 134273 -1654 134509
rect -1418 134273 19952 134509
rect 20188 134273 25882 134509
rect 26118 134273 31813 134509
rect 32049 134273 47952 134509
rect 48188 134273 53882 134509
rect 54118 134273 59813 134509
rect 60049 134273 75952 134509
rect 76188 134273 81882 134509
rect 82118 134273 87813 134509
rect 88049 134273 103952 134509
rect 104188 134273 109882 134509
rect 110118 134273 115813 134509
rect 116049 134273 131952 134509
rect 132188 134273 137882 134509
rect 138118 134273 143813 134509
rect 144049 134273 159952 134509
rect 160188 134273 165882 134509
rect 166118 134273 171813 134509
rect 172049 134273 187952 134509
rect 188188 134273 193882 134509
rect 194118 134273 199813 134509
rect 200049 134273 215952 134509
rect 216188 134273 221882 134509
rect 222118 134273 227813 134509
rect 228049 134273 243952 134509
rect 244188 134273 249882 134509
rect 250118 134273 255813 134509
rect 256049 134273 271952 134509
rect 272188 134273 277882 134509
rect 278118 134273 283813 134509
rect 284049 134273 299952 134509
rect 300188 134273 305882 134509
rect 306118 134273 311813 134509
rect 312049 134273 327952 134509
rect 328188 134273 333882 134509
rect 334118 134273 339813 134509
rect 340049 134273 355952 134509
rect 356188 134273 361882 134509
rect 362118 134273 367813 134509
rect 368049 134273 383952 134509
rect 384188 134273 389882 134509
rect 390118 134273 395813 134509
rect 396049 134273 411952 134509
rect 412188 134273 417882 134509
rect 418118 134273 423813 134509
rect 424049 134273 439952 134509
rect 440188 134273 445882 134509
rect 446118 134273 451813 134509
rect 452049 134273 467952 134509
rect 468188 134273 473882 134509
rect 474118 134273 479813 134509
rect 480049 134273 495952 134509
rect 496188 134273 501882 134509
rect 502118 134273 507813 134509
rect 508049 134273 523952 134509
rect 524188 134273 529882 134509
rect 530118 134273 535813 134509
rect 536049 134273 551952 134509
rect 552188 134273 557882 134509
rect 558118 134273 563813 134509
rect 564049 134273 573526 134509
rect 573762 134273 573846 134509
rect 574082 134273 585342 134509
rect 585578 134273 585662 134509
rect 585898 134273 592650 134509
rect -8726 134241 592650 134273
rect -8726 131454 592650 131486
rect -8726 131218 -2934 131454
rect -2698 131218 -2614 131454
rect -2378 131218 22916 131454
rect 23152 131218 28847 131454
rect 29083 131218 50916 131454
rect 51152 131218 56847 131454
rect 57083 131218 78916 131454
rect 79152 131218 84847 131454
rect 85083 131218 106916 131454
rect 107152 131218 112847 131454
rect 113083 131218 134916 131454
rect 135152 131218 140847 131454
rect 141083 131218 162916 131454
rect 163152 131218 168847 131454
rect 169083 131218 190916 131454
rect 191152 131218 196847 131454
rect 197083 131218 218916 131454
rect 219152 131218 224847 131454
rect 225083 131218 246916 131454
rect 247152 131218 252847 131454
rect 253083 131218 274916 131454
rect 275152 131218 280847 131454
rect 281083 131218 302916 131454
rect 303152 131218 308847 131454
rect 309083 131218 330916 131454
rect 331152 131218 336847 131454
rect 337083 131218 358916 131454
rect 359152 131218 364847 131454
rect 365083 131218 386916 131454
rect 387152 131218 392847 131454
rect 393083 131218 414916 131454
rect 415152 131218 420847 131454
rect 421083 131218 442916 131454
rect 443152 131218 448847 131454
rect 449083 131218 470916 131454
rect 471152 131218 476847 131454
rect 477083 131218 498916 131454
rect 499152 131218 504847 131454
rect 505083 131218 526916 131454
rect 527152 131218 532847 131454
rect 533083 131218 554916 131454
rect 555152 131218 560847 131454
rect 561083 131218 586302 131454
rect 586538 131218 586622 131454
rect 586858 131218 592650 131454
rect -8726 131134 592650 131218
rect -8726 130898 -2934 131134
rect -2698 130898 -2614 131134
rect -2378 130898 22916 131134
rect 23152 130898 28847 131134
rect 29083 130898 50916 131134
rect 51152 130898 56847 131134
rect 57083 130898 78916 131134
rect 79152 130898 84847 131134
rect 85083 130898 106916 131134
rect 107152 130898 112847 131134
rect 113083 130898 134916 131134
rect 135152 130898 140847 131134
rect 141083 130898 162916 131134
rect 163152 130898 168847 131134
rect 169083 130898 190916 131134
rect 191152 130898 196847 131134
rect 197083 130898 218916 131134
rect 219152 130898 224847 131134
rect 225083 130898 246916 131134
rect 247152 130898 252847 131134
rect 253083 130898 274916 131134
rect 275152 130898 280847 131134
rect 281083 130898 302916 131134
rect 303152 130898 308847 131134
rect 309083 130898 330916 131134
rect 331152 130898 336847 131134
rect 337083 130898 358916 131134
rect 359152 130898 364847 131134
rect 365083 130898 386916 131134
rect 387152 130898 392847 131134
rect 393083 130898 414916 131134
rect 415152 130898 420847 131134
rect 421083 130898 442916 131134
rect 443152 130898 448847 131134
rect 449083 130898 470916 131134
rect 471152 130898 476847 131134
rect 477083 130898 498916 131134
rect 499152 130898 504847 131134
rect 505083 130898 526916 131134
rect 527152 130898 532847 131134
rect 533083 130898 554916 131134
rect 555152 130898 560847 131134
rect 561083 130898 586302 131134
rect 586538 130898 586622 131134
rect 586858 130898 592650 131134
rect -8726 130866 592650 130898
rect -8726 107829 592650 107861
rect -8726 107593 -1974 107829
rect -1738 107593 -1654 107829
rect -1418 107593 19951 107829
rect 20187 107593 25882 107829
rect 26118 107593 31812 107829
rect 32048 107593 47951 107829
rect 48187 107593 53882 107829
rect 54118 107593 59812 107829
rect 60048 107593 75951 107829
rect 76187 107593 81882 107829
rect 82118 107593 87812 107829
rect 88048 107593 103951 107829
rect 104187 107593 109882 107829
rect 110118 107593 115812 107829
rect 116048 107593 131210 107829
rect 131446 107593 135658 107829
rect 135894 107593 140106 107829
rect 140342 107593 144554 107829
rect 144790 107593 159951 107829
rect 160187 107593 165882 107829
rect 166118 107593 171812 107829
rect 172048 107593 187951 107829
rect 188187 107593 193882 107829
rect 194118 107593 199812 107829
rect 200048 107593 215210 107829
rect 215446 107593 219658 107829
rect 219894 107593 224106 107829
rect 224342 107593 228554 107829
rect 228790 107593 243951 107829
rect 244187 107593 249882 107829
rect 250118 107593 255812 107829
rect 256048 107593 271951 107829
rect 272187 107593 277882 107829
rect 278118 107593 283812 107829
rect 284048 107593 299951 107829
rect 300187 107593 305882 107829
rect 306118 107593 311812 107829
rect 312048 107593 327951 107829
rect 328187 107593 333882 107829
rect 334118 107593 339812 107829
rect 340048 107593 355951 107829
rect 356187 107593 361882 107829
rect 362118 107593 367812 107829
rect 368048 107593 383951 107829
rect 384187 107593 389882 107829
rect 390118 107593 395812 107829
rect 396048 107593 411951 107829
rect 412187 107593 417882 107829
rect 418118 107593 423812 107829
rect 424048 107593 439951 107829
rect 440187 107593 445882 107829
rect 446118 107593 451812 107829
rect 452048 107593 467951 107829
rect 468187 107593 473882 107829
rect 474118 107593 479812 107829
rect 480048 107593 495951 107829
rect 496187 107593 501882 107829
rect 502118 107593 507812 107829
rect 508048 107593 523951 107829
rect 524187 107593 529882 107829
rect 530118 107593 535812 107829
rect 536048 107593 551951 107829
rect 552187 107593 557882 107829
rect 558118 107593 563812 107829
rect 564048 107593 573526 107829
rect 573762 107593 573846 107829
rect 574082 107593 585342 107829
rect 585578 107593 585662 107829
rect 585898 107593 592650 107829
rect -8726 107509 592650 107593
rect -8726 107273 -1974 107509
rect -1738 107273 -1654 107509
rect -1418 107273 19951 107509
rect 20187 107273 25882 107509
rect 26118 107273 31812 107509
rect 32048 107273 47951 107509
rect 48187 107273 53882 107509
rect 54118 107273 59812 107509
rect 60048 107273 75951 107509
rect 76187 107273 81882 107509
rect 82118 107273 87812 107509
rect 88048 107273 103951 107509
rect 104187 107273 109882 107509
rect 110118 107273 115812 107509
rect 116048 107273 131210 107509
rect 131446 107273 135658 107509
rect 135894 107273 140106 107509
rect 140342 107273 144554 107509
rect 144790 107273 159951 107509
rect 160187 107273 165882 107509
rect 166118 107273 171812 107509
rect 172048 107273 187951 107509
rect 188187 107273 193882 107509
rect 194118 107273 199812 107509
rect 200048 107273 215210 107509
rect 215446 107273 219658 107509
rect 219894 107273 224106 107509
rect 224342 107273 228554 107509
rect 228790 107273 243951 107509
rect 244187 107273 249882 107509
rect 250118 107273 255812 107509
rect 256048 107273 271951 107509
rect 272187 107273 277882 107509
rect 278118 107273 283812 107509
rect 284048 107273 299951 107509
rect 300187 107273 305882 107509
rect 306118 107273 311812 107509
rect 312048 107273 327951 107509
rect 328187 107273 333882 107509
rect 334118 107273 339812 107509
rect 340048 107273 355951 107509
rect 356187 107273 361882 107509
rect 362118 107273 367812 107509
rect 368048 107273 383951 107509
rect 384187 107273 389882 107509
rect 390118 107273 395812 107509
rect 396048 107273 411951 107509
rect 412187 107273 417882 107509
rect 418118 107273 423812 107509
rect 424048 107273 439951 107509
rect 440187 107273 445882 107509
rect 446118 107273 451812 107509
rect 452048 107273 467951 107509
rect 468187 107273 473882 107509
rect 474118 107273 479812 107509
rect 480048 107273 495951 107509
rect 496187 107273 501882 107509
rect 502118 107273 507812 107509
rect 508048 107273 523951 107509
rect 524187 107273 529882 107509
rect 530118 107273 535812 107509
rect 536048 107273 551951 107509
rect 552187 107273 557882 107509
rect 558118 107273 563812 107509
rect 564048 107273 573526 107509
rect 573762 107273 573846 107509
rect 574082 107273 585342 107509
rect 585578 107273 585662 107509
rect 585898 107273 592650 107509
rect -8726 107241 592650 107273
rect -8726 104454 592650 104486
rect -8726 104218 -2934 104454
rect -2698 104218 -2614 104454
rect -2378 104218 22917 104454
rect 23153 104218 28848 104454
rect 29084 104218 50917 104454
rect 51153 104218 56848 104454
rect 57084 104218 78917 104454
rect 79153 104218 84848 104454
rect 85084 104218 106917 104454
rect 107153 104218 112848 104454
rect 113084 104218 133434 104454
rect 133670 104218 137882 104454
rect 138118 104218 142330 104454
rect 142566 104218 162917 104454
rect 163153 104218 168848 104454
rect 169084 104218 190917 104454
rect 191153 104218 196848 104454
rect 197084 104218 217434 104454
rect 217670 104218 221882 104454
rect 222118 104218 226330 104454
rect 226566 104218 246917 104454
rect 247153 104218 252848 104454
rect 253084 104218 274917 104454
rect 275153 104218 280848 104454
rect 281084 104218 302917 104454
rect 303153 104218 308848 104454
rect 309084 104218 330917 104454
rect 331153 104218 336848 104454
rect 337084 104218 358917 104454
rect 359153 104218 364848 104454
rect 365084 104218 386917 104454
rect 387153 104218 392848 104454
rect 393084 104218 414917 104454
rect 415153 104218 420848 104454
rect 421084 104218 442917 104454
rect 443153 104218 448848 104454
rect 449084 104218 470917 104454
rect 471153 104218 476848 104454
rect 477084 104218 498917 104454
rect 499153 104218 504848 104454
rect 505084 104218 526917 104454
rect 527153 104218 532848 104454
rect 533084 104218 554917 104454
rect 555153 104218 560848 104454
rect 561084 104218 586302 104454
rect 586538 104218 586622 104454
rect 586858 104218 592650 104454
rect -8726 104134 592650 104218
rect -8726 103898 -2934 104134
rect -2698 103898 -2614 104134
rect -2378 103898 22917 104134
rect 23153 103898 28848 104134
rect 29084 103898 50917 104134
rect 51153 103898 56848 104134
rect 57084 103898 78917 104134
rect 79153 103898 84848 104134
rect 85084 103898 106917 104134
rect 107153 103898 112848 104134
rect 113084 103898 133434 104134
rect 133670 103898 137882 104134
rect 138118 103898 142330 104134
rect 142566 103898 162917 104134
rect 163153 103898 168848 104134
rect 169084 103898 190917 104134
rect 191153 103898 196848 104134
rect 197084 103898 217434 104134
rect 217670 103898 221882 104134
rect 222118 103898 226330 104134
rect 226566 103898 246917 104134
rect 247153 103898 252848 104134
rect 253084 103898 274917 104134
rect 275153 103898 280848 104134
rect 281084 103898 302917 104134
rect 303153 103898 308848 104134
rect 309084 103898 330917 104134
rect 331153 103898 336848 104134
rect 337084 103898 358917 104134
rect 359153 103898 364848 104134
rect 365084 103898 386917 104134
rect 387153 103898 392848 104134
rect 393084 103898 414917 104134
rect 415153 103898 420848 104134
rect 421084 103898 442917 104134
rect 443153 103898 448848 104134
rect 449084 103898 470917 104134
rect 471153 103898 476848 104134
rect 477084 103898 498917 104134
rect 499153 103898 504848 104134
rect 505084 103898 526917 104134
rect 527153 103898 532848 104134
rect 533084 103898 554917 104134
rect 555153 103898 560848 104134
rect 561084 103898 586302 104134
rect 586538 103898 586622 104134
rect 586858 103898 592650 104134
rect -8726 103866 592650 103898
rect -8726 80829 592650 80861
rect -8726 80593 -1974 80829
rect -1738 80593 -1654 80829
rect -1418 80593 19952 80829
rect 20188 80593 25882 80829
rect 26118 80593 31813 80829
rect 32049 80593 47952 80829
rect 48188 80593 53882 80829
rect 54118 80593 59813 80829
rect 60049 80593 75952 80829
rect 76188 80593 81882 80829
rect 82118 80593 87813 80829
rect 88049 80593 103952 80829
rect 104188 80593 109882 80829
rect 110118 80593 115813 80829
rect 116049 80593 131952 80829
rect 132188 80593 137882 80829
rect 138118 80593 143813 80829
rect 144049 80593 159952 80829
rect 160188 80593 165882 80829
rect 166118 80593 171813 80829
rect 172049 80593 187952 80829
rect 188188 80593 193882 80829
rect 194118 80593 199813 80829
rect 200049 80593 215952 80829
rect 216188 80593 221882 80829
rect 222118 80593 227813 80829
rect 228049 80593 243952 80829
rect 244188 80593 249882 80829
rect 250118 80593 255813 80829
rect 256049 80593 271952 80829
rect 272188 80593 277882 80829
rect 278118 80593 283813 80829
rect 284049 80593 299952 80829
rect 300188 80593 305882 80829
rect 306118 80593 311813 80829
rect 312049 80593 327952 80829
rect 328188 80593 333882 80829
rect 334118 80593 339813 80829
rect 340049 80593 355952 80829
rect 356188 80593 361882 80829
rect 362118 80593 367813 80829
rect 368049 80593 383952 80829
rect 384188 80593 389882 80829
rect 390118 80593 395813 80829
rect 396049 80593 411952 80829
rect 412188 80593 417882 80829
rect 418118 80593 423813 80829
rect 424049 80593 439952 80829
rect 440188 80593 445882 80829
rect 446118 80593 451813 80829
rect 452049 80593 467952 80829
rect 468188 80593 473882 80829
rect 474118 80593 479813 80829
rect 480049 80593 495952 80829
rect 496188 80593 501882 80829
rect 502118 80593 507813 80829
rect 508049 80593 523952 80829
rect 524188 80593 529882 80829
rect 530118 80593 535813 80829
rect 536049 80593 551952 80829
rect 552188 80593 557882 80829
rect 558118 80593 563813 80829
rect 564049 80593 573526 80829
rect 573762 80593 573846 80829
rect 574082 80593 585342 80829
rect 585578 80593 585662 80829
rect 585898 80593 592650 80829
rect -8726 80509 592650 80593
rect -8726 80273 -1974 80509
rect -1738 80273 -1654 80509
rect -1418 80273 19952 80509
rect 20188 80273 25882 80509
rect 26118 80273 31813 80509
rect 32049 80273 47952 80509
rect 48188 80273 53882 80509
rect 54118 80273 59813 80509
rect 60049 80273 75952 80509
rect 76188 80273 81882 80509
rect 82118 80273 87813 80509
rect 88049 80273 103952 80509
rect 104188 80273 109882 80509
rect 110118 80273 115813 80509
rect 116049 80273 131952 80509
rect 132188 80273 137882 80509
rect 138118 80273 143813 80509
rect 144049 80273 159952 80509
rect 160188 80273 165882 80509
rect 166118 80273 171813 80509
rect 172049 80273 187952 80509
rect 188188 80273 193882 80509
rect 194118 80273 199813 80509
rect 200049 80273 215952 80509
rect 216188 80273 221882 80509
rect 222118 80273 227813 80509
rect 228049 80273 243952 80509
rect 244188 80273 249882 80509
rect 250118 80273 255813 80509
rect 256049 80273 271952 80509
rect 272188 80273 277882 80509
rect 278118 80273 283813 80509
rect 284049 80273 299952 80509
rect 300188 80273 305882 80509
rect 306118 80273 311813 80509
rect 312049 80273 327952 80509
rect 328188 80273 333882 80509
rect 334118 80273 339813 80509
rect 340049 80273 355952 80509
rect 356188 80273 361882 80509
rect 362118 80273 367813 80509
rect 368049 80273 383952 80509
rect 384188 80273 389882 80509
rect 390118 80273 395813 80509
rect 396049 80273 411952 80509
rect 412188 80273 417882 80509
rect 418118 80273 423813 80509
rect 424049 80273 439952 80509
rect 440188 80273 445882 80509
rect 446118 80273 451813 80509
rect 452049 80273 467952 80509
rect 468188 80273 473882 80509
rect 474118 80273 479813 80509
rect 480049 80273 495952 80509
rect 496188 80273 501882 80509
rect 502118 80273 507813 80509
rect 508049 80273 523952 80509
rect 524188 80273 529882 80509
rect 530118 80273 535813 80509
rect 536049 80273 551952 80509
rect 552188 80273 557882 80509
rect 558118 80273 563813 80509
rect 564049 80273 573526 80509
rect 573762 80273 573846 80509
rect 574082 80273 585342 80509
rect 585578 80273 585662 80509
rect 585898 80273 592650 80509
rect -8726 80241 592650 80273
rect -8726 77454 592650 77486
rect -8726 77218 -2934 77454
rect -2698 77218 -2614 77454
rect -2378 77218 22916 77454
rect 23152 77218 28847 77454
rect 29083 77218 50916 77454
rect 51152 77218 56847 77454
rect 57083 77218 78916 77454
rect 79152 77218 84847 77454
rect 85083 77218 106916 77454
rect 107152 77218 112847 77454
rect 113083 77218 134916 77454
rect 135152 77218 140847 77454
rect 141083 77218 162916 77454
rect 163152 77218 168847 77454
rect 169083 77218 190916 77454
rect 191152 77218 196847 77454
rect 197083 77218 218916 77454
rect 219152 77218 224847 77454
rect 225083 77218 246916 77454
rect 247152 77218 252847 77454
rect 253083 77218 274916 77454
rect 275152 77218 280847 77454
rect 281083 77218 302916 77454
rect 303152 77218 308847 77454
rect 309083 77218 330916 77454
rect 331152 77218 336847 77454
rect 337083 77218 358916 77454
rect 359152 77218 364847 77454
rect 365083 77218 386916 77454
rect 387152 77218 392847 77454
rect 393083 77218 414916 77454
rect 415152 77218 420847 77454
rect 421083 77218 442916 77454
rect 443152 77218 448847 77454
rect 449083 77218 470916 77454
rect 471152 77218 476847 77454
rect 477083 77218 498916 77454
rect 499152 77218 504847 77454
rect 505083 77218 526916 77454
rect 527152 77218 532847 77454
rect 533083 77218 554916 77454
rect 555152 77218 560847 77454
rect 561083 77218 586302 77454
rect 586538 77218 586622 77454
rect 586858 77218 592650 77454
rect -8726 77134 592650 77218
rect -8726 76898 -2934 77134
rect -2698 76898 -2614 77134
rect -2378 76898 22916 77134
rect 23152 76898 28847 77134
rect 29083 76898 50916 77134
rect 51152 76898 56847 77134
rect 57083 76898 78916 77134
rect 79152 76898 84847 77134
rect 85083 76898 106916 77134
rect 107152 76898 112847 77134
rect 113083 76898 134916 77134
rect 135152 76898 140847 77134
rect 141083 76898 162916 77134
rect 163152 76898 168847 77134
rect 169083 76898 190916 77134
rect 191152 76898 196847 77134
rect 197083 76898 218916 77134
rect 219152 76898 224847 77134
rect 225083 76898 246916 77134
rect 247152 76898 252847 77134
rect 253083 76898 274916 77134
rect 275152 76898 280847 77134
rect 281083 76898 302916 77134
rect 303152 76898 308847 77134
rect 309083 76898 330916 77134
rect 331152 76898 336847 77134
rect 337083 76898 358916 77134
rect 359152 76898 364847 77134
rect 365083 76898 386916 77134
rect 387152 76898 392847 77134
rect 393083 76898 414916 77134
rect 415152 76898 420847 77134
rect 421083 76898 442916 77134
rect 443152 76898 448847 77134
rect 449083 76898 470916 77134
rect 471152 76898 476847 77134
rect 477083 76898 498916 77134
rect 499152 76898 504847 77134
rect 505083 76898 526916 77134
rect 527152 76898 532847 77134
rect 533083 76898 554916 77134
rect 555152 76898 560847 77134
rect 561083 76898 586302 77134
rect 586538 76898 586622 77134
rect 586858 76898 592650 77134
rect -8726 76866 592650 76898
rect -8726 53829 592650 53861
rect -8726 53593 -1974 53829
rect -1738 53593 -1654 53829
rect -1418 53593 19951 53829
rect 20187 53593 25882 53829
rect 26118 53593 31812 53829
rect 32048 53593 47951 53829
rect 48187 53593 53882 53829
rect 54118 53593 59812 53829
rect 60048 53593 75951 53829
rect 76187 53593 81882 53829
rect 82118 53593 87812 53829
rect 88048 53593 103951 53829
rect 104187 53593 109882 53829
rect 110118 53593 115812 53829
rect 116048 53593 131951 53829
rect 132187 53593 137882 53829
rect 138118 53593 143812 53829
rect 144048 53593 159951 53829
rect 160187 53593 165882 53829
rect 166118 53593 171812 53829
rect 172048 53593 187951 53829
rect 188187 53593 193882 53829
rect 194118 53593 199812 53829
rect 200048 53593 215951 53829
rect 216187 53593 221882 53829
rect 222118 53593 227812 53829
rect 228048 53593 243951 53829
rect 244187 53593 249882 53829
rect 250118 53593 255812 53829
rect 256048 53593 271951 53829
rect 272187 53593 277882 53829
rect 278118 53593 283812 53829
rect 284048 53593 299951 53829
rect 300187 53593 305882 53829
rect 306118 53593 311812 53829
rect 312048 53593 327951 53829
rect 328187 53593 333882 53829
rect 334118 53593 339812 53829
rect 340048 53593 355951 53829
rect 356187 53593 361882 53829
rect 362118 53593 367812 53829
rect 368048 53593 383951 53829
rect 384187 53593 389882 53829
rect 390118 53593 395812 53829
rect 396048 53593 411951 53829
rect 412187 53593 417882 53829
rect 418118 53593 423812 53829
rect 424048 53593 439951 53829
rect 440187 53593 445882 53829
rect 446118 53593 451812 53829
rect 452048 53593 467951 53829
rect 468187 53593 473882 53829
rect 474118 53593 479812 53829
rect 480048 53593 495951 53829
rect 496187 53593 501882 53829
rect 502118 53593 507812 53829
rect 508048 53593 523951 53829
rect 524187 53593 529882 53829
rect 530118 53593 535812 53829
rect 536048 53593 551951 53829
rect 552187 53593 557882 53829
rect 558118 53593 563812 53829
rect 564048 53593 573526 53829
rect 573762 53593 573846 53829
rect 574082 53593 585342 53829
rect 585578 53593 585662 53829
rect 585898 53593 592650 53829
rect -8726 53509 592650 53593
rect -8726 53273 -1974 53509
rect -1738 53273 -1654 53509
rect -1418 53273 19951 53509
rect 20187 53273 25882 53509
rect 26118 53273 31812 53509
rect 32048 53273 47951 53509
rect 48187 53273 53882 53509
rect 54118 53273 59812 53509
rect 60048 53273 75951 53509
rect 76187 53273 81882 53509
rect 82118 53273 87812 53509
rect 88048 53273 103951 53509
rect 104187 53273 109882 53509
rect 110118 53273 115812 53509
rect 116048 53273 131951 53509
rect 132187 53273 137882 53509
rect 138118 53273 143812 53509
rect 144048 53273 159951 53509
rect 160187 53273 165882 53509
rect 166118 53273 171812 53509
rect 172048 53273 187951 53509
rect 188187 53273 193882 53509
rect 194118 53273 199812 53509
rect 200048 53273 215951 53509
rect 216187 53273 221882 53509
rect 222118 53273 227812 53509
rect 228048 53273 243951 53509
rect 244187 53273 249882 53509
rect 250118 53273 255812 53509
rect 256048 53273 271951 53509
rect 272187 53273 277882 53509
rect 278118 53273 283812 53509
rect 284048 53273 299951 53509
rect 300187 53273 305882 53509
rect 306118 53273 311812 53509
rect 312048 53273 327951 53509
rect 328187 53273 333882 53509
rect 334118 53273 339812 53509
rect 340048 53273 355951 53509
rect 356187 53273 361882 53509
rect 362118 53273 367812 53509
rect 368048 53273 383951 53509
rect 384187 53273 389882 53509
rect 390118 53273 395812 53509
rect 396048 53273 411951 53509
rect 412187 53273 417882 53509
rect 418118 53273 423812 53509
rect 424048 53273 439951 53509
rect 440187 53273 445882 53509
rect 446118 53273 451812 53509
rect 452048 53273 467951 53509
rect 468187 53273 473882 53509
rect 474118 53273 479812 53509
rect 480048 53273 495951 53509
rect 496187 53273 501882 53509
rect 502118 53273 507812 53509
rect 508048 53273 523951 53509
rect 524187 53273 529882 53509
rect 530118 53273 535812 53509
rect 536048 53273 551951 53509
rect 552187 53273 557882 53509
rect 558118 53273 563812 53509
rect 564048 53273 573526 53509
rect 573762 53273 573846 53509
rect 574082 53273 585342 53509
rect 585578 53273 585662 53509
rect 585898 53273 592650 53509
rect -8726 53241 592650 53273
rect -8726 50454 592650 50486
rect -8726 50218 -2934 50454
rect -2698 50218 -2614 50454
rect -2378 50218 22917 50454
rect 23153 50218 28848 50454
rect 29084 50218 50917 50454
rect 51153 50218 56848 50454
rect 57084 50218 78917 50454
rect 79153 50218 84848 50454
rect 85084 50218 106917 50454
rect 107153 50218 112848 50454
rect 113084 50218 134917 50454
rect 135153 50218 140848 50454
rect 141084 50218 162917 50454
rect 163153 50218 168848 50454
rect 169084 50218 190917 50454
rect 191153 50218 196848 50454
rect 197084 50218 218917 50454
rect 219153 50218 224848 50454
rect 225084 50218 246917 50454
rect 247153 50218 252848 50454
rect 253084 50218 274917 50454
rect 275153 50218 280848 50454
rect 281084 50218 302917 50454
rect 303153 50218 308848 50454
rect 309084 50218 330917 50454
rect 331153 50218 336848 50454
rect 337084 50218 358917 50454
rect 359153 50218 364848 50454
rect 365084 50218 386917 50454
rect 387153 50218 392848 50454
rect 393084 50218 414917 50454
rect 415153 50218 420848 50454
rect 421084 50218 442917 50454
rect 443153 50218 448848 50454
rect 449084 50218 470917 50454
rect 471153 50218 476848 50454
rect 477084 50218 498917 50454
rect 499153 50218 504848 50454
rect 505084 50218 526917 50454
rect 527153 50218 532848 50454
rect 533084 50218 554917 50454
rect 555153 50218 560848 50454
rect 561084 50218 586302 50454
rect 586538 50218 586622 50454
rect 586858 50218 592650 50454
rect -8726 50134 592650 50218
rect -8726 49898 -2934 50134
rect -2698 49898 -2614 50134
rect -2378 49898 22917 50134
rect 23153 49898 28848 50134
rect 29084 49898 50917 50134
rect 51153 49898 56848 50134
rect 57084 49898 78917 50134
rect 79153 49898 84848 50134
rect 85084 49898 106917 50134
rect 107153 49898 112848 50134
rect 113084 49898 134917 50134
rect 135153 49898 140848 50134
rect 141084 49898 162917 50134
rect 163153 49898 168848 50134
rect 169084 49898 190917 50134
rect 191153 49898 196848 50134
rect 197084 49898 218917 50134
rect 219153 49898 224848 50134
rect 225084 49898 246917 50134
rect 247153 49898 252848 50134
rect 253084 49898 274917 50134
rect 275153 49898 280848 50134
rect 281084 49898 302917 50134
rect 303153 49898 308848 50134
rect 309084 49898 330917 50134
rect 331153 49898 336848 50134
rect 337084 49898 358917 50134
rect 359153 49898 364848 50134
rect 365084 49898 386917 50134
rect 387153 49898 392848 50134
rect 393084 49898 414917 50134
rect 415153 49898 420848 50134
rect 421084 49898 442917 50134
rect 443153 49898 448848 50134
rect 449084 49898 470917 50134
rect 471153 49898 476848 50134
rect 477084 49898 498917 50134
rect 499153 49898 504848 50134
rect 505084 49898 526917 50134
rect 527153 49898 532848 50134
rect 533084 49898 554917 50134
rect 555153 49898 560848 50134
rect 561084 49898 586302 50134
rect 586538 49898 586622 50134
rect 586858 49898 592650 50134
rect -8726 49866 592650 49898
rect -8726 26829 592650 26861
rect -8726 26593 -1974 26829
rect -1738 26593 -1654 26829
rect -1418 26593 22460 26829
rect 22696 26593 33408 26829
rect 33644 26593 44356 26829
rect 44592 26593 55304 26829
rect 55540 26593 75952 26829
rect 76188 26593 81882 26829
rect 82118 26593 87813 26829
rect 88049 26593 103952 26829
rect 104188 26593 109882 26829
rect 110118 26593 115813 26829
rect 116049 26593 131952 26829
rect 132188 26593 137882 26829
rect 138118 26593 143813 26829
rect 144049 26593 159952 26829
rect 160188 26593 165882 26829
rect 166118 26593 171813 26829
rect 172049 26593 187952 26829
rect 188188 26593 193882 26829
rect 194118 26593 199813 26829
rect 200049 26593 215952 26829
rect 216188 26593 221882 26829
rect 222118 26593 227813 26829
rect 228049 26593 243952 26829
rect 244188 26593 249882 26829
rect 250118 26593 255813 26829
rect 256049 26593 271952 26829
rect 272188 26593 277882 26829
rect 278118 26593 283813 26829
rect 284049 26593 299952 26829
rect 300188 26593 305882 26829
rect 306118 26593 311813 26829
rect 312049 26593 327952 26829
rect 328188 26593 333882 26829
rect 334118 26593 339813 26829
rect 340049 26593 355952 26829
rect 356188 26593 361882 26829
rect 362118 26593 367813 26829
rect 368049 26593 383952 26829
rect 384188 26593 389882 26829
rect 390118 26593 395813 26829
rect 396049 26593 411952 26829
rect 412188 26593 417882 26829
rect 418118 26593 423813 26829
rect 424049 26593 439952 26829
rect 440188 26593 445882 26829
rect 446118 26593 451813 26829
rect 452049 26593 467952 26829
rect 468188 26593 473882 26829
rect 474118 26593 479813 26829
rect 480049 26593 495952 26829
rect 496188 26593 501882 26829
rect 502118 26593 507813 26829
rect 508049 26593 523952 26829
rect 524188 26593 529882 26829
rect 530118 26593 535813 26829
rect 536049 26593 551952 26829
rect 552188 26593 557882 26829
rect 558118 26593 563813 26829
rect 564049 26593 573526 26829
rect 573762 26593 573846 26829
rect 574082 26593 585342 26829
rect 585578 26593 585662 26829
rect 585898 26593 592650 26829
rect -8726 26509 592650 26593
rect -8726 26273 -1974 26509
rect -1738 26273 -1654 26509
rect -1418 26273 22460 26509
rect 22696 26273 33408 26509
rect 33644 26273 44356 26509
rect 44592 26273 55304 26509
rect 55540 26273 75952 26509
rect 76188 26273 81882 26509
rect 82118 26273 87813 26509
rect 88049 26273 103952 26509
rect 104188 26273 109882 26509
rect 110118 26273 115813 26509
rect 116049 26273 131952 26509
rect 132188 26273 137882 26509
rect 138118 26273 143813 26509
rect 144049 26273 159952 26509
rect 160188 26273 165882 26509
rect 166118 26273 171813 26509
rect 172049 26273 187952 26509
rect 188188 26273 193882 26509
rect 194118 26273 199813 26509
rect 200049 26273 215952 26509
rect 216188 26273 221882 26509
rect 222118 26273 227813 26509
rect 228049 26273 243952 26509
rect 244188 26273 249882 26509
rect 250118 26273 255813 26509
rect 256049 26273 271952 26509
rect 272188 26273 277882 26509
rect 278118 26273 283813 26509
rect 284049 26273 299952 26509
rect 300188 26273 305882 26509
rect 306118 26273 311813 26509
rect 312049 26273 327952 26509
rect 328188 26273 333882 26509
rect 334118 26273 339813 26509
rect 340049 26273 355952 26509
rect 356188 26273 361882 26509
rect 362118 26273 367813 26509
rect 368049 26273 383952 26509
rect 384188 26273 389882 26509
rect 390118 26273 395813 26509
rect 396049 26273 411952 26509
rect 412188 26273 417882 26509
rect 418118 26273 423813 26509
rect 424049 26273 439952 26509
rect 440188 26273 445882 26509
rect 446118 26273 451813 26509
rect 452049 26273 467952 26509
rect 468188 26273 473882 26509
rect 474118 26273 479813 26509
rect 480049 26273 495952 26509
rect 496188 26273 501882 26509
rect 502118 26273 507813 26509
rect 508049 26273 523952 26509
rect 524188 26273 529882 26509
rect 530118 26273 535813 26509
rect 536049 26273 551952 26509
rect 552188 26273 557882 26509
rect 558118 26273 563813 26509
rect 564049 26273 573526 26509
rect 573762 26273 573846 26509
rect 574082 26273 585342 26509
rect 585578 26273 585662 26509
rect 585898 26273 592650 26509
rect -8726 26241 592650 26273
rect -8726 23454 592650 23486
rect -8726 23218 -2934 23454
rect -2698 23218 -2614 23454
rect -2378 23218 27934 23454
rect 28170 23218 38882 23454
rect 39118 23218 49830 23454
rect 50066 23218 60778 23454
rect 61014 23218 66026 23454
rect 66262 23218 66346 23454
rect 66582 23218 78916 23454
rect 79152 23218 84847 23454
rect 85083 23218 106916 23454
rect 107152 23218 112847 23454
rect 113083 23218 134916 23454
rect 135152 23218 140847 23454
rect 141083 23218 162916 23454
rect 163152 23218 168847 23454
rect 169083 23218 190916 23454
rect 191152 23218 196847 23454
rect 197083 23218 218916 23454
rect 219152 23218 224847 23454
rect 225083 23218 246916 23454
rect 247152 23218 252847 23454
rect 253083 23218 274916 23454
rect 275152 23218 280847 23454
rect 281083 23218 302916 23454
rect 303152 23218 308847 23454
rect 309083 23218 330916 23454
rect 331152 23218 336847 23454
rect 337083 23218 358916 23454
rect 359152 23218 364847 23454
rect 365083 23218 386916 23454
rect 387152 23218 392847 23454
rect 393083 23218 414916 23454
rect 415152 23218 420847 23454
rect 421083 23218 442916 23454
rect 443152 23218 448847 23454
rect 449083 23218 470916 23454
rect 471152 23218 476847 23454
rect 477083 23218 498916 23454
rect 499152 23218 504847 23454
rect 505083 23218 526916 23454
rect 527152 23218 532847 23454
rect 533083 23218 554916 23454
rect 555152 23218 560847 23454
rect 561083 23218 586302 23454
rect 586538 23218 586622 23454
rect 586858 23218 592650 23454
rect -8726 23134 592650 23218
rect -8726 22898 -2934 23134
rect -2698 22898 -2614 23134
rect -2378 22898 27934 23134
rect 28170 22898 38882 23134
rect 39118 22898 49830 23134
rect 50066 22898 60778 23134
rect 61014 22898 66026 23134
rect 66262 22898 66346 23134
rect 66582 22898 78916 23134
rect 79152 22898 84847 23134
rect 85083 22898 106916 23134
rect 107152 22898 112847 23134
rect 113083 22898 134916 23134
rect 135152 22898 140847 23134
rect 141083 22898 162916 23134
rect 163152 22898 168847 23134
rect 169083 22898 190916 23134
rect 191152 22898 196847 23134
rect 197083 22898 218916 23134
rect 219152 22898 224847 23134
rect 225083 22898 246916 23134
rect 247152 22898 252847 23134
rect 253083 22898 274916 23134
rect 275152 22898 280847 23134
rect 281083 22898 302916 23134
rect 303152 22898 308847 23134
rect 309083 22898 330916 23134
rect 331152 22898 336847 23134
rect 337083 22898 358916 23134
rect 359152 22898 364847 23134
rect 365083 22898 386916 23134
rect 387152 22898 392847 23134
rect 393083 22898 414916 23134
rect 415152 22898 420847 23134
rect 421083 22898 442916 23134
rect 443152 22898 448847 23134
rect 449083 22898 470916 23134
rect 471152 22898 476847 23134
rect 477083 22898 498916 23134
rect 499152 22898 504847 23134
rect 505083 22898 526916 23134
rect 527152 22898 532847 23134
rect 533083 22898 554916 23134
rect 555152 22898 560847 23134
rect 561083 22898 586302 23134
rect 586538 22898 586622 23134
rect 586858 22898 592650 23134
rect -8726 22866 592650 22898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 573526 -346
rect 573762 -582 573846 -346
rect 574082 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 573526 -666
rect 573762 -902 573846 -666
rect 574082 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 66026 -1306
rect 66262 -1542 66346 -1306
rect 66582 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 66026 -1626
rect 66262 -1862 66346 -1626
rect 66582 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use scan_controller  scan_controller
timestamp 0
transform 1 0 16000 0 1 16000
box -10 0 46000 20000
use scan_wrapper_1f985e14df1ed789231bb6e0189d6e39  scan_wrapper_1f985e14df1ed789231bb6e0189d6e39_51
timestamp 0
transform 1 0 380000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_019235602376235615  scan_wrapper_019235602376235615_84
timestamp 0
transform 1 0 184000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_334445762078310996  scan_wrapper_334445762078310996_1
timestamp 0
transform 1 0 100000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_335404063203000914  scan_wrapper_335404063203000914_2
timestamp 0
transform 1 0 128000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339439899388150354  scan_wrapper_339439899388150354_3
timestamp 0
transform 1 0 156000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_0
timestamp 0
transform 1 0 72000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_102
timestamp 0
transform -1 0 456000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_103
timestamp 0
transform -1 0 428000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_104
timestamp 0
transform -1 0 400000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_105
timestamp 0
transform -1 0 372000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_106
timestamp 0
transform -1 0 344000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_107
timestamp 0
transform -1 0 316000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_108
timestamp 0
transform -1 0 288000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_109
timestamp 0
transform -1 0 260000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_110
timestamp 0
transform -1 0 232000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_111
timestamp 0
transform -1 0 204000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_112
timestamp 0
transform -1 0 176000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_113
timestamp 0
transform -1 0 148000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_114
timestamp 0
transform -1 0 120000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_115
timestamp 0
transform -1 0 92000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_116
timestamp 0
transform -1 0 64000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_117
timestamp 0
transform -1 0 36000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_118
timestamp 0
transform 1 0 16000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_119
timestamp 0
transform 1 0 44000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_120
timestamp 0
transform 1 0 72000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_121
timestamp 0
transform 1 0 100000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_122
timestamp 0
transform 1 0 128000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_123
timestamp 0
transform 1 0 156000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_124
timestamp 0
transform 1 0 184000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_125
timestamp 0
transform 1 0 212000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_126
timestamp 0
transform 1 0 240000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_127
timestamp 0
transform 1 0 268000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_128
timestamp 0
transform 1 0 296000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_129
timestamp 0
transform 1 0 324000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_130
timestamp 0
transform 1 0 352000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_131
timestamp 0
transform 1 0 380000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_132
timestamp 0
transform 1 0 408000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_133
timestamp 0
transform 1 0 436000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_134
timestamp 0
transform 1 0 464000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_135
timestamp 0
transform 1 0 492000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_136
timestamp 0
transform 1 0 520000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_137
timestamp 0
transform 1 0 548000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_138
timestamp 0
transform -1 0 568000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_139
timestamp 0
transform -1 0 540000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_140
timestamp 0
transform -1 0 512000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_141
timestamp 0
transform -1 0 484000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_142
timestamp 0
transform -1 0 456000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_143
timestamp 0
transform -1 0 428000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_144
timestamp 0
transform -1 0 400000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_145
timestamp 0
transform -1 0 372000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_146
timestamp 0
transform -1 0 344000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_147
timestamp 0
transform -1 0 316000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_148
timestamp 0
transform -1 0 288000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_149
timestamp 0
transform -1 0 260000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_150
timestamp 0
transform -1 0 232000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_151
timestamp 0
transform -1 0 204000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_152
timestamp 0
transform -1 0 176000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_153
timestamp 0
transform -1 0 148000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_154
timestamp 0
transform -1 0 120000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_155
timestamp 0
transform -1 0 92000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_156
timestamp 0
transform -1 0 64000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_157
timestamp 0
transform -1 0 36000 0 -1 225000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_158
timestamp 0
transform 1 0 16000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_159
timestamp 0
transform 1 0 44000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_160
timestamp 0
transform 1 0 72000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_161
timestamp 0
transform 1 0 100000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_162
timestamp 0
transform 1 0 128000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_163
timestamp 0
transform 1 0 156000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_164
timestamp 0
transform 1 0 184000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_165
timestamp 0
transform 1 0 212000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_166
timestamp 0
transform 1 0 240000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_167
timestamp 0
transform 1 0 268000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_168
timestamp 0
transform 1 0 296000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_169
timestamp 0
transform 1 0 324000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_170
timestamp 0
transform 1 0 352000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_171
timestamp 0
transform 1 0 380000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_172
timestamp 0
transform 1 0 408000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_173
timestamp 0
transform 1 0 436000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_174
timestamp 0
transform 1 0 464000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_175
timestamp 0
transform 1 0 492000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_176
timestamp 0
transform 1 0 520000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_177
timestamp 0
transform 1 0 548000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_178
timestamp 0
transform -1 0 568000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_179
timestamp 0
transform -1 0 540000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_180
timestamp 0
transform -1 0 512000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_181
timestamp 0
transform -1 0 484000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_182
timestamp 0
transform -1 0 456000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_183
timestamp 0
transform -1 0 428000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_184
timestamp 0
transform -1 0 400000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_185
timestamp 0
transform -1 0 372000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_186
timestamp 0
transform -1 0 344000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_187
timestamp 0
transform -1 0 316000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_188
timestamp 0
transform -1 0 288000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_189
timestamp 0
transform -1 0 260000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_190
timestamp 0
transform -1 0 232000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_191
timestamp 0
transform -1 0 204000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_192
timestamp 0
transform -1 0 176000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_193
timestamp 0
transform -1 0 148000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_194
timestamp 0
transform -1 0 120000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_195
timestamp 0
transform -1 0 92000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_196
timestamp 0
transform -1 0 64000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_197
timestamp 0
transform -1 0 36000 0 -1 279000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_198
timestamp 0
transform 1 0 16000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_199
timestamp 0
transform 1 0 44000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_200
timestamp 0
transform 1 0 72000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_201
timestamp 0
transform 1 0 100000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_202
timestamp 0
transform 1 0 128000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_203
timestamp 0
transform 1 0 156000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_204
timestamp 0
transform 1 0 184000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_205
timestamp 0
transform 1 0 212000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_206
timestamp 0
transform 1 0 240000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_207
timestamp 0
transform 1 0 268000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_208
timestamp 0
transform 1 0 296000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_209
timestamp 0
transform 1 0 324000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_210
timestamp 0
transform 1 0 352000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_211
timestamp 0
transform 1 0 380000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_212
timestamp 0
transform 1 0 408000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_213
timestamp 0
transform 1 0 436000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_214
timestamp 0
transform 1 0 464000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_215
timestamp 0
transform 1 0 492000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_216
timestamp 0
transform 1 0 520000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_217
timestamp 0
transform 1 0 548000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_218
timestamp 0
transform -1 0 568000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_219
timestamp 0
transform -1 0 540000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_220
timestamp 0
transform -1 0 512000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_221
timestamp 0
transform -1 0 484000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_222
timestamp 0
transform -1 0 456000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_223
timestamp 0
transform -1 0 428000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_224
timestamp 0
transform -1 0 400000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_225
timestamp 0
transform -1 0 372000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_226
timestamp 0
transform -1 0 344000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_227
timestamp 0
transform -1 0 316000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_228
timestamp 0
transform -1 0 288000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_229
timestamp 0
transform -1 0 260000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_230
timestamp 0
transform -1 0 232000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_231
timestamp 0
transform -1 0 204000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_232
timestamp 0
transform -1 0 176000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_233
timestamp 0
transform -1 0 148000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_234
timestamp 0
transform -1 0 120000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_235
timestamp 0
transform -1 0 92000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_236
timestamp 0
transform -1 0 64000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_237
timestamp 0
transform -1 0 36000 0 -1 333000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_238
timestamp 0
transform 1 0 16000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_239
timestamp 0
transform 1 0 44000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_240
timestamp 0
transform 1 0 72000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_241
timestamp 0
transform 1 0 100000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_242
timestamp 0
transform 1 0 128000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_243
timestamp 0
transform 1 0 156000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_244
timestamp 0
transform 1 0 184000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_245
timestamp 0
transform 1 0 212000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_246
timestamp 0
transform 1 0 240000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_247
timestamp 0
transform 1 0 268000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_248
timestamp 0
transform 1 0 296000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_249
timestamp 0
transform 1 0 324000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_250
timestamp 0
transform 1 0 352000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_251
timestamp 0
transform 1 0 380000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_252
timestamp 0
transform 1 0 408000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_253
timestamp 0
transform 1 0 436000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_254
timestamp 0
transform 1 0 464000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_255
timestamp 0
transform 1 0 492000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_256
timestamp 0
transform 1 0 520000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_257
timestamp 0
transform 1 0 548000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_258
timestamp 0
transform -1 0 568000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_259
timestamp 0
transform -1 0 540000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_260
timestamp 0
transform -1 0 512000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_261
timestamp 0
transform -1 0 484000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_262
timestamp 0
transform -1 0 456000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_263
timestamp 0
transform -1 0 428000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_264
timestamp 0
transform -1 0 400000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_265
timestamp 0
transform -1 0 372000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_266
timestamp 0
transform -1 0 344000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_267
timestamp 0
transform -1 0 316000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_268
timestamp 0
transform -1 0 288000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_269
timestamp 0
transform -1 0 260000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_270
timestamp 0
transform -1 0 232000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_271
timestamp 0
transform -1 0 204000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_272
timestamp 0
transform -1 0 176000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_273
timestamp 0
transform -1 0 148000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_274
timestamp 0
transform -1 0 120000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_275
timestamp 0
transform -1 0 92000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_276
timestamp 0
transform -1 0 64000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_277
timestamp 0
transform -1 0 36000 0 -1 387000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_278
timestamp 0
transform 1 0 16000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_279
timestamp 0
transform 1 0 44000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_280
timestamp 0
transform 1 0 72000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_281
timestamp 0
transform 1 0 100000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_282
timestamp 0
transform 1 0 128000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_283
timestamp 0
transform 1 0 156000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_284
timestamp 0
transform 1 0 184000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_285
timestamp 0
transform 1 0 212000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_286
timestamp 0
transform 1 0 240000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_287
timestamp 0
transform 1 0 268000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_288
timestamp 0
transform 1 0 296000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_289
timestamp 0
transform 1 0 324000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_290
timestamp 0
transform 1 0 352000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_291
timestamp 0
transform 1 0 380000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_292
timestamp 0
transform 1 0 408000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_293
timestamp 0
transform 1 0 436000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_294
timestamp 0
transform 1 0 464000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_295
timestamp 0
transform 1 0 492000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_296
timestamp 0
transform 1 0 520000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_297
timestamp 0
transform 1 0 548000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_298
timestamp 0
transform -1 0 568000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_299
timestamp 0
transform -1 0 540000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_300
timestamp 0
transform -1 0 512000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_301
timestamp 0
transform -1 0 484000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_302
timestamp 0
transform -1 0 456000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_303
timestamp 0
transform -1 0 428000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_304
timestamp 0
transform -1 0 400000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_305
timestamp 0
transform -1 0 372000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_306
timestamp 0
transform -1 0 344000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_307
timestamp 0
transform -1 0 316000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_308
timestamp 0
transform -1 0 288000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_309
timestamp 0
transform -1 0 260000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_310
timestamp 0
transform -1 0 232000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_311
timestamp 0
transform -1 0 204000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_312
timestamp 0
transform -1 0 176000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_313
timestamp 0
transform -1 0 148000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_314
timestamp 0
transform -1 0 120000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_315
timestamp 0
transform -1 0 92000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_316
timestamp 0
transform -1 0 64000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_317
timestamp 0
transform -1 0 36000 0 -1 441000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_318
timestamp 0
transform 1 0 16000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_319
timestamp 0
transform 1 0 44000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_320
timestamp 0
transform 1 0 72000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_321
timestamp 0
transform 1 0 100000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_322
timestamp 0
transform 1 0 128000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_323
timestamp 0
transform 1 0 156000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_324
timestamp 0
transform 1 0 184000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_325
timestamp 0
transform 1 0 212000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_326
timestamp 0
transform 1 0 240000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_327
timestamp 0
transform 1 0 268000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_328
timestamp 0
transform 1 0 296000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_329
timestamp 0
transform 1 0 324000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_330
timestamp 0
transform 1 0 352000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_331
timestamp 0
transform 1 0 380000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_332
timestamp 0
transform 1 0 408000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_333
timestamp 0
transform 1 0 436000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_334
timestamp 0
transform 1 0 464000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_335
timestamp 0
transform 1 0 492000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_336
timestamp 0
transform 1 0 520000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_337
timestamp 0
transform 1 0 548000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_338
timestamp 0
transform -1 0 568000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_339
timestamp 0
transform -1 0 540000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_340
timestamp 0
transform -1 0 512000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_341
timestamp 0
transform -1 0 484000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_342
timestamp 0
transform -1 0 456000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_343
timestamp 0
transform -1 0 428000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_344
timestamp 0
transform -1 0 400000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_345
timestamp 0
transform -1 0 372000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_346
timestamp 0
transform -1 0 344000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_347
timestamp 0
transform -1 0 316000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_348
timestamp 0
transform -1 0 288000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_349
timestamp 0
transform -1 0 260000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_350
timestamp 0
transform -1 0 232000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_351
timestamp 0
transform -1 0 204000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_352
timestamp 0
transform -1 0 176000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_353
timestamp 0
transform -1 0 148000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_354
timestamp 0
transform -1 0 120000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_355
timestamp 0
transform -1 0 92000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_356
timestamp 0
transform -1 0 64000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_357
timestamp 0
transform -1 0 36000 0 -1 495000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_358
timestamp 0
transform 1 0 16000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_359
timestamp 0
transform 1 0 44000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_360
timestamp 0
transform 1 0 72000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_361
timestamp 0
transform 1 0 100000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_362
timestamp 0
transform 1 0 128000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_363
timestamp 0
transform 1 0 156000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_364
timestamp 0
transform 1 0 184000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_365
timestamp 0
transform 1 0 212000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_366
timestamp 0
transform 1 0 240000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_367
timestamp 0
transform 1 0 268000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_368
timestamp 0
transform 1 0 296000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_369
timestamp 0
transform 1 0 324000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_370
timestamp 0
transform 1 0 352000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_371
timestamp 0
transform 1 0 380000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_372
timestamp 0
transform 1 0 408000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_373
timestamp 0
transform 1 0 436000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_374
timestamp 0
transform 1 0 464000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_375
timestamp 0
transform 1 0 492000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_376
timestamp 0
transform 1 0 520000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_377
timestamp 0
transform 1 0 548000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_378
timestamp 0
transform -1 0 568000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_379
timestamp 0
transform -1 0 540000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_380
timestamp 0
transform -1 0 512000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_381
timestamp 0
transform -1 0 484000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_382
timestamp 0
transform -1 0 456000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_383
timestamp 0
transform -1 0 428000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_384
timestamp 0
transform -1 0 400000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_385
timestamp 0
transform -1 0 372000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_386
timestamp 0
transform -1 0 344000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_387
timestamp 0
transform -1 0 316000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_388
timestamp 0
transform -1 0 288000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_389
timestamp 0
transform -1 0 260000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_390
timestamp 0
transform -1 0 232000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_391
timestamp 0
transform -1 0 204000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_392
timestamp 0
transform -1 0 176000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_393
timestamp 0
transform -1 0 148000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_394
timestamp 0
transform -1 0 120000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_395
timestamp 0
transform -1 0 92000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_396
timestamp 0
transform -1 0 64000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_397
timestamp 0
transform -1 0 36000 0 -1 549000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_398
timestamp 0
transform 1 0 16000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_399
timestamp 0
transform 1 0 44000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_400
timestamp 0
transform 1 0 72000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_401
timestamp 0
transform 1 0 100000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_402
timestamp 0
transform 1 0 128000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_403
timestamp 0
transform 1 0 156000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_404
timestamp 0
transform 1 0 184000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_405
timestamp 0
transform 1 0 212000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_406
timestamp 0
transform 1 0 240000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_407
timestamp 0
transform 1 0 268000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_408
timestamp 0
transform 1 0 296000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_409
timestamp 0
transform 1 0 324000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_410
timestamp 0
transform 1 0 352000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_411
timestamp 0
transform 1 0 380000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_412
timestamp 0
transform 1 0 408000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_413
timestamp 0
transform 1 0 436000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_414
timestamp 0
transform 1 0 464000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_415
timestamp 0
transform 1 0 492000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_416
timestamp 0
transform 1 0 520000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_417
timestamp 0
transform 1 0 548000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_418
timestamp 0
transform -1 0 568000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_419
timestamp 0
transform -1 0 540000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_420
timestamp 0
transform -1 0 512000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_421
timestamp 0
transform -1 0 484000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_422
timestamp 0
transform -1 0 456000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_423
timestamp 0
transform -1 0 428000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_424
timestamp 0
transform -1 0 400000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_425
timestamp 0
transform -1 0 372000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_426
timestamp 0
transform -1 0 344000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_427
timestamp 0
transform -1 0 316000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_428
timestamp 0
transform -1 0 288000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_429
timestamp 0
transform -1 0 260000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_430
timestamp 0
transform -1 0 232000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_431
timestamp 0
transform -1 0 204000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_432
timestamp 0
transform -1 0 176000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_433
timestamp 0
transform -1 0 148000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_434
timestamp 0
transform -1 0 120000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_435
timestamp 0
transform -1 0 92000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_436
timestamp 0
transform -1 0 64000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_437
timestamp 0
transform -1 0 36000 0 -1 603000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_438
timestamp 0
transform 1 0 16000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_439
timestamp 0
transform 1 0 44000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_440
timestamp 0
transform 1 0 72000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_441
timestamp 0
transform 1 0 100000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_442
timestamp 0
transform 1 0 128000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_443
timestamp 0
transform 1 0 156000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_444
timestamp 0
transform 1 0 184000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_445
timestamp 0
transform 1 0 212000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_446
timestamp 0
transform 1 0 240000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_447
timestamp 0
transform 1 0 268000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_448
timestamp 0
transform 1 0 296000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_449
timestamp 0
transform 1 0 324000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_450
timestamp 0
transform 1 0 352000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_451
timestamp 0
transform 1 0 380000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_452
timestamp 0
transform 1 0 408000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_453
timestamp 0
transform 1 0 436000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_454
timestamp 0
transform 1 0 464000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_455
timestamp 0
transform 1 0 492000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_456
timestamp 0
transform 1 0 520000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_457
timestamp 0
transform 1 0 548000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_458
timestamp 0
transform -1 0 568000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_459
timestamp 0
transform -1 0 540000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_460
timestamp 0
transform -1 0 512000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_461
timestamp 0
transform -1 0 484000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_462
timestamp 0
transform -1 0 456000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_463
timestamp 0
transform -1 0 428000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_464
timestamp 0
transform -1 0 400000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_465
timestamp 0
transform -1 0 372000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_466
timestamp 0
transform -1 0 344000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_467
timestamp 0
transform -1 0 316000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_468
timestamp 0
transform -1 0 288000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_469
timestamp 0
transform -1 0 260000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_470
timestamp 0
transform -1 0 232000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_471
timestamp 0
transform -1 0 204000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_472
timestamp 0
transform -1 0 176000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_473
timestamp 0
transform -1 0 148000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_474
timestamp 0
transform -1 0 120000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_475
timestamp 0
transform -1 0 92000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_476
timestamp 0
transform -1 0 64000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_477
timestamp 0
transform -1 0 36000 0 -1 657000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_478
timestamp 0
transform 1 0 16000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_479
timestamp 0
transform 1 0 44000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_480
timestamp 0
transform 1 0 72000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_481
timestamp 0
transform 1 0 100000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_482
timestamp 0
transform 1 0 128000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_483
timestamp 0
transform 1 0 156000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_484
timestamp 0
transform 1 0 184000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_485
timestamp 0
transform 1 0 212000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_486
timestamp 0
transform 1 0 240000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_487
timestamp 0
transform 1 0 268000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_488
timestamp 0
transform 1 0 296000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_489
timestamp 0
transform 1 0 324000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_490
timestamp 0
transform 1 0 352000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_491
timestamp 0
transform 1 0 380000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_492
timestamp 0
transform 1 0 408000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_493
timestamp 0
transform 1 0 436000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_494
timestamp 0
transform 1 0 464000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_495
timestamp 0
transform 1 0 492000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_496
timestamp 0
transform 1 0 520000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_497
timestamp 0
transform 1 0 548000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339502597164499540  scan_wrapper_339502597164499540_4
timestamp 0
transform 1 0 184000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339732875283792466  scan_wrapper_339732875283792466_5
timestamp 0
transform 1 0 212000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339800239192932947  scan_wrapper_339800239192932947_14
timestamp 0
transform 1 0 464000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339865743461974612  scan_wrapper_339865743461974612_6
timestamp 0
transform 1 0 240000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339898704941023827  scan_wrapper_339898704941023827_7
timestamp 0
transform 1 0 268000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_340218629792465491  scan_wrapper_340218629792465491_8
timestamp 0
transform 1 0 296000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_340285391309374034  scan_wrapper_340285391309374034_10
timestamp 0
transform 1 0 352000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_340318610245288530  scan_wrapper_340318610245288530_9
timestamp 0
transform 1 0 324000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_340579111348994642  scan_wrapper_340579111348994642_37
timestamp 0
transform -1 0 36000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_340661930553246290  scan_wrapper_340661930553246290_11
timestamp 0
transform 1 0 380000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_340805072482992722  scan_wrapper_340805072482992722_12
timestamp 0
transform 1 0 408000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_341063825089364563  scan_wrapper_341063825089364563_75
timestamp 0
transform -1 0 92000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341136771628663380  scan_wrapper_341136771628663380_13
timestamp 0
transform 1 0 436000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_341152580068442706  scan_wrapper_341152580068442706_22
timestamp 0
transform -1 0 456000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341154068332282450  scan_wrapper_341154068332282450_17
timestamp 0
transform 1 0 548000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_341154161238213203  scan_wrapper_341154161238213203_15
timestamp 0
transform 1 0 492000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_341155178824598098  scan_wrapper_341155178824598098_23
timestamp 0
transform -1 0 428000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341159915403870803  scan_wrapper_341159915403870803_16
timestamp 0
transform 1 0 520000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_341160201697624660  scan_wrapper_341160201697624660_18
timestamp 0
transform -1 0 568000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341160271679586899  scan_wrapper_341160271679586899_20
timestamp 0
transform -1 0 512000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341161378978988626  scan_wrapper_341161378978988626_21
timestamp 0
transform -1 0 484000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341162950004834900  scan_wrapper_341162950004834900_32
timestamp 0
transform -1 0 176000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341163800289870419  scan_wrapper_341163800289870419_19
timestamp 0
transform -1 0 540000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341164228775772755  scan_wrapper_341164228775772755_45
timestamp 0
transform 1 0 212000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341164910646919762  scan_wrapper_341164910646919762_41
timestamp 0
transform 1 0 100000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341167691532337747  scan_wrapper_341167691532337747_24
timestamp 0
transform -1 0 400000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341174480471589458  scan_wrapper_341174480471589458_76
timestamp 0
transform -1 0 64000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341174563322724948  scan_wrapper_341174563322724948_47
timestamp 0
transform 1 0 268000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341176884318437971  scan_wrapper_341176884318437971_27
timestamp 0
transform -1 0 316000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341178154799333971  scan_wrapper_341178154799333971_25
timestamp 0
transform -1 0 372000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341178296293130834  scan_wrapper_341178296293130834_50
timestamp 0
transform 1 0 352000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341178481588044372  scan_wrapper_341178481588044372_26
timestamp 0
transform -1 0 344000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341182944314917460  scan_wrapper_341182944314917460_28
timestamp 0
transform -1 0 288000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341188777753969234  scan_wrapper_341188777753969234_29
timestamp 0
transform -1 0 260000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341191836498395731  scan_wrapper_341191836498395731_34
timestamp 0
transform -1 0 120000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341192113929585235  scan_wrapper_341192113929585235_35
timestamp 0
transform -1 0 92000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341192621088047698  scan_wrapper_341192621088047698_36
timestamp 0
transform -1 0 64000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341193419111006803  scan_wrapper_341193419111006803_63
timestamp 0
transform -1 0 428000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341194143598379604  scan_wrapper_341194143598379604_30
timestamp 0
transform -1 0 232000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341202178192441940  scan_wrapper_341202178192441940_33
timestamp 0
transform -1 0 148000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341205508016833108  scan_wrapper_341205508016833108_31
timestamp 0
transform -1 0 204000 0 -1 63000
box 0 0 20000 20000
use scan_wrapper_341224613878956628  scan_wrapper_341224613878956628_38
timestamp 0
transform 1 0 16000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341233739099013714  scan_wrapper_341233739099013714_42
timestamp 0
transform 1 0 128000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341235575572922964  scan_wrapper_341235575572922964_40
timestamp 0
transform 1 0 72000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341235973870322258  scan_wrapper_341235973870322258_39
timestamp 0
transform 1 0 44000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341240110454407762  scan_wrapper_341240110454407762_43
timestamp 0
transform 1 0 156000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341259651269001812  scan_wrapper_341259651269001812_60
timestamp 0
transform -1 0 512000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341262321634509394  scan_wrapper_341262321634509394_46
timestamp 0
transform 1 0 240000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341263346544149074  scan_wrapper_341263346544149074_53
timestamp 0
transform 1 0 436000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341264068701586004  scan_wrapper_341264068701586004_44
timestamp 0
transform 1 0 184000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341266732010177108  scan_wrapper_341266732010177108_64
timestamp 0
transform -1 0 400000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341271902949474898  scan_wrapper_341271902949474898_48
timestamp 0
transform 1 0 296000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341277789473735250  scan_wrapper_341277789473735250_52
timestamp 0
transform 1 0 408000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341279123277087315  scan_wrapper_341279123277087315_69
timestamp 0
transform -1 0 260000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341296149788885588  scan_wrapper_341296149788885588_54
timestamp 0
transform 1 0 464000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341315210433266259  scan_wrapper_341315210433266259_67
timestamp 0
transform -1 0 316000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341332847867462227  scan_wrapper_341332847867462227_55
timestamp 0
transform 1 0 492000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341337976625693266  scan_wrapper_341337976625693266_56
timestamp 0
transform 1 0 520000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341339883600609876  scan_wrapper_341339883600609876_57
timestamp 0
transform 1 0 548000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_341342096033055316  scan_wrapper_341342096033055316_59
timestamp 0
transform -1 0 540000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341344337258349139  scan_wrapper_341344337258349139_58
timestamp 0
transform -1 0 568000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341353777861755476  scan_wrapper_341353777861755476_65
timestamp 0
transform -1 0 372000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341353780122485332  scan_wrapper_341353780122485332_62
timestamp 0
transform -1 0 456000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341353928049295956  scan_wrapper_341353928049295956_61
timestamp 0
transform -1 0 484000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341359304823013970  scan_wrapper_341359304823013970_70
timestamp 0
transform -1 0 232000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341359404107432531  scan_wrapper_341359404107432531_66
timestamp 0
transform -1 0 344000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341364381657858642  scan_wrapper_341364381657858642_68
timestamp 0
transform -1 0 288000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341382703379120723  scan_wrapper_341382703379120723_71
timestamp 0
transform -1 0 204000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341389786199622227  scan_wrapper_341389786199622227_72
timestamp 0
transform -1 0 176000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341399568412312147  scan_wrapper_341399568412312147_89
timestamp 0
transform 1 0 324000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341404507891040852  scan_wrapper_341404507891040852_73
timestamp 0
transform -1 0 148000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341410909669818963  scan_wrapper_341410909669818963_74
timestamp 0
transform -1 0 120000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341419328215712339  scan_wrapper_341419328215712339_77
timestamp 0
transform -1 0 36000 0 -1 117000
box 0 0 20000 20000
use scan_wrapper_341431339142087251  scan_wrapper_341431339142087251_78
timestamp 0
transform 1 0 16000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341432030163108435  scan_wrapper_341432030163108435_79
timestamp 0
transform 1 0 44000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341432284947153491  scan_wrapper_341432284947153491_87
timestamp 0
transform 1 0 268000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341438392303616596  scan_wrapper_341438392303616596_86
timestamp 0
transform 1 0 240000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341440114308678227  scan_wrapper_341440114308678227_80
timestamp 0
transform 1 0 72000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341440781874102868  scan_wrapper_341440781874102868_82
timestamp 0
transform 1 0 128000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341444501414347346  scan_wrapper_341444501414347346_83
timestamp 0
transform 1 0 156000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341449297858921043  scan_wrapper_341449297858921043_101
timestamp 0
transform -1 0 484000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_341450853309219412  scan_wrapper_341450853309219412_85
timestamp 0
transform 1 0 212000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341452019534398035  scan_wrapper_341452019534398035_93
timestamp 0
transform 1 0 436000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341457971277988435  scan_wrapper_341457971277988435_88
timestamp 0
transform 1 0 296000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341464767397888596  scan_wrapper_341464767397888596_90
timestamp 0
transform 1 0 352000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341476989274686036  scan_wrapper_341476989274686036_91
timestamp 0
transform 1 0 380000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341482086419399252  scan_wrapper_341482086419399252_92
timestamp 0
transform 1 0 408000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341493393195532884  scan_wrapper_341493393195532884_99
timestamp 0
transform -1 0 540000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_341496918381167187  scan_wrapper_341496918381167187_81
timestamp 0
transform 1 0 100000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341497938559631956  scan_wrapper_341497938559631956_96
timestamp 0
transform 1 0 520000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341497964482527828  scan_wrapper_341497964482527828_95
timestamp 0
transform 1 0 492000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341497971083313748  scan_wrapper_341497971083313748_94
timestamp 0
transform 1 0 464000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341499976001520211  scan_wrapper_341499976001520211_97
timestamp 0
transform 1 0 548000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_341500800901579348  scan_wrapper_341500800901579348_98
timestamp 0
transform -1 0 568000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_341506274933867090  scan_wrapper_341506274933867090_100
timestamp 0
transform -1 0 512000 0 -1 171000
box 0 0 20000 20000
use scan_wrapper_bc4d7220e4fdbf20a574d56ea112a8e1  scan_wrapper_bc4d7220e4fdbf20a574d56ea112a8e1_49
timestamp 0
transform 1 0 324000 0 1 70000
box 0 0 20000 20000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 41494 686000 42114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 69494 686000 70114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 97494 686000 98114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 125494 686000 126114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 153494 686000 154114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181494 686000 182114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 209494 686000 210114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 237494 686000 238114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 265494 686000 266114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 293494 686000 294114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 321494 686000 322114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 349494 686000 350114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 377494 686000 378114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 405494 686000 406114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433494 686000 434114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 461494 686000 462114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 489494 686000 490114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 517494 686000 518114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 545494 686000 546114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 573494 -7654 574114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 26241 592650 26861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 53241 592650 53861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 80241 592650 80861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 107241 592650 107861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 134241 592650 134861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 161241 592650 161861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 188241 592650 188861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 215241 592650 215861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 242241 592650 242861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 269241 592650 269861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 296241 592650 296861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 323241 592650 323861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 350241 592650 350861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 377241 592650 377861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 404241 592650 404861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 431241 592650 431861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 458241 592650 458861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 485241 592650 485861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 512241 592650 512861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 539241 592650 539861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 566241 592650 566861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 593241 592650 593861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 620241 592650 620861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 647241 592650 647861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 674241 592650 674861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 701241 592650 701861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 37994 686000 38614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 65994 -7654 66614 41000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 65994 686000 66614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 93994 686000 94614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 121994 686000 122614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149994 686000 150614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 177994 686000 178614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 205994 686000 206614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 233994 686000 234614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 261994 686000 262614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 289994 686000 290614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 317994 686000 318614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 345994 686000 346614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 373994 686000 374614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401994 686000 402614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 429994 686000 430614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 457994 686000 458614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 485994 686000 486614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 513994 686000 514614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 541994 686000 542614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 569994 686000 570614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 22866 592650 23486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 49866 592650 50486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 76866 592650 77486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 103866 592650 104486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 130866 592650 131486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 157866 592650 158486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 184866 592650 185486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 211866 592650 212486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 238866 592650 239486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 265866 592650 266486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 292866 592650 293486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 319866 592650 320486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 346866 592650 347486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 373866 592650 374486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 400866 592650 401486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 427866 592650 428486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 454866 592650 455486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 481866 592650 482486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 508866 592650 509486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 535866 592650 536486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 562866 592650 563486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 589866 592650 590486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 616866 592650 617486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 643866 592650 644486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 670866 592650 671486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 697866 592650 698486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
