VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO scan_wrapper_341528610027340372
  CLASS BLOCK ;
  FOREIGN scan_wrapper_341528610027340372 ;
  ORIGIN 0.000 0.000 ;
  SIZE 105.000 BY 105.000 ;
  PIN clk_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 101.000 103.410 105.000 ;
    END
  END clk_in
  PIN clk_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END clk_out
  PIN data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.000 51.040 105.000 51.640 ;
    END
  END data_in
  PIN data_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END data_out
  PIN latch_enable_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END latch_enable_in
  PIN latch_enable_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 101.000 0.370 105.000 ;
    END
  END latch_enable_out
  PIN scan_select_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 101.000 51.890 105.000 ;
    END
  END scan_select_in
  PIN scan_select_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END scan_select_out
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 16.465 5.200 18.065 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.955 5.200 41.555 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.445 5.200 65.045 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 86.935 5.200 88.535 98.160 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 28.210 5.200 29.810 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.700 5.200 53.300 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.190 5.200 76.790 98.160 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 99.360 98.005 ;
      LAYER met1 ;
        RECT 0.070 3.440 103.430 98.160 ;
      LAYER met2 ;
        RECT 0.650 100.720 51.330 101.730 ;
        RECT 52.170 100.720 102.850 101.730 ;
        RECT 0.100 4.280 103.410 100.720 ;
        RECT 0.650 3.410 51.330 4.280 ;
        RECT 52.170 3.410 102.850 4.280 ;
      LAYER met3 ;
        RECT 4.000 52.040 103.435 98.085 ;
        RECT 4.400 50.640 100.600 52.040 ;
        RECT 4.000 4.255 103.435 50.640 ;
      LAYER met4 ;
        RECT 14.095 4.800 16.065 90.265 ;
        RECT 18.465 4.800 27.810 90.265 ;
        RECT 30.210 4.800 39.555 90.265 ;
        RECT 41.955 4.800 51.300 90.265 ;
        RECT 53.700 4.800 63.045 90.265 ;
        RECT 65.445 4.800 74.790 90.265 ;
        RECT 77.190 4.800 86.535 90.265 ;
        RECT 88.935 4.800 93.545 90.265 ;
        RECT 14.095 4.255 93.545 4.800 ;
  END
END scan_wrapper_341528610027340372
END LIBRARY

