/* Automatically generated from https://wokwi.com/projects/340596276030603858 */

`default_nettype none

module user_module_340596276030603858(
  input [7:0] io_in,
  output [7:0] io_out
);
  wire net1 = io_in[0];
  wire net2;
  wire net3 = 1'b1;
  wire net4 = 1'b1;
  wire net5 = 1'b0;
  wire net6 = 1'b0;
  wire net7 = 1'b0;
  wire net8 = 1'b0;
  wire net9 = 1'b0;
  wire net10 = 1'b0;
  wire net11 = 1'b0;
  wire net12 = 1'b0;
  wire net13 = 1'b0;
  wire net14 = 1'b0;
  wire net15 = 1'b0;
  wire net16 = 1'b0;
  wire net17 = 1'b0;
  wire net18 = 1'b0;
  wire net19 = 1'b0;
  wire net20 = 1'b0;
  wire net21 = 1'b0;
  wire net22 = 1'b0;
  wire net23 = 1'b0;
  wire net24 = 1'b0;
  wire net25 = 1'b0;
  wire net26 = 1'b0;
  wire net27 = 1'b0;
  wire net28 = 1'b0;
  wire net29 = 1'b0;
  wire net30 = 1'b0;
  wire net31 = 1'b0;
  wire net32 = 1'b0;
  wire net33 = 1'b0;
  wire net34 = 1'b0;
  wire net35 = 1'b0;
  wire net36 = 1'b0;
  wire net37 = 1'b0;
  wire net38 = 1'b0;
  wire net39 = 1'b0;
  wire net40 = 1'b0;
  wire net41 = 1'b0;
  wire net42 = 1'b0;
  wire net43 = 1'b0;
  wire net44 = 1'b0;
  wire net45 = 1'b0;
  wire net46 = 1'b0;
  wire net47 = 1'b0;
  wire net48 = 1'b0;
  wire net49 = 1'b0;
  wire net50 = 1'b0;
  wire net51 = 1'b0;
  wire net52 = 1'b0;

  assign io_out[0] = net2;

  and_cell gate1 (

  );
  or_cell gate2 (

  );
  xor_cell gate3 (

  );
  nand_cell gate4 (

  );
  not_cell gate5 (

  );
  mux_cell mux1 (

  );
  dff_cell flipflop1 (

  );
  buffer_cell gate7 (
    .in (net1),
    .out (net2)
  );
endmodule
